`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ww1cFCaKpEaygJUT+P6Z2OD0uzJ4IJG8iyHDm5UNlVWbTWS9KXjZ9jEg11wJmlv8lA2AVebHxIas
7nZJsy/GjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gy0/aj7fr+HoqiF2MKC2DdMRffpsNgkz3LCA0LoXsy3oP+ExvEwYs55sO8KAxVdJaUPMOFr+w6Gi
VDRBmTTzMTTD1KvHQEhDppUtYnGyL/2qAWb6xHvmSHDtiAjlHews7qZ26fM0sYgNx48H6LSqgFd4
hai7P1C8/gEiLdaec30=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hi2M/LxF9qgAZzAUuc501Ws9I83yzxDz1ea90Q5QjM7jLsFrH4fLD2d0WWY2wDTdG0Ih+QNnE4S7
Oq9DybBH0zvBRUhAQoExlvdlIfU3Jr1YKpM3lLPQTLIhhCp1eQgIZljQtMN1p0u0HDYYsZO5DBeb
LZHGhmPHPWGqNQ/iLmQ+PQu0B5Cb+1VKyvK7Ipxjf6wKC/NZlztCmWzwV4WC+jY2wHB2IofyzZfo
xRBIRCIpTb+tTiKgZ9oAjPNYVjgXC51YW/c8ZhnzF0gIdh/tD6GDSX/DdrrBN7Oz/gtduYw5jR0b
WsJx7lVGCa/mgRPb2+p2mjuutW8gGGnh6+Yo4A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X16goI57idQ5Yk2jq4rj0BhsplRtdzoYr8oOU2lBTTonp1Nx4fK7AS7KgGuzY4UqvPTHmPTfD5ww
0YcXmh8hr2Hk6aIz+aWFV8C8XcReGDrBhi5Np0Vi5hozuTfEPpWuDV7kTmarku7FYKZbPt+lsAsd
f8+cIo7ySKaxPnzoHbw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RA9GWDJZOdw/NASVbYOgehelK35X4QCDpOGKLkbLHbvCU34C5eqCOlazH25KMTrAHxM2lx7+fAsw
HHb2ZWqK4pB4ww23gPcOsgxVCyXs7Dx/H6E84snPbj5EBFAp1p9GZJoguz0skOVQzCSeso4vwekP
kvLqf3Ypkz4/BbGmeIV5O3MvxWppwuIHCb+NDzDYU2x9uQ7mLUtu7pYCzPfN1FeLiv9ttZaXRuYJ
ADExpcAMpFzH3bwg6Tm6wL+J1DzA4jLGZxI9jxK+L6xNTv2NtONryX7sLla9heWPJCSHR4TT8ow3
t3QklA4V7oRFEhlMh0Nv7QVOAHjukKSZ99LumA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12224)
`protect data_block
2JEuFaTgqghMsv5lmjCzRKFTRu9v2Bd7cfnnEymmK1IpMPqqHVgKVztK8UcvkN/cLu6meLkuW+GH
jEF+IasLsTsQoEbARf7iGoWy/qxr/Wx8iI4qK11niwKvKRzj3E/VIfcoFWMI7lDjskoNrB5ON374
xdQdL472o5haNrGgEzQCs124gMoZrq6ZZftrvXJyyhHqGqmNNfQbG065CYcPsuRjXxzPltG3oMhc
7n7pQE9F5O4ObyVFgYrFINih1IyuB6ga3CPJSEZRwp7Gz0bxN4RD0DBaR3vYvY1rH6jZ2As9bin/
g6/KlClzLL3bvhOha2ngCLKgz2aoAANC43Twjb4fUWJ67PFDf2GPtEf59dWM3VNyuNrEeNe6RWUg
jka4zLQP0zq2qshsXJQrae9LVhJ6szrSUvDOQAh3oT71FeB64AQ8gVISX1rm+woNgvHGbSKs7xZf
PBP7RqvUiS4Qazz5d0rzABAgtg35m+4/CZ6RQcd47z/v1puoo1bufBQHx73LzMGG/DN8vhbupjYA
svOqcQGNx9OB6DME6JsCHZsBHo8aI3x/a4hZHf41FqOiqyaqmjWc01kpYmeBfvzsPKZWMH8M7/bG
yW9X25BJeqxtOyeqdcRvqyQnEJ1HoishcB0BOSUa962dUzLqSDDUdDro7UpBLfafda9cVDS4XLbm
KBEIap5yL/BmCyInRk1GLXl2U/fOjGvBxrsmA9KuYhWFit/kiTe4yo9xZu90CDWCZ4O0JQa5IakH
bRCIdyuVLencac1svpY+HOynAZbmYpFgsLKUfER0UtkHhrvwQ7EebR1z8kAQ1EHeldFLTzrMcqke
GaF/TPfoe1hb2nFKWdyS0UJkpZI+u3UnW5oLYEi1eWSEb3nIu+pkTEFdD+NDeWyY7ooOUR9ukmJm
FbtSPJr4T6aXNoinEPe0BAAIEDnTtaWnygXYxUt5gLl9phRG7BhKf9pyhQxRhLaXv3dJm2z45lLW
t6hFppEp0o2lMyyEpTM/ADdb9E+ayxn24/aQWI57RXRXBLOjy81zJZYHrFlidSASB0CCEh2yC/wD
B5QfMrAMUIkaEsNKImtGoCZhoi8ZWl8cpvru2dtFWL2NYOSGChXVJTDw17BXMZ674am/KW0FNbNP
xJonGVPbVitbkX8OeFaJ7KZX5GgfEjccrXZbGLNsP0i48kwWL7OWQypCFGyh1VQ9E0Yg2t5OHpYL
mKuBnaRvMEKcW+vzC9YTkSw60mNXw0Tl0isvGZcgjnuGOvJbYzI0+tfsZjZhGrCFJgM6QwFkeAvu
i4tS/IgIp787GWG2VrpX/MyW6cWBJqtSS/VXG7edf3OKHn5BfLoILWkwkk9Ik1789H0M3dUtdVMn
1EsbD2HOTkQk6/uautsCMvJBTVpCUjdrfSGm10rIekn8RRYiWLpqHDBfjnvAElxsKSbxxkCFVqFl
Mft8QaEj/EkXo6mGBJR9FYtzGNZzY+hhzmDWJqGoaPALQuc+pukUZKLL4n40E40FY9fsCWRAsEtM
qN3O0NDIsaM1HXeaauf+s+No3eEnO2Rudm7JzhcUIafeH3aUBdbjif2yF2UZ2EJN0FTrtWj+T2l2
12GgMu8Kxib/0k7j5O4mGOfzdQLJUxZo4238IEgYqwOKZf3h3Mvl6jPtm8Kmb9TyRN9VOB8FZhAH
qnlvlJjq7TBULq61wc4zX8w3vYQXzAQjbYfJs2PW5y128zGprRL9hgVSOk8wNlWYlCt2VyU0cNmj
IC99Lw7c/En1+MaIMxzN46bmVZ6mb/00DRpuhR71e/ftn9nScJH9ut38geM9O8DDLavAPieUxJe0
E6KZ6dCOhk1Lt/S3Ye4aF33bEjg8gU4uzNJrLXnQ2hTDKCnNvB4n6JUcEDddAmAHzO7g8nVnoqBv
GieMtNsNaHKW8Y/KgqLV40lIb/HhBFQYDGAy528P5P3x4pMBKJHFuMfECLIAvirUczzGvqdUl4pU
Z54PyKT786VbzcnvGYwMFI/kWZQv+Iawx2Apx7YN9+6sOt5M+mq4molUTM51M8lMRe/ZS/4qy2nQ
iEJKIJ9J98iay67K0oPLYSLRJ7k7XK2nieGWNwACIwUeiixO6c+M7rTyyL/Fo9gV9LUck+s/9qEV
7nxjIVHvKSd4FI6kY9ZmsC8FX+LQZuqVl6P3WZUGAOkANctWA0MlQhcIPP3mwcqkYxqbhEAEcl+e
/r1lkS2nauEBRuheNUJeSY94VadNTUaFmeXwKU8SoMx9qRthN1FBl9c0yaGg+xsoYm3IkKeoCcFS
M6qwZwDXr0tblku+s9TQzIsTOKBHOgDPtHD/5l+RwS5BdGmpv0WRGDl/iGgrQarDS4ppeAHT6G04
fgzhb+l1xDB7yI3iJAJpc/I2jhxBckOofhua1zkq3xRpXqW9C5I+AZdFoToFroEuhElQ+nypFMm/
yH7fXEmSn0GyvMTdMm4qjUW+BgK64+n0IxIfvOceUBBzsfGLjADkHJ97T2cFuOD12zrU/WZlfgQc
7S7Rf2Pa/r4AoaOOcEw/ar/bM5rQ93nnPYLFKWBR3qbafJg2nsEKJv/O7i2pep0Y6q2WbFz3qGtW
AjyKvaR2mZZAFSqcDgFnGbWiS5zoJhF/5UI9Mkq0QlYYhSpdeDQZ4cp5Hsu04U4/9KnIxKnBhKZy
xRBEKrnPKVrx671lTzk1qMEWln53vvJio+DlDDg4tAKUBobJ5uuP6ckVqUifxunxKS5+3EIl+1Ea
LTbMkxG1oURsA+nG4ltGqvUwmcgVWhi1/VgWQ81XSfIlcA5eywDsxSqDfQ82FTS9kT92IGC5g2V6
bE/qfyPjHz2LQyvDqsnYZzHn83zCrHNd1P09JW2UphjZ3oHDVWVBSlI4Y+OF2pOOZqHhk01mggr3
dsiMild7YMtQVsSQR5IzD28G6e9qiUxB+vzh1IN9dPsLzib1GGmDqX+/620Mr0Ct4Qk9/cnaxFyb
FJe3p6/jtAYiGl4SxB6eBeZRgxNZJmu9SpEub6KGUg5VmGP/zs4rMzHjSEIoA26NhxIvEqG6qlAE
AqH9xwqFbYSoAcV+PYRzdRp1ejspFQqVM35ha+gL8QfTrXIs1yTFBm6kwErEjZ+x/Rz2ruAfVZ7x
0gjfMoxsUEIIeoCXTtEvwcI5PDxtQ1YJ3DMqPu/t15pCTImClfarE1Uf+ziz0duVqyM0g/E2J1on
xA7H7k27YJHv6Crj7nzFuZkH2oBAFL2O3r4wxy2PKiedp5GGxkNW/ba7oV+bVcPx+0PdzKUT+ZB0
nk0zQTGn7EqoWyGXhD5u6ll4pCZWvpDC95SN+jNUpNOBQKCzuPxWDsdRTb/E1voL/Qgsfp8nczSu
msXmc1TcQtOaCqRHbvHno8pPvMmPcQzwho47NkbmRsfPfzeREffQTtMs8IkA+Nd6GrLHBntCljph
0fzTge5maQwRp3YgE+hBuPD9MMK7+b2vWRpMw+4lvq4uuCBFh/wwIO57v3wVTO0SEC/C4bQRl91w
crs/Db7l9XIaUt9M02gHfjhnCIZnDwDJl59/Y7ELKRKMcO8v3YrYJr7n/boIp6GXdNRE83IL7kpy
xR75zI+tgayiYax8hZUumSk6xWWeV7GjH5tQm3LBBaaCasMtZuplOtC1Ltv2FQ2i3Lq7LWcySj55
eTZeYrHe9Uaoqc0jWQ0kpD/hh55h9SYqyeyhx0JNXmlI2oSmpZmAgyY4N7CPMXprFbsHjtwn8jVQ
2uYTk8f/rQPM/nPUIY73uxHmPlgdzQbJ+pUd/H15fVVvKA3NIcnbn7nxLsWQiLj1jpn1vZ3bn+U4
RDTCVSVTUsBwj9BXdi8ZhZnlM7MrraI5N7zdMrqJALFTxci3lCofYx4Ev9remJc4XHPvXb2EpGz7
3LL/TlQ/btolbnnfkOogOtssXtC9zOMyPwOKsz/HyFMMD5kWOo4pSG3k0G9VbFCcaimZkS6tPcL4
SiebA3clwC0lsDGCIx4RRlP6UGn+AajHYiNRoBH0SegcQ6TgEvy7M4oW9umnPnEX/c8bUVN9siAu
hrHPUt8XKlxzVcfvjDx7JxMYxugytW1k3IbQeLPvOyWVwYIX61WkNLrXYeSLPoEVDOIVyOvr8ICD
JxCAH21tnN5UQUpxlC4Wr0VX9OWD6h5NmcYOMW85jaOzcEn9a+bsZC/ZrY/KTrl4RiOmkPKCjeux
dWiYI3/6QGCe+r7GQnMPKwYmFhr/8X1RE8cwDS+9N+g2rlnTvT/AANR/miy4pr9TD8Hc9YblupMq
Bd6ROKAL0S7mxrWfNDAIx68wxu5KRnyT0/n3yM/0IK/NL0to/jtqcviBRhSqJymnR46XO3iHz8j0
jIuDtmYoaTAiqpcw8vvKJOc9I+n1kjknqtrWTIpX4njiWGTDvQPnYEKyTXZOsIGV9dw6OKtIEdNm
yHZ5Wjwc2vAYinnzvVV0LLpWl5D2hXddc5DF9dqANHY1eR4V8a+IaYej9iMDaibS2Cxp20U87xzN
6RZm4hl8UXLquUzc4xNo/6oIc3MLRtaB/bzCgNMzQ6FD85RvSd1a6GLr8YyT5u4za7oMUrzf+q8D
FP/5QSkagQjVt/ALmCj+H9nHaUfzuHslBrKBu8FaZ3aNzB89dYPV9BrQDPVHuFkuOTQOcwS4t4k4
QVYx9f0a8PygKs5ukZGuC2/fDXAjIo0yM29rHQpOwS6gjthWelaHQC0iqbd2kR9JiGm3/3JC9D1r
IjxeCQbAlJxla7q76xmsdM4jOd5jTedZIM+M1/s7KT1OOd+z+DJ7F4NBWtxqNTbSr+cL2kh22P92
VnEaysY6k1aB8aCVu3ceOd9F+Q5ZurTJG4Fh81W4a/Ux6pH2Oq39ndCz5a25p9iYQEclYNDGH004
GCOxyAlqbGVI9xl1V4mSVPEWYAHcSccDXw12/fUCWrttQhA4X7Adxbsk9WTT7rZGdy8q2vylGOtj
WmkQ781bjetd0mju3xO+eQN5873X7Pd3QO8CzCr5XqfwEwEvd4sx2UcegSFkZzNe8Il4p5yu1rZU
oC/WzdtWWjRJzQNEbk8NntIL/OHzHpYrzBGILt1R16qbSYbRrDcppV2LN51D68juYFt13et8VEp3
AXp9Ce0Na+bD8bNQJUllWFgwnSAJNtWk7dTcnhpPsi3eeG6NbTwU/iMtGZBbH3K+eOGEWex5iZ32
resqIejV8FY9r41tHaHFGOYnB3KrLjDGQx2oOvl65HnLfxc5KL43YZdmr57vi+sY1FSjurcFmrdf
zVazPZhtMPSqWwOVFroKANXxUAOFLXKSXm6SnCA+mDPe4wlm7KIsJmKL4mWKavXM/uKFjGB14UOd
K12vp9KI11MBIwOmGjFpyuf/FH7spawbEMGkMewEMrCfsT9buvU/Y+6ER+hylWLcNDH0Rv2m7ZTt
cbprmgBh91o3r2aNos62er8Hd0juQ53aWJTtKgHrrh+Ijzv5BNEcv06XhyBFeSRhqa9ygawLfRXg
n/ggX6fBhvWcOhIKcegP9WQimXfHy4Wxij3UppSMXmRpkYi3PyJBPD7HnF2ekrOQxgxLzhvd7IR0
6Gw5mcHRnwHVD7vQZ2zOyhZcBsKRkQYXj4byueZ5hzKAeazkj9OqbtWvaXkaPIzEOu6RMqa8C8Gz
WCputgmb/mvSOL0rNum/H3SaFUniQmd9sxZ8Pbe6vFKbkn9B9yyJYDh8dyPe8h+maa1/B/CW2mru
pgQ+rzJZaaVyDwCthsDuDNsBdK1Vq+nwLQYFO2rRRP2Mvm+iSDFEDcWdbFHOIvGKlwH8M91pMO4Q
LxskPD7QGIH77bUA95mreWiYIaG+/b8XlijpA0aDNUa7Y5a8sNIUkYjZGNZk6zYjBwSdEurkXAPX
LK4Pk8epJg5DDj+g7xiHPzKJeT4q47085kzC/e3kNr1vzXP0WuyJ4U6lEylSH9NshABcxpPs2RkM
ykQZI7tQeXFbW/HdP+OSjSlrLcw8ffZ0hVb6NYsRh5RnKabk8JXGdJbrk7MLsLZECvvfopVtGEdb
pb+qQl1aCl5bBUzQB9iq7kP30+o00wYQIVK95zPBY/Kzjjpf6oU3pYWshZ7Dn7CjTV21rd3V3RsK
ilKlmW0MwMMBj3aZwmu5m0F45CvlDc+TJ7xPp8JFC7z6suDHluqsihdvM8E6UwPZmEn1bPg4zkGm
IUa9gY9xoTTo0motKO5dowklfVCeiLa7yQLg/BUvuEwF4/nuEECosf0cOkOf1ea65GGY8XAzGLmM
6TtRt9GdScb/EgF/VDusda4f7qNAcQ5FBlShrwytRVwjc24nxYDvFujMR69NV2TiP0JvX/lKPJTu
g1mLVJWRpZmoIwM2cpAyFfWTHdfTcjxs9nX1DSb5Ql2am6P73V5ieFhA7g1Tt+HNfO002kKUFU6U
k40RpFe33a08g3FRbikv0t/1i8uNCeTlrr2M96GikPQCyyW6CUqu02XENgQVT0XUQkKrLQVDFXpN
GwRVAsw9gW1bnoYK1tOW7EzUWpBmt4yVVDbQjLXTs4wvB41qldVR8Sq99lM+ybwh7DgbprBlSAGv
1/Nvz2qnQLc2mPFxc6LmF3+2rYNMrjTYCe3svYTM0N208gHhD+cYMagiJhB0HGGxaNC4xWWq5nOl
Vs0JR08vR0Z2cQB+hhDxcpPDcNAtZ59wcMQcnQVkUA6tdK2drm/tucqEDdZoX07m8aP3CO69qIuP
9vfQhLaH361WyBJNJiIIVmQO1RRSHEBtWV+Jshk3l/JpkzQW9zZFMurh/uR9BbjTjGM6COtW57So
ukdLYKSUWWrt2R5b4AWrnaTQILrUMXDYA+c5RMOFbXp+kOBqpGAVninba8MymlN09SZ9UNL5BUMM
NWDs0/ppYgSiyVBo88fuPmkvAlVmg1ghgCkOHi+Zr5rtolWGEGfTYq3pyn+IgxulsD+/q7w57NRQ
eZrDQ32Vyre12tamY/Km8/vUe+LQ4+6+ONWtnwl0xtAOK5KA8KMSEEj2snUfQkYXuEBis2+TrDWY
CTAHqb6x+/ZrIRNMFUYZ5NCDZzvafXt98Un/8DcaK/TtUBBvcGL9Kf8nHmhTDZ1m3SlNLP12KBfX
VtWOg3aSf/blNaAq+RybdBDb0M4k4kx93SyDO9AI+qBff1MITDTqwTk3URX3Fbu+MfJ2WiUY1ORs
sTo4Bc7tX9Sl9YM2NepF8CQLOPgXAyD1g1alVr86t4bSG73GjyiVO+Lcp3/71zfdUdQZySyBR4x5
87i25Su1CrNCZHpp6Xffpcoeo/eNLVleeeySTStvE93fZlDB5Rha4VinSkI4LkfZyz/+4jrJ1RaO
gnSm8U48LILXc2DtMwC7cyW+8RYbf/wUXgw5iHwxyrNjIAfn9pI1Q4lSAkStDDJRnfi6p3bPEbdc
rEqpnUhW334hiK231285x81NmsXz4YT7C12tZJO/SHO0PP0LuLZv0Ee92k+hmn3AwveeVMz2Pvag
QMp3rpumxMqW6HEL2nM74MNheVbfI1jj1yOlCYpA0DePaIdB59zV3aokMqyq/YNoTRVkZJx7glPi
NA4/aez+giLxGvY8TxVVu+faeQCghzUMm8k+5oJlNNw1NTh19fkBmwf6Way7/saZhc2CGh5ggiwN
x2qswiI+m7vm/klEeR/rDW3OdLHOqi8WZUmHEuD3U9B837eGVLXa2wJsu0bIlmLOQna68uwr+Fp3
yh7x6qO/Hf0bQyidXoSopyt2EHJsPMNeJ2L3sZGTmTR87J1hA9u9ShVNvxPpupAMwqO0ytnuzGTy
aZSm2KUf2kzvykA1yBmHnPnWvaIzmHSMpmjM3+ydDoqATxhsKwyBxr7OtFOdyzU0Of2abbJCrgKx
8nmpetf+K742cnyCsJSfSHjfWdr6ZYFdGdayS7MqCCaA6McUqYRbkyNjTIKadyKMV/ovqqJXwmz5
u/+xpXENtfJ57TyL1KJ6lreCX6t13yncoiggB4gsR9Zsn9cEsi4V41oMATs8u1bTBRUeX2DjVulI
ZvaojP3VeA6U0/gWzzqX6XjSoR5t2+68LrJVFUCdELgQGwpO8zuhHikImd6V9lkD3Y8K1UwnySSu
ICUKzmAhW6ZAJM+nDUCRFYmOFA0ksgkbri5E1Q6IjFgv3rIj/N0Sdy9n9xPRI5nU7gAvTLvPrW0g
ekCxIhHtmNdkZE2aNUeh/BB2EXnHG/AQVHUcWT/ON0tR6idBDXOsfKfwNG0QUZrb4VTEeeHpNdaJ
L/Z3Y6qR3EjA6e0APDaOXA8YfcmzhqLOxI2U/mlE+54bbxbcFUOLul8QflpHo6zSJWOSIVOY/jc6
XCayjd960hu3QaK+1IARdd+/x9FbVBCWEgPkj1d5471X62arW1fgH8pQ1Mc6tQKYY72SufkdbxFE
1Ic7YebOhGeE+abk4lk76a2lXFk6/VRhvQG3WM0wll1fDXbPW0YI2WFdxsTxJdqYsDJkrQyB8KkU
JlyM6RLJSprC+pxF9tvUhpUC047IbQ6DDMWp+uapvnSRn/kx5ym+JsktK2DxX63ja20qqrWHJipe
4/+BzJHn17rcYUscxurxOn8bigmLNHuZAlOs7IpxO7vucUneNl3QknMia+3MXKA81UQcGuUAVjJi
8dtlhdjn6UzSmDomrJ/ITsr9KG7MSJN7tNqZ9pytsfvHNDGEAJ+orTdi6CL4GXFZhoBoc3bOxEEH
2WIYPkVpxPnJ8cE8llEsdfdINuinHEIwLfR+JBBHgPyz/IPoT+mjuUVcCQrPYjvqrIFwQzk4L0hC
EmRdGrDFyccPybivw7LLrEmerYDS3YgSVDBx4rpOtX5h3aTdUKcuryr6kQBgnbQ4Gl3SciegUmBF
TXVcJJWXsrEduZIOPpluoOEGMVozu354JlEUrlgNEJuXN3s0us3tIwIiPH8xKhAUM5bY+qS+Q/sL
5EKmRpKniMTmoUo2woQbccQAjgo5yFdGcTx5yQtNIhUHNaCzMxUawh11imwZ4Gww4H//02kKY7Yn
eD1OVXMXUuIooI725cTOvtPfZkr9+ALKt/qZcPlRHbUTpWelGiH9uc1kz1iUEwYyLlUn0bmOxPsJ
GOoIglAMd3auYSVzAyIN3rXx1P7lxgPj32OcZiQTkYo45EvJ1qyzXsNQoanrWKUNJQ29shmMlMD7
2CDJcG4UEr6d62CIwboHeEtS8bQUXrlD+OAvrX+4Zu4pk7oiduPH/hWSUjBv/UPS2V/4xVy22OZo
UAa9lRZdFCRnprvvTmg3QUZ5JSGIOiy/jAln5rRJYmBDXtAHl3mPmA/gOra17qH6snh6JHsIniAO
RvL+o4JUPDsJegxfe/OJqaOe+9ZhnEx6z3P6wi9sYEJjiDRiGkUL9pL0wLIjUs/tAFGW9GbFuysJ
rEDRRbSz/PEzi3h3yk7oGLL6sS7Bdzi3KR52UbJWwMGW94MYXqCJH4QN4vOZQqhFlM/HWkgCbqtb
Pj1GG2kNeNgH37xdR7WzA4fbRKspqcVdCK+FziI0FhxhGyh2xB59AwDceZiqyKRX9uAUedm0JmbN
HGDsA18UhcNbM4hOUC54iqJZ2aYAvvxTzg3+MmqsbWgql8PvAYE9FAGMKTW5lV8U+VUMAg2gAa4X
46uVWgeL9sE+6E8LG3Ad2nafHL+rOjQte+FCZOv1XMHt/MFR+nxJuZojinSOKSLc9oTihz4McvyG
Y0hu/tSb3I3Fjr24+VOFvVyAdVKtdla5bh5gLHsTBY75BY3iJVwzoWZ8rK9U+G58QzQ0UqMDjwss
VFGJ/ows2ldrjcy1SuhvEggLrqla8+yzkVoVAGZyXwUAaJMyNN2NylCxb0JTQjnHopHX719xP/wQ
R2c1qx5Xp3ILoEdBLxnGT0+RRxOOGFmPsr3B9TC/dIqTpqH2Qc9dULS1k3pPalspnEds33oekY0E
7wD7rrD8GFRAWMqUerpojwbaowXeM7Vncaba2eYxVJvc+moBPcgAvtnbWQf06LqJ2/7cUgXOzWmi
2nbs2hsENhwDW4UYL/Q5eIQiZ7iPQv1TMC5X3U9ttuY6jVoqXnxb2WVNyN4K2bgxaE0hGKttAOIl
skMgr4ZnwEzNmwZXI/v6A0y7EeDb7YnivLT4/KHuv4OmPAlshL3lku8ifv70TnfzKjYxzKuRA1Tj
KgiwUsUPe6ljgOBaooZ1dx6OTOgyKMLtw+p4/fWQCW1f0CgX2IcsQTUw1RVGOPxEj9dAkzxD0dyW
0fkSbHiuXmXz65KxwiPaJ6RNWbMMrKsMN9gi6PhfLd/fypnmSAtlHmx7Tcsv7iPrBrMqHPajlU+y
WzbK+7AAgOSJ9eG9/W91X4RAD+E3/Le0ReYlRd16/NzUB6bo7hNnux9oEocS2FpDjXUHZhnLvQf4
5OK2vpwNk+tRaQkyHeKGHStmPLUzbEEwH5AeGkzU/FIF6PzEOxymxK+q5NQNO22L8zs/0zf+vaHl
K9isUIS+8/SSEfQyEYWooh5/jpqejlLCxjOP5/lHLxHwVZ/G62wuIW3QDz6eK2ETQ5cNXqKTHIE1
VU8uOhKhpd/xlfg0IsG1yrxDWLmRaxmEw5m9mkeFZe7bVHtJsFu4c/5AEDvVTH9rfFTRxlE9NBx8
kLVAMxwyxUbgoA3omTt6GD22mTHh2GUSApOwacOGWvMlQ46xYxenncuWahrnB1NgCsTBiwqWu3QT
aa1jSD7aYNfQRHpax/OTfqwdAVQQyhZV4UDb56KGhERAEpjuhFztnQ8COP5x2vl70nSbOquubErg
Kdclkeg8921Z8kUtyp7CuM1SlWnyApe/J128d8HYzKte/IOyWTIL7QAVkGtjG97M/J66Bvfhjtz9
CgnA48wEBlumcV93puhSj6/M5t8/0MvN74Ieaa1kyx2rjMUGUp2oeN0KR+9n8bDE0wuqZeW36M+V
u6EGKxH6n7UcstGZF5sUwnUXDf9M1GfLhhAlVRBqTHDz/Vg87foAJcWP0dV0Gapajow1GXQ21xNv
JMj5FOX2JlQn7ss8QY+Ue6wirmjW3ydctedZV4TZLNtuPzKu8ZhytyMLDFqOW6/QDMR/J9kSzDSM
XreQ5LWaTLzUXxNfyxbpX38wOR+dtVaUsWamNtcqJynpweq6rULW6rFIOUt+DzhzGi0rHzUhV1Lw
p1o93Ks3DMMDWJ9AxJ1cSeuMcq6XamVgFCXxTx8JC5chHhdF2zQs+0nte8i0H6WAWwnmn94gmvia
BN52ZKCb30XJEn0Zt/j2BLuXptz6cYx4NP82aASNEjjiSGez1I1oY6DuKMRdD26G9kE+qpBSBRaZ
6QIBN/EreYIsxcRE65GEFJwxANjzvIgeBzLnYDdbGEAFctuir1WPq5PCpthkInGvS6gxh35T3SiL
1tEKG8xppNJYOp5EvDaDsbPv4QzdkiIkALHsd0eZ0srlN28a8nPfJB0WNN1CNXvJNwFIp+CPrA+3
NGjZtEbDnt4Di9tlRrMJ7sV7GtVitLxgLK/+o8QdSLTyoAYv/x7hXvv+bSlJMRXS5chyufVR85/8
P8RGgKaHFahNpeoyzY+euDjtjoheXJRUGVlsoksHM/KI1IozGHkw9vi1xLGMsczcsypl8xod1zxZ
1pvByXSRpXxO+4WAl4fR4ZVEhUeB0P4TpsiHwr67bG7TFbYg4m/7wRAmuWssXOzONvFWo8aLKrft
nN99p90gs7fSka3koBi/ilzdWoWNNLTyZgBs6889u8p/XEF+XXSGqPS+55fEMKjo8ysaMKbFkAnj
/f0t2m8jzm+M0f0CsBTL0podbZslyad+EU1CXjx6FRfZEjC0radDEuxsBDWG7ZkkLqSt0wWBue2E
0RYAMBm4dLVSWmpUoo0EM4EX/6O81jRk/vL1Z7hdz3jmifxdnU944nCMcq3V5myvgzXDtCBb0Ajk
oGQAoByOQJ1cgYnu8qAXVw4eoC56TyCZeQim+48l5mw2A6Vam1zPyqXg/U9HuQ/Jqz6Mte5c7nlJ
YZy4zOljnCRbWrrbPNE9wFWAyKrsr3LxZvtP0P01BKF+auBzcTtqFYunWAfs97G5RsV3rtd6j5y7
E3AAfUhAfdXM428qaYXh7vT74evg9QUKsaCa0N56n1SmwuqDVwieuzCZWlTjMZ/lOhPDr1M/dLVJ
mE3P1p0J0I3/tXjW6mmkdxYu2GLtoijpLTc9VK9TaqVOkJ31cDN87VMF3c8KHstTdtxeKI66egLP
kRzgWU75opDJofy05KsHK5VhDK8bfq4z99En6HhxrjNS5LHB2cxHqgKws7Ymb5ADDN8wd8nol7Ta
8LjOdEeo+Q00uQsbsaRbs6OrNT2AcOqF9hyF6rHPVuod859VTDtArZzYYdlIcO419MDZf6zGHmKp
liCAXqxyUUiqkuibxyHULpuzLYm+U1efzej9bOaviFZi15PP8ri8eUFEyyL1s4tk33gq5CXWohur
6W/lbU2B1KyrPvdWEHOFVZzOZkmSCRGl+CWCtD1w0X1Bgv96o+rQIq1J48Q1rbCxSoFF9rz7Au9/
MzIXDogrA6gRQiryYbMsRRqbu+xQgCrhWhCLToS6plcHVX6tymct7JPmZGVDW+8oMIEvVrpEK7g6
ovlh5o0uLuMdWwS7Kcw5r2JMx6YCly/BEebpAklh8UV+2kOs/H/t8CX1MF+8henmnTYrZpB89CKX
OADgxr86YS5x2um2ZyczPqzV6WNbCgmeccn5rQrH8tYJ7+PSDu3kYSBdPc7A/ofBDuy1xwneEncY
sYhYPVItbIvV5Ion2nTtQL/9hMXkk7QKBb2TwXM+b1KA9VD/Xy4bnDe1G+kXGjFs+7cIXtUTO5GR
ROLbnezu0aGuF7kcCWrP1UEsFYluhHc1T1mUmrKzwWdDeY282RMqH7nr1VfEicE28sLr1unG6zbH
SQzxi0F3OejAbJ6vd0abfXnATSSQZZoIiNnosf9WhBgxIBdKLj+qzyGHYlTI3vsXMqh1VTcsZLVd
Y3DGPn76XVTU3JIJSkWVH5KBUd5Dugztg62z0oYHKCLRsX6qcEhkyfKwXJpKY/fV5fS51rDex+0y
+Dz5c4aq0woQgMfHOVla8NMM9JuwXOdfGHaRLva4R6dmrOwtPExILwAPQUY8VHCt202bdP6VA2tF
X10P9aX1YfOFlq4PFwqMubwLi0fnz9/D7RyNk3gxeZhI2ZSCDrJoXaKEdGiWndO5SwBm36BVFb9N
wANhe+dtV4wPkxKaoJpjyCHSC5kWcg4h6oIsVJC9tKCN5rbmdUbK1Fza6pXzljpQqTHEbjGrP72G
qSiiWuKAdotOiPvx1MeQPayB2aSxm/p6tDpM1q8cVgmsJaCB3jVBK+EXkOIYNfCzpwWuZOeFe/vJ
GUyE6vKfeWwY/fA2HHs6d+1U00D/fbkU4F7FL4Dm0eiu/IkzjT8DClWxajHFvM+KYDUODfm8oNPJ
TyQ9ZfAYULemb8mAIlsHoCrhbFI+4MlXvVPLZ3fsmokQKEc5zyTW4B0LDxnD8Jay8GMZhjIhHNdH
ydHHU+jWPPsPXg8pNQvVvT2Y8YC4X5ib9KGObCdrRFzUVE4QqAUgh7IdRiDV8BOJHEIOTGSbTgtv
BqGmYEp2WWz+MqcjE1nvGumABwc5QTAIZD/1h9MI86Wt8CnBiV7AU26leazwP5OVhWS4T7R2pRwj
GLcUyUaIGIx2msvObXXG0QS1JM6uGYsVEilnU+0l38WeumfE7qoB1PRnHDRFDG6wFJE53wFjrQ6y
PvILrI6/M2/wISG666GCiq5bUhGLn39pPJvCKvSMs/Uxq5cQEdxI0PHw31BFKENzdvLVdSZxEkul
UULcq6LNPBGlD4/dtPXfouzpAnqCuJfzIgmqvSc/62x9Wl/MfRvxD3f2Dj9+Yh25wL2hlq5VQG+b
Ic61k42Zjd+JDLmQ/eLepC3Ni9HHYuQthw8WWuGwsMAd/CIsW3K/mtV/MAUc2JE2s8z2OMUGSAH6
zig+ndZVPLF8j+gRygx1jVYfL5GZi/7UVEQDSiK7n4Zezv7azfcNGQCkFQw3mj6L+d0uc9lYwFbj
+XIt87PvU3n1k3NSeISi2ShQGC33C7pTfYvsoIOz4fe7PvJfBVhoCVVSY+qY9qrhxzCC1uIq2C8S
FTEy6VfD3Rp2hrnKPIs3n7KAsFYVPdmjmaigC+m7xoObsSS8jaKiTnj7RBWqKlN3ctKDIVlg9SOa
p2o2y8EOS9/iGSaZXaXMLtWIxioX2kycD9ggxrHGwxMOpGdFPpC5AAVI4zJxEDbT5Kr1tph5U/9b
N2yOy23TssfGJDP16Leh30CymSltR3DoeN7Ocmch/xBoZp7+pSSeW+OsidCRoHpXfLNOXCqJ5kDw
TyS0b+LiG88mQuKjGaE55AsnWVjLqLyUDzNwv0L6g8s3yPPglShynSHrYyEMK+7Xt1r+9k8klp4V
zXN6JVGdBO+KGzismZburIYy+l+INIad7MlXUl/zD9IpZlEh5gn0MmMpiudq7yz6aeNsC0Vlmne0
LGC/h2YVQVR9BqoAdcdxSBdoiXP3WyGfjuLeMNaIO6j+5rqIP9RzoUpP2V7O9VgqhnVpkz8kUlxC
c3f1/xD4zIqAxsMPgKxu0rhwOTcai8m7yaskp7whwMVTzDr0LKpVWnrVXIp7drow5RQErILTtCJj
HLYRqctOvf0sopDzyjqVGOCBCy76mlW1JzXk63CbXQgonUemlvQD2qBkEEa5vlpD8np2QOumdtgc
dTDCuOTUIjd37EcpBGHuYBG8lEvUhA7Zwv07KGPGR4Be7bCFNB2TwwZPG75H9sA0qNhWLdinySSl
YebcXyLsEBT5wtixJOaXLWmK2VmBOzSPjaFaxDl1dz1IMEXn12V1yKausfG3foAK9fj+Fc5phK8P
q3YJADXCrX+FCa6hFCmoLIPdoizolml4+/5kTdrPlUuXXTH5uRIa9pomXrrf3DE5EkNevinH9zsr
q1wsoqyjJrXVF0EiEK50RV8isxNlR3d9cSPKmi2aM3+UnkIGhGLKIjWYWD+K1bWwH4yzHYjCharG
ALMWEwvZeWVzdMk7uq8YmqsPHS80LkHs283rdodfI+G2jC3YYvWinb9SHt91bdozH/BYN9Gpyc71
sIGSXHDKzbeMzcuYBYWDOCw3H3hBVBHFsN37FFclowBzq5ly67WnLeGYOBkWMOSKJwCgMNPG/opQ
LW4TmxqI/fNUeinuKKbXmjuTzDAWg8CUkzyvzAczWRJR0TS0ppdXQkGEsgGXrIOFBoNChiVPAB7e
NPw7g3XGt2ATxw41mS9e3PR0W1hxVQlxzhSTbCYRaSPUXxscg3XYjk9kcu905qDkmwMvck+iRI+H
LgqQx8Oc2Obv2BDZx/cqzy4fgeQw1REEFCkdIPrz17zLBfbbfjbSMNEv4YSIXb/dysZsaVhKZnix
I146HTlQ8LBtw7q1GNOkNKlgoBxBIdbqGMdZAssraoypShvcqpPDluHZba9ooXyqwUsW7CAVoU9k
UYLJtttVdlLetVpSi9mSPtmkSf9+p4YifizgK4kSC3VC6RpR9cIoLx1NKGUdnh4kxn8uoztFtl96
P7NASf6spKKN3CskDiavCwU66SABS7NbFhIQbaXIUp8vrgh4FskIFIF0+MpW7ghmph8MU9FI2yUu
xB8cc6/Cf67mqAPaJP+EWCK40o0ZHmSqyAA/LypLcqc2srIluUVqeGfVHMbS8K52/edU3P4ny5k+
nUqOfCy6M4zZrhiDGgeIXUA/E6kanmIhkLJhx5m4k5lpp7s3ZIYobhJlcXXH0VzxdwSXox0HJmah
mgvtSOD6gAzoiw8++cWwGRm7lNZmMcsFH8M5633UXC6joxzPcONRY8qrAy17oHX/X+65Y7E7m0pB
sS7eneHXZfYJgTyvZFOcwFJOsD/jA3yriHAQqy2U1WNapyPZBAcynMF1ppwuix0bi7GMvhV1AJFF
nm7ZUlMlseQ6mYAz8BG//0l8xafhQAlAZAktaZx/n8/CAjZmvKaBS4qVNY377TXJm35ggGOoUvc9
JyoWVHNvSVKNKFTy5Zh4ikgKWZsQbH32+eNGe9rh+NuImR/g7quS4x9Rrsb5GXBRTG+V6ALbIRfM
Y4QB18q8+dmPgzh3QdGDow9BGegB79TeItBdzdHjUpWCi/am3RQ+WpxKvF4TOB0NucFRyE9gMbBM
wDrMwtndGOXqlqr1yRs9V6/+tHHIyMlm8u+5EmH1CrdKS9+HEkElx4rerYh6k176CRhtOhLIv8FE
8nYCGWZY2WUR2fg/5E6TUJN59drkmX4DlBtg1PS9wKz5m1mmmhCaR09TvpcYqUnPcLL9/JySLNUj
EOCYuL3qMdXUcQ17ZZmhez7889u5P7p4oMY=
`protect end_protected
