`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57856)
`protect data_block
hTX64IeLyHzfa3tJyS5DfnCGfI2VwUPJSF+Bc54ckFz0mzldiRg8koOGfqr3Wv9n2pTtVUFRiQUr
inA2m+sGRHJyDdehqZ9sXmhUXWa6OLERayN7wMKbl0c9x/Wq6jOlfkiUAyCSTvtbAXfvPphQXaW6
/ykauj8UkQvGhXNBiLjiUYRcX7OC8vDWey/Uz84xCrRxDBq2pfIHwdDob/x6rG/fajiLKTCDijhu
mAFbKa3P2nZXMwI80e3OSrt4XaastRfLt6cvinqpYAXAJMIvyAkx8CeIICkAH3/AdU3lp4AY/mlU
a19fYXk9TVoDVA40gEd4eLM1gT46SVSeGqL4qpCBtr+RMNomfiotGev7g6DihQI7NL/40ZxSKsCn
cMFO9u25pZ8N+Rh4TzfZ+vGJODjjG87q8A95d0wIaFN9H2rtgDDAEHmDwgJaWdRDjpHalMOT2J4i
d8gU1elrq4z7Kmo3JmRtLdNQCFsIY1LvL6H4olBuCOzlGKfuPSp2yTvDuQI4H+I3pBfqJwfi0Q+l
qvTF6buq/5I4RvD/FtOIMNYOqVr0elwTNFmboY3JYsvZgSPXxCUVgkgDmUAvkhBDR64iuK28RdfS
tITa7YHNUChEOrdzrSUb1EmZN6s8zGWHMqqaqcQqjbwpnxj80c7A5TkAFEfrqACtkGH/BYxbKb0t
5W28tcpqpxect+7O/INvFQqrkpLsf/9lXsdETtfcJc3Stex39v8tEtAt08LB9D82OcXq/PkVr8bA
9nGb1+SiDddHGOirjkGDSCevcWnfvgtl+Daz0vqgshhwj2z9F+j8dcPkUabYHM+a2JfcLNJEvEZR
fesqmHBy3VwYo7//IXXH22lkc+t6WSok6lVhoCZ3tw4q6QM9unUg+G3Z00xkjc276TgywsdYzQ8j
gjbfUPftnBgqyqr8na4QV7zTmQCxctA2E4S4as/0ajcSnAnYv+SrU1Usi7arEIZcEZzQMbKoI37b
m7HaFIcfHY6Eiv0hLU0pXPlLGX5g1apP1tuHYs3u+sWK0iWs6EcyZb9ETLbS0TxntoAOs4f/EjUJ
c2XxhBi3Ahuak9FciSgrIDcYzsYMMKHfXIE2vs0LqYXW3hVd5yBfwHEBnUfmutrb9hh92GtU8cxU
yusgO0bJ1aabVmUWkYkDBRDt1Zou/LzdkXijfb2TrxqIwX6wrNOqNTMJdYKiRS7jU/ncMIqZJtdF
lNMRBBjFtNZN9CDDx7LKkyTV7Y017Fg5pRpMuqkPIqg1RmbBh94YZ9pm79CP/eVko+BXVq2im2Ro
BUH3WSbnqbE0Yp9GjG1jakmLmuvWg/+xDVq4CFTRr7ROFMM/eU2ZLOnKgTOTfwUK3SGFTXWCxkIy
JgdQJqN/7TuWVXYihoXlGRDaWF89ZGRBdltLgFJiTCCH5G7wu/Ie+8QmbxBmM0cj6VSDpZv2tRnU
WQ84xnRqhnN1QMCPqUWzFLJFVddr3/XQnV2nnzLcHFFACFJbYOwXO6UIzBiRuqfZJqv2MSov1w/O
KjnQmc/OK30SRK8g1E7APrIBHHUmxN4XCHdSGikPDKtV9lxa62F8l+h2TiDhvPguw3f/TWWTL/d2
D1QGibDMTK5F2tnJHkM2lO3rPGzOxuhkMdwRwlXWH/86u5uWAAzZc/d2acXU0zL9rKb6MVgsAp/u
t/rVGWq4+ZxqGRFX/SuRpwZB8xeOUCPZL2WVC1hyj6K+hDWFOyAMkIHR22nFrKFHAx+NKfxabtV4
qISWy86m/NtvD1w54LeVwGQULO7O4aw+CBjIvG1wMqVGwYwqNMS/o3XLu4IKMD0oatMaiFPzXRTj
upgEL52NxOP3+0wp7HZ5eCVLoTFthLC/Mar2IbjklYYpXAhxYDVl+fwEkG1EhePBw06bo+s03oqx
FX5dVDGxlIjlk6uHT7eXAtQ6jL5JWoxodsklekYcyJfFYnTph7D+82AshlOQJAIAdVmg2IEmuKLR
6LpLpPc/k5w+6nMdmvLsMuYCupe405YGZZs1JusxrLQH6q0iiXm3UhVHATCL2Qq5DT9lSI4lAT5w
Ofx/psHqi1UfBj76AVKkJ2nIYel+rmRfqslzuDtKxTwaCYq3WhRomGfewdisRvV2jNWg9kuAxHto
I+JlO3CjrCtTSXFFu/FDL9FdFKGOATFNFjoru3K+yDaIKwasN6unOU+zfuHW370c7JRMaps4VVMU
982TfNwF+pWZItYS7tgHMtyyHsV/tLSLwqLIQTstWNhv/aBlC5mgLvIK5hEMvlqfPDnvBtPxydk6
PMolNISUFez4+MgWtZ2W7pxGjXggbEoeHBylvCqhiBei20eNeQ1UfAULpUhfexrz46Axbpq9DJMy
Yl6qrTCXF1da0kIk4NqvrC4OnpqDib6uqClJ1e0C3fGXB7VJcXE8jq9g+q4jwLutgXTpaHFbOUX5
TVJFwn099SjPiX0rjTI/pN2viM3rusgtI53sV3JcNCMPpoq7lEc8Mafx17eEqysqJF9wYRbk0PBE
bKxepbHu2pFh/ZOziFkYo/+vRTmXWg2ytb5vHGI9cSOBWPlByWsPzvD93/eOLmIrkY5Iy2LkjjjH
QK8hqIQbL5lw5PNqIvCNlP0zNBxAvfqAfUfSm8xbym2RhU6vkARMojJjQuClF19cwKUBBkuo5k+Y
n/0NQdwCluY3qU44+WB+swLgObPtFuAYohiaFQHXQNytxuP+Xw/BPAAqOP/VLRHAd6YohaWQblk6
hzOGHHZ7iN+7cEzebspAD8DTl22pk5SVLe57uDW8enLm4kEHYDc+53eGS0Gjp1vfsI6YBYhFgHWI
muzCIpZ7iF//klcrnb9dYbCYjCkPKuWgN4/anjNlFjMmoH180w3QaaTl+ozPwgz7BlFADXlEMbdt
inC3RsWRTJB8+UHDtwi9Kacr4JTEO6HUoRY7P7KGmhCk2klEktfLbF0jf8+qqtpt38QA4XuLa1Fm
+mXndjZzN3SxVhHdxoPT7VECAGEKHG6DLu91j1gczZ0V7RCI0naD7501siqahGFWx6JKKHJC7tkb
1xkCfe2X7uQFYq+QwnVzkfGzj4iT0K+t7rmJPl9lOjRcnWOoTy3LS5vMK/QrKHC85EgH2+m4Ua9c
lTwof9pX0LqpfqRueI0iXcAuB3XzxgtvxxDdnQsqtwh1gQYhc7INRkmSlip1OL0mAaxb/JjyGgrS
i4ONPzWBZakf2zjC+o9NXcXIFGSBAFs52OmAXFnjTFMipe+oHAfqYBGxIDnvJXHgFiBLsV5GNRkV
NXgBGop+b/zCPaseOeGRQ2jhIHFJDIfqmK5OrB90MBcMADZcMtqAdzrtJ4YYPTguo1cyYkVDIMeb
CJ5iKx7BSWGlmZzQmo2KhcKwM3U2LddcDIaerT5w0XMZ4LRU3qP4mZTBmKrWUa2Kj12dv550j+Zd
1sjt6yZsYoJEeFsS9P8y9e7ABSvvGQPJXpJ82UTiqwOCXC7QXhoPsH2RJVKQH6wWfQQtqzAjdyNU
CzAsNDZpbna07lmV63bC2jDFARnShVvEfbe8Sthy6Rt+8bbqwcZDdraB21ZqfQSpMRFXKtHKvCXs
GDIM/r3RoPfLU91TbQC9y1D4gDk43QNgIV17Vmbt4HUDzLeFBZN6oYsA3vgWWroUskYYNcOgs4cT
JPmgUkG+FpAjFRMz9JPXf5c3B1hPfUyejLvNmvpmiAe9X/M8nNX3EroQToCOapY/LzXW2sHVVm4q
IrAOIXqFoPYVSjxPvWUzjDQBlUYXI6waYSZM/gAU7l7ZNg1Pr6Q2dLobPYlsHUmOrTGjixUNooVg
2MJ7e8FjRoidccE2PpYAOOEuS9WfMLuqvBlvvTx93fizC6Vtyffy3ZBobf1J6SiEmGvOUwx3VFul
vHVRdEvpHk0X7LAf0FQTe2Dg0x8U4+xRfrNxpBDZ68veB4wuBzM+ysqcjjLiJ3A2NlXjNdugrAEM
rrriOiZzYSV7xRXNO8jh9nNLhvIPUChVgk8Oq5zH4j123IafMpM03rWQMpXKSLvml/M7Kk5RZVUf
HEmbbmqQr5V9BNqcasGJBJpfFC8QX6/quAq4Ggsy7QkzZCdkwqmHpLffEfMN39OLdmceKHaGsctQ
pjgQtfMupyZc4O5e10uWYQzy0sYiuTVCA/eoKZgj8h/6nlxfP1b3GAP80az+375EpECpx+UNzwW2
fVdL9dDv3zX4pMNZp5dh/tGy6asQA7hAzdHSytzBsnZKc6tiYKouFQQ64FdxsZA1Y6AcjFt1OBIX
DI3hQtvX6FSqghGgekNY1dZaBRcbXVlxbL+zwpc3S1UX0I+ICBQsNOzJngIdQrhWencloWExDaH6
IjBFYMoVq62ex73aI9jT3+X1UpG9VBNTRioi8cfa4e/KakYpC2T3Bx+YOEttHpgq5jxBgsdRUh3Y
gwjFK9ANTmnPM/p0MKQBWFwCIe6n9r2tQYAvn/8mNatgtxei9kIYYKrKnurNl0Ceolhm/tvC7wLj
lOwIJa4LPM+sEyyOHmUfjsFSEqzWHMFI5vshxM1IH3+/NU43jqI5buHK+YWyaMiB9MBS6JAIp4p8
EMf16wiswvXpsMCm8uygx4B+rdwLu1b6b/N/8V6xokBQjknOQ83PDKSVM7i6AK+ODmptIMDXg8sR
zXPNQztBgh20GeCDb3dVPozGse7UX2vWgw0TeU4TFSGImbwYLnuxUdkmFzgSuUO7yLjljCpIBXng
8Bcs0APUFIOkKBpXxMU6/SY+CtVz6JcP4z0sDb30Yl2hRej0Yho1LDrIGgtp6i6iG1KU7nCMhEsN
uYBHaFVE3bVLuMWcgQe09lpGZMjs8UhnS1boeo/ffR4orW86VbaCI8Y4o5lR4fQvwhjsy8MwakeS
YdKy8vJSLiH1mdAVMwnUfHLmdQ2eYxWWQ83PUmufCKbtBjFzTBrYs95B55qjat/vggA2Zm0vTuTV
6bvrfw1/1QB+BrmXhq/YOyoDzMoVUnG3/+hLwxRKuXENDAxU1shKXt4Um7lHtotZZm/ZqZTndGMS
IVNPINFWLnoeYuZm5CztyvaL7e6qbX8zkRVr760ihkLE7LsDcR+Y/44BYyGJ7mfcNmzvioXgSrnC
FpgZPdKSeGPHcpc2Y4/afzHXEhr4bVvjMEX7ssOncG/Y0WXZPc3l662JYxE8kZR6wpClo3Ys/2b5
KgyBVTh6i1aeLbRefhDAyyr65G3IW4lt553xlYUlcMSXLeRcns+eBScg20V5ZCbMj/830NrqHQgQ
eGkO4qMLiUL/ZgSsTl0+Ku+HDbDADVDTRklyHYhoQSV4IQyAqE/A5xBlJvLo2ouGRDZwqOkiWLMt
jQeycbxf0z0H0TXS50bukeDO39rHtQVpaVl3WazyxcQ35+QI2eFPkHVGhG9t85855l/lpJ9ESLeM
FTLpJ7QYdOCKclcv7QNK0z4J9yuw+/TsseAaNVQJf1zG2UXWDC6KLbBv5L8xVeGuT2s1luFecvw3
UuN18ubJH1JGiU80kRwNnJiBlXyQQgF70Tk0k+my6/IRI44iE8veCw+mxqOUBeqRWq7XbsVjNZUS
F7n/DT7diiPqiU6uy+ipB+OynQcaZg/7SNwj+0X38UHjB6FTN+pIPRunr2jhFRUk9opNoKTc252C
SkmsG7DfDvdPLloG0UVM4N/bUWLXTqRxW5PPrfS9u3enYqhbg+MZUiuKo1fWKvHtKjXBBZLEkHqd
ZQz4G639F2/gkwfHwykWzxof9QY4k1EQdJSpoSfgIysCgF7GOHyi5MJmf/lPtaHPSGp+uaO+QUHF
YUXgyMre40f/nwo3z6JUY7m05xuFRUfKHzUcfLyFDFlk1n5JcN/gVnrJUO6MsOqQZ8R2pnBxLBBF
tdHaOd3/FimEJ41Me+v4bQO48ZDuRynux9IE8p+wt4I94q6+CYSCOVNBbhnu2txYe8w0gp8mZOqW
FIXcDmJCP5xxAWxUoKJKRDsiyFF8IRe0gDXIboaENDsDrj3HH47kOgpH8XOD2HU3cqj67ogimT/h
NRwI0SvqvZImim4Ac38s/BEjR5P49zmkZIC/abTQqrq3hhHSDnanMpgZk29sKvyI3j5d1KeSezvj
C5edxSSe9pWtQs7WNIlvNaQSk5pR04mc28IwCBBqgAk1WIq7YhoiKmLFx6ZyQ2ayFcshmzaBTgQR
E/Uv4N9OgLPvm9Ni0/4Sn8n2C8qwY1RmOAvRT7vScLt/y0tLRo2EsobDvMVsGfoIlyxlwiM+1DpV
hst9n+C2Ms95+nyaxOF6OZjCwsoeE81r6MXYvuB1nm9ssYq7Ke/UScCU//J6jjsIimCDjYIggc0e
I7/dA0P0vVyMYpZHSLhq2Z89Ca4iBf3pNBPvW4y6KwcP9wDh8y/K5P0kjsz0j3A4avSxJWURUN/d
5ecEg52omUQ/I47gUkOIKHSbd1g98jd6FZDD23CQIuzy3v6HIyQZTtDNVUKvsYhT9YXHdUHRFchP
YEiy/EvruSD72Zce5k+UFzVTHA2w6wlfCqFoLK5gSYLbZbhD0EBcQxAIatMTMUirxVBsvbH3gA9k
LMgZfOl65Jx7muXxFyGWYgCPNnbpvoy3FGHznUz4gE3tF6LTu/IGvky0qYoi0Ko++4VYWQmjQCbT
Mk54Sim9VCGdk4d2S391JujoyQR2xdLbhRnBwm0QhAs0TCGW8w91MCZTPuzq07HaE1vhciVeVZvM
TrgC5zcao4VshjIAgkkYuKzP7U9aG8epEOP45dRJq+QYq/FECHpLXf15YfOd/jmSYDPXnXz1Gr6M
nu9JItNdIpsDFmsJm43DKheFz9TjAwhcWID4Dri1iv+v86BfC0AUF4ZfS9voRGrOr7H/y1g3iP31
HscZC4U+0xOTmp71N899A91Nhm3GIqzR/IisEeyqAboS2vEIkoeygZvw/61fGC0VmchBd4ilD08k
PGMfRs4m1mYasZ7bxVI8mBLszS+VJSgmAzSE1OuZVBBZmFkRE4wx4DLZTjQl017UkLn6jCHdB2cH
ibzOUUSgsp4gB//SjCcVaOMo2hJMzU1HJs25aHWG0zUnggVuiIS4tXWhMr0lQKOax5e3JUj6KvSs
90zyq+emjingxn2EdS7KWeCZyqtWFWkpum/pa2+4HXWu9lLVJ+XW+xpUVp0NQWOYxKUd1ENmLUUd
PfomN4YMYRNhpiHfXX5EwemnQGtG65dlBtVFeTO/590rlfHVcxxoxJ6QwcKxuy/NTn45ofuTnrqJ
a4IbnUA2by2jbdpw0IsUiXbGhTHv7zN/IlmbGOAIx/Pl87HvP/fCVr3bKOQogeBobZOsl2mUpZQo
T38aDZlHb3Rtx4TZR1g6+SBO4R+rUnB/5KwpJI5pieBx5a5u4GGhXGuAkY7d8YUaTtWVv2sh+tEp
p7ZcvHH4jgXdch4KQ5QbKWLmxGNrXtMXX/moJ1QXcoCmTpBmX5OQtfTCjZcGEJ7p5r233EiN9Iqn
CYITOzOXI+sCeBgIoGz9OmNgV+Fc+BkO7rG0wNmbZC8rmk086a2i67jxMhIUT0jVm2NPNe+PoXNh
tVNoTMXowgauCV052u4U9mq9h8Nm1mfQzp2TAwO70jePxld4alzIbAhGgHkN5AweseZOLQC3Yigr
S6auQC8TtNuaXDUPVMIrA3O3G67Kf0/j7MtnMoUel7UsfOIDtHmxTaS//Et9MW6iccfQsBNdx3W+
938EmGkPxqyX+jhcJgqJB/w3IjTSl3fRHOAYoWGf5pisGmteir1isc9jLf8xSrjrLHn2AkHG2xAQ
LygzHJJRt7tyqq2XMczm3qKwJEz5QLLE2XlASCCpEMTjlWY0/6GH3qrgMfyEJMtFmbvXW/c8fU/v
S5grrBFMX1zSJqNftrGHqV6C71kIsQFpfc9GmPr74tuQ+TPH/8ajCbkwaHmmi9TP2QKwn7yZJtY+
fEgHfj1XFE606eO8p2ld2iuNh0/bnm0omdOaoTcMlA0Zz3lbyLmJVAMbucfegLnShgm1MX2Jabdt
Pg6GYKP1mgUn9E0LS/mXb7zp4qV/cMRrb2epbhJw6sAtJ/aTYzptF14Oe9GUAtDXjhixoiL+8A6P
MqwF92f0EGpjd9pkq7tng8c0EadW+RhIbQh9rZcHa5XwmMgse0qvLu0z8r1VIXXefjOLm/34Mnxg
eRt7jlnXjsP4HWdKbWm6jUUsUHAsYtcDFmM6tGBSw//LZ1cKKRTV0cni5P1ITM41QWGJArbKJvkD
9hfwKllT+g5uUlvHQxwmrX2dRl32TmeXd1yv/vjX+VoS5V1RyZraPOypIlG3Cav0tIG6KBDscVqx
1xf55ZR9z5ISd/+zv29rvB3mWvX05q0d0qp0bxzV8Tke1FtbrScRQbnDq1Cn2y8bobkv+rW/f/Nm
iyqKgw65xyDGRMs5olq7wmZC0sXOmsWC0pvaGHWT9+ek0mTil+Yf/DvC7j7aIcCsTj7rgR/vO0ow
2pMRa2wPPCRONareTOXSs9uwF1lYKBbcHmQTi6vyYURmMdCdBCqRjRNsduU7zhDcUeJfeSBpHsFk
UGuyGlVtwgGHAtr1jOrqja2ywa3AFkXn0G6bnmoWeYpXNy0HtIF2MS3O/WIDFFavMqFLw36W9gIM
FeLs0O4w2ZYtX3olgy2iuy72tFXx9cjlxftRLr8V8Xno2lWYFTW4z8roiyKDQqMBG2Uew4w904BL
UhSpHz/Y4TW3NeHDihTWUe7+2x5iY2s8sybboWGH2vRxa28YC+X9KqaS3BUNaCMP4+HxMmFyEuKh
S3+Xxxp98lllg2BD0+83QUFzkyUxYAEDTr1hGFES8ExlAXv1W2PS9B4ojLtlv7vDWvc2FWDAshDD
tDY9uSyA4mZfCZtHx15i9crh5P1xg+OowCvf4EiBXgJMYqoT8O7kTGualEVPDXF2uS0MRenwGAqw
qcCdeNNRdFoXOawajpInUb8IuLosT4hiNxS2ZFpty281nemIE3p+wgQ75DK6dUfKjMjkErlI5hYw
qCgQYTu/1jpkOSfObD/e8XU5nm1Evak4en9Sy6j3gOd4z2tr9sUTQQu7wyubPyb1K9eied8IVWUF
XGhok8miR8UwLTddPt2p9u4at1+Y1AjPBHD2r0wZSqn1cUZ9vQRVIfwSeEhAxm9yZD6tEQ8+rBg4
PxWM9mB2jzXxpqSbw4yq9VdqWek53OYKITRLKb9MEAkAMjeOXVVUJ2GCQM0wj/txC01u1jfv9pww
XUujECD8YFCGYkvPnUBAgSMS9ZJX83MoS54hv1zx8MeUvn8FqNwNabfJ5ykHJ70LRH3NElrTq6Ak
qeVNVQ6c1YLdqWdOQ0g0uZHV3wqpUc/2zSe422sgGDZNycpFy3BvzWPaQIEcmr9oBt8RGtxGsPak
/3Tkm3zlltEN70IGoOAnXb1ZH1WLoX7l60ldiT91N1mulJ9rZv0O8dzi80HtY5ndZfXur6MXS2hs
0d8uJQPCunbaHKDWVPoBiGJ3RxppHC6Le18TAEyz3hew4AmAmHMeVGFHFnWA6UA9xv10jZHHTbOW
6nLd6MWeiRe24gRLPq+u6Xo1Ma/UKV5abBZfRHE9Trm8uD5Ui99XqmH4i0bC+s6O/6/GZnVCKTBR
+o/2gQPt8xxvsthSG+4JySpwGnPkopl/oj3rblHjMf7v9pKo6VLq3N+P9G0BwCpvj11Jr98+9/gY
pvTrpCZQ8cRFHtvpiSOgGtoYtg+S7wnk1syPHu5DI8A6a5NwXp3htW9RtKHPdouKqlUYG67LTR0R
U+IjD9OSoON0UQv96qF2/nsBA1QM6N+yiXVJTXGTKaRO1/BVmU57eLYSeKsGe+OOTckFwg0ia/ET
3i2Uaz+tD+NK9dITd2lAivuh4naPHeFLjkeOGZe60Zk/rCwRKlnEgpOkMXGJ7DWhO/J+gddJxoIb
qu11aCxHBxuxWRhX8T/UNqGvIbN9h0TFShloJGL+wtA027e+8GEgmNAINcfGFZPIJrrO96Ewi+pK
6mvoyqziRI0GeZzEhqkHPEP1agf5jr+ug5wu0757vfr1ez3p9219Cu3fnt81UDiKHadu2dW+8flZ
4o0ulzHvILrqSfoXgMICtSNfZ8nRWQTdF6tBsrn/v9RLL1cmYfVyMn2fug3au9zexn88EpJAnr7q
u8H/ZgMpbGsIB1mRaMA92TY/i2ndYIpIPM66MfSGzYhFct0bpUdYeT/SFKdu37HK/cBAl+NuGWdc
ipS0Cho/kH0+HuaAF9sMlEPoyh4taYvUoa9mebZrHzJgSfidyuOCDfQbFmKtCZdKX76EW6cCol56
ypppMAk7snwdt/QmLEBivY/PqcWM4UvO6cv2yAw2oNvzgpY1ydqmKLI3bkxNDCHA+xs0UTnogVn5
Xgdinprwe9M8MrC3qmiWJSQLrbeu2t3rvFX1kKouK9sC9pdhfeecuSKhDJCOZ0sdjnDzlire54NC
bdzyIP0DN3Fv2fb1FbHAVE6gKuYfOjmw1Vk+s5CNBqQSb1tR7xOkeaDzq2TskzBObRMjnHMNq94g
XwWaPa3ta/EkjWZdmbcdQu138ZJcQMR1gkrKTkdX1K9d/lETLDmKN/AqitNjxibjiqmhqmIsQgVS
8lb4Vl1U4d8emtCpPZ0HTsrwPOVywt8GVk0P90yXU9or6127narkzkS5slqY9+kT1k8+3b8TFKbL
Umr7mM13PO1Zx47nhm5CIjT+8wQb5Bo7hqX5sHBijm0gkmgKEDfx1R1GntHzT99ojIC3jhBWAW+V
xgKo0dZHKNULW0A1a2vsCNqf1HnfzTPLMc3g38fCjjc4w1r12QxJ5pl2jL1SC3kLUDqyhdKeE03X
RCYGQREJKtzm0CFtgJQFGfcFXqHFkTjT/0Pi5W4q1frerpQF7JLQOOwLqu7+J+zRHeM835sqhgmr
gZIr0/W630BaAAkIlcqCLfZ0iNBZVFNPNo0zLTuAH01qBU/AwfXQS40cSibSpirXwhPZdUcUsBno
b+02YCdy7LkMTJRr5+SF2gScOsb6b826+D17FVrku9gKif00Wo0/0cLUlV7Qb97YOV6+nCMPdVJY
TmLIG3pXw13ZcAtsW/WZV6Jz7tkHXpLyDKFewmCSy+uSHbVJznW14Mi5fe+nyrViT21ErAggWY3Z
9Mwuv93l8flvUvw2kOLnYbWCBx+zlyPqJA0WCxBwlkS8LrXOebcIpInn8CvOdzuMOoiD/t/ZzHRT
/iR12y3rC3inwwIiRgdJZNC5iRNHcfI48m+Go36HJnTi2k6IjI3rff7qX/Xgk1heATEsoRKZGo4N
mYPNrjX43osM2U+DMiGCe1rLVGtnHrLXq3u+s9qWSUJ9CItpR3JbsgrogbuVe92Agepho5v2sKua
ZbVJTWNVVjQLoko5J7jIAjd1xwyMZkjYpCmK0YcFtlC1GLP9bCyvqtqmP2nY1UxdBkmkcHq3F7yW
nQoaYNR6pMsAVP0+yu1fCO9kcSZenJSC21Z/YLTIc304GgTDHw1befIN5GYumFK1jO1gERu9JoxI
smCAKXpttGRWoQxkkDmPjkmJuSDefktmE8R1sNC3cUuazfKMVeuXS38n8EtNjL7UgCdyJ8P6bEjK
VkEw1bgsuswmex5ahpfxo3IidQCfAAFIlyImoW984bwfep435SyTahyA3COwPothGkY9vwgIzGpH
d5eMivPHmQF+f3IvB0BEH27JyAT+c4hTvY4sbQdEKBjPK2xoN9r36uitbqUW8y0dcJi+sLxZL8ff
U9d4Dr2x9hV89zRnPYKQZYs/hMbbtSNdhNhi2o9MwBO8i9WvlOGGilBTdGqIsHk5avUnjDOxTmiM
LL2gAV7Y+iYbn+H/sDQTg63FVL5hNviwZrWmCw2yzDDAldh5QNh04dvZwkPAljuIrsHNP9Y0pE6v
R5BkjhdcVVHyo8RZlGGNy7I/oqah8rfWiEY/J+Jb7eawFbsxT66DyzvbWEbx1h0Q3bbnib3CgJji
+ScfjtZbVE/RZYLN2+o8ViVa1edUksaFe6e6R91C5QYHtEtLb+rJplrXdkIemt7E7JchBP68I/Vo
j/GKtrqzv2D+r/fCmh9bEqOmjiEPQYNfHUzmZvkoT8ErZFn7ASJHmoqyUqd6J4Ug07OPYuMQ/9gE
D2Ius7tuJEc0DEtWAM+lDsjVKk+4fpQWT5bD3Gr2vKORCjmqm05H2yU/zoWrFW25IEMQtW9IFvEX
AWNEOuazdwxhMPutPdbZ7Dg3BC0bI5UFRo5IY6WoI6XNYbgWO/5mgp3KrHu1Un+nO5YZ8bzeXMml
VKzhsb+P5IoOo0HIwVeOYku1Uupa1y3wMG2LCylQZDg2XhzExdJ42OPRsJPmiK2r42u7zWrZlRBL
cB7gPoWwTXNkLiZRIDZTA/MAA4YcmMdut3/bE0HTtkHw1JPT7/Ofi61H0HczIXtYEC/sDBe5Ou5B
Sl1j2gE51Jis0Xsid9DvjRLjoQu9o4qCgEYwBWgH7riIaqVO8ueLjmE3L/vbwYKwcvDNqicsHxzI
OWJAD6hyjv1IdSb8YoVBuIGo14kfjlkgEck3nVGttXlbHXSVi9G53tC3DOOSRcncEmo8w4xWcLV2
sVqC5F0+g8n5bqbZ/IozZK0ur9gJkvMIAR4a8V6BrKNQKV5hRc92018RtExV1Kz37ZsZ46w8E3Qq
IZxDlCym4QT8RoLm+uaGOkZNKglzRESbMMijV+91+JkAIj1D7jwNIBUGRiMXBTZYxqzTkcyzjFRm
s5TnCV9uqHfjZeUF6MuOoHg7Zfh9BFVT7IKibnBgz+RnOXuEaqsSmZVLPkl9NdGreFwSG2o98AlN
tL3PFK2G/pijAgrprRhdy8bbj13I5hb7sYwvQHiDoTaIMdD7fwwxKj9lqogHXP936LYqNILSxuBX
ImNv8XgvFOMJbm8YLDG/Yf6oqtOdudEbAMHCLc+5Dw7T+w96tMfqqM3rkjIdE8l0yfIl1nqg9niD
yVdclJya/5F4WLoclz/j5JXM1OyMeIMitI9FZFhxBt/4XnFPzBW7ciRuQ3Gs/B/UpV00U1geYf6f
jcw3LGiG/o/v0rmKyOOKGvG9HfKYjnOIUaylq5CnAE8ALB5akqyF8DEVNsJd5tgS8U1U522rS3D7
IjmM+cToEexKb6udfJIHktsMwsQPac5Ekonw4INOgeTdQfm+jsqmq+qJbmZzbO4cbYZFTY3/GAwT
i9jW/VDLDlFRW4MBnIuQI+Itukzzg14n6ywbGetOkfwKkDYVBbtv3GEu76iBwvTNSbDohpP2hknf
OyGkzXgSV2+lCZaCHRMP6Jhh30BWGZegMjnT0GU47LhWVuqgLrdaN4SnvlWvruStrTMqoKJqQ/kr
08B5nVR0oCVw7yRzdCHFqeFVzbZcZH0JV9+28Zr8eye+VdHaqlEeKouullo8wreIuoYThiwHcwQP
gLKtuwnZeRVxqD+mvsq9xYPIsZoapH2Wg+OHHvTXBBtU2Mo36PCp7AcHbOhMJUh/GU1+/69wm2Qu
rLR1GxPkIJgl7GNM0J8ty7m/6VR8znmJageQe4FncnzjxXJJD7tqJlizXFpIkiBSpMZ4PoQd4QL7
6Ubh4cmmqu5ZSJOALd8mRwFA9F0WtM1ZnrZiIQGHfb7+uOrqRGq4aFxE3zDBOftT12dlRExGv3S4
bnqbaSvfXptluS7mjJ5D/7mwgJRgS/D+XFjTgS1PQqPk71zYehv44uHDIFU50HpXzkRUQBeMDFAv
ExU+bigMiu16srbABtEECi8qAB3HAJBL8mT7Z0NoXgLlgIhzp93tC80EGn+XvSgQAlx6sXfyW1C4
qrtM22phhZmQ/Ii60y69+QWuifBfwxIarnYNsjCx8N3z0FuAtbkusWZh8VutuDqao/wAOqPXs2dw
2ASShaas/DqjERDuWXsRu20P0gzfTkmC3GRwsOgQhWrzRFWFZZ4R3tmTOFCMwyW1U7ToTDSwAhJS
eNdXpUdeZncRpZaOs50XL5zDKmWksQDbnP7MCTq1G4/lCXIDUh2nQQQ8EG1TePaPEai95m7Mx1uo
Ho+sbJq4CFAJZFzk1jtZobx/pJuo1NUg0shfVOFEu9n2ahmGKeNrAlh6hz3gbkhK0NmHmEYB2x54
u/PEhgT6HA2DdYks43w00wj7eDhslV3qxYpJr50dpZ2ydmERxH4yhS1PprP+l0QV7sn4WvMEslQ3
NdnYJeqQRh6F40zSncNIVGDuoVD/PLXy2jbRhGGD5dX0/9Wt/2KGJSNGebHdFW+tj3Gx+0E+6oPh
m2GJKvmJ+LkkwQMRV0/pMR4Qm7wlHL/7n+k9kFMQVj2Hutnz0z2sETjdKcpAGaByhbGLfgpgkiZW
TlEqm2b549IEFT/Fyr8Le+8y+U+yCMjVRsGjsDfdro2dOnQD98OJN/gxR1rLW0TEvNcUKi8drREw
FxOhXhPIPmzkhKMcb4YmzTzqPUOxEBeZADNPFZIQ7EeMEXOei/4T8KDo6Rs4awg0oIZcX+Es+tY8
Kz/KZN7A2SVG2whN7+cExGJmQsDGngzwk7xOtxrHKBnGKYqSGQVExCNDxLi1DbojISs8WhvV3TzE
UP49x4qo5OOOB9zGCIiqCIstgKXpH+Hac4RLE59i5LRwfiQzsK/8z8JGKfn7wcKes3fxPrfXAqZm
c4qf4H+7SHsS/rAU5OCFLR1aei+6L4UzsXTL32leyJiR+oGasXd7wfgMEnD/dBzXaGonLl+M39Vt
yQj/GcctVTm6Pe7/yES5cz3bmEI0vCpOrukvvJk7CQkg+2zc1KbIw9S56hUekEu9egu4FU9ppy4B
+zgS8ha7FFmTlHy94Y9XZvFA9u0JD5Me+r8KAzB8KAhehK0Ez/FP/uW7h0Kkzr7n2vyiA5xcuBut
miEoDATBOrrPHtNe/Bh6VJjh67dGCym11/2t5+XhA1z2PfnUhD6wW+pXJwcIcoF4Et2JCV+2sLNA
grP2C9n+uiQ9t2PdsiEtq9lGEv+jyBK/LjvkeQfgoBzo6dfnp6k2OprHddg9wWmCaB5Sl+5dmp4D
hdJ9YPu2AKVc9+2uzYdK/lNkNIEiF2it1W37JrLS/XbQ++f2AuZsjkVAKfecfkkv0MchHDIbuo5S
vvdqQDrhOh7y9dBHaul4u4IgxSJ5S0BGEb1r4TEuI/oxhsSPS3Sx8VNWWz7rYOVLdMMXbLpum0tp
38UrylFoJtzKxkt+rIn8FPKu1GHuEgUqxD6RLHAyuWi80tfu9PpeT69BqhYlJ+LGIax21L0PnMtH
qg6KEO8FaCpvW2ib+rGxXJYnxH/Oi79J5OWTKnsSOSak4vyFS9D70iLyssOGehE3yHlHdag1rOht
iBXDoT3AbmAxrbFdfqViVfaIbdkJIruRQHtGf/KHvfZMQ9wPbZExyKizWdq0JqyEdc9ns3SHd5E5
dBBOx6a9Uon+dLYWo5QD5ea0wAxXuP67iC43VVFbkdgbW0SMvDdPZPYVw+a01PufuW62f5RcieBG
iUafuavhIF/bkwm9piSeWVpwaAsZUCJOUOI4RK6An3kQVQ1HGu49KJbiYluBRVYuZZiCtdIJ2AZD
MUs06ND+rMkcDBh9Ru0DtX5RV43vh6d6SDBleqOUvZRWGLl0ajj9o1SN15iNvYSlLaKusoAsz2FI
d9Ze2XGZBzDyfOOM9jgfip5+zwgf268b7naXj7PTJxHelCFlHD1NE8YFabdUxUTKaT3Hr/BoJVvL
Pswqi/OUVi+8haab+t2efBtQefJWrZLh/iX0bggvXJjEB2TCAThiMKaQyHR1G/Stv1KJBBoxXK3/
j+kaP3bbcsOuHc9uDuEXOXaxLlzyCel7biHBV/Q/eFKmWhTi/aKhcsqpB+jHTawaz+mbb6CdsK4+
XMKCfqMLFTMe6kKPKnewzWaWRVGKSqJ9h4iVzv263/odyh0/SQO+oGY8KjvOvdixsGupRc4lnTFS
F8Vda9vkx4OBqmkcbms/y597FlR1kBjTREfxDptW72nacXa3PKdgPUyheCZITs+o7jFzTP9GoaBz
6pUqqfGsGQKDqSa/zjY4fCmsFYPd/u7oXDKt+GkyB+9vxD+VxR1TZs3tgADTXx4N8lKlVzDzeZM5
PXhTmDYACFf9jYSaezXWFW3NnsUnv77FmnryUPHVpRA+1vG3bUyTg+6P3IcJEeJH2Pnq4N21xE5i
EjiNlQnnyIaVEb+l3WjHux63vIYHXj1ANyTubmT9aYIFpaX7yTzHo+p6j3d5wWrDea0Gqw1dnzQ5
ZoSUqIzZkEqYDHNm1CiUf95R8nB1wUbOzFJka0hmKW5PFm1vxz0UzjQUhtg/UlKsLHesV7yN7QaF
mTs/a8ohuzT6aiqBxBIfUdKNHlv+Y6wqVsJQ52724+7T2mH8RKij4a07dgiROb9OkOA56XcQeNhf
wH6SuVNvKqKqGX7zHP5946GnrUd6lWXqntG88jcUfW7dd0o7w6JS8LAEpXdQJ442OvD9G1yFGNaJ
SULlI/wAN+B9qIcbMo/W/LHSP06O12jd2I6ccb8If9TthOsWYZxi0xwGB17mKdm7z6SEmRVg6wUl
A5Fx+aBvW3N6/5bmYeoDpEvRVUffiq4nmjyKelL6FaOEtQ08ICXL0mMS6IbYzr0wGY8kiFwZTsL3
maMEKJgYZ2AZ/oYNnVU0caOCW9vLD4vlwf8itlxrwukX/Kiro0t2vDdsKErDPwd84xnuJQzzyGOf
LSfSFO/5TMtIaUTF/VdMMuQarqrym+80Ln0B5ptvmxQXsJeCKE5AJWC+FrFRQMq3Euo3GKfZ+Yja
zUsGusA7GUoICaMhchN/fmk5gcNI23uV3OmvENxYX5DSOD6arXiJWOy4WGuuwF0PhU51RGXYspER
wyXyAbzZvPHO7LdXgzSpXyS4+6E4eJi6jCTsSruyTz0Rd66wQs5lUxMVMEwiA+7vHlbAUieBy+1m
19xlZFy6ifTinT2ICJ9Ietgg0gxdv4J2npVUDGOz5rL1tfo/xQANEeRhG/t6nI2pqXAFKXV8NaXu
n1Epstp+1DwyIcKoqO0g03tLSbZyYccHvU4/ej87jZ8IbV25bUXkZ7NJG+dTpPangYZ2KmRfsL4J
liKDbcAiS0GHhV+LCspWheQuOLwxhx0HWofUa6a3PPmcY/DD8vz50d4fEPK/CV6Z8TJjEkf/nyBy
bxkGgorJpiTHzbX9j+3Llws8bQFoo4Z2AnxiHf6+r8nKL9r9sAZIDtOAwrYNUHz7RBngeT3zynN7
pheLRBWv32Jd9uZ8nekKgDhrQOysUSSKUWoUYgVbLutt7SawT0iJsvE0+CttmiuR5DDD4p70XLwD
j/qp2kSWOj/gDJVuZMzatMmIWemIcqlTVEggxIEysKoHQC6qbX0z7WNvitHAeWgW1ALo3y1YPSro
I5Mi32ltOc2JvCTrJFU+Wi7f9HXs8Ira1PtRKbjv6BvHExBf0hHYFyQ6dAgNQS51cWPlO8tksTiG
C9O/xa0zsPrnuViX8RVQJCvhM8wZ5zFWceVxv5e/UXLD7Sh325+izabrVorovtFfnk68k6AbPA74
ugePxjZd9tMJdngwc8XPFKFHq0e5hvRXr61mvb4lvnnmOzRiHJOYaN3oehTo8Hn1wZXpaa/fqssw
roK0pj9y7VxTMpxHxCpvSlXNd6fdgySwuu9fTPYhsqbti///vDh53Fb3PG9e02t0uODxBdVd1ie1
pZXFvxEC+JRd6WpsPfEJBdqG2lFbyokcg/nligJlQfJdS9s0C9Ivi0J7N3sElg8aAfu9Yuq51r2F
7jj9dB3/EqW7mgiWCy9nQHyF/uzNTJr+0p7AUL/FrWRyxG2KTr7pSPEOKFXRHGYt55fBxMxOGfui
HitN1/mv7OiwGW4dW0whi00DkvF/xtyyOMA81b6wFFscyO7yk99eo3UyWqeiqaX8FrYGp67gj7Dt
z96djdBzmtfhxOWeQVY+1oDFmfjms+fwqh0+IMjOABjhKnPct2F1+OmKUsLxKw84SuHH/fgIlXex
7c4vDSnoqCakEebIe81BxRdNdjyntdC6MQNY3IBz9tEelDCDyYDAikuMnWN0174CyaYpW8zh2muG
gMaW8FIDLyRDnD1hzjYFyTLcTM9t9xMuOhcKO2tWSUIMIpzdZwVzavfoXMqiMLFmxdZc8+pqtNqU
/PwSEa4zN6N5jYoZ9aTycCxDTefl+5yCJ8nX01quB1WAxNU3mf+cF2Br8/ZrScRR5a8bLWS4sSIl
o7zHcLFiqDGTEdYOD7Ti7biPVHAG+wzl2/dkLEjgnOQdEZ81A8X5I0XhoXjzuHXec9+qcZC1WwHO
xq3v60qLA1ZWaSQIoxCg9O9Xwmgmp0hCCGDrshFtpTBkXGcPCOnZAyWuCWv4lrpJcwN+22uRA4E3
xSANNlefLjnb3tVQz76OFJbl0/BtNf8rzJ5v9kIBEF0WQGbBOkpnlO+iwBowp97fnqLgEtqWyO5h
S/gIKYntgC4QXdSp1e/07ohW6Gr7dX5cf4n3P3bVTX6ES0WoJRftXKYi95dqbefnqo3olFpC6ssY
NbWBQYStyA+6URrId8/gphLeTpx6dFyyP6ixEiXAnMjkcXJhdIdvR6iqJZSlr9zapeOmcdFoqJxU
KZe/9K0UYSHGabq13v21yjGL8IgeltOL9WWHmvcqFP9G65dvuLh0Ky+Ti15eNxc4FLJDABEm6K7Q
vpRWpa/OLxUCwxePsD037bb21N1JU2X0NhkFjno9vutRZT9s7qxxWhtg5Q274xQnOi3Qp+IHOjoX
8vd2mnpu03pTdeatspX7UPn8ruV5tUnsl78USWEThFsfb8NcINyyCX0sLOQc7fOvSJY7QsIYawjh
IjGyZwHz0xd6pwFii1VYEIifdF9usx490wM3ihvlshj2GsIfSX8al0p49pMMzJCO43v0081Vxn68
NwX+cbl/hDVuy4NgbOPy59N19quV2kHx8ZHE+VMC9AmtAtrtbIvo2tMKZdk0K2xRWaMs77WuRa+M
s3g7W8vPstShQ7K23JSvH0PQMcwvUT3MZvWlLKnDyG2TLcSAdjjY6PUG2sZ7qZ0HfmyuOif/eqir
Q9Q+ZwdMLBPsL9bQGWln/pu5eG5dzANOy8Yr3C3hQLXcTOu4iCeG0Fyb/mRK+co9jIaj43QGYJz+
3LCNuEgAciNbenSGBVTz81V5DsCEnbnbrxfLMk1MXNTmGgc8UQrJwBT8UigJ6wT5Z+Wyvr+dovrZ
yg/x/2aXK5nJ46L59WVlJwocWrAS1t22mJYQ0eicGstXI38uksJRk+GSpZE90LQnF8C0IzXEZIdl
8A7HLQjjVwbhrW0rTxzCsOfQoYxgeeov3iARfFV/vMUVxfIvnVk7UzKde4IlCPHyg44COgVvFdYi
/BEQhxcfQ2RBOV9pTj+SHjnnNgOto+nwaFvRyaHuYZQX339BGO4d5MlpcXZPGTnTFSzQznzDuzgj
XKu7tmJrB4RZhFmQew742a+hV5g6U/UvJZafHn4n4noAokDGxnzEjpwDcyD/s3E7D+wGuNfmGEgj
vteJGNN21IZ1O6F0fsroPmRPjLNuLLzRmQlQigtQFVZ50GQrZcDltopRku1rB5AHDq3Bi4o5sZbo
PNjS5k/2X5vRKwxE1pYN+vLpT2FU6Uop3iKgPLiLL6WKvZSk7AeAWU8++Ez+CgIYqgPlySojqgyC
tkHKRZHswzfQSYN02PSWGEsF9BfTrhdBniZR1MpeGK1Sx5juSk57bvc2KKDkuYGo2M5yykVtm2qo
/IPzfzDzmgyUW+jFL9sER0huxN7/AslBm8sRcHd9LC2HNNpJgYjutdWv+reTsNnyZ6RQ6chceSQA
38cdVnzL+Xdf0tBNxX0AJPLFcRr+SbMvpa7jB0iz6s1aHdRMTkAaloTAI2ypfRTcP6KWAZfc/IOU
SkERzJfLXBtu4v3mHiSuJ1ckt/XkBqGiWdAYPNm2d9HmE48wF5WZ7xsWCXeAxf7Bq5saHA6+m3fC
X5rFbapXZZ6MWBii2YEdqPGVmMpIMEBAJ6CC6+r8CMXMHVO6PfWGB2FzULpHiXQMNKMqriTOXGgs
YplB+Xr0Pax7lGPQgd9PuP3bVtM+GysiSPtn8wn/Djt/KxHJH/Azzt/g8WX2g7T8LKa0YDSdo+VA
z4sYOCw20dwE43a0FazaNCsYbb+53KCnX37fGFDreaq4GP+3THssuV/e5Pr2pdydb+AIk+Vr1C9J
B4vaugtpFt9vRsSLVETkusfm7MjzieSWyFPByf3Yf1xPbhAG7uKXAcHb0ABr/xrgnOcmRqoYrtyc
hg6pmev51jtNJ7AEu3ldU4eD6YMfIi5drys/jHRmuW4JyzYAZpZFEymiifnVc6V/6Uh9FHO6LGFQ
3n4EgwKG8B1b6SxDskj/TVxKOV8Cbe7sy5RIWDQqEAZy/2oi47O3B6jG7iPGunpmPLaZ4jMlViNW
+aqljox0Xb/aTOSHGzp75hybQfK2xRLmJ9w2B0APd4tJyIFe6uVq9liQiGatR67eiCaAwmYFEXAB
4KnhXEDcwzfPr3b9zSMlqmxFplFBXdmOgKR2zw0ZdF3OmZSh2gqkK7H/7vF4BP/EfyXNS5M2yt/Z
1WjVjPdBgX+N1wHvCuYTRsi4PdRsBZVBEDxO3v54JgwMO4dktFhuUTBeVULHjRVLzyL88rxjOERZ
be1TkveezbXNAoOpJldAIYv6CN1CDsPCMYjMIt2rw0/s+b83MeCi4CdCqlz5XZTQQDrzpEIHTc0H
wzY0XSkc3xXvk0csl9U2+U4MPW9qXKkr6qwd3GEFAepUjW2+64R0HMIdqSVXYdrgRTQDvuckkLBt
NBoGT8r8xUiioxZOlJIP/ck0sfauJ/A4Ulfy1+5vTKMt/JjwMkd5Lgv7X/VGf1N70lvJ5TkPihmY
JEG7nKI1GIJ+qhxANV28SPBY1TAjwSRwlCEDNevrGGp91NRHnggE3UQWiO7w1qq8O95MYkF7OS4W
gt1dlKGw5I1PANN8LeII/B57aoPw1jlx269yvb0E05n9g8/QgmXn6Gh2Q834Sda/c4Ulmvo+R+wU
SuBx/hIbieh75uc59E4TivRravc/b5gdbj8H8kxySZdqChyMxVBPE1AE5f7cHJ1kP+zBQDkp08sd
xyeltc3FRyw0ZoS6pS84GOicN0anpk0VIkd9gk/L0T3ptNWYQCSO87uoHlCDRjaqChBMcqlCF1LY
Sk9YGRcoSEihzB/dTQFJ7w1Vgi+LrYC4VdXM5Kanl4wLxpGMVyPuGajvByt8q1FsKSWMP4mWgt23
dhgHsW6pmtcEKB7Zg9plrm4BPcQw0SjehDkDAWttD8zjCUdFT7SbsW5CHHZVzixAxqUOg9A5QJot
N9AB3J9dr/5EQfRSu0o5hXs29Mqcr4M5fae+4ykmIuwR69cvLrdLjEcwOTUqAl7w6T6fD9C3nJ7h
4Hyyf1nd5DFB9mzG8qzwCTeGBRC5vql4G5GB28ZKA3u7bZDDJ5LUDgnK+WyYEhL5Sxq3LcO+8Y04
G7Cl3PVu5Q1CwVh2kr4IIWutCTxKvzF38CRO6Zxmyhb/260xg8aEfyvNf9yPLepjJU97WItF9UpV
Yl4gb94+slY2ZjE17xthXeLmdAYs7WzmzJ7BiN0uhon6pz6P6pYzHcyTvKWdqxSlfy0N5l60YxEi
yqwKSezW+Quv+pnM8H0iF7UGnFImyG3dVEX5WqwyOoQYDGW+v1/XqH1G2g1kF/Wu3iaq0UUUwkbD
+b0/amE/fho/QRmgg64Uq5h6vRpjM7xmGTayweRFjYZNSrYwu47h3Z+1ory2eTn6umXG284JIgoC
HyPfWePYL8wGE5Pg+w4mWVMMqYSmD2xGtgixwf9R8gC+7Aqgt27Kh88ga2SuGkVR8rx37fObq+fv
krpNuWHSJMbCytxUWKUTC2xkzuYSRHGvVMGtRCjCN6IVjYiyizVJA2JzgRepoixQS/EUPORU9siU
ssF6kKtphQRivfteffXGJpojLRaRCnohsG+9sHw5dWk5j8t0i2i22tI7gkqIDe1gMvsN2P5M5T95
tFdr5ShzBwkq7TlO9sg7m/6K96XgVpGB5OvkVCAxqcZna0qj9GuxnJLv7qvVUGUu00aqbchNmWTR
9CXt2ypKjesTAVzJkbnFC6VcpTZErq2EnQGEV0zH3cO6W3uvlXRMOFxDBxm2oVBvMYTC+d9K3vL4
cKfsEVO67UsKcAVFXUupM5QZYJYvmJOyqXV+7mA+VOmWBBZNyjxGbI8DTvIvS3G2jJri29xkYcEO
B3XOL/FXZs4udNbnbrNWr7xtROyo2vH1pDM0sTXzsi0b85UeNC0Nm36oA02QSXH3rjItKwA8LmZF
JMJRhRM4+vVhp+tJEA5ULfv/ErJpLcPNrsvkFyzWJV1WK0IFqHOQCJM1vNUb11UYFLLne56m1sge
3km3vBQmi2uTEUM9oPcRFlkXsrcfj80Egp7feg+1yE5I44pHWC/1vrCDGN2HtFJxvKFYWMgjwe41
ja02/PeM22Px4OX8fqGuB6hexdvdNe6C+h0paI7FjRMmGLxV3qdBNOR/f9VWDzXT5kqbPmgL0Fyi
EyW+zD/AAL6C8s0Ew3zZjW3FuLge5d3OJ6Cn7mETgEDSKoCsBB2AqArYeVc+2C2dzkmGR89UkGK1
OckKCraJIEbhVTxwhCTWyRsHHY43Skd0y8aPd1Rh3JVu0jUkThqvVfxvQl+C4IGWwwtAZfNKmNCq
EzsjXCvTN4lCVKS/U9iG5UlD035n6eDjR0gMkONX1kqXxvsF27vk3g3H6+P/KyiCvOwvUT90RAG4
EjU7dgX+QLhM4CUoI6xIf2hijDUs3RBBild+cKGyOYIvC0ySFE/GrEjOxc4GQzOxVczQOgY5fdAa
pJK/hecNn7y/DF0ZUFwjcp533g9Cdoih489XlmLcZfRr3OQgLpoAbkyEREE2lfpMU9Iq1Q2vLOOb
sB5oJmL4287MEFMfBEQjJc2usdI28/nEOSZBTmKhw0gwmHDvNt7zCDPZJi8amMRtlTGcuoKyHDf+
DzrSpqEchZ/0OQ3PFRQJKByZsvkR1cO5m9Ia7mRJMbRRv0T4Ffx75z59Esm6+YKFLi/vnNR0lEa0
Axcl7B7gFVPQKbGQDgbi6CyY2VdgPMCG9JWDhiCcITL7ivlGILS9cdwZ8Pnsmcfcg1s+ufhWLO73
pvt4APmXcwzzGv+uXWrJy4ayBxWFZlcnf/u0xJmKrFmr6/ET4GEj7Bqps0e4aQ/clQ3dqvhQp+xT
GUmJDO1kN6rsXgpht9Hdu/l0NXkpTb7PQ0Udsbb+iuUwp7NY/DC0ygDT1vTSOfx1hbXwBjlKljMH
Nrrlg1shcYagmVo5a6erWfRDGzalHbVrxwkDoxL1JL9zor9S9mpqEQ+FLiQmJJm4ZGAt5+EinkJ2
h4cOoo2E1i+k2OlIB8KSpp7pbPyOw7XhTkiM4Ddi9P6deQ96Z141S+oXexXLZ2o0f9P+l8lwZMje
8J1cXrDoxDWY6AdzQ2SeQHmHAGkmutixcNX2RG46EnwQVzHk/vA6gdqUG7tRjHwvmXQcJcXktAgk
f4GeCnX3eV2a4UOIUEa52YORn+8gnST242e0drdZIuCq8/1p4bsmXEKKnwQLDpwW4hOw18zNlc3w
MLT9se8Iia7a7wZXioQWJ/nwcVZ/b1X6syusyzEucOCnRhIMN+TMJFZIeu2WwEUMyHcSKDQ0655x
9vTOloAVzf7MBerVVkUUaNGJyQmhNjpSwPiACWrUyVD63/SIZrNFGN8gc2XxZgecjE5w1ttgtJx8
v60cVx5iEDSRULmGiS17nVnae1eNQTLcK+BUY+CVckj7f0rjRGwD4iBLUkFOm7WtlrohBUs078pG
tIZWXYGDAU7la3SxoL94Da3OLM/a1Oq/VO86Z8M5qJ74i4gEebEX3mNg6l/F0Xs8eu2z3KUXchXV
BY7gyB/h16xC7rHZo3Hxm6TwKZ5WJlCln+YWcq4/neaEZVI/gLUzzoUaYfOjhJwc/y7KmTHE7Nph
p+Hl1/SzsQPFXNrjyHdeWSHBRN8ba/RX1c+Fa50nKJWE8X7L+ga/yaW8D50ngXZZWY8U1dQQDeoQ
Mtq5BdRUqC2ywvVxRCOQlggfKDebXwqMFJhrznBQOCgfTLOr8vpZh8nl+2fBX2YjUJCe10of9G2r
PY9O9MBCVkKPO1yaS37UzQTuZbsN2V74EzusbKEP/rbaarysdriKVCG4S60FYpNvoJkWzrKsqxzE
tCrH/qvDcyrYEds8lLVJTpjUU7D4OhZ4/vv52w0Ad9OCDZeHT8YPnVsYP0vJFvoQNgxDCh3FRdib
X1pxgrFcAf37CU5n8JsRa8JJSx0zRYt73ugwsnB+KltbP1ncBLgXYKqudeI5CIu3ik2IHGwwHGFh
fxYtNH4DcEMMME+2XlHltW06bNqoEMMMtTRckKgVwUDySxUsmOyO/xem6DoN6+6m+eg3ULYq+Wo6
ZHBeFCmRuskxp8dce0ejgiqMf4N9biIT9B4RCAQ24cxkxGyStDcTGvw16T/aD2BlIclB9S1DW7XU
5Yq2aCSnaO2nWGRryWN36ez1iPZNDloQjgaZhcCXURl3YwPiM6BvCBCayNTKqLxis11TDv9hIzGo
md4JjrTPaDjRo1FbKt6/jh9fTxpEBeXM2ngBg8jtrQoeCXfDl40yPszR1oZSBUOQaWstbP4wNjc4
S1z9MoV85KEVMGHnkro50m7uykGef9NofabSxIJO517AM7v7xoPwZLsBNPtWfYa1Z/gm/5gqBag3
NSEgSabUL5PX5NBUdgzlc6qFY7yYXVlDkyB91UjVeqSFle5WgeE56FHlqQvZasPvo6FuySxDcVwE
w0r0qjMZP67DrRVugUA7YJTHUcoXpV/597zspxRHXqVJg3oVG/mu0S26ulxuk6a+9pfF3A1X6b/Q
/5CY9RzfD9PZIxnh+DD7fw4S9UaJ633im0y791AqXW1FD1eJuyVIJOwEz5LJrVKxEJE3Ktagr8sN
BKsKBjSbm6I+C31yTjOVuTSmMKVl9bBkGt9ruDwLTCoA4M3erHsKGmNv0FqmzcmTS51xFvfKDxbK
TOEv4LMJiwAjrBAvMy6Py5DcpOnO2H6FUR6tOfGo4BCgLB6og6JiWVpsNmx2C7R/UXtT1iT+RDIT
eKGCXYoTp3vnKqwXkNGUg5sDXLeTSyszKYZYN8djw3MFHAwEgdMD6XwZrZm43lQwHzisltxRKcvQ
J7WQW+/h2wPUMl89uN76qQcyzjHwtIMMHUwXSAh236sUaXk/k0R69i2Gs8cQLgW0vS5zvNTrm+eU
owM+szcdaz833lYt0Wdkpjm4Q0XCLz6shtcTThCHN0iGcs5YvHrMCU1Hii+PNVCfd5a2sRYvlJQJ
5oKLA1GAWboMYYt188xep3OXkBn0unpKcDi0vrfrKYi5zshwOcT2HsA5CWHj8rq6XJo67AI6gLbK
Gq9hPBNA0ZRbRzq0viWdcqSHq59ggja42ByAcEGjSFhnSs1kfnq7QvPel3y0tN2pveXn3OHRMden
BRyA9xlznjWBJRO21KSsphZ8CdWFo1y3Cn3nsbKeUUolFfRijkqCOGCcHStj9KGjzX8yuvb4xqo/
ypt3X7qiUCvEeoFVE2ufBDnJEKOh4jP91uinoKgTgbq4KvgFYKXAuA40+CYcM08bXCXp3hWSztTF
um45Q8bwPVFx7p+f0uK8BQoBMz7bRIJITwmOLNVSCcWW1LNKx+AoheEYpLyjCycHOYgqFELgQg0G
ZIRYm9TRQE1MwMrcN+8iIPrELEm1Z2vMa2YS1rZ81rEcuIPiYSMHnN3QUE0UO392SzsS9sC+7qCi
2MIuri+VW3WbOaRHpGKydCUwm4tZGI3WB+715H0jsb1eaSdU1XvVEF7VSkPkb57iEamHIQuQgAd4
Dfmnr4W2EZVo5iD0NG5FSjxDTMUv/0lFnBEaINKVyNsEpdhI8nPbo9hRCu+JQY3tFrRtpWo9vaco
3vzbo6hyYAozXQIWnsTaQ7XfzrPZni0e+aMZRQ0Mf7fBit4sX27bPYq+LI7kleZj/svx2o0HFD5h
LVOkSw349Z7uuIM5rnEr+93u15zb40rigsdU8q340RiEeOUIQLZ5djyIm/o2xYb57E3EHvJ8Gya9
wQKY5VulUjeFCbxp1tjW4TeH7tLNYNqdOpiAtQ7mMb78btiojLFVWXPrY2ri58hL6P4U/+GhZFFl
pA08cuM9Mp1ZXr1oarSV9LDjjRAPxkTEpVSSxlRH5Ea6pF6sjoLAD3dei9MCa6vZsRAwCPWt0GhU
u0LPKGFiDwg0yxeESgk/JF80vDb+Yu7/MoHk8s8TJzZSauMTmVlHa2z57BAZMxQ7Ibf4V16S08Ih
b2TLY4HqfZbaGBlGC0P6ZcMjbevGFkovJ8TOhG9ndhZ7yuM/xrJL/r5kbLjK9yeEx8AiRqnLcslC
XQRP1joF6ZxccQBeaQcY90QMXm1SpVPvJEMoCqn0cnVkea6eajx+fTwOzjx0/R9bs9TS4HdWS+de
OyEThSPuN3zX83KxofKzlx5+KATwR3iKF//YqbfZaF2Syt09agktb+tqTD+N4poumQu3/kndhgZB
AnxZMmkDRuDEe6RyGMCaJQFeQpVQGjQw4uBKQeX8T5t9CEr3RNw9CxoZKVupX0NVYuv6m28X5QL4
nxcqQeRHkZcdLiKHERDp8vrvd+yWxssXKPz/u1FVdNh2LJALrcksD2ipgtEDUmDaDTjnhAZOMzKX
ydu0i0YKnnxQa4IOWYLY+qO/evhqMAGUN5b8/edRpKhFHTIk0+FS0O13TtX1zMz9VlOpBZrjmWA9
qDq/L9E0TkrvawwiO3IFo/3FQVjRhgIEfdegK0YxI9BcKnxbqtTZo441mMbc3jFdoDX+oFiAj2EP
cyW/Hkb3CwIdBo2R0MxAT/sCIMcIEc3Nos4dGywx8gM2PyrOPqxvRDSz3AxnA+gBJcEPHfTBpkGq
ZMmfkZ4ZbLPKRntGEYnhRL2I6WIINJ31Ft5umrT6ZXMBfIImQnEMhZs18H2SZdx4gMK1FI6e0P2J
x/JgKGRgXvdtI02Ggs8ZGdWQoF4IUWlqN1uPsxP60UmNNFVWoyPDGVPZEsON1yVP9M9QJ1qShHYf
JPXmRW6ANXfwIrWPmbwitk9C07xX3AizeSylWd04rnT+JlPlYJGAKlIHKlVPLdeymng7skwD6d8I
iZnBBl2p/BNxjSXZAyXHUx8ggokHA+PKO9zcut7D9jfY3TwaOgQfmvoAmIMj2TYW/v5jGub6z9M4
o/IkcTAWaHP3DM9YGND8lBiseniHuG7odZ0d4yo0qEfa5Q/LZMkNTQTv2IauARb9NtoOk0JpEILO
t981Qt6U3hkqJ+6qHI1sWw+ec0G9osHELF6kcIQekXphxrKUm1XP0tXu4kz2fkPSQTTo+c3imdGM
jjHTMsBsXTh3P7j6u4Qeqa85/6HhRCUHr1s02C36NRVjVLGe5d1IAp2iFVoQcMQXWbfQmkmT0Pxm
lrzr5IJKWALvpu94qSS0VhfJOD7Zgsk1bIckDYyqStbT2BE/8u3mgXHSQyPbH1/VCXCc+rQTTOD8
FYpkfh9kSF4BBV8hvf7sTH1TLKNUvF3sZPSumJqzRQUqVuiupJkCWWAi9kgERMsdt7633Ou0omuE
c8IhOW6lQSHL9kEfkFC5ctwKARH1zYoyxdn+ez1bSwO80hqUxfUkDSED2sB12tuEwdbM3T1FcUkb
8xrIqfTawgh2rrHZzfW897bsHPf4++0KsEUBkeo7hOz53c8L5xLAQuLdpHmOz4GhkpVzywdq19u8
onF90FsKcFXEbOyvu6QwdZlL27MixCZEGesXw5XsGUO4gHJeKvp02/NK2rJUIrQVGHChGGsl0elu
OiLBuyubanxeL+OUhJ39aJKUpVXOZP4cjj3uh8ZYvl/CzID64byNPrud+QTPHlIAjKmeZyjjx1k6
BBuMUJ9z6It1/BmtNerOGct51VLW3L5Ms5WUoLdPSGKtbS7uaF64pE9TB6IbH2X/RBKEpAjKJ02f
WVYKoMnFHSRjN6V9m9jRD+SUFxm5wZb12RIcuEIXlmWhrH1CvV00lysqFvjLfDtOxD/YJBNicUtl
LTV949vuNGzua55+RO1WsZV9PnqTw0C1KiZbaluXojHyECPOiQJAWJVPAIMtKHe5qL6xEQ53/0uC
sRPtcwE0NpmUi2GGR6MCv+mRAmRYGP3nh611xfTjZ18YGwLkI5ybBJsoFkCrsWyzP/jnzVQVBlpk
jQ1u3o5hsdI9m5ebnkDk78hs5BYiohbbEP/OiNLc4N77aQhVhTrmnv7lo6LcbjbIw3KeQfbsmzfl
0E8dJx/WGqJ9Z463gmEOgIrBTZ8fseDTv/2xF4lpAHTEZm+QWKJtHiixCHwM8+QmCF9zv0KmViRG
MdHtzs80WUyynwuB+oFST6U6fe2eGDvYT++PGofyzlBZsCqIGOqSy3SwkGeCWsjbV57UMTaJQTD9
Bpqb036zi5PqUJeCP+3Q9Lr8FzGr8VnQDpvjRpBALjV4Avcyfw9iRS5ih4XsJjflweyGtZZ46GvT
aEDUuZB2AqTLVHIsPKZ2IElsI3qRduuezxSg0cCHG/iXMopw3LxmLfimyqNMIMdsxj8RYSDCjUe1
Psi982Xyu2ndL98XHma7RtinzAWv5Pg22/Tkid6dVkYhrZ+Uk4JsOAhED3j9hJR7g292nUnE6oWB
tdeeaVU3BsdxAObxU16JErMe7WbmGm8X5G9JAjdtNfB6cnl7KD+bvhgEQqOERUpg5TQjbTffVBxs
jEHvvVpUwl/FubwI0x6tNzE9VeufPlvgLVI22GO3U5ufH7vvHJMUajpZ1om844I39K+/Om+h0pKI
oz5B6oVFd4C90Xk0JK/fjvSS4m+Bvg+L7adexcKCqT7Hh1doky3r/4NDRjclQZ7UTIBDYMHECXVD
dDP4xySCs7OzKY8n/ntN//pgI8DjVoKGLQZgImU2O5vo+QxkF1iEL8YBKvZIbWT/ChpPWZMWbU6M
V+rgsdEWFYqnLCrx3KB/14tGgxxjYdbNjpXc5u+pg/AVXxVIbVhAG2/LOcyCGQ8G5fa/BUr+sNsJ
9FNbD2S/lNkcTKa4tP9HzNCH4dgfraHfo/+zwXA/bW9w/PJIhuxDLyuwq8DoZbasAFPLvP6PcFqT
AX0lHMuP/paDPiUA1qFs3KDM89xw8W47dvT5/bU/tSS8DKhCIT/U05iSxoH3Ga0dkU883UKsiQDG
VcLn55QuI3hUNjaFmtGP8OQV+zjjg8AqvY4V25aEt0JuH5LkX11zTAVb7DK+TFuS1QzG1zvyZ0zL
AcLAq+TWd7y/kCmoHsGzyO0mcCye/AgqymhyhK4m5t67uow9DgOigBAawa9gHwnTNRVFvdGFrXAQ
FD+gYiTolzskwsZQnMyGl5hqH7ET0cA75I/pzTd/J27CsJ2nxsg/nLpT2rsrX5NXhXqdkMwCsqPm
TLeHJIiUGuDDFmmoUUR5NlwpasfDAHqDTsJFsvBR8DSvDmZTETu5Nf9BHFWGum9Ayr6RZP8jTVrN
Rf5xSLcigxjxTSrUoEqMO6Drv5LlMDWrSR+ZTszxAIXBYhqPFUGIBrV/7b4rJHMXxwq/RIzKpzQM
HzR8ad9LUXtoJVdv23luSzNqlXRa5FvTtFksolrpbT6E041RTM+GD3zHQfYvNqFKQgczTZ8IOnvk
PU3frB0v7PlboMq7px+YSZDI19ejk7U0IKscsIbGigCx1t/oy76cc+kmp1khJXUoZ2aGRILt3/NP
0lZAtJacKFonWYM2mNOGEIRaVcxL4wvTWZw+8TOMVMLKwcP1HdqDVdh8w3fQwyCmIeqKLwkG/FRG
7k51k3AeGcTsX0vDLPmZR9ZC0Z/AOsQGIkGbTG/CVKcECyzSHUuOkdJKSnP+pWpb3ASK21QJIXzn
/ye5HKL3mUQE48Z1U0FoCf06fQq7S7IBqrKa6bGRL/wA1Ioplj8zzXxz5OBLxSyZc5RTibYlM0XC
7qKIgRiQDNFV0GuR1hcMQSwLZVaG6QrxD+PQUkplFNa5bvul4x1qV9bo3/KxAGLwvZ4yTyKowShl
Ppdxcj52angBAy1T4IXeuZxRfPuONEXngzSKIwGNZDGuL1LKHaZJDgrGXp6p+bSCmE6rLbBUv5KL
k81g5BhA+9z6AeUR98lJmUxp/UCju0Z2qvHBCCW2ZQzXRwdvzEBWpUAHHu7b4RXPP7XxLSbch6js
VGR34U8Yhf0VZiEsqlXVpbTjvbampT9+7zsGqZCvU6m2rHY9FaUqlemKTKi5ykE2HbkJQfnoeFZ5
n0MimOEWEY4MVK15W8evKCh0C/CTc9tok7rPIMNGp3+iSMgy1ZwOn1rCC9kFFfT5Q0RqPLyoG6DT
PmE7+8FONjcod/rWwiMVs2GRsotILIU9cbFRh23MtBpdl65zx9WM8EYr5kCSpGX/RbociNphJ8sS
KfYZZLbEa5y20cSrsdG3jlsQ/JGe3K13vZyU0Akdv/wpiSzWoIO70GOxiZJzSG8TIkWU/csABxau
Rs+e5syJH0dFx8sTn7SsyyTKuwHpuTObS9SkvoAGfIvljBUJQTqR3QINxKUo2D8J3QNdkOefSXJU
HCGYpE2njecdQsBjwxIB8O3oy/9dX5pts+FrHpVyf0IETerDzwhD1zHAc3uv7FtLiNz0ykKluD2S
8LAVayWceTUSxi1aOga7gwU5xYzi1Nt3mcS5hCtYwG1apWN7bE3AHl2nBVBnE8eAjr4/kiMwTO/Q
8HksVE2zdEBFDuJ5Yuk5ME0Z4wtAOA+c8RIko7KUHMpaF1W4XpYpdORhS5TOLXbkl6ZskhVWly4M
u74WF0np41qoZX7fxlpTMRqs5YBgxB8HRez8jS7OdxEVbZ2OI+oU6PvFP761ebOt0q8NwgbwSLoC
aq+K5rDP4PUGsCz7FXoTtaN99Ohp3DEHye1gCp8YKbdIJAjjfedysFvsNk9j1LgRQONkgcHx/Rmi
RSz3meec5EKHPgA5betpul5LL1Wf+dDfyQIq59vY0p9y0SYqf3m6M/a9UPGLlMwc/+PKO/3BIVJl
m4YRChsP/TelaE9XJ1VqvtzNumVFOP1IjmMNhz8rbxK71lsm6h0zLhq1ByKRbAYVZY8kMpVEyUvT
uZi3wR7oOV9ZIRXEXWQ14bIW++RMTESbFDd3eyNlSeLEwOaAjjyRceSKeuwpPqQtfI9EtPQMUkK7
n8GtDxO0OxVldb0wg28QcldIMFkB3skBojm0I/JnOEKewki+hOJdQvI2vCvlEd3HTSnk7pVELDkC
1HViiTgkhRKo0IZLYul6/8zKgohatoBFq02qYU2j8Yol+slOLL8GkRopYyL7XdEUn8Xd1+N2GCBb
pt3M7axS4VYcP7rSKnLQBCU5tSqDFJdC6xJzoW3XbN/IvYrpEcdLiFenVFS8mqda5R1PdkvKl9Zb
MZfOWJcQoSZEhtlZuDR94YDkjxh3tPocKC324+DsJntSBVtLwAZiHRfn+Dtspz8r1/AQwOT4EasK
GCCkL7EvczOIV0xickRaWxd1zkVuxEaYx/qNm1SxDlWLVPm6JdK2Seb9oxHsjbhlezsFBdv4gROt
g/r4CSNo9vz+bP/beJwr7C/AMQ73wZHXIVjIEbbPRkOMGkm4gSw+qha9NyhQb4KIJLNG1XjJ602g
Mgzfl/wgjDpzqgmP5n7iCff7j9JCTm0y4ppKRb3D5B08QQ9fYNeGzlhfV+RHn4Mg1LOip83cdpd2
eZF5E1O3Opgo6o6f7xQpTJY9hm0a8DHM+J18k9Eh+N4Xsa4OixNpo9hy80VHqUeoxXAFWaAF/qIt
+arhmtbN4aVMTNQzIG0qg17DQ1nVODq8alGfQsfiuNwPby7cwAb0saCK1rfrK6rfqpzcQqFmt0jV
9R0YeNQkQvdX3wOxZV0EhWJ/x8drpKWbpDlaErMBYMq1qQGABH74I+viN0PUn+sSks1m093XDw8t
jr3RNJjiOhrwHqkcJC7SEVza6x17kwIEgQLy30JET1M4rOH7nybI8RrhBvzVX2fnf8YhrUGsezx1
9k62rKH2P0ZRRHTHZMi7K05FCTj3A9HPvNUwRwS8In4xIHyEhub9zv1PlPkOiVzv4aO0G542SAXK
lRe9C8FjMXfY6d0ueHK54kiRpFbLGDMjLtZ8tmJ4erP4MfCdEYStv8vhYY44JPv9G9mkhPaMMgHW
tCBkd0tQ3/sSh9hAwcOQf3UnT1uDjsVUkd//M30oaHw1nZg639MLsf1qZSR4vneX7mBQgsbI51h0
UxbUpoZtuzuYR7KV9IGyVF1TfEgITBwpTs+vX9E3bG7w9L6j+MW5FvbvHvQsy9E9FEdvoZmpxkdG
Jq9jo5cY6zcUyFdFhovI2UXaDokv8KNnI0+MRmdgiHrlGjfednycWedhOVkdTCgDnEP5X/jUtG3h
j5kSmLAW2zLZqvJLCi2gEuxnBGgUSIPL7GxVy/Y0o4Sbu5ebBOxZ0RGFu3nP6MIfuY0jQZEpurTX
XZxrRqgUp4SaE9Mxz606NYaJHGTK3l35v6yGRtY6SfvlA6TRgPuRdhih+vzOntLO12ka6qmyp6Fx
lOEX/Zf/Vl5iFTG3R2QkKYaKN5YTBzu7rvmiLMB1n8Z+LuaAebYr10G28Q2hIQQgbnMu14b41vxV
p7KyqHGj1E7rHRPSVEFBfX7lVJfJ1AUQ8sZ+r3qM+EEAQgWk0CZ2YWg+ssRGLou47mAmgncYxMkl
aBhH4K5UlfCGk9QxdEgyWqHyL3Loyxyz/mKscWj1eozgFpLoAXxB8ECl6cvGqZ8LXnISMil7tMsq
jstf8Z76LdqgZfTTbe6edHUf2RhPfVyZbEMO+kb9QTTSs4WLyVAz0WpHxcEqU58l66uWuLPt3dE1
ZN2ELPtq250Ze3KyPsR58cOdm8aqeWYFjMkAUR0QUu+nDr75pHRaSmDFsNlu8ulT6XLdxE6BDTXY
j2ozhFBaDIRK3KORNYXb+svoDYw692B5JLifLz20B/OWT2dt9rfr3Xy+YL0qsTY2VZrWVYJkHVnB
PbeJOG6SWYMh7gtdEzbuagJVOG0Hi8Xl0o/YhdS4WZQzMYQEsbKbLQ84O9NAqiJUNyx9kLPmn6sB
RE7YPFSBs7lqUDJPt1MZPxtcsw6fw1Koiw8aOZUk0mu2yHugOQKZy9fahQy8ToCo2iAVL08fFk5+
H2wKl4XUagBxiVUKzyNT9BCWGFMFMb8+KXLYOQXt/UfUVyWoO878bJdztITGSC5iqiZercIMQly0
j8RaaqZ4cNk9OhVNXpRop8Ehf0oCeoNZJ+MZQFGo8szk24ucGoK1E4QKNT/ye0TRQbY/oDjlE/Fp
6dBN9Bb4rmpmEYtBhnyoH+wEl/du2JmFqGzFCfEAochX87bLi1jAbFL/EzHdhxuhOwG0vtTtLOuQ
56kYERWmEkWGhZifnoAJbX+DeKI4+uy8VoWpHB13UsuEF26DtOM5KEXgQySdMcm4MKNmy9fxpFsY
R22pu/5bkQODZHHYL9kz2GmVp6I30dvtauTzc+WbgZzqJ1EJi8t8jaZCgb9IR4c3zNq7l6h8eHUH
Vy1P1lxdab6PiTXm1yc1FSVT44Q9bYNHVSABw0RyTDOxrbJKJ930zQ9BWjspvxPM5lY6bYgfw8eo
aCDf2elET/hgIR/GSDvgg2LPbkyyb4OAObHU3OUeZwdeJz/cuJmBJpzyJyNgSXLFNR46yksoFx67
juGT9E4YeaRMMq5OHz6CoO+7Zaiw9d5e+QxKVXw8ufmAtmnyt8d507Kv9v/XmBW6zuIMdo8tPrLY
Az0TfHmkPalTOc8vWK+XNexbaG4XIZbbmO216CvfbCBppyeAjKrOTxO2h3iK9RjQjG9WSn8XObNs
xo12LCch7yARGgcJYDPslMuwnuxMqt4fmgD75fgo/wXAmpOOf+aKKpU21g67zqbl+Hs5H8tDRKVb
Yu5GsPb4uiJjOOLuPrrkEU5xOdTlNp+vDYu6Zzl3VMHzRcBIM0V85fhkjumVYjy5Vq0HYgQSPy+A
OBF/gxzdy84cVaRGJyn84commkK1wx1YD0okxwBqQNWKdCaX2Y3y6/WMj6Tj4GfAyTeV0teJ6So4
NvSS+UFSBWzncKXFJevDKkvLQOuRE9NZHkTihqpktGwXlx40tCbCjkbOzqxvKp89DSaTjJNTzdPS
ygwdP6RpPzlgHsYAe9cMqPwLnF9sW5oBmWUZ8MA7qlWxuzoVGkKcD5C9ydDKDb8ixRnam1NSFuyo
MDAtYLe9w/nh8mBRW/hfoLDrjZyM1uVGwjnvRAOGCDBHozGklu26OhwuwJtal/NTDM31Ciz9L0/y
vw5gdT3RsLinnzvKXRLsgCPGhtUhDRu/YVPX/aCqEJMbxeH3WaH9wZu67YVJdQhmKi2xtEFUOz7H
rPTcULYMNk6i+qA+FkCdu75Hr1lByhSPuFNZxoLHY64Au8pi0sUvCkCuSBIhAEvwQ823j6PqVrze
UbifyjG6E0Zt6e9miaXQuDfu7bXxXMHiJxtNRapunlYW5Q1uA8CbwFNgzCSmjMCtgwEdQkKR3NXE
s2bqe9FA+oGIgMihj+9ufN5oGwpBUfRVu1LHLaaoUuuK051JXwBFdGUFg2I3CLs6f165f3IZY27v
eQQ9+rW12ANL9I29h2vg8JMieNU1zhrAYlSoLKl6IRfnXP2Rmm5gyPPx0MqCrtUSlAItuGU0H065
9eDsGj96Sph2/g0fxr/uUuC/wmtfCM3t2O/hzWC155TpXzRKaeFA/pCaiUqh00taGclf9TXW8/mm
8LwX8O/zn0ObU5dhABTtMP3M73bqZ98xiUr043TVYqzkmhQFgaOkXH4R6M5tq62ufe/ZMuqgFVk9
ExvRJyZE0lDifIccE9Oek8MfxTK4nBnabosRBdJ94kg5ydW1Th+WBcj5gwauXAa4L5p2/YHl60Q0
PeQyK12YINm+RvWGST3WAYd/1QGIUUoQL7o51505cp6HA89kV1I/c8TRFC5ai+gst2Z5sGa3kH1a
A8oE//mf8SLvCPVvCqeJXB90RF7JDedI4z4iwHjGtVEZFiVyBvWPLJsWdmk9e6JmP8IwfQp7Zkj/
VKbjnFyVHAXECd/05IVfiVk3dYo91OVyWUlniW9zHii6cW7uuZhiijohTh3cHZVzdTW2w/35hEd+
6oBondTfACuTDL7A+F4Qpz7bMMtDnUOy3MlEr3GhNRUDcdniaXPgIPdR74bVeHADECOxFP4F2O34
ngxK/OhfFAvDBLeqq4aZ+3aPDybxz1GoIbdlJyY2HValau7WBQlUKu9L7zA1PKaOB44FIlNgyVi9
bJP6pMZavOLJxzVb67TyKyU7zbmhMRAFyrWPWeLaiM3gWmIQ12tlcy3e8AEJGzNSczlZjCNwhBQl
Vic6GVcCeCYlPnqyWlkLpARfV8/tlpfYUsnOvhdpg+HLvaSjvoh+Omfzzg5yvQWZxAVoyFIbWWyf
zm1Ovga0I7fD1S7y4T5RMQ4h8QhfzFTF/JT+r7xdLdf5q2Nx46rEil5FQ3nzRoExLUTRAWIaUQzz
ZA0mcAxSo7UZbkEeclTxdknRnZI9v58QAZWYMRre6CDGIucRYiLk0h7RssWgfo4/NxMDLWY5ucQl
FnBlullAfUu9Fv6ZqE2fGrgri7YI23pKKaHqVaQGb18cSTjvXQ2TNOt/m7Q5z0yhRN1DI30VMUSS
z/25PBnVCL7M6Uvs+FaDWATH8H/IPQnsjLAyOSphMbEdCNA47shh+mCIX8ewMrFXiaQ9Mo1bqP2g
vgdoigwKkzxaWtuZQ2C23NCGyFQWz2tHyQeKsKlR79f72lkY5lfMn3dOmZJ3KzpZHk2Uaow5AZCe
STIm1TQXLqUxb1O+IqYwYehOBd6wuoXztpfyDNIDN07NPtvCPrBlq+oNZFRWsaTsehn8UKNrYG9W
9qNW0kjouGgLfYv3nr70jlpNYCPl+TPam6mL8X1lmSAdArCLEt8KVH0guorHChg6AEB3yahTLqXq
iPO+ZGxJel0aYxCtsKnlrKaEyhBS4A3mdxMr3vzHgLlwlc4X9ElvBp0TLN1H/7Gxoqu0ZUFAtRa4
Szv+YndDi/d3IHanCj4NYu1VwaB71YAGI2C5CQWs9mzjoyKsYq4m7LpIIvy4iHKe925IyGgYmoK1
p6tXgVuIRZlYWQaCE5mS6cfIsgQteWhxeeT/XuzF91JLcs/EHCQEjG6w/NoAy+MiVxKyxyHQeuuJ
yUyvxR2gphmyr+GSxRDAWUg7XZH8IWAcyacvWpHEncEcLVzTXwJ62rfruxVyZL3fLaa3d0O2glWT
IHlAXW6a+O7eF4fLlcdTp0PHA1JG9RlU3nbPe4X8moCIx03XnEUMX9zZYg5xaNclvjeCdG25855Y
9x52Q0aP0afEg1WGSMbGi4/TTdmR3BlMirmf4VYY5EE+017kuDmT1XFzTvQn7Uriy8iOMXywzQjD
FwmLBfoyaiAjsoXVgJloDqh7gZjCPy1lZDRc4tNo+E9ryiqoXvk+QVul5N91prCvIHbJecABtEso
ahcMOk+PacEp5vjckJFAg8myj7OxKdSOBfrw3GTfdmpRNyaNKcqiz55KUPwWSLv2CLUFynPuYnBs
mMiEUqW3UcXQpZhLW6wuTltoxnqXFqZne6PxX6Rg6aH5AZMOWhsVDzSHMOgsd8IN7A1QPub7Vu2h
KzB9llRT4z31KC9OBJ6vgcjtSiz45zOTEGjEaEWDP895L1OMJ8/rB5vplk+TOZD7gA20zgoArPad
StH+mGmrxPUMhYvSSN3IePbkiyJNtXZsGWz/bSkHOdwm5Li9yX2WfMd8QcbE+5Ld2O757LLp4LvT
1WO0M1mcBlWuseCCVdqOPgoUl7vFbNSlLAX39cLit5pKy/F2dsVXyZAaXGbIl9+m8JorSDpJa8OE
znT2t04QArs2Wtlfd5whrIYsL4MLjo6DFrz70yHHpYtdwlX/4myiLRuOSrBgFY+RTxfb/Rmh6gj7
TqbkxNJxe9ITxwtUTAJrgdlZghy0NUlegL7Pe5U+lilzmDZBgYe1dqahSxLHZ4RXQEbqLlb5Dant
TUfTr5hS100KxFjoolQXiRHMm15aqbZq7W0D/pU8oJCNldOY5cY+3rg2O579YlJ57UhjdaZj57Dq
UbJRhqd/T03x5+959jmw3sEzO22qeBVYBeLIlI87HuOEWdDovxTUV/Wxnd+NXmD+hseiO6pX8gvL
vyTUMmGdFB32CgMCzF0m+8f1GhB/wRnL8x2B7cDogZzTC0FZBwdcNXv1uH7BwDvuD+FYQTE/Nlbe
zhnTTu2tV2zhozckABYr2D/eYfSF6/mu6nl6q5TTg2c0YAqj8z3h78SEpju+DgoTTdPCRAMeKeuD
DSs+pdRiIahHrZfhGKqpt1kx0IQP/nWoYTrkEk/T2sJPkSuVsI3j5LA6uqwrN2cVK0wacsu0l4SO
6aGwSIJyCCopcFQdu2ofcb/IAFf9Z+hFc+as0mLpCQ+k+uKsgdk2xXjzxnf6t7LN9KiFobkfsQ+s
XnLODcb73s2XcqewlQpIejOWk+osnFoBDmlQaSp/TMml9d81mjz9kqH848w33Tm997WtNTMLyM1H
996WUlcwefKy/Lbz2sITg8Il6uAhX9lgBKi4Vw0xscy3ZEs/h63Plszdj9RvgEQkeaqNuQD6MhhC
QPzd27RYqL8qmXOfr8lzrEjlLGwCIp6+lQ+XywPYFNysrXGDUEia0yZMvTuq5yqUdruZn7pz99kE
mnO+eVWsbGTEA3Ivm8ZFlyaCLl5WA9htlJhBZzRVQZbgzs1UDLC1K/XhjDbFn6YS6h3ip48IrrXz
V87R2HawE748H3f4NbqhSVa2YpNq0r4QMWd9+grfwHd0yirK+ghx3+Nw0kiSTuLXbrj4ewu+AVSR
HLKKTiFURv3bcfcpB8OJW6A4WIq06V0CxBQMMNhguMJOKhGBT+cxeVEUJgoIv91+n41AmC+uedgD
gEdbQI6Alyt7Pt8iwvQNsbswgQ6xLbOksT5RGES0tKGBs/bnhTN2LxCTkaUNRaVmaE3bq1p4Qvsy
hDcqIl/NgwWCLEEkSSg5hcEh/o34y1yNG3cicGprWFN3ZiJcy5eTxl5qFWPebEFOzQ36eElisJfI
fMxp8h5ms1CKIPBzpnvdfSyYjTTRVaHJL04CHL2MxgNT/t/bNe+pDohWV/AHuZai4n1wxJG/2dMc
U0g2MnHZYINCX49s1eMyxfl4KHUNwwtWKzhQ+GnGYQ5tZuHU0soQn6nDFBnUknSj2Oqq0gUp/Zh3
BXoycMiMNQd2qXArvHmp731W406dUPgQZRUpSjM7L4/IjU6D3wqziAr0G2BasrKGnvPVWzkLT/mP
CjITdyw6gIJqG9tyLEWp/cvSdgFnU9tUZjHXMUQ2YVXF4T6ZEReuxa5VPkILpENgpiRMbnCzG6sc
tO0wwpxpgIzJnEV91H0pw2HeEOlLOVzBp6W4JIMiLZ3Dk+USPAOOAXykMNVuUy8I3wWmRpajhNfw
bDdhJYegUEwxObzz+cP8wgk58qK5Zguw3rFa5UEfgHuCI51If8yl8yJ++BaNC+QJjBmLpfp4HMFd
TIIkc96djdUzKQWVUwADRtrIhkPvHzo0pNRTTe2IpEN2EuD55UZhcp3oQA4fpVmNhB1gy1waiIKy
AMT2b7gvb5uAfbLFqJk7hG7pVONHN5CxvaXXp8lGRaPJ1sKQAgR0Ni8MEHcWO+MWPg0dAMT3cEwA
7MchSFojj7V2SJ/wt+SV8dp3m0jlpUESqgpsOz/z/qFZUkjnwl0kNLjFpHrrF8r7zUKDZCyJrZFx
OAjc+jhPl/l4/vuxfFDIYbmLiwd6L4SpGL5M28k0IRoaLlg6tAi/2+nqcxsf7Q1tHKu9pTzXyJvF
eEw9+carEzWg2uMnxtN3vIVQYrytoz+sw6FFtNvwsWJokSq71XV/RSDJPB4su5Ho42corXAqgqCz
1i7tzmZhn2B8K7QnExnYsmw14avCh4AhyL8RGEdxkw7dh4a9w1FcLR9taBkVIeAKvJNmA2mNif1/
kyhJEFmOTxwkqT9gtROedgF908iyFbw/tYK7bSCi7e0mO9y5AERb6nSYeqO0qW11o7FoNsGVHFiF
FCUjClJeEBj4GFN66Lw4k5fhYCBY1l1hQlXLlr49ieWNGbynvyHrl8KGYnbESd4iBFQSiwq6mgfv
iodFnAyylPZgdrmRRPhBygB8g1wYagfAacMqXD5h07Vkjsf53D0OK2/xipsI6PSySlidMTOLmdaB
blPBNTn0cJIIhrWmQ8Bip54nIEH12J3BX70zKvq+8U22ySFngCwek+wXQzeqwQKsTlXkTTH7WglE
2rgiCzsJiyOu/GwFJgNpj402t7sXpRFQczwOptCKDFF07XjIptIJTN1CFWrEPJ3G+AMeHVi2Oacm
7axaMaeXnPyjkOkAL7Sw59ZPZmf48IpeTR1Ai820lKlnIR8OyVgL+bQxIOeDZDN3FYhWlcr8R+pl
J6PmhvbsDaBxqzv/+jb0EpPWb/I3fmLS9paTeHttdfVhZMFOiPiAKu0TXIzbniHsZ4JNEC3OTOvW
FRW/tWL15bxTw+bRqdrdfNI8KgysRw++bopxrm//Hf6hWAQaHRgoCIHAx3UtYQu+Oiw3AxXb/LYZ
qDXCV/09HD+AhvndQubUt3vgmLPl+M8bMP7WQRqd2pIOiy9HCBIMpS9Lh6HdjrEBe8AP4ytZ3iZR
Cz4Shjuwkr/b4zyigbyR/8go8yjVnlTX1Y6/zFdmafqhueUd6BAqQ8CEf3pmRRcfL182FHInuGXG
+wRSNeyCVbe2DfhbOjNPZVkUCcSTxKgBDOumnN8uAcbttGMvbjRsrgKh1xxUQWvfd+ni5ysM0z/4
uw/JyFd944VKkTmQoheT3wz053eD1hg6vjeGn8cfQ+LszEkwDRgbzrdOJlfCb16TSlQDZ+OVn6wf
V6L6sFVbKfDunm9i30KkyREgJxwhvsgkK17HTLDnqM4ZdPAcIkcnR/YnZMczuMflXA5BdzfN1u32
WcPDdmhkt1UFzG/CPPmC55t8gg51K3eC7pNNsZ9MsQ9b18N7N9ZdtfxYs6+wXzpOePZRjL4mapYy
Ny25OJe6GoqW7mWm95vOj43OZIsJZU5ESRr7Hqi1j1D20yddBghZoNjFLzLha3nG4zu6SZXQ5DM5
SvbpWXMxxsFUUdixCxn8/uXUTqHGIWyeZV9sc/6Sbef6lh0YNLElLJI+VD8qMChfckonu2GxVpjr
OsHjmjugJf7m/zsXXTTx7PiZh70sjmwgM858zmkz5f/R+g8YenR7vBv6Pz7BZFqgnCyfwVuoVjPV
TdFZu1ncbNbE2Luo8HXUpCgt4SbwtATuMWuQT6d0lA2sadx8cF6tu9phjIrtCiEIR28MzGuCMYGf
YXC83qHhxskFEwl2dlChVsJGPqQaQpoBTRtLyeGvikwshf2y5ky3Izf4lfsp/ighpuVzG7tqvVRZ
BBUCk5wwEvfjVEGK08QHsWbLg9yNiPQr0SOJwCdD/G2PpS/CL+o1YlGlwmR2bSHZYazmJyrACkkv
5xuz/XbVIbFpcwtrZimXawlv/h99JMebgYgVNeZVNM+rb1Sc+n5pnFmBRyN33oGURBwWtH+j2Ady
+v7teUNGu52PacrAEQwiZd2C1hGR3jkJ1bCs5WkjmLgPJutpzwED1sxeK0JTDN0hZcSevTHLAff/
pzmGWNK/YadXiOvv+bZ8V1g7SPbq4dWxnGC4oJ1bA8608be0+VdIkF4DnOk+NKF+e2ypVAYLV7O6
yiDdVqgp7OZjgrHtU/Rsw/KuiFzLArClEetL3d5ihNcwov62G2SRDsBcDdNBnLYYcgt8etCq6myx
AP+NyLnxObwv9oVK8D+sox5ffxveteaZGcKkgMiSM/bCMO+awF96lpmg5KUvRD9UlaQkAA+31Unl
AcvDmr+TQgds30XsMlYPrJnWPbrbpdSAK4OKVL3kx4pn0ONhDR+O7Ab1EdMtL/rR8euXTx2QsgiQ
0Ma+JtEhHLfZxPDRnG8vfB2OVHR+52TbX0PMSBQDhqL9meTdLrUIIoZMon22NGlaBTNmKXXLCvCn
gnnWBlathLpR21ZNnrJfkJ6ZsVGFr8517K0dCA9JcCq2EDZkRd3mxlLO0ylBglBtrQyMJyFhgGGu
MZcZvtBCEsn1fnYDf3moCaO2bffk5jnWhi/1R4WAEteiyt0D3HRyTkezKIaEeXN4BsMLTBd+FLCQ
v/jXcftZPMiMutzelL3I2ziv/uZsJnZa6uZwO29y8zACAJX96mQexFSjY3C8djBqfQ0Z9LzAwZRo
JQuo0HQOOWmbYithsBtYMKuyQiiVLlrf5tvB9I4mQrkc8S07JOhQdyzmzfTmu4IF2rhk4SjHvUzd
pOWNMVQGE4Ld2f0WqNj1FRBzfD3GcCI/TS9tXJDSLETXvjn4EgND7UwBlmGDTXk9WQt0UoytefJJ
qV9uN9shPShajjgaYhLht4udlcIq0ojBOo7r3iPwYAqS8YANGTr9BGC3taaD5F+NVf4PsVybm/hD
/O4gohD9N4/V91FLXVixn1algihwEGtC7W9upaDtByxuzD2yAO75H7x7PLcYNPraKWTHHc+9CUBU
IkjniQC0wh0FgoKTKzLURquVY6sB9Trlk8U/Z1S4i3tOw3ViKR8PBmVJb4M3+dv7wTRXZHs+C+F+
N0PgpbnJXXSuDpf8MWg/sUaedRuxtP8RbOYaJjzVzHCXSYi8ZAAIJhm2VxSLdVFK5bCm6ontJ/g8
R+o/taiGn8yV4dbJughQumlkxkVFeMTGwXgPrJZwHuIR61aB6ERewCZ4hdFcDf4nQQZwA/YJLRsd
XMvvQczJJF5jJfPcU8t0LfQTYDVaDzOh2xZDZOY8CE5GUep1H6je9CQsvv9mpyRQlAK0JVLTouyq
/eTaDOLiL2Mm7q9brhWjDZytQ1zFC7ERiJtlXb9KzaFlI0M/LDoqyrtRAOrTAmtBpfHawNZpG+ux
GWqyulMC1HT5TYL/u+IN/ggAuny4hmfNPBCWpFL9pu1R6DsAknXuj+NrLu9yOHrb6pGO+Xwox31X
nEtbyKKfABYYUg50rHI2SnN36Zf9ENBFPtn9375MfP86EOxacp2NMl1dYSWOYSauGBAVq5y1OtYs
m6HzREJMn2dRssFkafdMYVJjJVn/5YO7Dh2wU2/TZnwUH98gGFR6cRNe6jXhIbaZgaOgiHNq3tDM
QTACoDeq583NKOFqpTZIUPTcpIwega7GkZHzdIaxhpBBQqSZtf4L4ZS/YwBiCwKRimVerFbSEObl
9dY0NFa/zGZ/GVEKdjnlAdY2z6uSHNN5+Pf7aNYOLZe5ZgrGMO6kNwzGnTaCFrf38sYhvm/GYiJf
i3Ti5H9+zowk5p8YuDReAjjgRoGCKlqdXXbf/CO4EikVHyQEMSlXMz4lVBoNZ39TyXFoanB50fdw
tQbN7Tj0PCPTTHANk0XSOYegsW+4LWCVIpjMVkPuIg5XloeAk18tD1H/9yVgsy3SO2JbZIOm/LPU
+nlqgO+DACpvhf4BRPBsqB7KqkGbUexXFdQxilUkE5l5S5kTT3IJLTHRsrHfSkcqUxOdDw6TGr/E
yFbF5KzDkwkLia6P3Q19vnLOBD2Ac47N+3d4LBSaFj64ypUetMPqeO3lvbpewEBZCOsHhSgzMkEy
ra5t138CoO5ci2tsXf0okC4qNeGnbzmB4Q1LVeIlAA+p0WMdjemEDZZinPbNA5gTLH7ATyKflJtn
BrvN4HKtIdALeJjJcdxyuQz6EBAuo19+B4V6RbePq0f8FwYEa1U5NBsKrlXsqXx2c36dfnlblSSq
yEDHW/B7QowDX5Qm2vjflw54phzgeQcJ9/HkX7+ZoKpgAl7ZkLC2yzGRFYlZyua4YWsnm6vZ/10f
95BhEImh4XcARPIwf+NcRZSbW0tAHddbLquLFVE4Ohr9lZqvR6y6ekDU37joAJelDsZ/t4aphsmB
tnJHmGa0YDWKoFti+Tp1him12og2Q0+YnbH5zyRmETF/mqcyFwGAiXarIoprniW7zTEsaPMTu92S
YDrMxmHdUkJBg3wG4axBtb2ROKEE6CvhWrPzSGTEuZDvyk8CRRbvpI2DZ37mw5WVU2cf3sNNoquE
2q6I0V8tB745xdKSZeSpANuDn34EbwM4ZH+NJHA2ftvP05FTXW35t/QovG3iz8Q6Q6ev6jZucHJy
q65La97b+YkuaNDf7bno4lToLMIf/830E1iZU/FhLsClYUfKvAagM9lDh0F63An0pzZ7rZvVbTFU
ar726RGVYtWhvCmhWJNRXK9mPXe31lZ6fcNh2jnVa9dQOtviZe1RFUs3Hxl/FobjmmJXPD1aJejn
hiLLIUrB6pKZxZRa1ybYmK9ZsWCMhYdWwTJyvmvpIZb+XELpgQ+tERPi+EhCEj8SfWSgD9d3blmd
NpYaqAbay3mECWzUisDzIpsmpempa46yRHFvazKxqivbhHAg1Y7wxcR3iqasM33fe0/+EwtVFGsW
mRQGs/bvDGcEIRmigJDE9LsldS91YPkBMIdVOySwpXUuh6SQaJex06855TQ8GY2E4a/rFghSYH2c
AfEDFDtrePSpB7r3uUW2Ovjw5GAXd5VHKXrAoLitXGPe9rg5VrMX9U5OeX4ggEby48mZ3hLkN/fm
Uc/0Z9BS2DVNY8XVC4b28jEj01aO+f591q7HP6dN9cZAhHPbgCKdE9XL2p92QZPSd/rCjk0UwrA1
9eszLE+S/WRH4wiPqY4fJ7veINihh8cwGA/a+8HL5p39AB8Nw7YKMzgz9gdJMfxUQlVmscCnMcbz
RhKggvHWL8vTKGhz4dNTC/mw2e0rls5WDlPJ1BFVY0cw5xsrl3dWz3XocloyAbN6nDA/mCWqPlgD
z0Ut0mX976BeMoom5yhylZKM/6iSFw8cnwFpeeQu+8MfXptx/x2aGLhzDB+UEmJxqewNtzqbZYem
xO86ShnDC9y7onH/LTEqLbMbD6QHT8Ryn7JqpVx0YHAulBd6P+FO8OTERGzOLw5sARfPG0kZIKw6
jRG1bH3Dv2VFcoveCS5hKK+FazV+BdJ+5n2J6oSVNZXAZhOwtL2+3YfKBk4mij/Nl9bujxqz3vlK
fUy1Zj4hXo/bInzpcjFUYztm/rfacGG9VRcMAdjJJ1kHKflpzngwJL+XIEI3W+RNI9ydy3rI1ctJ
S8EYlYXGhWv6ikjAZsHDv0r+ScQ/fOqF7WxJSUP7SDqiYbediZUEUtm+mL6/dmtiAbBQJ/OrE98T
RzdS6AD9OgvRYg3d82M8K5yj89CRhJBGixdkxv8k/98sjRbTelXv26rSC/ANyhTmm9V1hP83k9EI
JhL1E8indHHXnL0Hghh4MGlmFgsVH2FUA8oLW4rN0xnpPVIpGRE1frQ6CgIrw5m7jjGWmFo4hpnY
oHYzviRTzeEF/IAdGS9q+pdmnyohJigt+ZY2JBQfPFjFcU+belBClti9pmxt7IK9GXgZruJT8MbO
orTi4xjuOj4WsG5L72Dh4P033eSqC2Ei/O4xRUEbk/DItxhq9qR5ZWfqLdnk2Sg8IWGnxRQiO8HU
TtvETXis8DtrvlEjJ3hgbD2RZLVMkDeQuSABDUrkJy0jOreAyav/fzj+uf7egHOJ/auuPCw9O2bQ
qXC6a7QdLRR/SFezR8kfCVNW9XCwfyruchKZx5I8eFdhB/5B15MT40CH3za2xsevw7wwWN8qR2ov
q/5CS2xjZsFGMuk6PqSFF74D0fbRgqjoqaU0KlKA2UUo80OEnS97AhAnY1uHgp+HF5EjhF1p/kVw
jVOXKn+HnJ+Dv7o/3fnuwzBG8GakPGgMoGrN0IwZFncdvlGjRJke21sp6WZ8kCumwKKVRl7iibQK
d4lguskHxCoQdviQ9kLjhMVBZTUpg5KA0+5ozmnLRK7OwgdDarofmMlkG+7QorBops6PiuwOdFdU
9qpmuPZW5ar/pamUuEDOV9zuMe/5E3CuOKWzpPGUyDadP7xxlwXrhWAdzU7j+w2zguoWhX/cwQcO
sv6bJPRrV6fIYf4q7AXnYnGpC7RlIggBXutXQgXFgW/zfTUkaJDtzY8SuCClY6xsJ8rZkltR0QXB
7MFBej/9KzntqkP68JYe9yPfRZRfdGih2LkkqgU5b2D1O6QSi7cm3X1L8Wf7Eqz5HES3wLJfk8v9
nDHZjmT3aZwq8DNca/safXb7ihlzKXExGzx6N1d654NIwXjPToNlQ6EYrgttS4u6NdSsfm0VV0e1
YshFSPWiL87Myykfx6G4nRilmV6u869faxKC6wGRkMWbQTJ7zVLIAzWoCoKu8llx8nVum5k2CpWI
dFMTcHKGh0hYns6Jl5dRcvFnaeRAJ6XdrjrqLNKwNsbVlqNXmmQf7fRSiqhqMUYvdrVOgiFYnb4m
59KI363AyusWKm6Wz7gyusVAkTcvzlk8/4ZMZhTpQVubLu//mVDpxEYlHiVmXJYTuMQU6BUJpw3i
6E8q38Dw77GmvAaJhi+o+sbACZ5UwkWsUpBTD2RhHANMouUxSx/leOpfk92TKrhsLSC1srBxM9pP
JyXoIGOWBXesR9ZIU17YKLGPd0BtDVShUU0l+RHBNpYtaWm60jXeJm0qCGLl6t7pOGg2KncB33H5
jCX7tat6sFN/I6iYU52QIy5yfFWDsYXGzAX5nszbYCZ2YlK8EftuIwljS/MAmQNYflL70si23aOs
ME/axthxsGSYW9nN1dP5M/nEdwJLLhGqN2B5oJmC+gy3TeeLmNC6urSFy58RNfykTsXYSqV5++bE
8NOiivxQLwpn/y7x06TLluS+j6iMjqmS5+jyzeRIwZlG/s8JpSqDKTc5xGLDWX+zAnYojWvtHetl
8VgAZPjm3P3AYD8KxAUyygB8Zyl6GWoPfUdt2Mx7gTceSDvgqQ/ZhFI+zv/ywoQ73kU3FmD3rzvD
5pRxtD/2T1iYCd4+aswg0iW9Rs0zQojuyY8aD+tB0n7VtHaAKR+lJUufyiqRaTmbXsR4q6QzfxH1
yWaG68oP5aTp4j0dUNVv6eWHAUgGsSWNmaJEDyUI3E3TsvCcG9Ro/5D5ZEpBRyxX2DDbdhp8DqRD
DAnQAuVtR0nPpHYrJU5cY540deAiOHF5p0ZPv7JIAukSgXrIkN0Sc061mkW1FZ15+f8JNuD9bNgt
4usc8XxAKNHoxzkQVbNZwdsdyUUjaln764OBuHH+wBcgqBJMnOhaApPKS19EDOy1GCM+ewIWifG8
bQYbCKhYH0FPP4NH+4iHNboxzzaN5AHhu4hUwKP9NP19HX7aim5Ekpr5yKTTKxAXOw5obSiNO3T8
nalAw4lDVYKqd4kLkEKs5mrVs5mai5xXj0+B1cf6xS0km55TET+S6egry1Q2LmssL6TJWS/pPquA
DinMrHSPiKrjqcqxFyxEWgUKEfB6H2327vNY1GFX4a0jRuVYgrwoAEbq6Bi8a9OJQ6Bu3Ym8YtsT
QdCVDIz9R5wwt/R6mxQ73C/mAq7xou4MZB/UmklPPtjxulhLBth3/Q5pnVxDVtJPw8QpcAWPpXWX
6VfoL709ETgBjPn/ZcNi6Zov/wD5rgJAOn/QysTXwsOvx8MR0qzHPQaduXt0PavcKZd4y56irVrI
GBQZT+6aUG5RkYFWe4daVo43pk/ZymgCiFv9tqVnmKWkM+9Adk3CC8/GwnpDbG92TCcGPjWOAnLr
byyNKJc8DDlihE/gwcSlXX+T/zwBVoYthSGWHis4ftRW8NvjFRuTENuSLYnMAi39nGgilgI+G9YZ
sQ8Jw2QAAxqdInhX2mpXVvxoKzOZo03CLqTnVmXKmTZdT8V0Y3HI7Nn1NK8ZD2V7XBH5qp2dz3sY
FM0y5yVWTo7RoQA4+jMSYhBUvafYbAHmVj/MRsCfqaYnWGuGlgmjwg0gm4BImGzssQ5rVanrBRT4
nD4mYeUDw6Msai0oQnZaUff82iXPD5XU6Jb3nhI6IKIYe5OeRUBywj2vN1eMxHRMHKueLHa4FadL
cWm2ibbCamTzyBA+/TeaqoHFAwJi4Ub77hLaZxNxlejK6PAaYxrrcNcj9GaLzALfJ1JjyXE9Ki5L
xfFPh4FTvDmMffTQBI5IFpdPEv7+jAl3GKS44UubRwP0Fq61+RWS+26w1BgXSsNdiOEbNMHtMeGR
i2cy6ne9ZkG8Yfj3fPWDJVW4YhRJPL8LA00pD+XeFKDYlzA5TCuiHKKLtn3w5igsa9vzMmn6no/0
qKVVcZ+DrW6+T7bNiir3KaSGprXPqpEo2xiuZFF3Zc6CEChUkbrr6iFzHgcANi1VXbZjXS+NgESi
DtaKhEMCSYBBlTyzx178odYZewdIMDD1pocn20q+gOoLWIiojEXCH2wq4+e4f4Q6mSBTSoAwTJq+
6FwKccAvY6tSxpoC3QiPGl6fCBd62pNztLzu3s1q2RWYelAKN7rtc716Qk3zCLH7RloLeZpdeKgQ
d/QdzOd12vQLn4nxA4Gb3QbHrpfTm4cmizf84OKl+S420Kf8fLcTP86bN1uLksoLyzAXEHLhvHWa
D8HnwZNWqp6OdsHQ4EbptKROS8AuDdTLiJ02CBu8nImPIYYfBXEfeMarjairBESbMisTTpEMOExk
u49HURd41YiPT51HDy3TUs+/FVZ9HixIS2AUDw3Ob6k+XHEdJFPDk8qn8QbPnIgK0hfsqfk3i3ek
DuK0r4PMjkNNGjxzXTqNlTIWVyN2byLTJGoCQJv0rYJfxKPwfV88gCIZS7a/OFhOKVwZ+YlbKTgh
7llD8zvhAwrdcVdY6RnHxP72AVIRywwwe5fh9jhX//oBiJyJqVkWLif6jCf09AmPuxB5FxM2TknF
EzPrbR22V+i5PaBtiloeNvD8sYv1gcveswSsS38FavJAVNC4nPU9QYlHOcUypgnoxUNih7uqUiSM
VH4Lf4AfDA3QnILOG8iobgIikA6jmEifsu2drdmEPoG7ofoSeuMEwqcNKwj+83Y6D05c9u4xugk0
JGnOsNQEV7BUAmWpAcTyP3F+KwIIwZUx2v/0EZMm8X+xYZPRGxvzJ9P7lM3h2BB7oBQj215kBtuH
sAtXc0ot2HjGbJWSwjV2BN0lnp1ZxNWXGReOHI0jF4rFsn+WsqnfHq9T13SyCA+EkOiSpyQ4Zjla
JCC/Y2uN3NWIuYpeOiQdOsaVpFbezPsb8Z2NWPLsbRlA78I93GB1g/VeYA+XdYk/a62oWyr7yAkq
8b/j67AGbkIdcSE04dLbEFTiRK7cANbaB0aaLDJCMPJyBt8XPb+JG58NSGcXfOBsFpeQ2Rw0KcdD
Qi75cHDL+Im2jRbrHVwZK9ZeGSueyFb350AoNUDI1yUdR72NWtpGlg8HgPMHx47w1jBTnHPrMwG2
/TQ/vz4o08qLN4xnBd/lQSaovI38yHjL9TMxieuXw5hCe5HDK7S43XheEPYFthYy+E7oyf/acCJ4
wdL5ghwJ+AV54mZXU3CfXOpjecl+AVFMHNvW+XymmpnS+smUod085JWP32XNBl2mFYipU28yfHat
MuB0zsAf8xdNZvX0DreMMjyBg4Ca1J49l+zZGiT6qQdfip75uQ2dr4vUDjTHOfEO3Pusp4S2caru
MRlWB/AOjcDM/TnVvwwbtLnaVku8EDJgBPLmXjMkSFVANseMeknMjUlDgkqsJcxw1vmp+hFh6QpC
lcyC9+hbI/X4IijYd3ZlpUM9er5zT2aPFJtn0iaxGF5IVrluN6rycumvtquifYK4rY8EI2fDvCHR
XBcwM//tlPD1bjHgYaCrAenlw1iWFy4ufKEPg/D0WAeioK9cM1/QNaXh7Tmx6Bug6BHHOcMDgN6j
N0reXJg7HagAvPOa+kmr+66q1jy9j2LtAYsElBrtNIgljJfCMJdERMUITtgo7jc71Q9n0bU2l4yB
1nF4k2T+DH/Gs4GbYtmzBrf0zvpE3eRfttZA3woe8WXOptuG/5zJMW6qoPv63d22HonkJpstdqm8
3fSxO78hIoa3l9FlKrHfNLm56cZn9yQeKPdKBP5znPcS6v+d9kIhYG1wb1mrZt9weXl6X2Ei0Hv3
uDu8L9bigU94oFvE4JynjSKvb5O5/iF2JX4FB4+QMgCVXYzBcTN83QDgs34BOOSXpqhM0mf6E88l
4T7viWRdYuFZYN3nGvnLBecMptbauNBPGnWNlovtphH+/M5E8WGzZApOXORGThF9/SdGcOcZKpeW
AJrJZr4rkl5QqXzDuA+n8ZAtQOohD1qPTG5x3iXty9twzqsVXTTTUF5/BKEvxf/DHYW/qlemEIvx
hx5IIgMkA3NcdW6fjLIx+5KFUJMrxIjxWnYFoP/bay1wWvp7Q4Z1PHesvFMEOg6ju21qlfUyqZwp
gRn9SfnXdYxP80PCT0TNhIJM8LfeufiVcdFWEZv2Ftwz7p/oy1M/WVIpPFy/xBQb/mu0sV3i+g9C
iDltCeMfZAx+KzH9p6cy7jRYnGbiyisLMpIf8RMp4Ddcz6C2eE581CdPoDwSAcQYQG36WZbxrWjN
tQmI0LLKMfawK/vM+63bjgHLFknJSi/Bx3vWxyFnyn5AGw/TzSlibCBjjZBDM0zEuZpJsseb/FpN
Hle0e2sAD3J6CdvvzZTBlumeEFC0pYL5EjQFzRaleY80Y34oO2KDhfWCOvO5e1DXJJj8wtJHml4t
m6GBTBR484Q7LtfcKPY6Q9BtYoq0hXaVPC0WTFiqpvoA+Ks7/PJ1wfqRsX7+BuqCKXHRM+e3WS8z
thXP/Fac7ZRDUjD6SbEgoy07mKVik4bxdGjF9/FT7009StVvmvZG/QMPc/23uL5ELC1Q/bSjgZG+
OgSZn1tkftTdqEwqQtPhxS2eILOH6/tf3BVimTEDkQ4vPVC2acStGcxTRvmeCISaa9Rf4n9d533v
PUNg2c49f3CmYB4AY0ckY8YuLX+JkR8+zjSwkXY/dFxVDCgffdEOWKzONwiU8LVPnYfrtU6+TjIz
1xNhfxxwCJQKXHLdg7yT3Eyu2McCdFUPx6ODUolnNlpfY+gScBvIvasVcOrzQlxtmFL/6hxMo3zj
D9jqyLT/ZLLcsWgR5z/9sEBNVEML7M5POD1L3X7VDLs2mo8/sY8bYrZKERdITgvh2lH+VJ5ybG81
y9Uh4WJ4slBBh4g26H2/AQ1t3DnMchu54E2OTLmmrwbyukuAKv6s7YfK8QzFciaZwrPnYcTn3GR8
k7wY4mpc6xfAlrr5XhOE6DBqPNmLMPfXTEKa5uUNDr5wDdHN6414yKsFOvrtGsLuG0gMqRgnhddn
Vi+764EmiJbymXY1Yb42vuiVPUTcIdu/eaU/yHNEDvn5P6ceSNTp//H/dHSnuvsyKUOgA5pkA8ke
DZZ2lTT4mEJAD7Lpk5h1cK9iaytUt0qntYch37zYqWysQj6KRFa2KsxchmwQP6ScLI5RidZGLwwf
EGQqI0fOrt2VTFdgntVS6ECX5vWTGjawBD9UOrcqJpN7x0x4BOqT6/mYUjWxe1lq6X8xJaLxr392
m7HpVFI517A9S0qYPgUK45HZyqxHgqyw9knwUvlotbhCLZsYuE3yjsrRdOq7Tx9N3UED5l2iN2tM
ALeBuwWiZEAjI+bqVbP6/jjRuoz7ECxfJ3DrEXPG3loN+Oo06pVNk6qhZGqiwOO42fjrzz9hTGWn
OJ7+oVrYhYjBoI56Gt2vqhyaP5jLgB7atq3R3gWt2f8X82KjDYbfQeIngDDIkeQ/wChPFc63OOYx
k1FA8zSirp9j9uSJF1c7hJTE/QuAaPALKmy2dvIh3iSwqXFDt466sbMU7IjRaLgG+EntcTbMj26D
lHBpmO+PHMYIRpwf8TWGCXyyXpJ4ZOoLtC6O9zZrj4ysC8PMR9WomiFPj3lPitgLFPvvyQCIbWza
gwHWrAM3sSZ4PFHXKzYq0Nab3JlxKYj4ddHF8OQc/zAQ8G/XOi3RcExpKikAE9XPD2wDXt3E1kWL
9C+HFFLTz25LSMK8qPPTYIoS3GIcve7NmEZjrXUKrhE+zI9axnjs0OT9CHfSxKWFnaeSEEVHfwaR
yKuDrgN16uyJSHa60XwpY5DiSaze6PoHRsYwBx8XzH3M26L+//ncRIYLszT6Uw6cWI9JpC+m4NXn
EVYFIfJRzsylBvK5/T5rmA0atcqkRS+rYIUJ97u+G1up+enTdOhqrQlTaeqOZ5EQoA6GbYYIjQjQ
PfpIuKrn3az7YxmM6bR+5paAaBieuQXEY1ihUCNQT5EiwfYweZoobUl5svH69y6xcfA1Qp9Dv6GG
7YRWmFVdfvQoFizvRswCYYarGHb+/4oc1tThFEutb6PNcMtvlnC/k031TlqeFHkMLaYVg/WvTEF1
oFxc8infc3He67Gyvvizw8Q8ah3fdRvSi4N11Sz+z+5B8Kg7eugd+bRn/f8s66QWVqKjr8CqA/Im
wp2OebiMdvqUke7kknmZZH2piVC0Hd//BppFq4u5SLIUFhTM93S2ckgtzCYynKcqZUiUd6i8g4P+
02lRFtDn6z/GF7r3ByysHP7injgCloJ5RmdZzXAAffyRAPUCvNwQ2SYBwl4L7z4P+pRz4sn2xo0i
IuVmB/4wDjHO8XboHeiLPHn+UF22twnC6IyOOkk9v4Forc8wYSSG9do8vfFt0UuiSSKQQ7bJv5QC
klKtA52TyYIKEDWBynzEJvXEJILdfLRGWerWgxq8eLIA/hZ6iGBXrSL50lcI8AhDN4plKSrx2g5C
+TuiEQH4+oJFywe+3b57wsZYiPSTWmcsFlbU/fTCtxiF5HETDsKaDTTbpRQA9DCHL4t2l4cD626d
UoAafr1vU6BD/RIhTTveWhuShTsGfcYXoqNN/IBOKKbllc079smXdTlkeWGcnqicX/UWmAWyMG4Y
/1LBQ9/BGKw7jYbSaqw+wEICMal3EhXEKGtUwvPWfKKAH2OgGt0a5MTg4wkBNngaYC778xD5KOYW
igdnynax+eeSpZAHguT+CINf217c4dJnkpdLXbohhmUgHQ3vEe42AjImv4XokRmsBOj4vWQmozbs
W8awhxP15T78NwZWbKHbHs4JZ8pHvMoxaJ+MaTRXOQMlefgA64Hh0eJ4P39N8x5tLhEtlwwu+thd
01qEQ0X2CzJ+0uwDCl7GwN/SbXu4pzLZ52E4qa/gLTQDfGkqcRDAbOuMGSPf++qGlcWmhfcOEaZw
aDpvtX12iUa1T6k2dm/pMo6oLQrzRbtRRTMmtBH0B+0JW1KNOSd70omoaEfGYGkm/yrH7X1iDjp3
9sFbZPrytUzyE+1fri1IcnV8A1CDvE/UT6n/wkdr0qS5UavQwRytHjkYWVs/kf79a0lovlGQ6WpF
/PaIGNHPUDkFdKNvvrgH4QYB6PJc/PSBTnwg1OZr0ghJY92zbDnxKxp/aptf+P7jPRRTVj6UMLA6
XuCH6kJNRlkApaK2dP8poQDoRBStcDfuvIXvALSDWe91Y3eNtOs56Kg9NhBShQl0MPo7P2AoBCHQ
BN25EskLk2b+Q2KjKAU3WkHlXwTEn/HDQFvvvjWblyla2Wd9ZnFA2FFxcUbzUEMWGPnIaNQRWJxs
lyYgBAKkrCf8OZb64Gyy2ekvIoLzeH4DAqahx4ZVFpxLrRIQg0sJ85KkyUi6FW4T2F2fJU9AwRix
w3bJAjFZYVyGRN4Oww2VbevYkG+faVqSnRcigqLJjYVvA57z/51w5otTWXIx2e5G7s83Kbnajogm
/3djV52oAi7f390F05QxyDDPB4K8Uav02BZVF3T1QY5lwDk2qPp0HIEsJFCU6wKw+Wm68MVH+MN1
tqaQjh+QgFK6S52aErsjoOARhN8nVQMMa9u7pvjWi7VQEt6ppJoPgdIZ1NDDmY1vfMgDxFw/xZND
XLT4mH1mI815eScGMtRtpviZPNxoECoUk2fjnCRkyEh4mrcF4lmtVM68/5SjxLG6kZBRvhkaoip2
RsmqyLAEGEWLsD9ONos3cdWy/0lgvuhpwRZk0fg+9nhpytZ5Gl/Rt6r6M8PQir6tjjHzyQOujEX/
O7XNBAqHno9SAsWNlFUJYj5VBA4PbvVLVTU9RtZ+cGz3Fc6ZSfoRfYuiW5RBJMgHJshfel0FGq+p
UYrA2LlRDebvBcdm8Jg2U1aQi6rwqJ0tITAcacXe3bkaxyTiH8ln4J9PZ10f+4ip7Ci0fbNjYWhP
z2BCHv/A3LpeexZH/Am6LS3htK0MAmH3eu55wwED9R4A+l2MHXleZpJCRQs+1K4jBYU//QZYW7mk
HVW04cQUXQ8KXXKuNbxS+OVk1VvwPgcThGTMijW/7rXU8/0M/AgKxqOO2ii3KaxVMmnvpNfvFy0C
zHeXNPLrgE/l1S0Diga93EhzPiTskfXuaa/ocQVih1SPtpFEN6QWGRyqilJPbePy8M6/UMcRVonJ
6lZirocNyxQxXBo51X4y7i5SYcHUaf3CvPBcwH6fZQH20fMVP/IWwTgWH74fJhPIf9o46qsSxzKf
czxBhttP3axxjwGWh4/isBODYsVhd3zglrj7naOHLAU9Zqc4w7ilOWi7pK67wHmOEFY3mdLwzIOb
WtjEWh1QrqORI6MzDDXFa40iJitGJh+/tYtZqJ2P3NU1LkTToKuIBm9EXYvTE1XOzLtOqTUFtCrx
U1zrrMlp14tR3x+A5m6km9tOdsc4QwGaPvI4jf0PcTNsjz8mhy582zys0govpBa8wCWEHGaaT4vS
+X86cxonxdzO7jnlMKv/2sE0M3aCbGO6OEBEh2ZoUkug/I2feM+FUC6sZzFADCzlm99sxzcn6V2P
adBMxMcYJR9l3o33uk8tzdkNKkRbxQzk1CX5Ji8wBr3LBoiQLYSdt+TDtNBHe7MMHdH5ce4ThDMN
F7TMfJHb38kiujHd4MIjrNO2SyOeHNfyQDMo19qLfLRRI48A+zmHjb2Q0wKk/ftTH2c+COefOgbK
ZOjlOXpck7Iz77WmtHUsgv8dl6NEOlwcioRXrOlcd85c+N0FJU5bYWwiJOEnBHfBc0hUGOuSCIm7
oLPF1h6DkOpC2efTtvRvMJiOGt58ktfypG6ni1BHQTQilGY7KbE+ySVlJjrX+jL8gRSmbEilwWxF
YkqTjIJQfCKfw2/ECpXG7lfPzoJ7JyoqEcLO3zuZI47byhNsu/CsKI6mqCFAlvhnxO62WQilT4Ai
5VkD2dPmQkm1/4wrxtiBMAUVMQFcaFa4j1DptU1nDQkzU6e5gHVh6Xturmx9X71vopPo2NUqVXF8
EnEck9dEpir8hXvTbTcapga9x5746OlMKhzaH5XfYH6VECfUKe4l22ccDG0Tp4ChSDO4WzJCCYZV
HWXFe0VsQx7pX46fCpJD2PN5Ua+a46faAG0RWKeGcku5L+3UIXYrktlriC6LqL6yUGPMTFyDtkWc
FERfA1r1b7qXYr1RisHlyAKeEMqXdmuvoOeFrwqYwUAU+Q87sK7xqZQRBe2t9RqMiB061UPf6XvL
BPRL7l/Z3D0MSv5Nw7QIoz+ugTZk8YUe0qRv/wPrtTpO2Ge+1zMYhG8ejkD1zzkdG/GSDoZUQ6rD
AIduHjsVo4fqEurU4delOugSv9aIG2UEvmUdKCAS92kB/zSVIeR1roxJhClTaLmfxeq+KREth27O
Z7bzCcsu2w1KRqra8m6iXZcoueauhLWSgvLUD9GDAIxncw0PsGiiIA+/atw5zM0wlmHIJCUftE/Q
ZJyz/oeXPnePtbXSE13eB7Lse2UYMNi7TJR5b9ZTWXMywnagnrkQIifMSio5v847Ea7XqCWNejr0
wIVasMDx7/C1DlKTqXPixI4Z7gqysbZHgMGUGdUxG0fxZyyRS6071SshylYC3aPPNHowFQfUiPns
SU18WNUnjEYi+UR9DoerlwKVEucaTdu0FWEEly53waYGDmWzPlZi76yzKODfirlz4kCEcOEBO+RQ
NRV3GtJAZaIWs4tzaS5lp5092AK1TNi3bluGEjxLV0nAQPwn7l9OwCub6feHiV0XMg9mGbgKcu3S
b395uKuEm7zOySRPND+qubB02BrzXxRyY2h7qoPV7Kg2N3U7udlX2ER2tAQ5K/POjOBfGPylWFFF
y9kIWbJFhtDPJdxsfxa5IPW2Q++dSz/mZglCCokmgQHPvJYbuRAHQYUYAlWmjn8nkXCN2Q8nsRmF
kWIOs8esLEZKwqeni3/kbMVo80rWmoKQ15Einnkw2N2mPV5cloPyKlvPNx6Yha3dChYjy0UW13Mt
ePoqpbbXnjkd1prKeY6CoQas7dX/DFS6qIqesggcYZL8KXI+CgLanP4YlK3D01vtJm5L0/9K3RRP
FyJeOb0nOlnEjohHQtb6nJtO/1WFhQnh86qlgSlMUoD6cMFbp/vkoFB/wCwzJBYAOeTt9pyA2+r1
5PUXtMbWnr46KGbQk7WumGQnP0JdARRltbMVPhIM+kgmoA+wTR6TSPR27jBPUvxCbD8pmDJpdIjD
r/3vr5ssONtStVev0tjp4+bt+Pt6x1I3UHbz/AVy98fvXvcMl/NliVjA/Cul5Bu4bd1Ob8wVLr5/
EOjloWPItfn2h+BqpgmgmKf9yZ4Hv/hN4kxIhx2m7MJOk3zFnMfna2sSltt+ljCCsTEHElb9F2qv
HzMHQxmYJG2t6sfn821Ysv9UpwQotqqIFhLWiozxHM2sIJmPUuWZ5PPF+tfICqy/pvP/W/qEuPmm
d1qCxV7VILIMqUvJtvr2Md5JJMGwQRMCnu7yUHj0NrpxRzTf3QvEoNt4tkvO7nhqmtsNIxDUmV2L
rrdWsAi6ZkTqDvUouWc/JMw176t4Qbp3kAW9U4a4YHHaG998rq6Ul7/o5bkbjHj9tClIRSTIG1Mj
yEczaCtTmTaZFMjiUIoyZxk0MTEDpiksNDijsSSj90fEmXX66CEsqlstHMy8Xug1PBwpPyDr4QGY
MmkEkuQr1aiVSdLeg/RbmdG89XgdOivn79ycgFObIOJkpLRySPDhXkiL+rwPqw9VUEfQeEeGTZy2
chZGu78d4Fkf3Z5yFQBNhzp6yoGWtXn8ZGoa81shAHOlnrAtil4QxjZe8pBjKRyqrZAPtYPZMtlf
QeqYMjzEaVIjRFrhamOqhW4TaAUM93ZtNuWip9wzdmtuvzTP4hMJvBwCL2A/nwJA5jDhp5mU6MtF
aQ9mV2LRNtygnZ2ATatFcDb9cL89/bYpL1O58pMB/oH4pdtjlu7xdwQNXxUMy/YyA+5tyVWkFwRk
nib6YbKMpsaKU28YW7potNWKsW4J36HDbDTlBjtkddKR6o++E3zhow04Yz5GdbhAp2H4vxuvmDGA
hmDokFsDWR9AowcfCTQg5qnOKe97lt3Hq2S7UlW6TK0aVgHkDYtUdpeQYOUFf+sPtQUM9490MCbN
HvtNeZZZUCZfLxOVi7C3LBiT2DHMRSd/urM7TAiRehsSqBY9yRUcDW2RxglxPTQGJtNH9S8ruNH6
vqJQkyAvF6vBnzhiOeQfzaOeOFiCcNtGayVNahKiephf6UtB0NaXFTLiPQ3zNpZT6I3p67PMCndI
xN5KsGnqwkvP8CpiURkseP1lz2lcO2SURhDJvFBVQEHs/boxrfwG/qL7yVBDCxutbEkoeyc/HzKk
KSJj75BJiCvwB66xPiFBJXjcQ1fqUrVCr69HAPW31tVrw3mYbISm3we4nPUmM1W0o4mDkbTUP28s
eky6QyecaO734iJylNPAHTWpfRlGeATxJOo+V4FjqwxfOBL01dtswYn+hHPDUC7+9EuVSOenPLrN
57omdLKI+g2wdcuqwc035XTP01tTEzvM7efOSxeyVPxZPlsjxm6FdKnmwk11Mxfk/x1Rao/aLVmr
uOCk3AKtAg+azxn9StQZXw6+E/ZgiPoQv2YU+8Z6grsFlcDMSbz/CO2W75e90RwZU0uZ1dMtsjRG
FzYBUxYhyyy736tFryW9tUuNeoyDhPQGFPXFbUF3Hm3X7iJKS0p/4E2JaXm1RyIuaMP4C/YVNiSw
UuyH5jS6o12fTb/Y4KcFMAN98jagwDPhcW2XSc3gPhl1UiCaCE7Kxhp2/tb4mAqrDm0gG+HF3vXM
IgRZXoyn3eOs3iK1OZclig934XXIuKerbVMiYBO/a7XYhQ1RsI4vwJ+YPYqWzd7nHvJyqZ0FD7Wl
nxxF3b6QUT+JoiiaxS4KeM+QMPtd0JEMRvXHXb2Gbbs2vxZv4ae9ytC5gVWN2zivIfRuWwUUmes+
VdUp8hJaq0FENPYXA2U/lzVXpLkwzxmwbQF8A656CDd26iasQT+hCNAxVN1HzdmOuNHGSDtDgJ1b
JEHFNd2wRkdYQCLI+f6flT5ufH3+FHfQYg+6HwQdYHfV/g6KopXMLFsl9A/71DvTPesC7NhLwz8+
MfrseUipchlCSeO5pFs1oWBfkrmXUJUYdbDuMlcUz6tC6KCubipefkvSlSnDMjK7dxU+uwna0+WJ
+PBb1pQezk5KQ9bS93pPcMyTbOHbQsp0QMwgI0YGlUIthZdIcm9wwfFy6Pxfy5ZlRcBPiSEt1jA1
38nMOEiwDtxmTXTgEef1NrKE3Yk/xtUlzb72Rap8eg+U0pa741qzYX43sqzlx9UZq9XSnsK7uVdO
QCqFO3/Lyuj9kBms4DecHvDqmj3VodlHb6ThC+CuQCuGkcfVKYkaHdnatwdkTO4H9D16S49iVYow
AYC2K1gFSMjoAyukN8EjGxvPcbsjRGeItR8qVi9j3iy+bZNliRbtzddrwZ3HGUeE2YC1VL/gT8w2
Ujl2UGVMRWTgICDtxhC/e3jSMHAlS23fE+Z8PD6jbafVZDFIBC2OMLr0Tnhpyay5MvQS5LkvqSIa
GtwavutUMfylkGXFTuc5LCVyFYGbSOOUQnE9505zcgNBhvL0kRak8yRbEnowcsyuqtSOCrXioZbi
0dYs4wIcZlwug+pVq7rjGwHUNIPPzxt2OFNFEG3OLdxbCJV2bDfWlylqMrKdH1XX+weANZjGq2Az
QWwb/4Lq7FN2EGrON6RxEjGPgzcTcfpgVfhYa4BmT/pqJgb/bLI52IA2nC2b5Tn4E5wxuXbSFdqM
rQNUopLYv8sRV1PDeKPVvccFjQ3br71EvGZlQ9EfFUcTyAHXMup/s0rljGGo+vZ8IswZrAZqEh6c
3SrNoPsVx0gMAUz1ULJIhsdX32koAWlgbCif1NP6Jj+qCrprjGbDaGfVH1BtjogiLEb0A2zeucKI
sdwERZUTWHEYdj9BseaA3Kmsu30gBZinBcxCkJEHgH2SzAV9m5gVtXaybdfopPSKl1kHFdmjlvfb
9tCbZ5Wt+ST/QHR4zuALVAI/UFPP/mJBgp1erhNcYVdCxb8H9UpxGtt6GSttGqQGc372zxGdCZuD
tqwZslwwrw2e8LtGfysvmPAMUmF8+INzCdBJ97CUEoxpNryVOaPUIAPatWB4s57SgKhB3B5DMfRF
l03+5v1hEcpbcmCkNXCwQLPvA3s2Tmd8H6liD9JowuM+qMr6xZrX2NypqpTC3lzg6SZKJwIFsmZO
Nj1eu++RzW4h9Opf7h4RZLkTWFv8ztGnf+i8QpPZlzoQr0seC5A0W5DVXUAgWF3Z+cdzIau0gThv
hl2bswdJEG3vv7j9DWK2Iu0a482otJSgrQEiO5xL6wWxoWQ3HeYsubzb6MALUyzkoMZTyWDfyW1G
X/f4tynN0w0wRD9rHFcp3vmttn+/c3wph3RMB95ij9mHRKN8+IWZO5y2SAh+j+y4rG9tfgXOYr/V
Jjk/v30KYWrd7LW9mASWhtE3kOZ4bJrT/dppZ/Jy9qfDf/jXUQ/UydaMO4r+xPYNKky91uxQBnMe
2YKGH8w/Cjs/mJTYhOWi2jniLtbb50dv3OOct11YmFqjCkicyHUZ0tPZk4fqMkBzWm0sGHXd+HDk
dksWnZvuvFoY9KP71sY1KymoSsWp5o559kDeCmZRE/ju6MKJPXRvRKjBTTLO518uNsZ7+vS/Hk+V
UrxnVnA1tNu6b7htHfOIHoXCPxr2ThI2J+NXHjOzVe3ExY26MjveWKBi91JavW9lJXH4pCFaQKJf
74W+sDSmKbJzPRVRQfMKoeJ835zezvrMPs0sMrQKYaJLnTFcKEgnOAnVgr2lukGARtUthV5jc4nJ
A6NnUN8u+bDCI75U05ccNrQO6canE9F3zq66iFycWiDuHr9Y5Pf8toTUdO0E/Vja+PToA0W1klFF
twNa0TlW7zS/KCA6Ufuc/PuNO9g/XxY7E5P0QFYNNYAir07kE5MvgII5bQOyRW2uvBBeZOo6QaZC
IbpXrBM2I4Yywr+OtrflN1A96YIZZYs/59+7noiZIFESkuntwk85nXAME4lv/Ku9XrU2fGZEk/p3
LB+uQ2pV3lUZkXksPbT739QxQYZYLVnkpQbAZNDwugURD8ySHhGkJBHA3p4GJnxf4vteup2UJ26s
tjLO0MdbbnlEOuB6mQ8jlBCBfxiiDm04jxagzPGxhm0Zldm1xr9KUpf064CNB+IKjbqVjWXpPB0e
XlNlOV9JI56wcC5cq/pBOJlNEm2mX7t1rM/xk0a7lIqW3RIOye5zN8PP17gcFj0lAwRepVx8N68V
AVI/v4l/VaD2skV0AbJ2oF7VeGsyw892hyY8wVtPn+srp/KjTMvODYHyksHJxA47XsxGIeudCK0q
8zsDbokuCpc9E+YGBGlBnSkJizPcr+llBBNKKkLQemPNfhI4akXMLEHe/Z10c/L7S1FyvKnHT0q4
Pz1yf44RoWw9ldNOzFUavAiHnlsGG+uBaoFZ02b4Ng+h7u8d5kCU9NY3F2yobeRGCAgDp88kNw6q
+vtZKq1N6tCRxAlaoTdx40lDSAwJ6utcIr3MxruCFJ1ZGiNWxSL9M8CznrtXCq4lkxDa60wk59/w
auX7K6/xKYQdaAMd1pHu+l/gI8uDfambNOfFTOwQE9/+669F+TZHUDc8ctHDA44YV03Eo9kR+Rx5
8HVcDQiOfwwdu6g2m7kW5JC/ZWLSZekGfkeHKvU3NZuF6qHgSieHQ9k9JbMtxIA+EfFPk5zKlSbi
4/uv6T7NGAszpYaOA96mu9OwJC5LGH7Bzxrz1MSWI/qtYFfqwOhIvMEOB329MsFbMN+n1dQs4Myg
ITNx0nGwrAzVbPCp6GF+a6okw2JIuc7KMsQ+Rf6M5WchT6TC9q33h9ABzBLUFCFGcB3X/R3D/K2Q
EaIIEAyr6xUQVDdoxf1odp37zWv1WmwIQBac8mI0Nt1EF8oL1etg/yNXt39ZPiU4/AxRUjbYLpmZ
+iEjd83puuskdcbo4yypLPVIvbhux/GkyYY3EPCXVmRKYfPIm72TS4QQVwyJ+XuS0ahwRPCDMKLP
NdJrs/BHzUhESrWd/e0pR+c1gT9Lp67MALCNYOwsx58o3g+GZ2C8Vi2UzhynRkwb4zvw1G1dX1Zl
QyFQ4SFC7IiJHSaj+S9VzkexH4BJ5BxJnTHWarNev6xuEJkYb1MOQcdtK7gQK97D74Jh/FnUPmLz
DnTvAIyj5E6y1YHbwhJfGHF6S5I8lLSXSIT1eGg8P27B7pW/I18voJwsNfiT2sn1vv8bMmpHH7HG
Y51nX7Skc0uSPPrGhw2GjPz45L2xQMWnsb7CxuQos6iZ2ugTLXBFRlOs6m2gBv6kcv4PF0CJ2Ddv
6p1EXQYUx0QJXA0iQaKlvWvXr7rt8ynMF2U6j5kisLuj2F1W4Qkpo9phVgsZmk0oIzIUdAbP86O2
cj2fgUoONcd5e9Lr1oELYvAFttTF0rjEH5hBeuXtadARDebVs87gEjQrU7Jd+ojpLJ8RjDu6sQkd
umt2dYmjvEcDSFBPFxowPbzjU7SoFpr2fFcro8GUQ8sqfniSed5TgCvQPOaez/gR38nfL4HdRDLo
eQRwJQN0VYsMRaUzWK2Vj1YVAimJtA4XGIENWfTnIwLJkwsCRl1nKBhgpSm9lsA5i8WWNHF9fOmQ
C6sXOaJpvCBBIaVN12NzSexsyUy1zadLaGYtvAy0OVipVvSPF8fzG77/G2jqwGu48NSFyNG8BQ7I
KjrSjtjGQA14huSy5GeFIb+kfViS5ijqilYfJlSdR0BqahXJ5HNiLFMhI+WME/O9FVkicMFarbSk
qFA8/gXw4U1pbXl884JUKgC+jFSNjQz9GLhQAMI9jGcLM6EtRFZi10x1osJeIQoJSASMZjBsL5kq
cbtd6YUjmUYThoSFU3hNqHRWWjDqO3vAc/KjMYRaIzSPsPBNzxfQaxg1NOxCEDku2Z0+zdfXweUR
GPFCZh0PCsdfi4Q8zby0JORDhwuROjO49H9OmtzhqkiNoGXRpY0V/e1padGj+izKyhnDoytKMfb/
JSZnjFBftkLPGw+BvlKtLbKyP8rfAQ6O39gaw/tfKpdkQ8H8z+stMCxl9BRnulQ5D26IYNNySzLO
dHMfYupPRYs5wGIOE5+NW9mbJkPThC+Z2+OnQY1LTojcBoUkALnIIrMDCOLnOEOA7kHD95gOFxM7
mBj3y7uvnmObaXi222pH38O9CTbq5kDG9nIJ9nnLmuG2TGm/L4vVmCk/WXGk9Iey7Zw1AjIoFP41
JNhUksFrJEUZIsOx+6C/tzWqufsyLQGA0LC5yL0Un7HFM4oqKeLdWh7HIi8l3bq93FhRUWifq+6V
YJubFgDl9qh+e1d9CwJtp4pSBaIFel4toWNZNoaG+Aj+BvDmQGJGuINYOBCREQgflaDFCgGUqwjf
5rW29jwrplom4G0H+T+BhacQ/eagHpgEJ/4AJHJ2OszSOJUEt2+jI/5WtUX6dBpmgrd4wJiUIKtc
FBY6eF0sMrhBXtzQgoKh7S7x1Hr0hgiTCPu7GwCZSiTg1A4oJ7YYEbpZ+MIn0pHy1lXH0/PT6/xv
u73PnS/x5WJ3KfbKeBxKTv/eJ0HXgSNfFVytP78rR66o65FHM8BT/ml8fv3pUMSFgmoRZP6kAehK
nUeqbPYMTcAnL4TvAcCDIIUCRfvGkeMKcqWwjBRw5DLLocdAITyYlPwFM+nL/MEavyQ4ojlzgbga
jZubcH7NtC3vhS6Wj17tH6hkPKqSoluFw/dzAwnonUrbucFoRiXhsFGrETT1xQj6VBpSToQWOIKL
eJd3A/pbZ5HkHjmvgecvmDHldVZX/Pup40PlsYF0lFAQA/ms+65LurL09aRNZSAEsEDeZFAYTEZd
46WorLIGmb/vUinXj3yTUaQwMug6Web06VdxzV8rbzSnDtyImxTmpeKYYeeLWgE7X8VI4ONjzuD6
BVIbK9SNAav34AU5OPM5zpUKSWAY5XZ/FxoKs0Y5NCCe1B8woMMFpYCqo2FZXGOCvVrn3/6GH0Pi
KJe05f+GA5kDKs3hSQJaPGb0yV0/vkOoq0jN5b9YfzmPzZQjWNKKdFpEiXo5P1ZC3HWQuymPx0Bt
FbBV1B2FrDP9uVl62mF8o5yuhDc6kVdXvl3o2c0FE7Zsxm6t5nCnr/J80rUW2YuG5UAe1siFVV82
I8hKneU68cCTFzGcV8ZuENj3rIcMe513h57/vbbjqh02+Nhyml4VD9I3r84MBRxtSvvx4bpqt12e
y3VQKJhFFg8maRSe+Ccqb4LSkc51BOzkPn4C0ArPjOiR8SQjqpIEwdO1/5wz4cA0X1ToaltIUOM6
KB0lx0+DCL8TC4FkslPAtWCSxJf/dTi1ly+qygkby5Wnw/fVBRKzTcQPtty5c0/psxWwoMviV1QY
TTien8ecoebjfdlWT7edU9iD/JR4oNVw4btlMq5kvzkuNo5WEkZ2+Gn+FUntlVwCRPCPNoc4XM2Z
UiCyPPnGcUdRVHAuWXURe5cwmK6yqJsUmtEp2ShyZ9wZ1jczYy6sPH3qz7cyk81E0HKmWev4A+9X
+AjyKTZYZCPwoyG23Os7hhsmVOCAcUYSVSCReHdkTMS/ACFvNt8czt7oTEx9gadE1QIahJ28jMPH
YNjjChLM9CRlZh7lcbcMlS82B1E33HcquML7l7ZE0MSvcBRV8TzvYPLsaSBcQpub6IILa20v3+WU
+ry8u88eSLS8KaT3Y4danT61Wt2tRvPfU8ke+4o5JXc0i5x4lLeRDcxmwr1oTx95bslcv6ggQBs9
pGab0Lk9D+uv1PzMGFa1rRNmxWmOXzSPYbvycMmrEm0hyl/iO6mhhUKf08WPxHqZijRvSpfx6Huc
2M8CSAMck4ODpQrF1admSBWcG45w4egk1Sj343GDeUwJ5/U2OGwYbN+JIEp2d4m9nhXT7q/TXTuN
ZCmDZjk3laFmwt/KOeALp73G/LSuni+5NVCH9Cf4mv+0G3aaH0nDhfiD9B8ug9fcyRxyHl5N/zLV
4o9WQMVXkdy3xjKA/+nbLYkrXOaF2P6hHOf1yK0MAGbZirGLgs+ZQKWmVc7GZ1+QKzQDQwrE0mns
7BSlvwF+AqD1OiltPsCDi/mbeLQcp9bErOX69S5GDmkb37ZrtMCtvWooZw4AcR5q4YLCfzHGkiom
v9PpUMFK7qzKlfYh7bLdr0u5VmIqfWn2is1Nz2Hb4q/pgCPCytVsj8TRJ7xpzGpnvhiVnMMCCT/J
136K5BWLBsFl4eYcD60SbP+P9xD8mqlqCTeFgseZczFuFoI8lXetEcvby9OvXWPXyvmkbzLgqTmL
0XzrN5VF8aBs0uR8JmMMzWpprHlEfuk0J4oJW4k3b4DKObGq+bMw0RmSghUln4hBzO9DH2j18xCn
d2hdFcFbNE8vMb3D9isID2U2bmotOkfO8NX6A8HyoUphNg9so9IICNHYrLlFRdRiUs2dZzKn/Olm
+tRRdkKR0ZyJoC6+fU7nrbPTVduBRWW2FukNOe8m00qrVksaD7SD+mj1k8saKRgcxGmKu9ZlGt75
ujbHQwqE3LSWF7weiIVhrGuGQxtjfk0KJdstxFsyjIOtzWpul6/BHc2GmgqqjU/vXpWRoJqXsoKR
4Db0u+Hlpbhz1yDEFI+hmN4I0HCoAGz1f5yCFAxIabumrA+PMyXXjC9AxCTm9hMoEdHFBByhD304
nmu6eSV5SIOVvM2az+Gwtl7xkf2I5eAHPA8jhlpGTMg3TpNndIWm1TjDnC5TDg4lG7LO8c87QhFb
UWbCzB9OAXea7c5jfsoLgy/SK0jY6g6XEp8/zCyaq7OWeAHd7U+UIaDMCSJMxlXbp4B50C8mBWRc
SEhE8HKrKqVNfW4ojLGLQ58IyuClXXD0mhEA8vobAVnUlvQLb+EDwDBt1tSIN/JuxQECyDzUDSWG
Eq1Bx7vZFbBtSWO0KJNpy+Lfujk+uy1ELt6gRavrhs72vEdm6lHKlIhhlhJ13eHkC1wxWuDt95Gh
+LzKuKocYXDfQxSld7zOILo4Th3d+l2b6b/oJ+zc85SHN+d8Lowv/XMGcGD+WQPGa3e8ADMGtKX3
wZaca2ExbouxNBTqPgH7HaC6fkjYgFKkodvD0nWfGeK+WWuxzkLHKWsmnbJjJlrtbjhondqxAmCV
j4ZEBIzc0URjHcrHOWONwCM+WxW+wlXfYQT7KxueLuMncOnUXaIHXes3GdBqm4LIsXXN0daOdpzB
ad3JZEo83c4zLNencnkBLa7cuxksxiOYPqHZauGTIZnW/tr+k3X6id5LIAjfFi56zt99toOPKQK7
6V6ozr0otXk+PSLd0T39bNCcvMAmYoVicY3nUTvpCodgF7Dkg8OBcZTnyDMa10Llja97hojY/twS
QpiR+JjmSMxYrcYwsSyChokAyH85LmJ5SUg8fzrWKHTdg0yue6JuimFkYDrCCeu+vVXS9oNiKU7E
9HfzVPC3GhLAyjxIn6BwyXCN5DdkAO4Wc6Z0DkKf52kQ23U4DdnsNyQ1vnIaefIVmzAUzZkEqon9
zrqppCyBUwsf0c3zWTVDnFZHgSnwwBOFNu2Pkzyddj7WfEOUEPbYFlikvCdA1IIvHfni6anpuReb
ZHIAC7uv6QI8DashSsk8DEo6cSYsJOO2At3HbYto9Nic5c0SZeuci+ANAsY5yuXjURcLJYu7Nd/B
U3HAoubtxm3LMRnjlHWF6eIJkWx5+zBXNHZLgXk81RYNaLvp8szI8JTK84WIMI1eP2FSP7rkeTQf
i/ZCt6JH6WydGf4Pjcm0tsRWdXcHNSST2gWwGcjk2lgQ9+kzyfJyUAm6Pb02+2Yah8KrKv5ZofQp
uwfDoIznhJF9HOz1wZMb7zgx5zEdP60WUO+NgWVY3wnIbWKl4qy+0mIO1tuoI66pYaRRsm49CPMI
iC4sSo7IgOmi39EXN7rl82qHxWRB39PxGVZe/w1w8ORjWxn1i/m4j37D7xWZ1hD4X/Q7iXAIhonC
spfDyKuVwDP6X3lkdqmjNs9Rls0AV52NSdQGO+Vks/WK0/pm+HGqPBGIHVWEB1BKpTuNfzvligUW
MpzGijQpZbziBM6N8vF6Xmv2AvbP9k6hJtTTy4pkU5M87dSQjpJh0vF29VgFbSmzwA3zDlaIhUwY
ds7usQITT8KPU6ylE810eOnV1JvgE3/dGaYQLSd6mhhecxvE1jz6nntGVHWh9u0WLFJ2jBMoCv1k
uImeCFB2fs0gXi1moj8MV9nnnUb0hnYd/uQDSF7F8En5pYzKGa6tECJuCRu0tJDccR4dDzu8PNB4
kr4cDjw0+g4rDG9iFZl+p6NjwWgYOjjViL5XbRyDsp0Vc5MPMHmCR0oHD9UKPvD1sw9TIfp9lHRL
0FF6A2MlO7yKw2z/vA10od5I5EaFh+ZiZrYDYNE/TWq6FYnP+RPVjr7FOf+iM8a6GHYkOtqK2Hc0
k9c1sKvNZ83R5hOssXXGAy5eHhZMIuEUrNePPBXPmtGw01F/N4t+yWkYjTczgd5Tt15FGHoPSXYv
m88d0umWGtu3U6a7WIwkuzpWHU2SlUwDfztv50M7x3DE4iCaOVkG2jNRBewJusvjf+YMtksxTNN2
Vi/ilihGdCH2PCUDZU0/mHhEcsRIcKjBB+0lcidWgwxMr1cPAT54Ke94eto397Nh+Lc41cSpE/Mc
zWjO2MJrv1pi2umVD6v2NljL2ZYQt85HA6Yg0adL9t2sVc0pRJl6AM3u20oeS9cKIiZ1mPNY3H2T
1bDSyWh6Vci7xoiiBbhCKNdbik8Jbp05aHmZvo0kkMk9A5mKVNELAg3QhmX54HQcTySm8w5RMVP7
mLZdxTrSmgtED2hDujSy9/dywLnRzME+Luiyrfkc0fAPtmBwhgfrQxIgJbG7jGENHbA4xER1ipQt
SC851Eyncr9m4+1WhWM1gSujRkS597uPM2e3hEvlYU8sTbCNNLCgguCTXKyWtC0Tk2yHqc7g1MoB
3WMXwmZepNiiCNT3vL7V/za5KhmSsod0G+OpKwB4cpxKULsWeamwtoD4QcnmmRfAYFWYVr0SiDeC
VR/DFtsWpF2R3GoQlhyFJgn+53efpDzsaoH4MGOmsWWIZpOdjaDp2bKtPHUUMbExEqy2kXmWn4JW
jxu1vndsqlAQ38mtOvnWVJlP4tDOuZ+fphD2MUQZuexLzQnZlUYySIuezktPyKZI062uB/liW/ju
W/HtIhMIO332X7uI9acuCMM1rEikkmeGHuwWCgI42JZJZM/JFLdnOc++6AToGo69Sk0kNtJQpOQl
2YrUYYu1R/i/FjmA4XUlEUvixoQ5M1GycTu882EyhwDPVamxClumYB/7yXYTLWZ6arBHqNlYIuRn
n5rWQOf3elL971SYyiKpbfeWm9TkdTYNpSVCY8Fvj7Xqsw/1zipgzLndMwvfok0oFrM2MqRbUyVK
vQk0CtDmGpMUJR/eQfQimgTeKh+CKsJ7kx9aaJuHn/ntNrUaPzBCCGnZ4CgbY2RPA+ZBqUGD82sB
huJkhWTfx+2RbNLWX9B2YOmlo3Mvay1ZFlO/QNr2zFaRm+Mx7C+IZtD2St05wrDzTe3o8jEKeZ20
fApJec40LMZ8NaN0lM0wKiPWSBCjT30J+qJL4cU4EaHXz5UWh4clqHETQDD1ZlEUAd0RiUEb0Byd
wCCgB+/hceaWhWM+L04oySDGcKmeik2tTHSwc/vRr31KgO41C5stHE2CW88PP6lKl7fmes+h2wrN
aR1qPEIiZX+nTtHfa4pcnWKVGipLsGKF9GJxLkO5R83dIaT7+EGsoZREC6UlBNSTzTnSzTMz1Oce
SPuL5DM8kPF0M67xvx7KBg/ihhiADkWGptpySwUDeeASUkr27ik8PqIGXgfM5sIv++7Y4b3a0+rl
wZqwKxwncPmQMbWsj811PxHfBbrnMXyv5dmKK5zWkv0UtGF/cZapqjgWFtzvDPtvRKuSlmUhLxyU
vI+dAh3FeAo97P9bHWl6NLU6RlxSnVqJVgswJOyEmu+FK8BMeEYAzgF+6XjxvM9HPNfFBLwso3UL
n+gE/V4VSB9vYK4VIuDhj+xZ4Bd5Xk77L3KDrde48Ccf/aw8rS35FlZuLCFeq5lFGW4JEXmLzcZf
aQBweKr98+iOublqjloTR9hDTEHUzlqboyRICi0++K37D3f3b1oLk6RxFAthZylTcoK5TrVDVh9t
Tyig+4LF22H1qkfnDiISq4s7Pm7P/H9Vc/s5GjHWJi5GLDQWCt2NkpRoqrWai43hGHNHa/zg9qnJ
8runQLfEq3E/SL+5I/i/ieDDMX/LzP+LKnRQIyvvxxTqIlhuK7HXbl3FFq113naL8H0L47bXVMzH
tz+xftnHtMaBHrCMgiM4snSS1LTP5PSmodUrG4Ua+CM/ffjn3uTS3tn6CY3sfar6h9jS7rkulkMO
HLfrHqH29c+vFcbzh8d0KcmejoIXj54kOaf07uzdu2CYPyHIOKPjCPZ4qUcaL9JxVDqSUCMrEtwL
efZRymAG6i+jvqOvxZnShPzsTsCwGls60pakGU9LAlSCtbngXr8lj+3CZZFvby9eXGPzyg5Aw5Mg
tl6cf76p7QqIMTBU0Uy1HF8oEPpB84zzb4WEX2NDsJKiKgDCoPIU12PE1B87SuLjqIsi4PuDQ3Mw
uZLte3sHXPdn6tGikWhrwJxN5gB0t8RyBF9EWXcXrHAjtAozKXJ3uOv0JhL2rVTUWr3a2bJuvgqz
JK8Npcj1XEqmWD/N2XEm7H+ciMIVdREi2p6iVp8tOb27kDQItGcaLdaqgq2K2BbYQDVRfq+z7m2n
qu8AEQDXEwvTG6cqEE3YjVu3FJYnRXM31A7x7EGWyWvtj+klzBodKMSYBlqrv454STtmzdDZbOAv
E8SGfrglWRPlKs5NO1zgoiJkwYqHtEGjWwgSfQGlQZxfoGvDbOGFiRop109BZ7eGhBBAy58mm9jX
bHuUcMQla450zacUDCAlQG2H18696aracnKUgoDIEJkGCt4niKawrsRae/P7SvVvdtzYzPppgHAk
5IEbVDjLvYTS1DL1fbl7X1NhwoJSJ2QbYBe07ymTezjg/x2th151R1F+30l8KxFwd1KN/XebjAko
/dwdTXy3VmN7dsim4jXk91I3MwnYZJgHO5rwvDBq07MtUOXVDuuIy29YK8gKPVbcEU0+s50SRs94
yvpaA0t+5xl7yvkYEo07NoTJdVW9883j0dfOnUb+c54mNYXP60uV1DdIHv4jT0Br+dOA9Z7pBd3n
iDhvsa8XIa7neGGyNmELvGeyBTB9y5HMjTrxdqP5L27jwr7O5l+dxFylZ1bmxPeTBRlkseu2+xps
nIhSfppGcMQEWBcTTf1XTW5s7FBS92Cq1mq385mSzdrCDFgvwaOxHyOmG+4WTHMH782P36PQL3xG
vPv9KasDEO6iZKMQHZHuxyyS+CL14kh250LxWkjwgdBc1hWXv9BrFj2XMh16MkP6Nq0AV/uhbISA
z8tbwLxgb4hWpxeRvUx66RstK+UvY1Xh+4ktVIigfghSTsnoCw+xhX6GFZXhUXzTbOBdCZICWSCA
nFtn+kbCtvaVJg8sp8k+WVul1jgy5f9ZLngNceeUOsUHAyBcSyVDay34ICEDXkYzaXB2/TipShCY
3WwpHsCbp38E5XTV35/7XvGUb2mzmiJjTy8v3rSV5aNWbCugBvRtQC8o49gioHLRU5C+UPuE3cKJ
X/pOaJC947H2FlRwkGxzKAESx/LuugxFXbReieUgBnDN7ioDjl6G2tu1X//FtY76mTZq1P6XTi0+
JtpXpeJjp2XurjRf7WTbd2/L/2zwQMxQYvDnUgwhgvZEgeEnA+jLwRBUshOQaszc6BZBqwXA7keO
TkNOU3UUhbKelGs5ev9xRYj/wQQ5kn9t04g0bKtfNQGqLFOJVaPGyBhMGW8gBjoyVa9mXazDFKNx
VNml4yCdqeSxBsVRZNectF+ZIEr6ojaAENLGKjbvc+ncaa5/Ax7+L+d2CFcE3C2ncx3Krwr3LOiu
SgjySevrJNx4Qe8c0boZnRmFgP20DAB3KjZ3JXVX8FaHmnRoI4jFEKCRpYpr6vQOcYsl8yHMrFWG
OGPqnDRqtPN+bTudgmM/LODfbXnLQkYrIRAywy0RVYiTMo0VGqIdjrvPdpRFVVpud49o/S2HXCmQ
F95p7i0vpCUH1zo+3JRFLeTsDvqIIasfcKtlmUUnm89XUHf12E3F23FZgqROxcPdO4QUkpkgkkVs
reY3s+YggBBEbt0SdoqaoUW0k2/LR07Isv0sLm9sNE4DjLp9vonBciWL3knv7mOB5ZL0SChXLCZ4
mY5mzpDLJpweVnPzYMr3CFEYZ6U9kok1YGdE8+rA8pGGSMqJx+xSxoTLYHgpV0cNEXYrQlUOxPkQ
ud51cZ40DBKVo0MmPEZPx5CJ2eQiaiCA/A25ZFT9/PZEK66ah/OgDFmen2gSKnpbmO7GXvyjFr9z
XUWaQI4XPjeqdiOPRGIVejz+d8xem2fz2Ln/ba3ARbo8jlVqu2Bfd1rnQ4DuFiMEbCCMYHk/NzJB
7gpdo6lgxsI1KjhUWmrlLv7GOEhLxe7BRXpGxOaVjI5DzXkq/jZ7fGZoiDie6SM2YmfQwjnSfg6+
d3CNcdYhJ3E8yvzq2U/Eq97//j75VhxN24JIqsYII5mrdT07yxAV3/46rGv5COyM26XRQZ19Qi8H
KPbTGWK5/7Y/deixEtEUm8vdqD5jbtj1rIamAnZ2w7O8ii25rih3EUub92UhKNe2OP91oFmMKFP4
P68if/NOjJDs6BO6hjvKUm+s5I74jnT5FJXqgpsafDemFtxfxsgqNHREQzSvkw+nh7N2PORpNmE8
hEBrzQRRYwIpiltNyq80VIkL2vPseRmt1+lfbFoQd5yrWTvMQ9bWfpwMlK09/0zUodhqMYEFQ9tY
6SiAGgLz5m+OHJIrnGIYbHXHlzXpKzfdJhjiOycgYkWPKH4Ja/RBnGeSQ7qrTGTy+uRD7x5wpg+4
E0QqXQ6KtqcTlpl8olpXhQ+tJtsX98womj3n5BH7PoPq86xVJeYCsc2emAq9YK6mEjRfW76G0U4a
J/gvhPWCaVBZPPfw3jPv2QPXwt/syZwRMNw2HKOXwxwKJ2knWy7JjkkJsD5K0GL5T3db3sXYmSLj
Po34ZYxruQ71k1jN/7j1jUhixljOBk8ooNffuQW8eXCd2By8IOSgPgLjXXbLy5rvP4TL5ydrk/Cu
ck6q2zqaczta4c1YW4KgoBoKy3YLlBFBhIvHGqtj89vtr67WSXQZSE7bsMp1TAzn1n+Fm2JGHmG9
HXJuH3mFgJhKgoVDEwP0Gpxbp7Bn/IM510gGQsySnHpdgaCNVPDm2/9C7mrZP3jxljEX0nR6E9Oc
Lz0xuso7A2Nl4Et7n2d5pAhdmrS+LOzJcgA2Cp9KOjU5bNgG+YLePrFcMVyIX1rtPfcflTFeG9el
y7yOLbplxqx/cXDMMIBerwlpB0HCdfhMznEhwInw+LFZPLqtpb2ZaVx7MuYXznxfudEsoPXmk3/Y
BoDDrJPhtyCxuRPpzQJVcNOFusNKWFlcBe3+XBMpLM9oToTgUntqsIRJAZS62lWnnmjc2PrpFqhk
MU6fisLcQYdfsFHpxwof1P8g/anOT8UAkoaC+D9mOvMgigj1gz589LyUgSmnfLUZPLaKjBHeeTEW
B9tFnS5slp1+DyMX4e0izd/MI0OyjsahzSBMeZUKvc9M1sVljQ2spWGTO9FHu/pTBnkSJ6b+v/XF
oA8LFBRVUN9nlOWN10rIMWuDbtaw0UBNeAYzIsDBwMvl86PPPcR0kC/rZrL3vPR2MYFJ5AFE+BbN
p/BIWbHmFxzHK3c+QlToUDP7dTCJ/9jB2xVyqDSmJ12G9fe/OEAE8vwG28bBdNu2DrCH6VbgJDHK
0KWvbB8wOWnnBhhDUP+ln/4SKIQ2ljIAHEyBeZPzkcDk5+SE3AU+wpc5P7XtkN+aK/H5UMBRE24D
iHhngOKskWFmcrupJKIsSLVY88hPT+CmarTgJ03DkXlc2AJSpHwYGfRZsqpX6C7Cw0fk03niti0s
cZn8FXywFkzC9fGEx89ypSMN+S8ieSJ9Axzd35cKLoDZepzA1Q0IXGnexyRlHbk+pI83p+F/cuTz
JQXjJhy5CljAaxudXIXgXG/Uyl6N+KDDvIPLhxZQ1V/N6+5du0gifu6o10+li7fv3o7Tx5ue3ntn
tspuIFnMPtYDxx0BByZOQ5TUJQDqrskcB7ZxWprkhF23bUihgUkDROuBR/TClXIyUV8bscIaJjAu
ESb8u027lsZScJ8pD1sBznO3cNdUBUUQPJUJwJzBzZT/nL2AH3ZSolBEpOsStnyMy0HHjS26EUil
feEX20gKIxw4VIaAXRa5Tj12w3+6V4WNx6YZoXadItqX+JaRvNbYRtvvucE89SXkbW1/BFqUbrcS
8nThseC0k7Hbwy9EKqo2fO/JoFxLThUYb56zpgOMqm9arRUwOJneoGC6jBQ3KmVBs8t9K6EtSB75
GMZIhkdP8vlFpOV/cxQCdHshmkc/W/D+uTmKKR7wDTpIIAA2a1/SFqgqmHRTc+behxSg4sLLv5KA
DB9GJW4ITvLgIvcnrN69koLNXM+mkysFKKUsEElgxNy/Mik5DgI6dnUQzUajG8rq2uLuzeoM3GIP
VI5UAFqAyLEHx36WBr32Grji23tjpjaW7LJGFJFiB13DlXV0o5Yz3KgNB7PKZUyBbpwpOhEd7dBO
TWyYl8V1cWlmu9HjKr4V8IUNfcTdqR5gApSllL2obtg3PEU/nSjOGB43C2QeltkNoyFi3wSBTKbn
3Cqd7UsswBH4UXEDQWopI8TdVohOEIQYQSZQw9hvvAxe3hjAsfa7ICbPdoO1UL6gx1LpLGa1VcdW
S8kutfNzR3FoKeyo4g/f+9wbFQtOOD9johyIWekL8F9C3SygtMEa9if4iLDJaay23Fb4Z3KPGCbV
cmK70O2JwxPw4TVuviT5NNhJje4/dxxa9paTNhcFU7hl4pgUfKLpdxVhVZ4zAkziaIquybI3rNGH
TyNUOywg0p4Z0wTG4Jm44muGqdkcx+yMGRY1pmXaLfiPo/4epFSCx1emrSwIEyPW7SQr4EznyeE1
FmfF3MlOQmYvEGcencvF+1xPZOS85hrrH5HzqK9KIgTjVf4asE7sJoTzmXU7Pt+jfeRTsrd56lr+
79Q2QJX8UYa7rukn7YR4wECddr3otzP3rI5EjtDj3LLUmZVJ47JA1Odfx15/7SgvFxWGKBQyqD1e
MTxCEsCNdx5/Qg8xlvtS+wO5/rKsiU2KcSg9QUsoWdzUXmlVU3xRuH3OnvKGc0RWbWgo57vQECD1
5qAQvF/buFKPaO8w3mtWcTa52Ms8MIWfVf4Y449bka94osjDr5kUBHdj7nb4G3KnzlD7jucgqjoj
rT3aqaszMgZ+1KFLxIKfRsTeD2rPERB0iqOQO/a+YBn8/kIeSSOU2NXkpQjp3sNSqiEpxIcTgY0V
Dyv+lJeCVQXUR2P1G4KlShNGSn550lNHYKDpNnBYOXwp7NvI5H54kEkxcU4PM2pzThaQX3YrMSc5
ndQzZpWtKabpjaix53tMv4YBgUZYWo0zbbMAEFwZNWrbkqtv1mnkN/OJpPH0cQzeMggM4ahn9xW0
9oi8cc4v9Xsc5TUO9oyfadB4MBwsye6NO9rWyKM+PA8R3Et/jsuNAwXJ/HBgsgw8OwemiFfh8e16
oVmcQ0T6hB96nd9yoOBd/1HzobI7xr9aW/4yeVXRI6GT1cAIwsRo/43qQEg3IqhCdYR7IsPCBF47
2VNQLaAm4U5P2isKq8a5C23va35i4dZMUKVWO6jBtW+SqQG9Q1y9ttFiVlSyHYyER06EHxz8rtYc
twjNC79bhfFMEN4VNvH2dbUAHTDT2VDLYoXSV7WP2j2f3lHuwaTGol3eEtMj0tjOgDA9YgTppcVp
5hbC8f2gyFZVh+wVih3JG+xhvrGC4Vh907ZfxDrY8O8shLklPDY3o2eXn6zfAm0JlLFs3GhOjak3
e2olZ24PfS1ooZTKcvzNCi9CY3ai10XcnUE1f5ST1lVkDa08M7n6L2WD1XJeb70oLOfJIWPqVKE5
V9Iuc44blS/oehBGf3LXwbP0ldlf8M6YfbF91nNMIc3CC272S6z1yMuCk3d5pMA163zqw99VA4dl
iDyUj09/JNRiCisT2UdzjCvMEeualEW4pGWw57e/9RpsNBoT8zkAPlRKqpsaoVHuxllCX9RbXxui
I/TgXVQ+qG/L8/a/Gnej9q2QiAfLcwr9ZnaeM+HjBqpEBCMSw4NkTl5yA/3jKy3xjgLk1ur+spoq
4t28GECgUojpVAtuQxFXi5ywVWGOpJ+ya7NLVSQTdR4B5o8hv28xsaNsQltxsHZPUyP5XIWZDtso
eKVbG1G/0wTmW+A+HXnb/1b5y74UZLKpFVnUfxyGqrWA072N8jnv+MsVfMRHYtiHxyQ5gmsIyn10
Nqo2jm4kFr7en6HoZ9Kzfq2ewyUtnez0oz/L07tJatAXIfWjgAahtsemjLALs/x75iIIpDeOJkUM
g8Kf3FrRFnZ3cviXtZlmxAnwxfw/Uhwn4MkZW3UYPybeUW36Zwp3fcIunkyvJJ1YXoGNawQz002b
sv/21Pap07FBFKmP2AEWxAkkEeO2Q5j3iD+EilRVoehS3BHfonWLEjgJDJQB+msjMcfmwejsKBUC
YXnU/V/ZIYeU/VFYDTbIE2ngUrsXo63rbz0W6+rps3EJrzhwfp3E5lUkxkgYPEoqggvu3A5OFZwD
ansyMxNDCmpbasrW/eppnzk2q9KmdpKCYfUXtv4GHdMgZqIhom34SEHhmA6i6Kl4+aOfUu7eEbN1
ZK2jJZFDKRovG7e4D00hbAD5nbzuCsfpQSyHoaQZGXtBlKT/V5xeAIV4goxfu7dlwCZSANVjnMSN
nTTlK9UghPTZlccxpdhc6zy54gG5b/rGywhSI47xn230sZ68J3ynPoK7RgZpoe08bq5IMTHwIi59
GX6ni65AQd0zS28Csk8MwqvABxH9JL0LMl5i8PzDiCuAr1K98YHRGDWuCtFynNVKkcSoC+wqW9RL
5CRiaDoc1+Io+H5fyfQNNMSqrggvMKLyWE8NReNAgD0Oo3F2XUKFupv26FpVyGygc5XnDv6j/IVh
lLu82JnapFXv6NmdayFtu5exVNrN54shomToPfY/58veQvQKCz5uX8mcDpTMUebr/wuEMrP2DXpo
D/slyxZW5YCDldgsxW6Vp85OVmoEn/4rCOX8Y55uLHCbHrSHY0kTAM5XE+Kx1kd0nCtCHIyRYl9x
BEecXtNbCVI0QK0/Q6QmMhJ54AU2oAKuO/qa+jGdomD0TfkQgoVJVgXhjGCdB++qNvy1bVO1fL8X
ZZhSe5zOImm8eyt0xMGsQwdyMsexsi3inkq6LGAe/GM1bPlNnv25urN2EldMO7dFao62VW69XJQK
N011uJcIyi1RSnQMmkfFEgWkHp6mxd+xmNe5G7GN7djkVZ47azQvHynrjgecgwDcfgLdUpwBXBeN
7FP4ePGFJj1GPFX4eNe+/LyK+m+/OTcoMbs37cYXU5AO4/uDR07aceCUO9nEgUkUgXpylYk/yg6u
bHMFDBkwF1A+k2HQPOLhlJthVw1Ccsh/IaqG2++26joIwLMg3hxgFAbmIpebJwvbGrEfPR0WIkLv
avmbS6Qyqnqhz8t9JtFEFUwjcIk/7sUdnZpyN3jmtVkQ0U57VPlwSKg/evJZepN92rn2olB//jfP
QBiXRu/+z0+OjuGjJeWepMaK0SO8uY3TKBNaG5zLDDEEVOqhWmbHcBEGBnbWVPanjX9q9G9phxjW
ezuLRHtJuGuYQjn/F35BofY4GCs+hRBsjuo7hjYa7kzDly6fd3WsQwrv5S3NNHiBxnciSPee0zrF
QNMd9SxeXgb0qflCpY1TL8n5w4XvD8ZghYlVHN+Yt1q4qbYM+EmXNr6T1uqq8JM2eGD47/aXWVmW
yiU9KysvGbKsGvQcqpPBV/XUFB0pmnDZwYDgPYTzrpb3esXQSu1wF2WyHH0+t5wTVrSy24LB9xYO
lH8grIWFlW/1ajeXc+57We/dbcLzS48aJN7n8LkP3aLqbHrLJHQP/Cq37BU57MMagPb5uw5I/MTC
Z/6bQwFeRrL6eAKQXkjKEsQhxSl7/sFOjxC6HDoxl5xy8KkhDCfXBf1UB0m4NZFH1Y6f80KPIFCJ
n6NVVS/IF7gjv8kKSFOLSfO1TbG49cyoY4+6d1JsKq++41OiOro9jwLoAtGkuoT3IWeZsst4L86h
pF5WfdSvlaoQ2UgAg4RQZu03S6wSYw4eMOnNqQ/0VVbSSZmpbwQrlvmxxg4AI2t/wo8qsZcDH4lh
VyKX/EM5MyOM7mDaTlU/rymDHhmDfr2tUWEEjNkRemxk9elaWnEG9vjFB395bnkCJGLIIM+ilIf3
I89z3D/6X6NFsGv/T3O77xhx517c3IQuAJ30G3JVql3mSzaZNbbBzWhxMwiCebqALc1mxfpYGLkw
APJbXdhH1svvx9jTfyIp3jqcvfzi/N83qn6HNiDF5E2mH+ZoC9CZsillCvpIBxqOHGSOh5FuV+zM
aUxiAk2KGZjqwcwGyH7wOU1Z4rd6Gq2ciVNMzFlZYO0GnsJwf2N0Bz0cgNn9qxwEmIct0tVYmDP4
z6avH3yQ6Ovb1aDi5E7d/I9EvUeH6jwW33feChXi5tI521d4EqSgAcSeBBCr9VuuEcUIZHitZ6oU
ssIIaCfQyqO+gv3eK6eWMT4NNfPEJ9aQzGbTHsrYl1F4+EjdfEo7Z1pNR+ybw04flfQTLmoMbNE6
F7/yqEKk0ng0TTUAO2bgznpUDSfEHY1Laq568odpoEkFQmCqJWK8wRCG1xYmO2LGhEYGLmLisw4t
ijeFdxYmWClsd7Rdb28J7XNEtsh+Dedv43jadz+lt3hGR6tEW3eEk8Ygn/zBFzCUZiMckq3zMBLa
kbN700u1LybhOQyTBzhWiYplAxpmHXQFi58iL4WOnG6Pen1z9V5TdRRQL2/ILX4h1ok1HW42ijvz
t9CbMU18sv4/phUxh9LRTB6n8c15Gt5gMGtShE7iV0ga5at+EczUcyv39earXHicapkjZs28N0KH
Bjo8ezI76/Eka4GwTAngePoH6pPkHyOnA89PMksghHsFh9iBh4ycV7MF9RceF90FyLOh7/tm4IS3
pACkMkf8oVSSCf6YRNtF1clmZFkp+KNnLrpI8s5oQTfhVdyBDGRFyPNKNeUaiwIWbTdLyuRkie64
7Pl9eQ1pci/0XnVRTq+bsr8LYiuSjqwNSvGSxdzKTOGnRGcH0UxnroeYDSi5+LJs03+wh2KV9aIW
jYbPcJCUCMXCzOiwZICl6FWQ/rF5PC1n5gnXdHCiJch8Mr6Uy7vJHJDvQa46cB72IBymmkuKp40z
uRP5LicFi9XotA7cqaQjFQGxBvmebh2dtQMTDhPcv299XNHokVH0C+H4YWDFyEhsDcICAwGA0DbF
rmglAxxP3qjHxsDyfXZ+YtxNI+iWebtHVITD4VGqNyQ00SIbWnOYj7F9XdtrcX3Klkq17iVCZoJz
ZZGFoKSeb/LnSOXzmN3bXSeqeeGZFGAi/lbjk3wVuQC2AToteqMDcyfwT6gvZ8CX/t2Aquz7kE0l
BqVc6j7xyUkqDlFtFzeluCiA1CcfVqVN8M/iu1UOnw1aYXXzjmnm0m73HwklGWQutrVWq0cbdohM
S184IVAPm9BrQq5I3oOC3ddQyfYhWydsC1DdSg1f9Lk9RT3eRKnzkxWmJ0GMyNnUQh6RXtz2bO7s
E+2etSIafs5ZmeB2zHrbE64TfieoIhxoWR3yuE1byYJgc3zisoVDLyvpb2kktishdZKs6FpdGoCz
5Q==
`protect end_protected
