`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 107920)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf+kF
201k+6QR2npVEY+494p8x3Y/iVMzNwQUtTTNrheBLY9h8bbdcsKyZaY7KuUU5K6Dirm5yCA5/cKy
fVLBS9aoQtd0++VTEa8JiZ53ivfBgt7O4dPUrWryf2eOg6vahaqyDuI7QijBHrtM0mffeC4icvET
5KSC073iVZMgw0Z2so1EQzosT66HOudBmWfbcElxS81rk1QZh5OjzgLSlSqxFjzcvu5rHGpQcO1w
qnaGuoQFnWjNoSBKSrzae7L5Ftf920LUqRwwTBzn5W+l+2DkbVEJZz+vOcY+z2jFD7aZSVSIIL1O
wK252YqFpZjDOVCgaCNjmWl+wBEtjhptK5mkqHrYNArkesBAdxwMDfhRCjabFv1GWh70PaPBrtHy
xtLHhcUEyGt7Uj8Fmi1Mn8xu3J5AduHH4kLys8MzyD4ej8sIYC5BhdMOlb3/CzY98m/4CPoSQwyu
sjIOavnwCGYLV7tPkxqjoNPcVUVBnlzeyaty8mR4fTzgT7pn8Wxz+qWAsToBbfvrc6yc3ULGX4ku
9dE8qpMOurf+tzHgL53mUigT6wTpjyH7LRseYHKs/I+f4A64mNXBs+C+wg33fvDl3yxwqkT2ylHS
f+8vkTjh4OjxEX5/khVWDowb9+oeSWkSBf4yBU+yZl1lgHPXI1ZIZFq/JuAqi0csPmmmU0/RT7BQ
su8VulrppPO/YlAIDcVi3KwVtCkmaV09z+FEup4VbeRipyEVpAB9DUNaFCyjAUcVbbvJfBU2hA8w
HKD59tiRvlwDA3gepVbAXFmrkujLlH+Nnk9ev18QubE6mC6zPq5jlIseDA0AissvrVnHro3KFS2v
ILX2Knnz2mrAqF+/AuP+pK4wC5wObPpcPfDhW9v+4Qh/+NZ3GaxrSNtd1aIP5WeTh5n/KNnyzEdq
JvW8IbWoCTAtpP72fQ5ubQmM+3KfXOWRsb5Xu7TDPcqv98ppvoHv65QPJE3xuZo+GzG88l5+rwzY
E2XAaZTXdlPaRovahkaex4mC4sueHo80tLZsZ1tHoxfyfLMWvexPlKcMrUozBrZguFUFFh1H8JmW
z1TQVNjaFSbB2iUtYLi6+jAmgI46p02Td7f9qHQ5mLtxNTVRDsm7xin92m3Zuw7FssYfS3C5CeVJ
7JWLzWONg3oX3DvDQTDMciBVFD/eXOQaLRSWHGlUcAClcE3sRjGND5xHwdAjY2dn9ZfSds6CMCpp
aHMRUs7bR+Y5x3bYi5TKR5XRBJZWQ0oYN6fvPU44XM1m9b/TiTjmDDgMPcpEs5NHbvThp5RTBTFF
fyxRkc3sBJ8sQmnDvexsmuqMF+YOcYItTvRQbUQ7InN8lFxYOBgrqCCcw4pQ/tgilsEvLlp0NUH8
lzyIqDiO11W6qDj+0TG65cgOIp5J6WDm0wh9lRHAez61adh+TsBGO34N+Wa0eULto2Bi9S8cP7iV
KzghSp41zR0YAxhhP39z5N0TEgC3bPkARRPcm9KNf8YhvMZ33qzUb65iGTTNiH429Bdg3+7W44YY
JUsGdF/N0qh76zCkeOItivpfI3qRuK64rYBQhJs5qpWKC1qhfgemW9wpuLZiO2ISTipGXEi1DtsD
BZGzbv+0eG3Hhu+BhVG+ueDD7ssTYjddtmu28zMhuPAPSGdff9v+fwDBAW4jktWT+BWp6+F1MnZi
0zUrt1GZJzUHb6T0BTKaaJS8GoASN63u7d3ceXypFY/BWQfC9G0y3j0AgC6eODj5OdkMlf/HwCDE
QrEGgBOY3qDVkwLNKIkqElL9ECuoTDqOsrCf71a5gYiyVPBVv8w3d415XWHlIg3mSyCbnMrR7ZcM
EIvNSIWsDlbbrLA47zF6C/JwQIJeZjsns+yf9HZQE41iFnhB9XOOTP3iUeP6U1IpO+AYBRhFRTif
ih6P2IqINzPQ4AkVcpJ04F8fgcRJ3j6b00Ts9jVOF1hwDeEWN4EvTDk8Wn3xGOpTDFATHiotto+R
2J4nAQFAJqUY9GF/zah0t8zAecoPynXYV1hDZ540oC0Go/Ohl2fYhLi1ONmJjKbZ+6SIGzwj4+pw
+ULkBGGKQT3NbktDjus7X1kWFzMA89LH6uSwFnqSL2o3r6nAlj4rPKvwzgl2x6uLdZnE/aT2DgLX
yWe9P8AdsgXhOQWdqlf3I40K+2/bnxLT/T41QVADtaeHw2h8sq4FYkOb4l7hqjwLik1eVW4ypnaF
x+iN/m3AcHvoiUoTR3RIfwfx9YukCYBnW15YMKn6/+0BIc5gzoAFryIayPpuNOIueIDTJNrUoerE
NhwjENn2KmulgrzcNP/DU8U2zUq83AkE3Pief3wL0mcIYb2WVKC4wgRAR1E5H0CIFy2q6Cj3tb8F
xx1cV+8hRwH6Tsu3oHaBXs2boydZf2Gp9jisG3qH2i69+p5ffs4aM6JVlu86aICxso4qcTbrxaIH
iG9zSm61JOEU/D0wiZUmIAx3wcBIsyDBoIX06XbsYmgCZnlv0w4MrBG2g4nIOyW3qRSBzryOo9xy
3f3rTjnb43onJ0z4J7TfcPCg+LWv2KA1SOQOa1Lnj2/HkAFpeeW5Xh3B65m0D4o5PCUYZwfKPYLm
x/7uucCYzenRnlPVRoSD+5YVU6VRxOd3pgMLdv0nGgfGxW3/PE3yrMdT/PuZBw5rV5l7zXog4ZCQ
tKlm1okizwuS5r3Ni20wp2MgtTE5Bbql/UErzda3ClTEHn/atSfu8OZbib3IhhLMqgsoNdvXPbXn
tT6lRL4nj3pOry6uqHJWRRquoDzUo9apJgiM7+/CG4yaJieQ9NeyI/0QpcQHzvykvD6Up0J3xPOR
uGXKX7FpVzNgH3P5hHjsW6JjKgKXKviLzLcntIaTb4plmXfXuH18oMrG1QbppJxboG+rbp8KzO6I
+UpmQ1WcvYPI0yB/5PcQ2VWpZrS3kUVRpdCJc/v+csn7fAXzl3ckdieC5ci20tPa7Er5PncqVi7f
2fD8wm0OezWs+veTNzzbqO2SOpgMp4QKZPKVsS05k5YhEY2uXPGe7bN470go0n0leFbQqyjN9vL3
Ba/0Kbi/VwQ3MSLXr9BR66apvnqF1M7+SVzxCs/slP+4ILqzCWV336TqJAU2wt0DyvbiPwZgViy/
ROTa7nUxJUyLyDw3zAVjR5HGPST5eiDZZc9KeQeDGtonnBoRFaFreqDHFd5hyhtE0u7Cdg/ZIDxo
EAqb3Subz7E0d51KhixfA/Xvd4xnuuImH+Xg/tbJHsamdC4K5WJ7iALxx0QEgkNR8TZZ/lDBr6RE
iSsD+s+6kGXCJsR/R84WnzRjqbZNxoEqAU/k3KRYDDlBDG9p8Me4NQpLxCgiVIxlVeCb/TKx2JVQ
X1CbHHBYmkQXuiJKja5ovU+De7LbHxtIbBQ+4ZbD/w2IswN0yt6wzvVk4e8PMqG76SzIaZNbDc6W
TYrPJ09DYyLVA5Aehxq2JwjQsNTVjU+Na55PfXtcrMdM0yhM6FcRiTBwAnSzJ7GK3dJZxzbKMyfp
uSFQdqDN81+o00HFRMs07ZQlXe9KUMEdQjyiZqS2vm/QsXXlfMuCREwvMj9bz+f8uEKBp6m8H6Ts
S/51vIW7e5SXF6Fed5bbTXBlg4t49QwGQ0G+OzoibcM9YP6MDHgX4bjYiO0xOP9HcqtaxBOhyOoD
5Hfm6McUrfCqPjpGlf3K3U0DIVTd49iHztbwGWGu/stWMVzEEYlWlK2FavP6sbzTcPegWSNUiIF8
N8Jad1oNgyw4GVbnMevMdgkMmUvRvu3GGS9P3xa961kdOqT6j1dMjgRXim+mlvO/RkTDsxuvB5ck
YSL1fIkF7z+v2ILvZlGDaQEtL/X9g/8bpwymv4G5cP/AJguUHxCkT5eNt0oCa5IMOOhpClHrabAi
JSSw4HJGuQheaKhZREWAr8i6aMX/EguS5/s/CYgqUKmewdFbo0rLIEn1h1YtmTEEaEPTd29f9E3A
LQraEz3mv/miTOHJUlStQiKdixMGMDEzVce3tkchIQHIlbb3uXa7EO5+DsfON25L6vNaIv8BSooj
0LeydNnvar8vaxRiUlZ/sF3/ygLibYd5e+4Nfgxq/85m/9LK1Dt21YGBeBy6mXYDx2U9EAdPXNso
oedxLcoYyxN8bjjwUm7Rra+nbdOt5tvN5KEHGxG1O/o8LFoZH9lQx2MSZQJHXNKH1c6IDQgo6eHn
8I/vRAYCOMt1cJyUxBJSIYzhf9ZP4g+F+MMj9buHn1rXnQLVe2NPs7MthGNPgx0jwOjQ+28TFUWL
cNSS1sKKN8TznKjHBOdhQzQQS+oECMYPJopknTaRJJ2I9QtFnG10bwm9KCve1EbKTPz6zdfYVNuE
zQNtIQDyYJOW8o4lrp7hW/q4XrzOFPXCpRt+qd2/A/ZIDe2ZDf0S4zT+QmDhJAjkMkin6xJpNSjF
HMMoAun8YyZIsVXagWDULgj6zMtOhIuB9YNA1Sz5e7tnj7Mmf0GFxHUURTFwDoNfW3k8aj7C6pvF
6RXQN98K77/kRKk661YfjiIPiTpN1jDW4Mypg2aAEBnb4QFcw5C1q0gZ4gZa9SbdHQEEangLNHzU
d7lqe1FSTs3a1sEtEQ6TsGrtfeC5w74ELHwhNA0ktybzr9Ay2CyWFnhivBqJslHGO2rKTe1JYlre
H086/nkJlrO9eCfjKKYGZqIuEin8YuwsuczQi/20OOEucJvnneEBgX0uYuZITPHptdR9zGIUoijJ
g+X4cDheLYrHzxVbvCcMcfRJZJ6GWs/eODvLgOkoTBbzk98/otS5SyOrWdJFCaAH3/OI7Q9+4x20
vnQq8FcyX/2pijB4a1qFJlsWMGsa+W0AtiXH9iRg91pYqHqYXOTxHOm1Ykok5wesMOHHQUAmmzbm
/pB/EQbT+L4Ed6AwBKZvjdptBw1fwYQP60H+gJ7kb5ELc3YVV6B2Xg2+QzmGXpFUmAgyxmN8G6rK
blEC8hwZ5xvSR0EMci3VO/gy7emv0UDx/uG9MikPKeMmn7sz/9crGJTZknXJAzsGdPg9Fk4BN9++
8uK10BSj3Use1zSLcp3DclZ8BumHsbKCfAlaZhyaj6A8ZwvXBEkhRKSDUuhPzgPVvQ426mL3gbJV
PnuUGy0koqt5/EsQuq043AOapzl+GKPunJmxEkB/T9IIfRKldEr10nMzZ3Df5G2Z/42PgOIjV8V4
/vGQ0mVEmhyNPcusQFjTyEF6e4aMupLwzdDAvrjazDqmIbkHWxQASGiVQ7jekGHO4IReH5uz9Bkp
SHOFjeF14/QB9MySlhJpeWdfHoZ2zUP8ZrNR89hyRRNqwZcov1QQe6deRfSCtAuQSdKO95hBFPUG
1KaDmiX9eM+X+sfU/7YewT1LXe7cUTxWd6qbeFcUAUQqGtJrQEz9Qs2DTUDLzrcQaPgZiAttazN+
c0Go5gL9f+RQ3v9piNwVab5ywwIOHjlyPgiz0kjpWHGbeEZi1hg6qb1NacVFyr3F8hz8RZzc1ro0
iStTfq6qPe8UwySMq6eDyD33HYFd7gKwTUZoHwiJ0xmlOVzoxq06l6jQBYgf0zQCGmEMMDgmGDDE
LEdBVnuFV+dVyrla6+gkdXT3OzBDfZc6lfz65o5hC1IBWr4fsQ0ErP1elckl6QvcqHfVfNSFN6Yy
X5r/HSKBgY6DW/z+Q6TmcQ3G6XpYjIvyYuAVKfswTEj0vyKdBnyrBm5amOmtvSN6dfaGukXliPaa
4r1q2YnVy0bNB1pGEZ+sog7gwlAih26butW0D+OodktqXctjz9v+u2JYamCr6TkGw1HT4PWd6gsO
7pA7OeidcKYeyLoRAsDX1lhnmmMxbtWLld2igsKKrRpxEKfLynO5Nz9ABBMGtpHNBxaCey3NJO5j
8lqgdTE+xxBRM9obl2m/XWwI5FM9yo2U69BI68mcZ6NVAhHtg0xbB7rhqWELiE1fZsH1Fi3Qv6lj
UsYfokG8TGQtEi86WjGACyVsEH7OXWNQxbo3mIES8rbxar/0yBAQsO7jgbbqGd97OvrheaSo4sTA
LrNY0WjpbTdco8lMqai/PJbsVpI9gOMeo7guhb4ZdCgs5Y6edbiG565biJArCecBKcq0J91DpUbW
iaa9iRM+25BVilNvRPTqsQucwrYJm307HFWFmEnEihPzxsYDanWVanKyhSrVR/Ggy8KOT6QTaVj2
Y3a30xyaifOcH3BcSJqRQqsaGHVx7XceqniYh+1bcQzXvRXyc6r5+4zktiouTINq6w/NbXszR+IB
nryA2sG9bOjnVkDJqbA7dz1JJZhRsEEo+JpJjDQkNhP6sHHQgcreZiTJxoEsoRY4PgQI6K6u6rhK
YAQa5hixoLz9dv4KbukvgwH6Do5xyUsgcpnjDxVaLitOlox+heP6mId/sXICfCojczams+18MliS
kMfw0An7PDx05UZt5rUbM3fXa5kvz89ubiGw/5afjbeYdYi4MTDjt8MvEzVDGAM6bzLMoSKYw21V
JnE4JUWvKp4Yr+0F+L14UXeaCZXbDCHbJ74ujQovAf08ycE7AxL8tJqPXTf1UgUzavJNBK7+kOzB
x9ek6pCCsdy3zOdBf10DF35ZrfQ5BZ9/DW9+l3kGbTgAg4qo043QpE4ljmMuR14qN7qayMNclAOq
zLTobcqEPFYJLiTpU/jzV02UAHUEB22NOhXgKxDndZuwIKbw63KoFyv7HnbV3ircpawNczT1wpD5
7vfFn5wqiIqXs+PlWyr74LiM6w1cCNEwuoWChjgWF69m9F3MxGYgrtTgqvkGhsVxCI8jTVK01uYp
WeyaD0z205oeFJbdwkiiqcfNe1W8aMxxYz5XDTtcY1JodZfv8ajRKpVZMFeAOZgIKYqM5yHV6SYm
7w8nFGILmBwvOrKO8YHHHPo0DMQrdZuOFsqeqyIZLaqwdDs5U3R0Hk9ryz39/e1bVHgcR3No9MaS
iSBrx4djIoowrwl4k5iF1c1PhwxvBJTrbD8L6Z12fops/3zZMkrPOocXqJHjHcOb3EBypPlHSjgE
3Ia1kXU1bldxtj9t8t7UEz7cHTeN5ZHNYjKoYKOzcvKnn5ST2e4nKt/CA5BhEcIktjObuNFEiVUp
9FXaP+5ZDB8B46QgwxE6q4o0dxUZ3stP1s+Oaqgt+eHDOqqcyVrYc4Jp65pwo6CE8pddf+LCPaBB
tYQDozoIDJJi0P+JL3VnubTe2esqW3c3D7pfL4IeaevuuC/52BKMH0AOY/8fvwMwq+4PyYr0ja5O
GVLrMOLEQZNygKuJbK0frnPKqU0SAmU4Fqf+Ils5KNZ/YV6Z+6ZVpXW5awmu+REsLnDAdhAyVnuF
281gXC/anVGmHCWboiqyi3LxXStS0C8R9qRbKhdfJq3pcWNIXeXvvIQmSqghgRcpJ66bH2dHucsw
DKwRWiA0PKMJ4S5bgc4C4P5M7dqg+CGfW5yzdyq5wg7Q7Zm/7QbINVA+SKlU8LgtoqA2MvLqBPu4
4e6fD5aBPLi72Vgb82QjJQrwwEu6bzVmfVOsZDRGX5/LB0PLv3nHMCCkY43Z/NKJE5xosvIipCEc
/qR+vlWUK3MP1E/0VQ12YXdsZH6+HCFdjZIzmP3BVFZ3MLLfmDA1lOYW6TmKzJQIRzAdD5QVmLK+
bAP4KgmZJ7WLxS20cpcG3Ww5Yvz31RjNqbu7jBOqRJf42PID4J0CaDnbLyIjK+NY+tjAF6FqYqs6
xmsyEzfBZ4Hcolt1BCBvoZrdk/U3P4bcKlORTmrCUZZj+4SmuuSJl8RB0MCwvoVjg2Ui01KYxJ9w
YzPvOxpMautwBJTuzX7Xb1qPJdfrvnxDtbgG2bAGFtQ9QdDHyaExmLI4QYGSe8IX13PvEYf/dacC
uSpQd1XMRjXHz4jvbnUQ39PUAgx4jct4GRY3YkQ/gopfyS4lloPXXcDdUvRn//pg8ROu+BJXO02c
oGo5JjM4uHjHcNnE85K5xvxY4tfsRyYSAHUpp/YJ6krXtn1D1jAba4c6HI4oEV+rrVLan+pUhW6C
h2nIzhb1Vh04bj/Ha2hDrZl8dl5nf1XL15JWpG8F7B0sdw7ESRiLCztQQDiNXzVTKFsGK77AlE+d
vGwuXpEAfbfp/HoIACjxkQ7fEklLaCLkD51RxVkiYKQUIiL/wLAl8Aj0WnoElReZzoBOjbLcOlJL
LQnjXqTfe+N+7Encb6G4SE0env+LkKQr5c85tj1PTTzH7xPtV3+krcwbrNTY8Q1RopfFRrM71LDo
8IkrbKJ+vUAgb/zYI8DSc5HToDKFWuJA9IJvHybMldQJzNIXsH/2pKzxO+LByw66LNQvfWZpTSbl
o8ctO2/02Gx0wUfp00gkZ2c6pAWgMBUqXfSVZodTmyvNbCGruM4szNu00XDBYPmtTUQpTUBX7+XW
hOMUuDz1DsY1gwSDFD3f0+uOg2mCTYTOZiuJRbmRyLJvrVMah7Gvy/Vd9CBVNrDnMJ77Z1jR+vSC
mFZVm4HTFIcKab5eNCB55UN6pcFLsXEnxtwsrflXH1GAEG6G/xGHzwAwSr+dEZp/yur8whGCSaxr
tezEQjodI94swZMKGcbl1MuyotaF9UkjOx1ewCKOLtNOgkntxPpw6/NcjuICu5dNHvog5RxhTfLi
OEzPkRZ78StjloiPh+7ChJA5Alv0mSa4P1gORHt1CCJdufwOAnw7GgvzF43La/TMjePjFlA0s5w/
lgwrsntICaE+BewYtD91XNEIb4e92tIRj8Y1EZem3cvSfpZTN68BEt0uzGSHuqqLGUS4EClf2owu
NXBo/vlwSEA0ZB9EHrCIcSgMKs9Q6Tt7MdBJl2CasZTbxpKJJNY9Zs4gSnwGjD+3qIIhDHQBpZDY
ZKCv73fJSPiSgh8G9ZHc21SHGqscQnoQucdjLgXcPNug6Q7SfTQBAITNqaSDAQjH1tNfY07hyC62
0Ej5vBg6QerWgxHa+fU7+90BtaPc3OOwpAID4BV4FlwmtSruqE0xBYMMRe688DGR6eGxw4OF1Zkt
4CnPHJk4pjF2uoxufyARO/19c3q0NP2QuHxmLXK7xexJJQfAJGxpMDRNFTaq013ftMXWaKZNg9zg
gTuo2XoYyKo9D5YX4ZbTrELHKHy4wT5PSYaFhBZHno3vi3bjO/EFwlOnpNyEHNatKKWwepXWZZAk
Ay8CLEdYuGhYKhq4kWL20VBQZU/i079PNq32rqZ9i1TmgfHYHuyQjolCuTrVuZMs8uou2mT3Mmkt
85v0uskjA02vPSIpnSWyQBmn+cK5HUp8y/C2j+tkSu2pU3rlbluCbMy5v8/mXinqVD0jnNP7KqQK
jf8X9Hj0CX80Duc226TBBzNW00KGzckuvKQ70suUCkwRA4AL1z2etAAt00Fb/RSbhw/lJtxBwSvq
SiZpB5VYGjdlzrB6pBc4QPM9OAQsoF2qfJYVinUdAodRb755jqiEgDrOlTd29dYaLfPcz1sLuyeM
D+hop3e6NGADSaMYzWFut1IsPOXBSIhqIudFT7Y70CU8Djflt6B3nrx8+FeIoGH/XR52htI/N+qZ
pu1HThETFhVgh/dEaZW/ZrvjWQ1NVlVaXLyGgbT7ZrE2UiUBVH1Y3514tPN/TreRglMsLutvU/Al
uNZa2MeLAK60bWv/gLw7lol5A12o2l8vDChbJRfO6Rv8BOj5vbaiCKoEDiZavc7GDJJFHEhq0nH5
U5eYUKnsEPEo6UuVlizdsq3p2/LHeG+uJRVFsxZfUhNNwYctKW+NPJqlS72OFwIcGXLzu/jsxmId
rVCdTpKplfIumiod1U7oTnNI/lOoMB05kDEvo/X0WAD30Jyt1JIjJgjhvDZXI58Rr2jyJqGsnc3k
mWXN+TRWB1ydnxrVPAJxAgSVtDv20n/Qj2Y4g2WLC2z8wEvNha1PbvoFCoHfu8EFgLl8ue0xSNWo
A1PoSrNO/oPqoyjj6/poxMgNJgS8EvSarbIUC3Y6aLO98Buic7Lj4LXL85PqgrbWMk5yjbBscl9w
mOp6XdFOC+WX9DVaAvslBqXGwCk4UNjECMjC5tmikeJUcXMKjeWlJl8Ai97rCmdXSfdO2OSf9i/E
88IId+4Xz40hAoHHNegZwm9nli9XUutNQYmhp7xCK/D46VDZi3+KktQxkTUJanuYrf3hsfYFQqoi
b5/dmTykcas48igOdhPJ8laRPUxGJ+owJwx/5px8nAKUItTPTop6sHyGn1bMX2O4HRQ2ibBeLQQk
1++LNSGSSLY41Jh88A12GdGDoxHZa7ItMCzTdZXYL1+PaZegrXa3Shi5ybhXxXs5XpWi1vhu7BsN
EWUbfCKDmNPCplT3Y293XHZEDFomXs1QMzoqkZeOyg5JXR11Zh+8N2xl876FsGtsncOI5zv6VFuB
UyPxWkfX+GTa9pJJ6RyQpQumSoLM7lYDwaqnijbVem96T+qNwE90WnppWotBqDtWgcZ4JmYu6ms8
sMcNAfRvmyhOepZ2UmEJDuEpZMurJ6IoVIv0iBoUb91f9BbkU+hr4hmIGBO/9wD2PuPz5fvRGocw
MFRPahjzAQUm6u7+HBpgDo3xLmPWDGTzMXlylWek+q0vW+Ioqi3Pq0/44jatynsuCi3kmO2X6a62
pcY+rJLhYWlS3ki6CDYZqqrVcIJM5Ve81kimjNuuBqo5PV57N/h60saz3J2IR3Im6kWiH8cpDwcq
DW8pOoqVf9QE7HUibC8ZEoOpR2ZqxycdtvJ2nTB6g5Gkgt4thpNaIM+CYey9FptQ9tuhPPKDU3wK
OhIBnwc7J5BZxvoiwYBLSipyCGFbwRsbviFS8XdeQUp+vh7u/25Z7LU6mbpm5M/7EL9UdDMEygfT
ar/z8QsUbr63l08oZRx9FWAQFQ/EHMmrhX8k+8Q2LOpY7/pbnVWgK7f6JaCR72o7eREHRKFKoCD5
3ONai9zTugftTLv9l7MAAljeWcEgK6F0N/Efh8MnY5RhavJW2LhsUqXsbZNZqk2hV0M5QCkWTTPE
wMoROoTPIH0nGyuSjban+H/u59KWc8ApfVmtOBwhJPvNh+Cam6DSCLOFh780DuEMVUnIlsMDPR5u
nFi9ZYPaIeiIV9/sPq/ZMiUaXHZlrkppq2zSMf3WpuqLVv+6D+LfEvpzsaK0HePaNxo33nXTgCKc
Q8FuHlXncQ6EX1/Mfpt/TdjmS8SxSi5m5DKhvUzbbXihRPYBcViImi0XnLVVtfTokI+v1yU1SdZq
hd/z3sU/8tfG6R3S3W+uHnYCBnIFxvHZ+VKXQdrGJTrndMV8/YDbZN3NtEPjvOPnX5AcN/zK42Zz
PyFJGH/bPuMWT/tDE8fnv5xEPqKb21yuhFZoDrrnQ9K6RWHBHEOeHY0sRJKcqYtmqQ5gFAJqaAcU
ye8KBshaWcRhsxPxVnxQvAKzlo8PfuqqlFOmIzWBT5xmXaH8hvCVg7A7T/Cw9tIM4/DwaSmk0YkY
hkh9NGe/RmbffiFgwTy2cW5T80B46a6gX62ew3nVH5Sdp2hoB+oER7gO03gWwC+97d+urfHN1nds
sWp/6BViMKJfgIpkV9mEYHA/Y2N8yg9x9090I1oBCXEyD5Ny7j4hoD+HjM0kBLLdQRrwGYD6A01u
5YXZj972eeMm8d1zOW9Xkl8xsEa5rX3sv7mCSliMHkzWoBSRa5mkS885LJABtDKI+q46tIO1VLoU
ksryiMVc6UPzn9J8OPXhLhPOieG7sTp0o7K3uW77lcQUGsKtMCQhjQqApXE0sB/KrM0p0SxendTW
eLcx66bCwKSowRyZgeRhpgDn71qW4Gc9bxBWkKQTOG352EckcQrUlpMsL93OG52TfwHAvoQgpxN8
WAtApxVmyBZkeR7A+YZacCY1AcJtSo2uFlmMyDHj7i/BQ73rCe5LBZuvR8RRK313KHkJvTyc73Cv
mN/uWiDXZ3QyPnfluGFyFLjgEJ/9d+rp532W/BTB2vO8jD5p/7WItJdQPL4vHfNSD5SXhYAfQgzE
Ri9WiCnHl4JVmGRkbwwf/ub0iDnb5qFZd6IYSMFDfPgoHfyb0IDL/c3fI69AzaKXAtuDnbAfh5px
seb4MJfeU1OoQfnAbyleu1P+MbClbdL2hJlM1MP8IGKAXpb0WD8MbT5jiQtjc4h9RoEUWuZXcKcJ
mHa+hSplY9+TOiAULV7FPHHIkg2jPzCTS+/KhotFPl/nmMM7aQyIrnrY6NBSRS4P9iHo0OIAYITq
o4BcHoOZnexpsISd5E1eRw+n+hekxSvIZ39BrznyaoxgLQg3UbtB+8DqfLhxFPO0RzfrGYVBEUqE
/zw1tkSjTJSZsiVoVC+Bm2dbrUVQo+CFtI8VCHX8uncsfQgpNCInXLeg779gOQDqSWiE9LhFelu5
Vn1WwK9rS7Xxo9cwH/BgvF18UjTeCfxMo9dRforvfQHW3f2qaVhFyJ/IxmCR5n+AX9+J8GvLd1Cu
6gF+t3LY3KCAlKq1ryEPlejFaoNgtJMv4E8DUwbg8+psduo0Nn5w2tDerUM7VdlX2h9E/6JF1ntf
x6bz+QJVwq6HpasIMo3xT/sKTuipEl94TQ8a3uuhBHHJ3Clb6JqkaHb3JOJl3FF/+/UDAczkTbLS
TVZasUrdJWLP+zE1nbdO+ftZySWnj/g860bYJQeIxeZX+Hjrv+qdrG8SjFRP8m3U7ZUhTumcPJk5
DOR34i6UtNSSl+24+8Y7VPk58MWZxaRgcn3MmfqlvsmTwpen8KAm8faawNB4Voup4j7AlBD/z+TS
PC7qgBZ+70MJUDd1GdGNoi4/5c+b8BL4JYuTkzNPQb0mAUa+g5cKFvQamKwSbkI2PYDpmEQ030aM
lf1knxiuxQD3w6o8Brc2mfHO6EQRBA9xs5JMh2VUfj1Dq/FWlrLCQ65azKf0xc2PY+FeurzZNOkQ
Vwg1OtrdPD50dnLshDNULDAfbVo3jVJl5mVDHKvJ8nVbymTJeKXngppe5GqEQLqzZWyY8xD7C+D5
vBgaJpTtyBfIjkwOgchjOQ5nQQ2SBoIRrowz6cLS7vdxUBkba0XfCim7fhQ6WSpbzSnTpoDC10J4
WfwE5tbawnI2YA/TCJ68xQ9k6DeogQyZcm637sSOVdVe0iVf/Feblg5/Z1LDmTIjzUb191sfXJ18
U3m7YXzj0lzdEztyqIH4INerunjIiBYV2mI19al70Ai5nLJAipUdIfnQ0k5PyITcgS0plju3leoD
CBXdiy39Y23LUMoacVXahoY/D5mCrWL/ihIwZecN1adR05NIld18ehHmJJExE6d3JGVLQZzCR31s
mv+jSYs2HFM06cz5uv4dIX74Q2p6SC7nGfghKGypAdk00oZar9o29TwbM4xdqPMNUnuiQFJcVF8t
9m0vypZwCFrwO4PxPl4bfYRQiaeiiSkFn4smX3R50609IfCWY5xdkfIG3mOEHzXSAAFBVn2lClMb
8gpo2Z8Mlfvko68PDASeFGOhU1Qb6phHt8SXB8Ye2OccwYIr1Pas8EameIsI29kFsQ9sHtbkoFA1
PZL8cChxJw7djcSJQgUkGUnK9n+oL3cW01/SlGm4Zilb9cpJbdOtLZqfc7iDqUMnaNP1D52SthiY
a8+mO3ICDPdRgYJY2paGaj0nhD7GARZBDAeNhDUpAF8NCSZF9mxOBag6+iD5VTaFaJ5tz/79V+XG
c1LVDCzVuHJMkxFkDvAU6EFZyFeWqeDZvuRks5467XRWQs5Av+lhHXznQECLfjrrvLmoICbj2jzC
sTiivz9rf4mSfpdbJl0BakeIOYFrDppoqxsy81emXesZM5vBmFkxLumEfv2w6cVd11ISio5Jr56E
jY9gqUqVHVKe4d3s13YcTkKEonQz2rJlhzVka/e5ccFn9RY1mN5kJDWK9V5SyuI27dnr5T+FMoWe
rSkBMKoM0H/+v9M8RQYe4AtFFj92zshNlY5axravN1nJVZZaDMPZ65VkziITJ9bzGWTBbxIGvBcE
wWwLsFkhUZ7EU41LVD/DBK5VIIbrp8u4BeWe8ARl9CoN1zZuQdePVBB3bL4dIkOKmED2zW61rIdv
kFuW6Y1Ajt3/NaTQ5PFBd679wD0BlzUOsibE9HiPdzHRt+18t/dWtQwcM78z18WELcfRnDfQeM+T
Kt4pQ49o8rxdoNKZL9rYbD+s+Q8gKagpb1JKBvCxApk6VEdp9T/wSjFiJkJrV38e8qS/LA87+Eii
nKPMgzkuuYoKj0nfXFwWmWHj5id/i9FaCURgOX1t2qoeTpW0nEM+MhLvBH1gi1PGq20RLR76BNx5
iIYcGvVNHIEkLebP8oBlD3Mbr+M4fa4/39/k3PnVVycVdEACcSwTKhJ7+qprstlZbwE2FS2hYBIx
uNDJYlJoKfyWChfYNnvPVb2jy7vF0TADcBVAyMxMLcQidnI/+yslkRv4hEbv8RKM9iAVNMd2EdwL
dtJbXo7M7biVBiQKXvzTq9CnqQRfHW1StP02uMAlHgyST0cHkPtIF0VfRcBCO4s//+BQxiVm6ZDL
rEanxYYI12kPfS6N0obmXz7m97N+bINB88btK4HRiEfGEef53Wmla8JpZrZqKkaVEGvGe7D4I+yv
mKxOKePizzJYLDAHpU+HWtM+rjgkNyr4vT4VaSN15lGJ+ZU7dMI2ftustL9V8ItVcoqxeLq7KzDB
OMLtRGtJh4f/d/pCil/7QME6BXTpK1X8WEbzdwZBT7PdLEe0V6hlY/UbcBK3f/5clgSvygUN+E0U
kVaGQuXiieaPWafvldtSHxIahL47cJDqozOaHxeyeHDHvqgdirUHHXsZ3z7PlwThqGl1qdCEkIJd
2XAtfd8sLFWHMT1bTEHFxSFOCitmvvHXniQZikrJmmSs5EJLZgEVipR1t1KMwglLdA9YdkY6mvp8
faq9pK/WL6x1mffIs/1RNIR6kHRwxDqvwICyJdvFJ57Gt1Sdnf1qKkiueFHLGhZMgJCc7UYsfLsH
dOdn6FyxlA1RzMXNt/Rt94n11yg9Jnccc7iP01pLvXb4BQxmwQ5tksYMhZzkd7ujZl/2vOOn6cel
0nSyfpCPFps7bUiC5wlYwW88/GwEpZ2t1QdJddQKWXs3gSHJl5RE+NoHoOAKabXHczhu0RTQolMP
7lgwqZoJZKLRFHwEnGQlh3VEp5YBVa9Nhd5HWFxd9OmrwEBUD5qEsrt8KkW4xqMh9k9N753l4VyW
bS2QRqBvwdWcIQmFeeZBs1mhIh3AloG4XyB0kHtw79FK0zLCmtoCrfEuSGMRhX5AGlYHkKVGPCOI
x7bN/3k4nRzgfAVWfCyPScHjN8x8qQCvBUwrc9zZKyB68uJSe4xRSDQZhtgmFj1uAKIkaPVf2/2a
SWA3ZFkXADAlDr6bb6xzCxugG9htgW+aHAS7+9vUSnvIR+kMya4yVCJarG/fxNOrAIRHmOwz374f
FV4sbFDVLV7Xj6RczCLjCGcRVqx02i0f/RFpjb/XNHJfwf7Fa4nK2exf7EmmYuPF6LVzqpvKxycr
LFO9oVviro/NS7Z9tRX0K3TTgVGhdS/9Q4ah2Zfaj9WmByS2QYrXS+5wwpSLA9hMtoJOuEGUOL0R
cuavWatIMUCkxRrloYQPjqJgLP9xcu4auPfj1xBbmFh3j43IsD8vmYAO03xcryDMAgNIzAUrA6Vx
LlfyAMNjSedZDrDSXCyM/S8tSIFqC/4zzOzLWucWD/HJphKUnrvibDdOLFLAlvn2Rd82KyFTv+zC
kyv+gPGcm/iuSvpemcQItqN2T7tr9ha1C3MTtvDXaRdRRLS4EPR2iMO4gMG+GuEy+Lg75qQKDpCO
uLn8NXJAr88gT83fYLwowI0VxumkYYilHXZnmUPa9jPAySYy4KuTjCaGfmqTKVthXcLA0lTZ4e7M
0+7RAw/GqGNtpllbR3FwqlBN/4jptw46tONnaXD5C4qPTKSffPzy2qyWU/EpiEfH+RszFkOPcpLG
vOZXDgkdPxdap0LCkwxnPjPCpbc4u+zLZtwZefWVz4Be6KbfUTYfvI7W9nkw+qgl3FKRuD5A/03d
HyMREli8jJhO9oJZuAylQ8glMdJKaaNzSI7YXkzCCny0z9VtlLnsoWvM1Wto+qP3oh7CG5Mw2UOd
faJU2ArdwxtsDdu/nDa2D56GigZjPbEOlq960wvVCGZJ+7t01GeGFlIzdktbMnWZ64mo0ts++Ku+
l4GfyW3hqg3em9MCzxBd9qof8ijSfHVReivYCpPazvU1ua4wrwLZBq1ZrTETOAD9QAy/ZvDrmYJs
EXakkCpfs5J2ki24U70JnJQsjn2EuxIcysPhzIjmv79LsFqMoqtvj8B2+mQroIAtzNq85VzVxuQp
zetUnqQtza7SWAl4R8J7SnHTcspfB3A+k0GPuuhMMkm11Y7GNA4evZL03ilnnCpWFZL6SUXwvdTF
r7RYldq61qDUNj57ciHcE42ZJ0Y9SJNcXlmPfrULTG2ql7a1eGSz8X4f51VLLBe2Z/vvZBRX1n3a
9TDXQI+B4iuQ0yfikDKFTetiA93WIYOXG1r46O4nkNiKdew2oIgHCH8MnxfRfSc6HB0ZMujRey25
CEXZK6QBCgGOWN6vrAoAOM0COJupmprhBWADY+UlAWq2R/WVALrbrSnwe50svVh3Xy9IOMPCUr/r
0iM2I1d9e6GxvUR5iAWaL89hj8vwsBkzVPG+QbpiJG3KBp7XJ9RlQiis76jejcYfEI5fGVwT+bLR
IdGex+5ZD1sACxh5Ui700kM3+ljuD2K30MsKbq1lM/kYk5Ftsa0wAUuccQhM/EOnPaKjn/nno73h
SsoscmOCRwDPh4z5v2NSHS7TekFGTiISb+t52EKI57zC77Cl8NspniokLTHgadSHgiFW8kyIVTCV
+0BKaB9b2S87VrcxpuFpRAfSCisJa0yLRE1zvL/UaM4JpKjiiYlwy/7mRKo6GzRd9nsJmix09LdL
DEZodDi1SUXFwIzlqX6MXAvZZtYL1+Hpm35FMqCIVEOWab+t28CEftgO9YTDaTDDF3oFzHgpMeg1
ZfOkHlBLxRjB0eCdAXArLnzmLt/4UqKCrTBrOy6emkANTLwKgYROb6w0tVRIlRJ7MublZ3nUQIlA
7OGD19SEk3aKrsMTJcFZ1PpOjV9HtLBu/JjGe+vhcc5zm/4VFPJV1FuADrVSZY9z6SjPmU/Z+BG9
pYAZAANdtHquwjty+ao4CHqgMDJD5ac/NwC2+CaSfaxwtEbGWj0A+NlzChzPfidzAgQv7z3Zrj/t
hZyGyE//tlAkOj7eV5hAeAPB/6xIB7ZdwsOIrn7QNo2mqHln5RSUQZDcW+3wnwAesGl/jHvBFOKZ
txpqO1vdZxLiGwoAGp2qmhdb0+9POaC6T4osIkCQjAC6B/UaRvy6+Qr1/4f50mGqzVOU2vl6nJU7
wclDyJ1PWO6+J8Dzo4BVbDR0wkHa7D5jBOOuWuY86D3gcjXC3mHoaDNhQg1Qfj9hI+z1uw1sjQ+x
tiBQIDsCcsFLxYjnqNWqKQPUIej4haUIYPyIUAyJ8KfBGUOzl89kq8G3my3IIX5HRccbWQQXGcWO
CxOqFzE0VAQrTG4HwU9KXfsYrl6182txG2vDNOJHsGwvNgSXrHN14A6QdLFgDheZg+PJ1QrcctEo
dV84MvVdyBGSLn4zQsRBp+Dd3z5dH21KxZbhz5Hl9XStThWaJ9iu6AQpg9flP/OsZd75BzaKJ4iM
4qH6NLflwX1wzL3WOafE7wO4pUdTE3T3epqinP9P+7T8gcnhVcoID+jl+Oc8N4KuvwHSvi9jIkSy
NcuVkOtJ4eElTdBu6OKhqoBtaDQyC7nc8iDsDl7puhAypUPKZq0ewFVu5EA70wWbxqilMoWscdvB
wdngdtRswJdQhEba3bgDGVL4G+DD797vYK2VFJ5u2Ash1vWOdj5M14vw19xyrrJdmhjse6SmyCn/
IpVLF4qGuoLbCsiDTliRHguJXuzWT2gmV5wZTMNyCqvzntWlzxIoRuhstyNVfgO/4Ao7SdC/sx+R
d53SHuuGCAgEMKn3po9j8pEptaRvIS136a5YGt113lqv9v+zaBU47He9y+QDPFYa62Hzxq0mZoRY
gMiwsTaHPI2xQYNkhX8O2HsOYYW56y9nDo779o+VpToPQWipn6B3BKctXr+8ogM3VxpvhDRTFAW6
i6Sl7kWWdDoaTHRGwpj1KgVRg+Xh7VZuXT91ruc6SKvwAPtqRMUKMRVuezgdStQHHQHw2HYivQb9
ILioCawTannVcrpHrj19RD3M4TxPtfXhASWh1POWPa8JBCPTq+PTCqv8npDWffwtOaqjMqcuT4u8
4pxKKd0VGEgQm74yF9kmTr8Tn4MbnBrmlVoVUwCrNLt6iUsppYg/amt3SL4GeYflXUjUbfZpYOYi
yti7PVv4235eKG7zzmHReMXYrlpf1dxuhA64dgRSzKCl346DYMW4v2MzMUvy402W0sS4qbMxYZcy
ZXyDTezi+a8Fi9pGz73tFAqfZPGiQnagGw7LmYU0Zp4Zz9/L41qFMi1ToRit1kkXpNLD0b2Jgfwm
5s5GD9jb0P6ranwJnYJMXl2r6SEAwz6Dxxjb+JJ9SBH/tmaUWFbSLKQo2dA/Tq33vTDrFumnaFM/
PYV0kH6QvIxfL49lUjza2SckVPARqj8G8LJ09cMBpyUdVNqOQb2VasbcnvNSbHMwKHVDvFZflmtX
II2yEwIZ+3XRrt8wua6bVvePcR136j6w0YvWCI+Ve17MmKz8TYHHdxubU+/tZr9PatCYwrReEhB0
6aYjchC3HzvELrMWT9Uhbiy6CFB0xjeJZtmm4hHbIg/lwG6OXiAWtxKXP6lw1un+DanrIBM6lOU8
l8V5CbclVBYYS5mYRoQfoWJLQj617ho5FvcGmRmdpIgE/u5seY4t3D7amMCRmPT12PTUmwKoDB7v
pxYN856YKEoMHHuDi4C+1L2yaAwKjp6pjGXxzipw3GIssiVOsrMzs6LGw7IAK/GCgs6YJUKdIJ0M
YvqoMjuqKegayGWJHyp/kcIUKPw8/TL2eAZgSXbV13g1uy5bFRUHPpsNdtMYrOnjcA/jin06w50G
EaT/a9hGQ0O5al6lrOkRZkaeYozqQdyZMK5JR8qbAW2JYGW8JwJbQbnf282+T4BztSwuxgVeXWrr
NfFM5CpxKpJleXJ7+sdCiZFSUar/ApFXWHvMHjhwEuqvKCAWJYLS3ukNAm64WqDG3R70mvKxIOjz
RLFxqvXufsuAhJ+H1z/nXXIEZxxkBXDISD7WrndXBrGUWs54bpo7jbYNeuYoPkhQdBkAUo7Vtgo3
n/joCeni9QVQDcSX9yYDzWCWv5bJ4tQ53otJhdQm2YMUDMcwIgpr1zsvJbRzf5pJ1ghYqKQ0T/GI
Snawf78nsV8+N3AxVbILwyw4WZE3vqG7NSr4DEWPhNil/vw9d9aVQav6/tLZnj35+u5WO+zeitXx
t3m+8D4uUT2MqkhL2ikzNkUU+nyglvchPHOoyRHsGY600GU4lSWNFUDqBXOZ1K0DaDOvFkw2VkAk
N3K6WarHEVhgZRMg/+P6gtzt0jVtY4yI0EwK6anjlOpvrReKo2gipuG6g3826ZnSvcAbOmJAoZHx
KXxDnocrcxoGP/qQEITUYPVc93e6Lz5Jg+saBXEqhc9Th8376lynJWh+VDU74w6+FFfgApeTGc64
Xekwl+znJcsq/q3WSElczzjhsZjFKioRR+1BAVsBw/ydaKvbDdefCL8wCm49f7pQ11q8ck7AsOSj
5Jvo5D/c0uiUHRMOEJ1h31Zv+NhMhXMz8dZgX1uWmXdVTxDD6URUEs2D17yIW/t3nxMxTiNZtlI6
beNIvCOXUh2/UySRNi3KDzV3pMfAm3gDZ2ebatnimV32WaaeDqXJKbg4FOC/Rgo7PWaL5sZri09c
QZTctwyQcYsSWuok11bGvJ46XRGog0WlfJ2PtSe+sN+CTSYoyzhOuHeeq91b01QUb75ojuFVC9fY
mjxjIVP9K4qMFuImrjNW1CRTpkUUQd3htlo3FE6X6L0x4ELLaktoKyEWG9VFzLgKGymHEdnoB7Sv
ewS1K9WFAn8sGrRffbMV/NtSsLCUxtqfTmQVI17k0cLPg90Ou7Cw0uGo9YdC59Dtut9KpoPaqyrK
L6KvCWtCYbW1C78kxQX1rdI22vSlB9oPLIuk4DB8Y0SUcmOj9M9FGg9BCZvcjPQv3GMmBGj3OAFO
tdx5Z6r/YhMj62tovbPE0NC/Dx8nC2OM9nKfUdsOKM/Wlx/qUAjwmNxrVSln3ig7q3Pfl3kFDExW
3P/qok2opozlLI/7W1tIt2CzLFkHjJDscUVRwPEz3UTILpeoKTWV/Wjf6jWilV7vT+vQQNnZAUJq
eWmG3fM2+siqFkYMHt7u7wLCCbotrh/P51gNZTlXbgxVAiLCmLaJ6fUaiPd+bXGJdsv70QjpiMpr
l0bBV9qC2izZUlj0xTGDJcW7pY/3aSIs5y7z3oNEWnYobw2wetn2QUzLep4bC8lFJSlQ2ypZfdy1
nsJvi3++soL7RovCxUl3ibAdFxs30aEHB1qtuENbAOqiH82oQvCbmwVZbanRSC6Rdn8VR9QxfLKn
2F8WAbwGWJJQ7E86lKA2gvEho0WlPKiRaSWc2U1ID7w5FaVtL7vH2jstdh+tFIpqqspbxN4PUwI9
IRmKqm6jQ7C4MWUEqKs3FVwxSQzw6ua4jEibEBudK8B3COsZV5kVCQdEcomYqoPMEGX+L6VSQOM/
5TS3mU7Uf7IcitCTNRoCoWfAVl2Rg0PCfZ84sQroaYs2/19OfYmYgRO2apMzZke8H0hAmbKCVgOi
n0tZT1/0Iy5otK40Jj7PzSRhuSCokStNgHE7UrPqL+twDBxLHthyjb6i5nfKGdh0Hdf8zGmyf84B
RhuE1OMBH55XVxpieHfnNk9+m3BnXa1mDdjC0eWgtbK0L5hdM9uMdk5lvsYGO+obCmkbBeBGZGND
UA7Fhu6OvIfWBkugsvcC0rezwxMuEt5W14fZl4uqhwP+qEDqdJ3cFVURpsmwFF8GU3EcHIVivepX
WWyvqgBDe9udFhQfrq9TiliGibI2vskGU1ypmCuROwKzDiJtZypTnzcI6F50ZigLj/gYK0pR3Nu4
Dp/PEPpg9mCDSug6QD/Xs7Cgkr8gqH/GGhkM57AicScjfVAumU/5OVWNI5RqILzR94RqbetJY+F0
+7EzTXOq+/aXLpTH7GJqPx3+Wb9qKRlqmkv6ju5eqZmkDba/xnxn0darD5+mpVnuGElHuCrt0+NN
dD1iA84tnViFidG1RBBLDe24qx3rpTU5wSsNVLnUVTuG7Uffp8dBo4JaPKjgKf6WrbG7NgMGr2Tq
PpkbRzmYW9qtQThoGBbOm+s3NfyXQm7dcyuJZgC1RBYP0JH1ibZtzurYKSxSVTETOBjRzDkcOrn4
qWUYNoXdCF7kgmLIIp5kk9i3IQvBvv4QVR2m7i7UvDRTAsU0gPDoBlG96RMCiV2XXCgwt8zQqpCq
8Dqk3VomlWpwwj5CF9mdZdk9VWI5zJhFeZWc7mPq+wVTsv6U7snnXoHqsPuB0lgFUNxYAuF8tZaU
sTd4uWftubmtZH8K6ou+BFrubWAiqLPmg9HEvd1fWnxtI6BR6KlgIfnN3Hm8HxXhtw16rQ6gMabL
O36g+ujVYlxJ+1yNSXMoI+wc8IAuXEgSSXaTVbourffdxuO7Kl2lybiQiOXSZkoQgmHCNWnIqyc5
pVe2CnlPla5a//7/reRTRgmUD/PqalyPJp4yNxqTvBgoAI4QOV6yFWBBK58hT3hUnG6CYMKpSds9
uRlV+9zBiJzcOEtmmuYy31HM2YWguCgSGYzA1oFXK6cp5cq1X3kwJo3d0PnMDt2ObAgI8MAsOOZK
mqO1HE0GLGwR73lZO1V8giqUH4SRnsI3dlnqcANcd5UScuHx9uUyKrP8kI2ii9MXpPdhI71r8z2S
x0aKiDoX/Eq6sAE3ZNn9orF9AWgZbUKkKom8qElv1t9ESMkq8OxAj5N8mZTG6n9PjlbgvhsiYRQ7
xUoDEHJaUgd1ZQQ2EHfmFpE0eeHMszh9EE4yUap5xgiPkpuGuG4bbN2GaXxgI0rn7KUfRsMOvqJy
vCjiMfuLdTGEc1Wdn7g6C0UPgXcfFjFGwfD760iijqwA8ndh5RlXfI5rIvoCTQExU3x3Z377onsN
FV5NohTEbJPzZemaUoUAHflTpJex/MKaW6DqdezhNOhvSNAp9sdA3YyGjM6LH75RG7zuJoBEMUMh
2W88qnIQYkScQYcgW+CEv46kM9bWT8Rd6x6zFDXkBlktmGoBp/sex59s+eAhVDqPUN1qteDeTs6n
pSHXk9vBf2GsfcD2tE7Dtuq8fYuxZzMk/fUeBGWmMcqWv8JpFBqbGtzVTZngD/pO1HgMQY2J2SjC
Qwy+FbLc325gofdRjlHo3ekNmFGUMeI/BgeUc3KmaENbp8iLAwKlTmjRWZv1VAjYJNS/o/SqOaC3
fVQUjPvqr44VPT4Wig3rOdIYvFgZa1hcpHvCWEAgjeocUYOGm3VavhNXUiL3yWXxd8yvgwzs2ywJ
g6fcWyCi4kd0+Vasu8Vk6BtfxuMmYzSPcgIpE6IfKoqFzWQVF9H0Sreo8U/TFSSU5ZjCkPWlBmRf
jKCqx9I+FyjClYX5MnmH3JZHKemhLw8G3vDRchJOP96KmjC5GhnOUVUCC3TSCVhzjel+7zUJw9LU
TeqbNUJnjoOl53pYxmAufqrwTcN1jYscC/W80OalyEOY0AWukcUqvhZ3bZrrLAWYb28q8CheU6cE
BCmtoxwONGp46oj2EzZpldG+3o/SoiESnY8uk4VrOClMMAJK9tzZ//fpvGzkDciUMD1gOmA5OxSs
YxfbuP46IOHzFfOL/YqZHT7KySjd99qGXJwuHZ58j43wdlXF2QKuanOa8s9/EeUMZadZQhCs/SqH
En+JzvuoCagW++WQNvWbFN9Kc45AGoa7BeX9yZL9xVj3wXWfFZTsLWRto1qksXAabSY81Ao/wfPl
+5c00IEzeMpb2kMOuXJ114JlNYnq4zLSfnBPxQABrgdPUm+8He3uWtnF++jsK94deNZzOlQ73m9l
eV5qaVN7X5C6Z/5jbKc8apvAKlQU8C9e0FlP3WFm6oxgQT5cYjYdINRA5pkUCe5XUlumxNleiIxC
s9xA5IGyqeSHmXoTxU41TwTVKMSDjNU7AgJi+V7D1/ypecfkvM/XbsAyATMIpVJu9+sjxtWtnzFy
yCUJt4fMC/Z9SbgQatnM/PvRbQPsCxvM0cVcKEiiPoN901/HqFT+eGhzU4T44XBu9O9102cfSijN
aM5gleTx2qpXHmpyUilwowr4Yf5W/YEodjy5Jsg6pviMPC6dsdU3msQHtpbFnZzlnJqFzC9yKwaK
qBDoGo3M54H98FNn0Ve5SQg1vZqnf4bCiABaFeH9+xkHnUFrVm9aGdN3Z/NBzqH9Mcj11CQ8hC+b
R/B4Wng59+Ug2GqdO8WTPCbNHAtVnTO+0sHX9oN/y9NFVg4CnaN99Y0tycKIVFIXSAIiBvNPZMca
OkffwGJuOYNprocymNl2fQ2wEuXQZgiLAnJwwgnQ9y47dqh73OnAMZfjLjQJPLXV5Zd8IsXew5wk
H0CTHnpG82OfKitW8XWuEtFK9+Yv1r7wIhrftTdR7gx4jctOg/Qp6wNfUqVVL7hjFIvkCv8ctHdW
7Q/LLeEUsjac4c582+fEl3YmTA2cplmwKN8xQlayAltH1KRwWjL3zpLUvHFAIz99KCJBDjgSTen+
6JhBySae2QELpbtXcr7jaWVqcZNUunNJ5dpl7doaEPJuKmY3y9EPvn+8mn8ujbfN9K5ZdmMGfLpk
vm7kZ82Z//EznDLd2zNxlRP7567dMVSJ/NVBHc0IUVclPreY9b/dmFXqOwFRdyVYCbyhUsElAGQD
iX2WOVvzuKmEdne6vygWryEr/y+4Lz4GHY7SrvHMfUbkFW1k/cmCP4A8EhinWHREwsg7kzQjhqkz
qZaamszrH6SGedWz/kKsdvjOL814Rwxn8DVx5GagCZi08GYEIbHOjb7UHAhsC42Cbvnqe+O4V/dn
CsxLqG9JIkT4bFeZIvNzKVod8fdZwu4VJAatM30oDbrMKF50WZk+R3ekJtU9Jk/4frPeQMat6hcz
XRbW+D3oSYlMwh9QW0TOtqBaDjO+4plCkVVwn8NlLqZQifl2MnUJ5YlY2uxs8QJwJUzrN9eEN0t0
FwSpA0alDfWXs5AvAk/RHGmFIHPNwVV0bBSP21bVm42t2ZhyDvr7r7c9XbqLq/zRc4UzEPKW/w6p
FyMiqdlaowvzp3m1imNzCjlS5ceIGdGXJc41DwYaktDF3WjNM/3uvp0mOGUtnemsnZyLQiJwl6yv
ipvgYhf8NZCD5m2YrG8OiwES5xSE1SneA2iXGq5uJAQKS4WcqgTryzMd9c4gExuaNefiTFm4oPHx
aSZVPzXRaHHqjgYbXsEYBQm9OfncuxXHuiJltQcAZMl/p3fuzO2/do0q+CXQNU7/1G7MO4UJ+5p6
/rQpfT9hpMc6vjBUliZKxa9ve3XwtSEGUK05++AjMcHszRxY2U03IU2vRFWOta+MZs8xWruYsK9j
uxEISFfH/QPSXTXvA5UqkicxmzEFedA3p9Gln09ETPw6r2S6NMCpvD+iKpsodJM8NZ+RXybQkYJL
Ec/Wd33eDbuVj4BN2IeRmaL7fhzjL5NH1utOo9GcglT9BiJ6AwszF4iYqRzcN5PZSdtHCQKeQtJS
GznhJsIWS6eob1l6muvCa/qufuX7PpveYS1fXc1dSQj/BhlqdVZBUloDH3FFMoChDRTXHRkCLZx3
jYBy6asMUGMFGFDUCL8YE9EN1zRjyLVyjo5dduoQgxdQrCakihcS4giXnrTUbLz5TokpmPNhqw3i
Q6fj7XnYlQTKWAsinExx+4fgRh+9iv3S1vQJfN1yMxwDdVhqjPOssrQ0rV2f6WupHFx6IWwEFujx
hb7RqnMuoBzgTcjX7dL7PoF2kRvGEp2ulP3LhQQLoi0cSx/YjUhYBtNGelOo3K29fCSdR6qYENt0
TsPivlpS0hFO+m7ZFJHfUn1y8EDEjRRZWP4XU/CdiOru6ZMzVdUV/xVtsSJ0QCGNVMJAHoHs/xQD
3kNI2dU3cbnwsvofyVx+haNsCKHFqdAXESNDc2E6KUtM7Rj3TbXXE+k+DK8obcezgE5YjeEJnNeR
W5pTi7oGgrXQvCXAY22ouqHcKhempFmeBPSKWKejaWkcxDZMOyV82IVuUvrm7ftY1ImIVCUt25Cm
WgP6sO12r8A9fMg0uhsPQIb5OfWMhCRzZPhjMMfBZB2AOMLs7ukOPNDKi7JzbBbPn1rRQEtZIGFF
GSQjHFVwd2rlKzF9dbypWW+X3KX12OZZNI5HoZei8ajqLdzscOZfvIyybRFwUR82apLaG3pmSAjV
VHkOpuJDm4Uje2LxkPhu5fuDO53tWkQ1hUsilI8Ayr6FPlvQnOYrvFvJyCjW/Xm/t0iFarlZ4ET8
fLai5thPiP9bMTx7cyix4Y92fPr5zpPyPCKw4+SAk4BZ3pH+kY1mngekMbKpLw3NGHm8bCJH0u4S
jejJ9drzjZdn5pgeKkqNdQqrMyirQQrTMrfZG+1t8AzD3gv9V3s/8094jxs8rtmwQi9zYeraHtUN
GotIVuGwWoYWTiMGg9iMOuMW4zAcqakPrUodknwwpOh06mA1TnFhQUgzfMZQnDciIw6Dgl5IvdOW
kpx6Gewd5iGrP25NbMnwK+9J4tR41od/Do/MzhSNeHqYwkBueJiXN9pyA4wCszhNpeMaaH6kSopI
8eqWXH3+S29lnJD0ooJU/o9BrtZwtilDUquqe9L2Tx/pYwnkEGmbJu01W5CS9HBYuMaXTSDv7Y18
mClu2xRWKzLpYFKtiyOzp5k6fezwsGIjKAnvahCYo3kUmKs3rrsXw5UiLDUXKjyech9Fr/vHRavq
yA/S24ygO61oyZ7ywvp4vbEtiEFvT3OYFawxGxJ7xqPCbmNTEuWVwR8kaQtbrIxbovkjr76/RTTu
e3DNF4IQe/K/6AK6YDQE5D7WyE1PbmyHl7qM/gxNaDboFlQ+zPeyvitpNoBifCZI4V05H7+2qNRv
eJeoqKVj+Hy8HQXMIp/uZBFVioFe1t3UX/XgOUX0IbAdb3oUtKwCkYm6AhgfB/7D0nUC6hUlF78G
9btP/JBy2NTl6G+W1Gng51HkrNnI3RYf9/QfJDlU/mcNMdgmtIGNkNEKvyJ9yOeUN/qRHLH/3cgI
Cj2pCVyKdEbUbfXvqa9HozkmUG+WBSN9w4hM3+Ss9vjQPHWlEiUOpgwjiO5puA7g3j+kN2FuHBo+
BSE8LBisM5LgBaKrr66e9eC9gtE79ukuDjFLrdZ0Fvb9N7QRzGzElGoTl8cwAw3U5Nvp0p88tEyH
iE6YrW5wyXCEqGHCnBHJf7b1RdPsMCyhgcOpypLqD2RPAM53ZY1/s3sxvN6qUzDpvk6QaEh8fcg1
Cuvirk5Jp4IdZBt4KHcL6xMvsdGwruEPfUw+GhR4m0NsTaZY4rj73UTife0E4Gcu+a5ZjASxg9VV
H7+SnCjCmJ4MTiE97Z2GbbLg3BZviihJ3CQ/33rr7umAPDG1fNQfjqLc/P4cLGOtA7c0h3a2xm1k
oPSRWeyjiLs51WA/jwCVUGa519hrMiKGwhKe/luHKkwRfQw1P1ap8TPTRLuo7enZcjyjvUUeV0H/
2Z1bJ1L1fdzGPTAyxzkotGApSQrsFynGf8KTIquv23rN/r5QpokUDzcpDtUiirtbolz8y5+I7drE
qskvPMPG+2c5OszGYifJRMEuap4mvSdijvwTIf61UdMwfL9jzjuX93VxGESaMxjoEqidWoCPsocf
fn1X33xw9KsoHUZYCmtFqXKaPXEzQbJe+owQbL7eF2D5PakGrgmo55l9sTSqxHihO1MmWGAS10hM
WKaLZUsMozl3Vy4iak08oWQjxQj7GKNKAzrhDzxGq8l+osl6v4VLaZUUUzSsqT3+L4lChfDDgZv9
HC0Iz8gJVdKKc+kH2PKL3idUGmlGQQ5bhGz5gNxeAjNuEcnyJmhOG/hUw5BNlNoBrZklmTHUElnC
jy6aGKeIZJYsaT3D2hDUBC5scaKhukyWDLJ3mvlPufn7BsT67pkiLkJnJvka3eI+7J2bJiWPYwJF
Ru9B+n7LhxFHS8XDlxIYT0jbdOWIDWTDKmewiKJ39lP9k68i0y3gm0jq/Ybx4r8vy5Mw89ezmg/r
4424lYR3Ww9Wv1KT+TgkmMhkzBuSFbYFuS0fQWxJMrXilcx5m0xXI+bVYgzbsywRdR1khdBssQcD
kWuYdYR1DcOVtx/GAqmJEaBQewFBfxiuJFA8Q14P84kFEEgsKjq0vwq9kazCZESjVXKvdktjGPDM
7l9LduufBZG5l2KbPq8E/XC6veeAbYroTb1kzsdbGvpmKPDF11Db0N0+u8SeEcLq01cMqSNw+FyO
H/QE7QOBDEBcXTtgoQTUFYjewV+9STELc5Yw5nfMlU93iw5Lp5WweQfco3jJzHFjtw3c+Tqpboy0
V9gpCoi09Va9HdYTMMcMEMp08JXMKWeFVdih8ewbAPOvL1UkjIPu4lLEFOXDt56Od8ZdAFvKwGhJ
wk8+a7JUQ3U/zl3FCsZnk3vckMIQApaGxSk4Itl3hG5n8oku2ss0PrRnGLnvJSbZhekLLKs/pydi
U9euxNyEAwCdMw72CxyG7z+N2P03OwWvhcQM0W3QkuAOloLtdVxAKJY1N4NU51uwAS1/rYu2ZW8U
KHfmTKU/g64NTbAea3CtsrYt8B49rZtvpSaUtCwU6KjqPzyVirM0c2YkpRvQNJ/GUnAsGWDWUfAK
Wzk5sdo/qeKE6mafI7wnhdmurMfV8UPYOOjL4QWdg0kHcpHMuZhxH8FVY5WWSSU55RDtQk14Jnpa
QvhUkqWEopCPAADraBHsY/AFUcubr3D7Ar0/VjGgRBz+9AOOX+w4hEUqjryaiJoh4tDjsnLpEaJU
Z/pTENv1l/KihESEXgs6DPclV3hQYM95x4MaVzodpf1Yf79kY80HyHVsErCbLcUjXK6OVU1DNfIx
kkb37qfD9xUxQ8UHiRHrOKDuhyjYdO1gfIg6njN5FNhO1hXraHLp+0gquv+QWmORIHlYlse3TRV4
ey45ot8rfkQKR0hMLA8rz3HZ6moXWASgLnl/w7lxRQn6Fo14g8as0sKey4kg56dufm0Dly1AwFAz
rv2wJ3IYQMbaQCXuwhVNzESU0UILnNtryzVPwNjltF1Cx37F9go4TZxi/My/SEKCmZgPyZrIvqPD
ciUPEGrd/20FTApPvk3oqmeYrfmiqCLn3Po9kEHn5HJf3YJo9bXwKcEGuZstUjdMyVIiNTRaxnDv
CGqG2DOajZR+SGD/6+NNLDY2xMjfCb538gubtI4ULjo7xuMiEMhiyg/xLzER7B5ny187U4FUa3i2
Uf9x86EudrhiwqpyXdZ18EmEQHdju+jR/bsxxgTA+2JY/yT3cp6F1ZubplppKMf57BQf/Oat0Abj
hfVYRHnhN1D4IlPImUi3szgdgbSWfdhTuAY2Jsrc+veC6PWxFnN4IcZe9uf1coajo30Zypf5W/+Z
zJm++beHvCdbQnzy7h/6VM0ruKMQxcZs9FWsTIB2sUF2FgHHxa+KSuix5G30L9xKTXnlHjTUjmAe
HrSCTh7kiBWZ4lzgPLD6MoMrZZ8FcIIZwJ/yNrNpS+7+OW/T+ZzzlRujM0nCNcrCZPp91oNf7J/B
hNh5jXgnIlhm6dlzyK7shkqx9dAO271lHwkiJfWFohWrfHfXK1gT9PsxxVYYDHDd+pussbm6NkcO
1XiZnWF8mrsF8qVDLhfUcBC1mhu1sbWlkwwESWuijZqBir7qculDcIYay0nD523PSzKpFs5HJJNl
77GmpGP+76VAiS10zicDPg0M84heRFYNGGGtBTgaYGjlF6oFncHw9fN3MEaCNv9sq+4K+kqzDaHp
1tYk8cZlKW3zlM9ZEC4w5hNWEutnS9javSlhUIH6yjyEmFaV4wYvDr6V0+awLQFH0gXR2OlsaeWd
+oOmt5l6+IvUcOmsqsYWjp0+pGl9UMdkO8kXgZAvlgg+cRqRxeQV6WwypRoxDRXn5QPHlHgEG2M8
OAjCLGOojLYaahhFYB7X22iqR6epnix9EVsZuJlOQMj+iU7FEJvYbt7wpBMf2AT/NOnf/ERwtEdI
2G8tEJYRsEi9MUKv9OAe+PRmpNZW5bv6Yfw8Vbhcg1SsLIsQfUz4OcxmlYKxRY44ytwtloyD/wBx
Vee5zcsmTHYNsyvfD7thf/WwqqQmQzIJCm2Mk8EPwrs5Ro/PnjwB2OtQYWrL6Quzj2fZ6UgnBnqZ
MTbTCgXEdNmuqNUD7jMvF6EB/7GALIBMR8hETsSNjncN/ox3W7Zny+IDsJ4RGVutACEzmVsZm65i
StwW663/teqg3pTcnoU2xTTtPalI+RZxH0I2EgTHxuLcWk4FaUK144PQ5me9veknLe2Cfr8ImNpH
zcMpPBsrlM1WOgiFuzGBOlfFChebfxGe3DRBhlPQ04pJtOxU40zxH+vOc+2M5RZBBuUZh9FK8vCy
uV0LSGqkWy+0hYNPTQCwwz3C9L5Gce7UY8K9FdgTSDTfFNnkZJp32sTGvWSqA9ufGmlGFaBrp1Ho
hrN4xkZ61JEKjVHoOM0/sBtUvLz8pJjlwX+J6c2ctL/t3Y5bSZsuNTahofCQguvrvjksBkQp5wEq
rBNjpAIPuF80+Ao3agRrv05siZwXeFLlKJMjWJSwq/ckxVZ1tMTv1rJHoenUASI+3bJUyMH9n2lE
d5bEYlr47s/CjqHYJ0MKfVk41T7mVVaptW0UxggAh7mwP2Sl69MSWrH5JHKe3KIdu2SjzuaUEYrg
VxhLdfQak20KEqnN2APxmMS9unNUUtvIWyEhxxAJyxdCZtNv1iDtXRueyQqW9TXd4oPdrRBpaBGr
kM+9oyNzyFTXg1cSzCTfj887JzisdUiMd0SMfHYUqf93M9B85vimrB2x+XGiYiJHy8oMg72ORsXc
5q90V6ct2RIhkDlHq7RIHxEY6MeE+ZQTOXbA1TaywpKnXkDU5VB19X3HS4v6Los4PdalYct26vfJ
uGwM5p5eVpcPaKumCofiXmkPjk4uA3Mho9HIpz/mllTS89h4daiOXldzI4C99P/clpPAEOlaj4dK
0tn8kV1FLJQM71rDqhwWSWqqIZ3QGfwxI6GjN/b7CSLXFPKsdu+AZnEIHA584gsaey7nG0/P+cvr
bKPKJKZnMc0wvWc2EIIORvRSdINb9lvM9mXHTeDZgORWbJ5LcwVYwH1HA3xyIhHXaFfR1Zl9DT2Z
p3a/yjXQSdlq8xyWM3/SiuBWM7+u5roJlJJDXHahTsE0LzRHKK9+4zqbeZbSwr0noKT45pBXX9yw
c0Fgk4ADscZO3L0yvhFpbZnJ+5him4cDNFvbLXKE/Mpe9BJ8rQAVebQVLDDqavIGkyPkQtdD5kEY
SSsT7UH6uzrAG5KEuf3jpOJT8TvwCY3xX4v7rWmfg3dvSA0dpzgPx6cGXaGd6Wrn4bdDbqnHcNTp
vynlNRIqEn/74P7DZUMgcFWR6lPeVOZcwNNZJXxq9bzbBx/QzMtn3OP4u/aUN6wcDp6aiOwmDEUn
sOkQSr3Y2FOjlcfjfKJnICiF7z7DB8VTwXMe/0cQuSnD5xn8q8owjiovF1Mv967a7pf2M86UDgKk
xMZX/qHoBbTaNJsV1ZbaLnSAjDerUMA8/eA0JvDtO1+sSpjrVvmGZTGCJE6f3zKBFnT+W2KUkNY+
QCjUaUCHE54+5tJPBx3qakeBxINpxakZH/Jd95gdK4bo4++xUEnUKQgUic5HKkLxmDvFZjpZ1B7w
/nzWmixNjctR3CD26RnkdT4NUN/DKFFtRPCRcm7IL37YIGrsnR5wW1F7zmJglTUDNJ9WL4qUfMGI
tYrP0AcOKVihQ1VdmL+chwYV1jRwCDetJK5uJB9KawJEIMsY2cjWPgsIESCApRR0FfZnB3MmYSQF
jHPgmfxZl78B7K+DtDC2+zCyT+7oH1/cLeSRecQz6OH/olDrMCNpse2flCnW0sJ52GDbyPrYRDcv
YlC6SaX4KqqiBcbycZnLaAzyL9YmWexRGP3ZPOTLZjaC8Xk76iAily44Y/FX5l5zh9D+5WLyLX6Y
GR4TW7oOxNNtUUNSCQYBm+jeGgLF5bEx9yIgtD51Ce9cRtTCeRHhcQAZDqviHcD6BpPFaXpcu5FU
uhHnuO5VXpyGP5stj/BNFJnDemgdUYGFYFEsNR5G0/JCoecrews/gDPu2WQXsFSbBdELKbLfyPYJ
agaBFuJo2HcFg01+IMMRDRhNCSVRl0tnLVlUAJTy5/LFzM/FkmLiP38qSdys+AhamRh98pao1Zge
7EhHDhtFKbClD675kthUjLajhDweitQEtWyRpmc4Zpo7HbbB/Tk+tNOMgpfRY7afZENBWuJCxDCv
7s/hM2SibgRKYOJGyHhEx3Ii0pQYHtb8UV308CyPcG9QiP/Ofy6bGtArEpUeQJfEE2Ex8ugYYSJm
w/X6KNLn5cxnwCw58elWvrYAUczdKhRAV/TNw0B8l1yzIrk52lWxXYZgheXEbOA6UChHgV834h2r
iRNYRpvEOTSh+Uk813ZnqRBCk97A1lC2HYcpCAZPvAJO7yyn1aQ35LyHx6BAd5O89u3o8JEvVmLl
puZehZ3SQY0gHhrDDs/ITaHMXGsNS3eUZOlt4Mxcsmq8bTBHP6cEbledzKJi9qnN2iBYnvtT9BZ5
EO3ta1yDp9uXhzktP5Xb3qUeuiALEyE22w2J45sRjy6ojWnobS5MRyEjIHP9fXOTpx2NrZvG4+qg
guzRtwKT+9xLFSxRkt4iz/TRR4TbmiAw1d9LAkvjL/HljkOLf9wHGet2s4TkA+ibFHSMViVv7IcF
CW/uH4gYVk48QKMddaQ7yilJdmq3xvKhx8mZOe2gtyxdzqlH11NSSm7BUhXu3CqWrdwYoWoMYiPx
hlX5i1a1r+siAqUXMxDKc+rKVqf+PevsexbW8zljJ/4o6HTFegm1RLKwO3TajGe28mH8Smh9Bu1O
Zw7BUC2ostx7sDReuk6Vs/wzAQ3tlPa8wwmSC7XqtGvInKNI/FM+GYuhxwhjgw41JC+zhEjsYDSe
+Oo8BaImxYLNAIfUE/TLC7HuaWvVxaxHG72AUcr0HC/ttAdLDzR9VDfTOkTlMeZWnB61KNGjtwiT
ZMWq9FoErZ7YpVreybF0HZXaTSOvzoNGr1TY01C2MWPRshCrlX1gWZQl8PfKtq94cQHe66XB+nw4
MkX2XyEkEE9BrQC6Mu6rAo10Tb+CMyLrpBAI55vTVylA8xQ2+VsP9plTmGkN63m82Oazw21YZyIt
244SWtbczGwHCkSno9jjjcoHn4nEN4yJbYFKh6YD0e1FQywvam09BPmGTm1XbdZ5ISBzkmM1QqAX
ce5xlGI8QpKALVzuXi2iwWyb0o9A1nHPfhRsEyLTbZGC4BlNUiRJr4yl9B0+apO822S+lRN4rEqr
u2jaw7WIdRI4pMB7LP/fIzmjCG/hdsec34pH9MJB2LssPyD2Wri1++90bKOUcve7gTRWhvWMPq8q
tZ/8D0Qr/Qz6Oi9/iR5zHA3dDZGv4w9WfXsiN+kvhgmK4qBA0Je+BI8pxuQPd9MFkuHysvyzSLxn
KtZ3cc7nuOXUYvnzQ5Srm/E8pKONmS6VkkxzQgPJmbxAReL02BTNHdJSXySqPPKOkJ82U5R0s1z1
KtuYs/iUSWz3WUrLvGhM/5ulgsXd0fFLscVxOxZe2B/vGvRsTrPryyhy960XSeJhZk9wvHgDzs1m
vV7gp8uaJcsSWQMj3cgyJXHP8h++VUwsNYnwbVdLKiXbKjJy19sC+f15RqZHdp66ydDDUgcgO+nd
saGE83eVrSbo5UM36AHap5K1wMa4BbyxoFIrrsCO+K+YusfwyoSMW29XTABTlhokOOuMbtnfbh56
kZr8+uFRHU1dzkem73tP+XtdOnsnNSmdctZdJsBcLSCwDKvF/ohlcubS859YSH84ARyGvIec54Ae
qUDwRS0DEB9iTrveTUrUyURpFYbcqiKQXmsmRpGhXwFq6K6aKoQ3gaUe9wYNe3MAOW49vH//1iLg
tLjQchNojFFjy3Wd8LhQ+silA5Nfg737NXO3fk9rXfkzBZmvlunKXS9wbDgFIlbbrG5AKcRbcU+T
SFh7j3pGVApdIG6hZGt/uMtxzd20wYPuCmWWNfQB0f+V+vLdNbdudJobn/SxqKlL4v4hAF87ZYhU
z+x2H0En9LV1rawQRIUmr8r39zsctx+MKsggTzDEoKhu38f5fhE65+7uaZ8SRvM8gsRkISx017Os
wq4+RK1tB/0rU5sqslhnk792mISQ1D0NJwaH/hUXM7hv6dkIAE4F2H1a2GYIo+JXZL4ldSyHrCou
CQSnmyC7sOBVsn18lkUbpIjSmrXdR+F87SDdeOqWOf8Il2aj/N701tBDCpLvZBC92Bt2CdKcwBhe
W1O0uRL5zpnI/OgfVNxE4CPvDy1cTcOlK1qgAEgsTwET3usw7UvL3Sp+RuTd3lmt9+t1odzWsHfn
RsYYxR8GVnFasOet4VFkpVaDc9rLiL4ajdFOqGTmcALPcLLq0cRLtlhZ1VGlWwoZa1aZs32jMj1B
HeZuZSMSSc3erRl42AAEfSL0ksDszIVehL85oDjnMxFSqw017seirQqQNNx42iNvDqUbCKk/lJiS
9fuLDs61VfcJzWBq80ewjNwS11EhY/IbbO1fSC9z918ZU9NQGTgAVeXhK5ZlS8WMvPJDzZzApgqS
mPQmWzqYaoeYjSu0k1VlUl5khJ5IEVv0j5ak0hhCmwoE0Auf1Xpm7ZYZjLF8dCPz8j7yQ+lZOLw3
ERqKjaVmXEaSPXZ7a9NRYyPPrlCjDakcQY3oc7HWMnSl9+rj5uv3A2kDwqkAVlwwq7lhsR+85OcP
xNIGhkBX9yIEtj0QUqOs5csDcG2Z1BzolwA7KUxhSIeMBOWGJ+IshglMKOOUazANJKjvnEQYvJ87
STQqLbHSPDomF4ARVl2WHuTQ9HmKhZldkGQbBN3Nk6DT7IoZD1ambogAV0mn9dv3ALb2yifHPMnI
flFdVscuWZ59QW0R8pwYmZIIweI5ouBtcyl2X2QLIYAQEmTNZDq3OPT10aArJ7RHcmBSU0trr0pf
rAKdGCRZ1EDp1iki7pWpKZDita7v3Q08vB6MSna/kCHMi6Y1S+AiZafPkPXaNauXaGwZNofUpPDs
6vCFk/LU+A2bYVhzRiduRtCfFb+E471DzV0X+CVSL6jHd5jOqs9Z2ZvXUHHj/ufA44M4sqQ9cucd
4PLcNQoHd/oRAL6/SngOYQC6KER+ffiViDGfD59u1HW1WoaooJTn/b0jRnny0qN4Nl4Z6je9LquD
nsdazbJlOO2jAM6ti5/NFv8TUKb/krH7LOmosJ7mOZuAvDXdVPMelzLbNfoDzEphCV74MW8g1X2s
+QIHe1dKa+pr8FholhEGT8DPfpeflmDo+J6zM9+KTpfElX/02GRntHqRRGBcUOAQQ/TYFBIexz1H
YeB1l1jhp4o+St7lUK9PcXHBb5KBXc5u8To+3jXs/gJZqKgJ0e3xUB4W/NKXXmABTVO4s6pUNyyK
z9r/idcOGmh8vT7Ku7JBrZm3VG0rhlVH/TkaR2Y3zRLp+vyVGmVc4mV1/tr3qur/1T0D0p4OxHC+
BcmcrLaDRlfTuyqHwdHKH9FGZpyqh/AsfUAqamk1Aki1J+qfWx/+6utk71n53OKELbHutCL4LTe5
wr0jO7kyVs3OMVeTiRIcfK2RlEq8NJxEmwGqpu3aBTxR8CS4Be4zibAMwKMH7cmc+APEiVNGrOXw
HKkMtXVZSwUlVpeGAzO+kRluj5UXCx4WqtLI74+GDelz7/4El8x/EuiVKnMVpH5/l8Cb12TGAviA
znN9XBF1CDEXXT7rKYK94xHgDHtVVAx/cfeKkpo5SUr2AUHkARaDowL7q1sQXu2aXJZYCEpwdOph
hNG0RdFD7F1f108pnap8/sKHky+NzJR1Y2G2S63ISbyWUBs/rNQAFfIYPG9nLEPWKduVzteJVwbu
3mi7GNvYlJfuqnavxw+G6r49+f9XKzd7Tbgr3fSY01GF2RjDPG0QL+sortploVIk/3g7vgI71ufm
DKWV2Zm+zKVyuE8Mu3ScPqwRvKOfiVTgHCClV7ecKDOlhOlh3wq0NApETVejoC44eCzReolXDbdn
keYsMhqGj9Wg2ocbcAnQyoCbqgNTCjH1jM9L52L2F78PLuKmNDr7rSc9LUlqwIP6KP5hXvwEKVID
m61Nt4hdltP8Ez+RF6d9tk/Lx+6i5qE5T8kiX4Yifv0sUDP8zNp8X/jYoY/zIfeqsELv3mK3Cu2r
/q3ZF0aXNiiINLLo2ptSPVGQFK0UvfC1aXww85UWlt95xTjJKQGKlVqKbhoyWSfr8JieTH4/bJ8Y
5o8FkyrYRt14KVbIcI2tT6JJeUBQ0qUODIfgMOSSkEIO9PS3zkuMDw8tT2lu2WsYudJjR1nd1rgW
93TvgM86eoQtIeSewplvb7qOlxyRof5FUcKZ0OIiDBQSBFBC3EApIhd5fcdVQut73XeqvZ7eSlF8
euv8LS0+NDkQu8uvR2ett5v1G3VfAjE4E3NdshfgxuBSMF0XljCb7lNk4x8n7IMANKF0nVDvwizk
JSVGjaOwMKTUWp82//MA/H5JTs7lIpZ30awo+fEfZNov+/bmk95TP7V/4oxTQqNV5iBVrr6LqX96
prpAOmAWdjVm5R7iy6uMuZ/qri7q/bXjDj7JGQTfTOloeg/uA1ftxTmFrmxj4+56tt9/rdmzdKhr
eGMNlLWdnjEIi76uPybYZPe0MgOcrjRsyCvEB+B5ibVZkYCN8hVyPLk6V5DupjgFr3fjjVj/yJS0
zokICw/AkZIxc+lGPY8ZKj69bSqJ4VauBGZplAZGnSmFF7nLVlDGbDAc6IuyRbvViOPS2qM6qqRT
x1OkmajJxnRor7B1GOZghSfEc7HlUFp7nGKbOkOfMfbsLhvqLbFhJm5KXhCNWIwm+yPKGzYVKYa3
6dqINxfQ+Ls0bKQGzOx7m3AeGnW20O1sql+ci4jfVg+qLs/EEIyTsn9DnavzPTqCtaEMIsccu0rv
i6qqLYbBPiDGrsFDpLdHY3eTeBaJni5r+U5/0NCSf6hHTZZy4D4i2cpLHPkoklvtlgUlazuA5pKp
Q4wdddv9Bmb9j5ojqspn/Gx0oTgUTrWsQyLS3sOl3mKHHLch8hSkuLtWq+D4DEngPIoZTZXYnFwL
r4e0fmO4vRVpImoSXApv+ycnBfME1fP9n2NFgQn66X/4dRYHmdctdiuURvDY/x0Yq5Oip3YAFZHW
/74OZsaFuj32U9CMLKQZPYlCxg07xTuKTA3RHVDV/BsKfYi0waxKj9fhDvId7ycI8giMMrM8LWC9
OfH29JPyVWc3yQqo9EujhhUw5agQXrs/aO87pZWDSPRPZ/XOJLS74cbptgLDp4mwL4SA28aEi0Jt
7pRIAONtjnjyzTDby6T81A6v2ExvKFkCGzhyad7nXyaqPAKSIBYjflRlLbFhUAmh5fGbLFovwyDo
yfq0ewB/ssPotBc3QUlF8rcun5cnfKIZxk7zZGSiJNN3gckxdIKBb6+rUZbboHyGWg+BaYGOTgqL
0NFErTVX5bBOKZ0X1uDXvgOAFpxjvi3aXmyFCFZ1w5J0ZN/khx964+pzRczj7WWrTuhqdIfHpe/x
TKoh9W8lqu1O6x4SJP4iPJ5TloOT7USkiivp3+PBouyU+RUa6/V9NuMi4rbHET9uyhmBD7Wj+Eav
kNb0kanntGQa6YBrNdFhEJQBaV9Z+eQbMbkFnYFJm3Y16KsEWRwpdrYssgZ66myBeibJM2COBcaP
TdUbJ/fYPyOg0nTWr0q6k0lbIGqNuQW9rhtEVd2X21wIb9sJcc6Ek797sab9zHoHr6e6RPySsOw0
XWkyrwbTkzAtChQkYCInRQQo762AigXzEvxM481ROvAyH/AqFwjXM8r+4gLiRC8utu9m+rS0a14J
rjrmPEipNqZ57ihBrk/f5eqDJohr4nIcP4+yuGlU0YU7lQUo/nP1aC28ax84RR9LTEds5OuQ8+HA
K37mPivc/JmXz5DZy+jCHAuCClG2x2pDDDpzoM/U7+roiBh+PsY6iw14plJfQoZTa24VoyU3iuT2
mVuOFkiNjruik5oGz0pWQpyulWpeemZEcblyfeUMTovEO6OKkAJuIXrtZm/DyqvWPG91N3TzCkU1
G+QPbfzjxtusuKvwt7zx3W+h7N09WNHUnsDKg/KfxXfI4N5yet72UNo8TTRVfX4pJt1s3hIeyz22
02h1fNwgCwo81zsIZhqEOYSQACs5qTfkTC1yKJ5uNfc6K1X4Re7c3qP2jJdQPML7/GT7c1jrCmYK
rigeUUioZzVJ4LfXF4qBY9wUCu4Ymvc7fBOQ4ZE/Ql7IYwuXVF6GD1CTcc2KIDJPWuYpFhCUuRBD
cMGS+xlu/8Jr0XT/k2x+7sTnml2avVEf6AAw4TkIWZgfyizJNIz2YPL29gr1I4YW9u9sP8rsumue
lSlAmdrHJ5YU/43A3oZ1bPhalPAS1/7J+wyK2OoBhBS3ooz74Zke/LqHXue5Ap60f4Vr9k5BJ/wi
Yz25AYmpXkRd3vdHcdvI5fOsZ7wQiv2xwcV/jW1EvrbGVfoSl8pt86GB7HlrM9aj2SomzMQdYQDW
x64gnDUFMtSA3t2701PuJE9+fSSGsR49ckedj/Znag6+wAXNHnidC3d0gnxE7J74MuALC0o1EeiU
7emXWpZMZfNnVTyf7Ws+bv+VcNsAKZfMtky56i8y3m/e9B/EHbM3L+o5lx6AMXG37Brg+a4Kc+Cm
uurATeoJ4mVq1BogOey1tt0Sxq4Gm8trIWM+pApMtBuv3C+1i3m9rs7Sa1m7Rix/LCw/ekciYifc
Nx9lPhqezRTbg/f542clmlLaPjZ+btjTdguY6NvNhOiz56jeW7F0L6vkSYCCqUBgUrnSuJmY4wCQ
sLSEzhsPjNkQ2aZk/rt1X0AoTEkkpeccRZdciq8SCPmkviVE9Z7/aZvn6LPi6duXrBBqb/1D79Wq
dmf5144kDxEBPST6tzFewZo+dFkvYhHTrsKCmvfBb9s6NkApIdM8Ems9CHH1se9sTB6XBrnlGra9
ZLLcB/p7B4LD2NqSGpdtyjNS3ADuwHcTVLKY9HLN5xXp7grFbluireV8fpON15QWmwlkIyhVMgTp
hGaxQ1Rsf/9F7Pb6j2EyVlHnflwK6LR3ACiBibB6DGhA3bBnqyHtsLHJ9XoG6OsXJOkCd29wL56R
shUR9SYU4ytx8Bd0HECOmyp7xTFxL0BMkFuLOJdhh9tC6lxKozPsqwudNQqAFfJudzmmQ1uSO9hc
+kBph6GZ+Kdpf6BCVI9aoW7Xc46CWWoiyBQuIILCDuNZhgJJ4v6HGVQaMvvopf3ChEfyjH+a23E5
4HHuvpfIn1Xga00km2c5PO07JGuqxJ6gFrm5+FsT5nVqcB4Brtjaf7ArWROYeKM29v06XHXuAU4g
IrO5/WfkL+zfA2DlaWSbaW8IF9giZFyEeRh0FiCT431KpaCQnwxv+Mtg/hVEJd9ki8teNp54t2Cx
rHotY26kbYICcfBbVeRvWnCoEypsahhx9NuOjQpdgB6YVcgY29aplaXXTSDBdCTDEf+LiqtkKuCP
G8J0Jr9cR6mq45XJF3+3bclTMDjDuI4ho0ec7/eIEir6GTBnAUxbtKyPxAj+i58YVB8oTa+JcW8d
NC4wKdxxBBQmWgroPi1WiKP/moGix7M3Jlh/IOjCirSmfSS0WzttwXRB4ekI7lCFpPjEVzKe2uEG
YQVcmxBQnIFwXgjst5rZYp4wucAYgWndIBzVEuZncDuFmvZFH5KHc1uqejt/f7QTfLM/DZwdsGxZ
eP4Mce3vI19cARmx4L639M2ir2DwfLZU4LJA1EsP261HPSDQXreFx7GnhBZ2lh6U0dfPcTfVNX0H
hlszojNx97IAXESeks62RmQ/N/ONL5WNdL+0sbElGFT5yDKDZE0R7i8fVvOnVosI5X76YmRScKcr
kQcg5ucWedIacpvTlhmEYSFeCyRrHvVDHRI3YyXqD08BXFJAewWgfyk5m6G/TV+AbFhkHwbsgnHu
LOkfcSF6zwD55QHySbBMYwf/txs+u1eeXzwL3Ugv1iLuBxrl+jO8pqv9UBkJbgaVy8ux/REUjNrF
c/+8ibCGGZpeda2xJjrtHjuW8ytgqQ3vtlnpRYc2HlPzztjgj5Al6jGQlXuDzliTvffjvOZzfO0W
Gy0U4RPvdlh1kMuc+Po8LYA0KQKPtibPs0wyMMxFgBhNo7oKFZhRasdA181v7IUa3x0KZGmVMc1F
3Ek43JTkmqPebki2xY3LAphzG0ywTfqaSYE4kIq228lAJ1EjZgmgPSLi4DdaFDsE0nesBIwAeA0r
AbaFP9dmo/BmEeZqtCp9gZg7mXDhsW/8ITdfGqM0IwuJyhJRKOWwQXo51pLmCMCc6Zu2l4QOtQIp
XysbUN0CUX7dNvwoJRPZk0opx6fFbNH5f5yG6kk86uUJCdeJhWZICaWVrm2a4Us9mfqChmydG2EP
3DFz3nG7whpJSLnZIDghpwyoQNjlYYU7scQmcpiYjbt6pRbtYTp4MpN8xseb2Zh0Qs8DTE4pXS5c
n6PQpR5Bk3a7g7B8Mkd3lw1RH1Ejcvb6nWCBEN3N47YAxiczLA5o19ZJ/t5/ayjc8ixZ+qaNU0in
tFgSRKnToetZrCJuy/Idl/DVZBXU1il8insdy/k0keyrX1YhSipgGFXjEp/mM+a6ddDzCId9HNIP
5vB3+BXjXJsO9qjmzAPUTE1E6HilCcx0JdZ3ECGxd7qRtgAyVO/Jl5vUb1ts+TNtnnJQ56rLyH3b
M03c1dva4tVzmQJ+j0cXeecOCHqO0STXy0XOQFI61j9FQ2l/YxRzVXWYYMY71d2cX6gSr9Yg6UhC
fcm3sfXn2+W2ceBsf3nalbYIJJAewPeV8ZhJ5y7Nxc87ba4NGJfPtIvkyjXBxk80m7NGHrREgZ5/
fGgpeg/VBaZIDXrjI+58U9f0Li9Rhvh6vheTGP9v9qTbWARPFqXBHtbGr7JqInr5FsohV3FbU0Cf
yP8TNJ2/V3RTAe0dpIjbBjiWKRpmy0P/kpP80SLt6tvt2vhML/QMNII6kBq6H6oG9tY2iGnIk0Vk
Z3mKFEEccWJJg5wafsjofS7Part3yIPahuAuTyX0ZH8asrq1ghx+OMSJ9Ji3YocE/jHFhgmPJdyw
CCTwHiIg/a93efRvT/mUXuc1m5NYzzSEcCKv7xye+xGySaTGKWkT/TrZEO+eTptEh3E3vRFwRTPz
l/iMtBIA1CzuG5CB5EWy1HxhEiVy8MMv72AN2uCZnF88US7b0NyixjJ11Ni0txpPRdKIwssLoy/c
o7ZNAqwcLP/HplG61P2SZwncnjnfs6hXha1f9Dho0JjxsAr9Q7dUdQR6rkrS8tZw+v+I8Is/deDy
u+D8BnmAuErkrrRpyNKNN9gZgpos6zYD1jvoTN6/uHJxzkCPiWyn6++d9jXcDfubNmv12rY2+j+7
q2xaGIetEIMaNUxX4ulB3SzvOFW00UC58zFycRhjpMTFJlAqi4OJVITMo6yGSHGO8QpZh22AsakZ
GBxklSMUfZJWH0dIkL8NSKRs3m8hlfFlHfaufCNbKUXwgXkKW7vn4EZrQJ0Meyfgsy9Sv/WJGeir
+Izaz6u4y5P7GtTIE3PhgEoHfLCqelcGbqz44Y4bd4A0KEXHmruGfETAKJ5BPimhaKUzASpguCFf
Tm6A8GUiHH9Lz7AoNTQi2ptn1YbeF5RQQzg7qVimQ8vIUr9vRXC9bqj3Uew1VVdkzsXeN1bnu3zF
IwSzkVbj1NwSJ1A7smHNL9haZ4XfRrtFDCABuOBKC6CQtLqVuiPb4WLRLxDmbuXqSMZSayXFnnyk
BItExsnwj6AFtSjAbzXjlPFb58DdtWicA5ASvVEpIpV+m6mjRuMemhasGpqX3VwCPsAZa5tLtR0a
bs2AdeQTinUHLhn97x4DURiCoYAhaHz3GaL9QQanILc80MJHJfXN4o2LO8vcZVzmiSjH6UlUElfe
Wu5AUrq+AGyUVYuMRMygwt7agz4cr9WvoetpSk5Our4Cp3IBQ029+3rjEYBdaI4SmnZNKkPXlQtw
ziFXkiNSnc9ZPVWH4GdaxTLZbv07v6/88Dd/zp8ZhZ0xNwzdFZyuMDbLyKUc60J6mGyOZgw1eWTy
fqgS2PEGvMD35eoqnu2xOwWHv042r3WTQhGjTdnR28nof8F+ECXouUuP8w2OYCyotWYcjFNQOOgt
BpJITzxwqV2tjri1eIlEcZlx+x5PuLFBGpPYUP4ledDCzZ48xdEY7KPlavIPB/viCzd06BpK6+ad
3EDQUI/xEJU4lSiWq8aRZ6TrEM7G3RiVma5Uzfbplo/W8IlnlCK5aOrQSYr+XmR6g2r1XqodRbJD
XHqws2v05zfblS6UiU9NBYvH0nmgKFrwTiuSiLuj7NDttFHe4fMQpKIag6x/yxxnVlFzwkv9Ahk/
XvEKhoraomjni92pDB4vI5vjdKEaazoXVef2fOinrxznsutVRq4iRP4eD2jv2cXZdXytP3VOzT5N
si+RUzg9fkxswGvPfkS/KsefZR9pR0K1JpUt4xrQMwPlbm3PgXcJPO/FzKxSd0x1Hcw6ZKNcuIfN
pUZ9Qd6/ZeGAeYdgaVhrCyBT6Cku1CufSgrvlsSXxWTs6/8Hm4uQ9zBFzESNMp8us1djgvCGgA7D
qm2lQDSblwP2VA7AnKm7TX8bD/iDRY5TjIQ4sjGBkiYiZRoIQRuMwG1+89tD6A/UxSdr0ndr8JXu
QXTxmrYg0KnhjdG/3d4o4SgvrDdrU+qc9FnB3ydTtctPNRApus+6HDfJWmIV8hd7n9rQnnx8AFMP
Y8tmLEgK7gPR8N8lXh5YdCSM6UvctXmsBNaXC01qUtAfzui05m6vaw2Kj8ZF4hCycWlIaXQWFsrc
SyKk8hbo6Rr1agUIL2rqhDBUSZEYXh9rEaafM+pGaRRyIFz/iDwQ7TxR5YV0f7Z9QsCIkspmlmNJ
Xbi9+U3VCl7YRPs+QxAzGLKTHKD8VQJZHF+RKYN1W0wCwTt8yWvi4MIObjc898uRzPyH2F6p06kP
ORB8A5lkGywEWgxRNHxN47nt/PWo/2dzlRXq5Y6aIsGeR/5N/ICfXuqAEBho2atlRZbaOTtUAWyo
dKPZp4AFidpNL/EJhEGij4ATB/S4DyERbM5a87LayDQ0ZOiolH0Roa8rDnae6Yi15mRdyjV/33g3
NVKU0JXwVVWSyITdXQEpT33XaYS1HxwFOz7GhJgxu40cpJBmWfabG6VwtL15ZL4aH4COq7GzObas
xg1ZIxB2Xo9nvLG3CBqURrdkYlOjRfEyS/oFRvsN1aHlSXZy8m/YEl0nfcr9K/QWiBFlkIfRiylH
2T1Wzx4nkn+YDgJKF0qhltoytGeW3y5UVZGEEDSajkVNzhC9P4hPQvtiW0T7xv2KsFR6TBUjCAvA
j/KauIWw37TxJSl5515QahjNeRYaHHc6YTaBQeD4imttxVHs4O6Cy0W8nvf5/0qWLl9MBO0aUiQl
eGAkuo1xqIiM6HNh3P+vSWsc9uo+8JOerOPzIn1PGIvpsjcn4iZZejccIzhImgwH3HVQgbi0Xjkw
a3hITUrIB8ZSam0ch/bhRKZA/AHMGxGqBGt72lELDxjSdQ3puyPSN/ItyAmiXCDY3mlwMEuQnztl
rpeUX01K1EGisEF8YlRqk8PCsRAef5etq4mU8xvlm4nlVoZId54BgaKu7SnlwBEOcnh8noPNwdoz
E7+sL5y696ejVIYUAVXaPC6HXsy4BiQdOrOnBQBl58oteRhBmSqb/4DgG1SG37esiWDIL47joIXZ
M7XYKKmECdIwLJJWJIr28vCrQ3sOpHughKZnfAa12FKFgCEJfD6rPAAkoZUMzx1vUq5h+faULoWt
4B5Q3i5Kan2ziiaWXQl477Aqzu3L9X9fF1r5bmoS/XK9GQZf2Tn6BcFZNv1JxJT54zuwv+pKaqzg
cWxXaf+ybjMpvU+fDIbGVhHd8P+CH7QRlZ2uTKB39VqAcxByYfxZORWsRw4SnFkpxvREIZyjbJrX
7vrgleTZ9cXv6JJ9N5JxSdoJPwglgWSJrQylK10SDhsCuGjqwP9hX5lxU0oY8YrTEGoEZM3RtxuC
HqHJRcztBqzWsGsijhXZE0o3lS1ZxqENdrWoRB8//RcC/XafWd5KCXHn2FzXdYkdGgDwJ2kdFY5A
aO82lBFuxN0t2PrQ7LVFT4Yqd31BsH2o0fpC6tJnVUJ1OkG5EpnhQd6/OgzFNW8wY/qtuYksbq5y
TXIOiybQp/BkSqdzbNRlA0NDj+6QoscGBFtSSgu0HK+i7wrn7y6arZgV8/ITiV7x7nkYaozoWzBp
lwPBX5i3uWomAZTedrZWTZJtzw5eSmDagaHbibB4sI7tfiDBjL1lFPbcA/JF/UUI9VYhoePHeTs8
r8sv793DcWTp7nTD2JdNRDIXLJDmVqIopW4oAtECSw5rFYZUAt2nh1QRPbhAh4hZ3zjdx8lmbVdD
d3bSXf84tqGlGpLIa4rjKCgO9Q+LTHsYKnInvOlRtTnTsjHKuysVOSlgF3Cf/wumyOPIFWz9gxdJ
AR+88sLTr4lyDG9qs3RvKGzYQcZ3zERNK9SkMXeNhJ4iL3AmEg0XrcYUaRGZAC5VfOYutTW6Spht
UB5m0K3oRY7z5PbP6njktwAPi/UgdKDIdvX2yAa327z8H5vK4lf87WSIzh+A1BKPwK+UifoehP3B
UPomQL4C6zpewWqSYX3M/xUAbQHJk5iiEDQEf9CYSsDI+lb7zcvydMryTb+gQqUr7AsVbKicqWJc
yNE2l7/shdVdCJ6FuMeo2/XQck5LTrjjnLJUO4Vqw6SnR66+JqCvIAbEEO4wB4VFIWzt64ms/iNS
CnoarHzq7B1HpKAP/fKixgj1B30Kbs9KeIMmx3k/qssO6S7l1PBcrbsBttnHSkAgXdewuak2NVXg
ejXqpkjh9ywodFvSmSy+6Oc7O7SmBC5rvx1cr2DbxWmwfb8Md96WFJm/DPE2m47cK+/RbK/jjHm0
9PbI7zNgnVM2ugzjsTPE8B7kY68Kh6tJUIH+mn9ORmstF6XuOJhlUY8fqafNjHobPSIiHNXZB8wh
VOTKKr1BztnXK88suhR6An7c/dYvg1CnoZpdJzLEDD39C2MT2y2phXrZ6TRS0d4QyjM/ARt4Iys3
V1DMw+51485Rc15m2j/oD7kZc1rKPOjYIjYUKFHg2MJ6DTCXbM7OFnQD7GlvJQGvJLZ5Evdv0CHY
ZgQrckv94WDP28pXtntFMeq9ipNvK2RdsCOpz8GiCH/C/S/LwoHdk90FYyihZ0un4MSoGih7YukC
1iHrOrSqqUASv38K9xVf28Ix2hybevnjFl2kNjJp9XqoVqTHH6bYCxsauURaUPOjrnueNOMLfjJy
6XdOUfG/p9k7bQCjlfEH/tT6OopWTZV1LsN5kIfNFI9XO2krq8FHoAvP651qqRpzw9OLRyvRq1AP
EUW5lkE6LgByuGEbcFDeywuv/EBdoDBrCZMRnNJ2Aqjdp0va1tO9eD9htay4moHJKjbDp/+UxLKE
X4TXlnX4EGkzY7sImnzKxq30ItyESOQSw6pXYBNqySxE83y9h0afQeged2W6VLrYZ4hWkpZEbqqN
3RDfmyF8doM2n3wvxG7ZsyjOkRSpnc9O+ZRoKRbNve/3JBX1dK9xX7fpc5KcberMzJy/K3w2HeG4
k9AhAImPrk847Djhp9JET0h+zjnhBwDTEFuiOySBUDB0ctv/WFKOXUm/FFx+wuhOYFyANMpfyTOK
PSoFHO6vVveJIyeWt0puxLZLvXXRvagfKeIf3rrloVeidF17ADUcJvQ7ytPa6jGYuDxiJaiAT1QJ
72Ag9s0wrUklKhRG6WZTPNSDr8rJ3kNYOeJLKl9UAtJXQ21MPJfgVrF0vaq/4g3+wM3aMkIJc6zA
2AV4/iCYCMOuR+ZBsTKHNDO/novsLd7MRvk1gvQleCMmCJyoPaIsls8GsiJtuIzS42rUIi/SvBof
7UMxaopIjpF5Yhj9sDjqTAzHyKlTYuhVeN0SCcvvNe2q0uHzt/9g3a6FgeYjYhnTX51X30v8vMbE
2kHvZix/5gPbL/CIAw+c2LzDX54hfZajL3kRWZHBt95065QXTQr4bRD8+XSSdbpZdFnbn0vYdaFF
XjZzT7rQNTW6ILq30Sok0a6vG4TLkIMTgcmDFrO8KOZt/IfrBlWLzEIPwGpaLzL9zhahiqTmH531
S2uT81Qsc2kviDMSHX/ymkdWDTm4HQr1EtkWdIhfijFUox7WT0MJot0yFyR2kY8rMzujcc6wAfAr
u9mCDYNrdM4tpaIJFGL7pOlhQhMcjrXYfd+DCZvvP5pQlZnmtEGWq9+wWIN7wSSKaXIgNJ1Ol4Rf
olUqie2GNXzklCVgB76vZec/nLKp8sJK4kl+8Cn2FHPwXlaE36hx1YtPOKnKYYjdoeqq+R3G50S6
fs/iFwL7FewW3tZXVaIP4m2deIj11iRIVe0bjVlh3MWI+zesl1Ejx5+0eDL3B1/ESCa5Mpk89LWl
sAQqbL9szlxI55MGFu1kTcaXQ8krD+KAcQzfnl4bjQjmQ2Ffbzvy15y2TEOZalqXTujsUPm46cCG
PX0s5+6jgZQV1+F8xrNZAtvCDC4zui6LOCAUCRy5mKr7Yq17LAalb5jcxBI7UMJXOph3Fu2x8ja4
IuZYNLqGTPhWph2Zs6lA20SnPIke7+dF6UuIHR2K1ldHbJGQyZj3f5EbagtDP/+1xBXKabb2bu/k
98tWxqRVH40GPvu4ilX9/CvYDeN9shsqirYCsTXuF61qSd6vciLrj//Kk4MOgbURK/ju7Y01aN9L
et9VC1y7nscOIG+gmqVm+WJ420sMMvsTRvGRlSAT6+OXTJ0MeJsYlYHGJKbptRUKq+820Z/D5aXM
EThJVaXyLROAbUaiUSDzznvNb404W4Ty7o8DHHTdzQKX1xj5I26F3yMFdRbiW2A5yetj/uvYcPHB
OIOKD57qBDLQIKfO8iQKUsaDwCq+m+dG7n7F/hIAyLBGl9oWUczykgd/hfAJVNgRlJ5ClaS9lMnv
ilXmEjLsuldP1mmOAU+jZFl3iNwLxof9xUJ8XMGbysogQ3OxUizlSv/PlxCCONMMXIV1M2B+XSX7
eY/9o/RcBetaz/NXhYCdNMkGajp3ML9l18cOgaFtS68PLM2STG9n4sTDmBevjsEctXVv2dIX5fVB
EbsFh1N7DE3iN4YEyRd5xKz+8SWTMACFFkk455gwdWUBQma2c6PIRT+htT3L/2OYTVrtdz/gNEpw
cs5/CoKNr+JnJgJdp2pC/I2mD0KtS+GJP08OSb5sOzqDjOmKXIz2ZedQBZyDnt/EeW/B4ni3MXyR
H/fYJawt5X6J9loDeL+GKZ1ot+w+z4VodDIwFWkmmdv8Lnoou8+w4MiXNgYMxL/1xSBTw+9nRd22
EhndmvxUwsmJYkciWTWJDw78GLovphow0XZlOH2pv1vmczzzzuDywblt4vqlrjvv1CHX7zIO3EvP
uzpmVisjA9d67G1Hmo3/RNktPG/ADtAnSheKf95m5oGPQSMMDLMvLRAWlgIodAXjGW13hL6rAGiK
76HZlChx3SugB1y3sbXdFWlzcmx3H2Xlby/bT2gkPqt6fAyS3rP8H/J9FLC+2rFnNKcSwTw5DVHy
17432rLZNjsMe01iJyfSsnUMZZO6NPicyR9ZpQbqRgfuMeYsaZYYzte8irvEAMsfV4oa/Rb61i0W
u2yxxzM9nT/uxNhbKs9omnPiJvG95LDBIGLdoySLukckmJHeSIhV6VmweqXa8JUVGZlZnSgjnUsD
6oCcb9dyIQQPUXCnKg2dKUTsIKFuTLkuZHRy1OzAIYhkLX+jkVGGqKNQDR3l/iAe30VLyK1i6LIi
iLy1oVWocILcUwSZeXZhnSXWwmPNVech0s0hl+3pvyylY7YoVw4KsgrwinHE90b0IOSbjQoBzsiG
RatQtaih5+WJz1bwML0YHkau+AFAPAR7oaWxRPIE+xVupbmWHkTWWBP6T3Zea+9pVpZzITZMrrz8
TozwNBGPL6eKA5h29rusq3lPIjFzU31IP6VC6Ef7PNo3c1eKTkcr1JGNvgMi0uw+jbnBbCczF+Vd
k2ByLYcoiSi1FERljlZhMtTBcAEQGgGWeQCB0BMYqhgSn4ldiDSwi/lm+uXeltMhMLngy9KiCQb9
YTCoWVkaKD2fjEi3IB2dICHOnyyHcZ9S87aAYyLip2gqcNOiiqqWLDDmsMCSVe1fQsUWseUoRQGW
PaEWjMnoS47NbTqqH23fiu/sNcBMCmF78fxqDh1kZEahaezpAQ23HMfhE28ct3ZGnnOhBdxJp/xK
LBKFSPcKJGAhXolEOXrq2LOyCT6y+HKBJc6DyYns7dEwuCBdK2gCXNNW+i3rJVvC5f2wQPA6SH/n
yy1W6KEj5dg9e1Boh1QENIfp7T84k47BfqNWAATUIi0cs5+VMbYS9KZlCVY9EXAF76HPfWjc68x3
xSUinApU8N9RRXZHrF70qCWx6aKt2fmMhzP284veyI5L6iBOJY+A1vjnGWbzcL50FpP5t0xWBb6u
RdTnTQuSVcGVY9A5Hks0Fuh2sp0KIqKOjBmFJpbRgg3dauZU/8vqon22zrXeYhpSSRwWV5Xy+UAG
hhFNEx7uKoG6P9UszWb/2HBnftb70hYG4tXLSkdKcfgqqFghEdC1nKDGa/BEybvo8Jx7pAqGPciK
UP7V6yp09bFrEgelt9DaV2/48Vb5YhPyQQ6ChShEYD2aTgJPGvBcTMtFNGgEluLcen80FvIqNcWW
CDVCf39wu0zkNXPccRlj4yLlIwNUzNinC3F64BrFQ9QfAzRyXYECtuUj+NGL9TSGlID5YA2QAuMn
jI+peWpbqztYiefg/Cm2tVP2iwjJGDJ/8XdH+c0uEZykuosMnnpbvvcUOVu4PpdTesz+Wj9CSsBC
4Cql5jNXIQza82GCj5JFmNaiT632cJxufvnxChEvlMM/YHZI7onoPB6ML3aw98J/b5VYm7dgt7KB
mu2fymNkHDCWsmeDBwlt4BwmqvQ96lprp+q6Ri4YGIHMgM2CHeCKrof3q4HA5wM+HlnupgmFiSfg
0VoldJLj0QhuZjqCd0KJS5vC4cPJbS6l5HswH/To5UxzTCcOTS930BSMDRcakSTq4ERWMhNNskvz
oWj4vfwWziHWMuEHERH6zXsi65N2FEyqsjWR0i8G/n024SmVoDJ4cEIhLIGd/XmhUsAgNtM+oTVE
SeQlMFnpIPxJmGIX1QcVollzwi/fRcLVACZS1WWIuE6hOZYKXtDGijIkp4wkjdQlTjk7sFiygem5
dTLtos7DLBQxFcoN32IOuFqvS3N4pKRBYXYCAkV87fCjo4/t71lfNrhTpXObr2uighkzrtG+I+iR
6aN0F7VPlOk4TJINwGHxs/NWy2EFV/mUUOrjMtUSxZilmStRItQMku8u2kMhJ/wqbi8YREn7c7DI
aWS7OC3ZsHhWj7eUux0taEOnpBhuIP3/wgei+OEMA68Ux69MGd4m+L21hNOKvOzJYk9wkYCeBfKe
YibsTeVx4qQVgJ/pCu9WZYw4nxkbTyMfrKwAqJiTpn4kM/8X0JEqiiwyzgRr9LdaoyIs9iNkUJ6k
A8B+s5TK/xThXRyX9tHSz/XfJg9GX1wihCz+LCr3TKUNR6MbeA84fMUhSvaIqWuqUqEGL2/k8XAg
pp3wcukEwaMKTFzG1C1/qv8hHNsCAYp6sYejUXAkjB8+ik4R1YXwZl+eoUgA7h0ljzv82ljTD6rf
0HSyugvo5p2g+mS9TPkVCdopdabnCqla3fVSS/zdm6yDy4FRwjCLP4gcyK8JV6uKmYx9Z3yYDHSd
awb0kTMjH67idbUKyleVem2XnaxrGzTq3WxGd1BUQo5VQgBnRpDek+PJ7JuuMBk3NHHnSSpJm9oX
OHpHTyT/n+c4r/5wLVztI/z1aT4LzSuBI6WQeo/+F0I2cmF5XjCxf7fTc+JjAruWDndXp0XEqwEV
ARxDbNu1MxOQ9wk0EAc1Xx+RZZN45x2ZJtmPao3GtDLafws8HVBbaMEs6YHA2krZg47yJqxZnyFO
6D12iV16JrWT7XUvfyT5FMUL36T5O+LuchCo2eARa1xRTbq4M/VjpXwsuv89urNFAoRgbvzxousz
4P3iTaQzcrO+hcCsM8+HMjERTXo3c3n8C8qywrLS44M7c5ELiZmPlC4e4AnninYXxVhIpAgKZI1q
bgJZvmKbtcn//peMQ24pYza6HL+wcoN3pj2f0pJZyiLf5SZJnlRTVeJfd3xQfKGyFtCYMD5SnyrB
JYsOE39SbV+gAmuJy+z9lsOpd91e76cgPpVNOEO3VyhnwL6cq/35upRJJ4zeMbAv99dfN3x9TKeM
fSHg8rvFElXFVvCjka7leq02zOI/4lJtogpuyMk3qACHRCaDkyGmPpQiwCPmd+fx0ShS8ix2PkJe
BY6Knb6Qk42b7z0DKrt2wQANKV4gXiqBBQaxvNFJP16GWkSCIihfKDzW5GaWtLBsGvxb5vy7oxnL
n4R3o6pTgBusjP4CD66Bl0HmBDv30UTS79fn7p741KUEJdzWkKEujNmkT+9qWacKpGy9A+fHXp9m
7AgDcjDZ8h9QoRIYuklUMpk4mrBqdjt/qndIMVgNYaI04mE4amSCN8PKslW7l3wU8Q5u6EwL6ESp
VvRzBuVUIROZmItIiRECPHqTtylhBh3zOVsfkatMncB+csefbLtqCLQZDrSn7392xu9iemiCA/7p
FYRtYciuEI+ZcfLcodTIIWWIJCmvdMl3RzfQwbnwNQj4KITccROKbAR/oiaSX3oQ98IxfDxCWbRW
7XqeWysWCfZ1WYfyyoPBzHiUv38M2dQEdBCKiZdv0rQG2Oeo9zAEAxUwtP+2K+jwyngwLLv85T2/
toKR9PqRgBHGfSxaKnyfqxZkwzIlWaRRyhlSNjCBU+PFsGGQ5SLLCArm0CiO7FvJR2KL2OG7Wrlm
LFm1CvSEsJ4PBdgSe1Fw4nkp76rFuFnkCxSUQBs2yoDj8iDHYSiIDZAqhlt+iyOAyiXPh5l5poRW
EICuJpJAZ43sg6NyUOzKu5MY/NuEdCUAjV8kNA+wM0R+LKBii5rbzSEH0LyL5tZ4T8GOdSENZla7
c0XaF8umlF1qXlhOIY+Rb93lWBSHGfWetxTh00jl8+fZlvwx99wu0IMwNw6wNlg6RlfaXglStU0F
fuNfbU6E2VaS999rM2QqA70sgz7BfMCX3+qFfBy1Ij39huOJU5Camw4Z9OB/4Ok9Jjy5yMO91E/x
k4QPa7lBk9LgwE3uR9SmWHnQEMvl/1CpvzjEOWOFQYC9F+NYHxyXR9Bg8viAVrwItM2RTo/hEzl7
iOgEKx5SKu6J0GlUp9rBm3HEePKxEEt3VjsDNPtwFTFH+xzWIogEOw33Zro9EwIY3l3y+pnSZzh9
y1xZYZaLb5sanpWMgUEf7YA3xgnvjHZG9wdGaR9AkOj8CHeas3RK1GC8/uL3S8pEKISPfP3cIDUH
Grxns5JtPBV82Dd13+AEqoJ1p6N0+dGa12uZxwsti+m/yqq/wodebtT17cSZs5NjfhgXE4FSC8Xj
C4iWMUzi7qts2O4LfYhviQWYmqgSXwOdchrrNBlPWjD7oYmDwbkTsbakobcnf6U08/PHQv3qmlIH
qOKwVMNbMiWajs4ku4uJTArWEWfmkJYnczu/8H+CJPJeFk4FmswshzGZIhZyLyFNShqCxVQ/o5Rj
PjrGjjFLKiCL9w0U8/M4WmnAmhN03avUVLAYNte8pG4jLfEqXOgXRa8NOkA4RC+ZT/dr8pa/i85L
pTCvZTUOFACjwUYCkwfPuPZc8GNuyJvbhdVsvVp/YuddECRpJiSSQrDJnrv99SAWhbf+SSsEmFqQ
1ohPRDp7GnDkNS+crU7Ac3l3pznpHt0GuwtnUUnjnG+XpcO0unOVjHglHxElADHQfNisFpG8G4LM
swq25c7FajrYz5Zd8cKAOL5biYBqzXNiokVIUvvcr9kUvja+QBx3QBJZiqfljj0vMTE92tnxdkUE
xqz4oeRFmnBsCM8o5MzgAKc8B0k0JONgQiSsf8FcOcTZboavP81vaCoG+ETkK6MnXoJThzcr4EgH
akjwedZiuNYunmjUInsmhh2/7XFdyOWOD+b7KcAIMY7OzRTd8oTXuzaSFkGW5uuddNw0kwGF90BX
XKPXea/xKede1itL8am89qiGKBnkX0m7Onhr8abObYaNoWxRKUXleaSjeSm/DvWHPA6fU3fc35QW
JQdLOqgG0MZtFX2TJPFGzEnV5bc78s6+PIL6nu/TUCD5IU4w2P4/TyrR3Z/i2A0fLo1GrfG/VuYf
f/oP2K9stsS9UG1vGHzBkew6Q4P37iVOJaarDMDBt9tUsLKpfaitRAK5m5zHTu7xIV/j3DkOvzlq
X7qB1Ag5J228OX9k9OLYfUaqx6uL+ev1EzCgQ+FeSS65woJiW1a/X6FND7LmhlOkPgIdeJJBX5H5
yKLXk7xOGQLFz0GIB9QrkswPSOWickOlG9KkAL2kxbu0oKfkB1jMX7PIoHwXdCthPFf6BgtskKCf
ECk2f9wBqf4Amq2msrrfSdI2n3MWWIC8uJlCRH4Vctu7D5XjVfoXAkS0Kx3FAZyPJWu6KmbQHcV5
phW6cyLFvQza917y0f4vAMplWboprLxrQ7iJZhkHch66SWvkHPX4NVpq61/p1J5yymaHPMNqbt1E
8weRQ29JuicMGrKRJwAP1amhwTpD/E4nrk1rpHHcyiK9hJEAz2yDAlDJnVUwby0fxe8O0hCOm4f1
QHI/4si6GZo3XpRUe+mQWX3gichDAlo6q9XLELr/JhOzuU6bYFJbMGie1GzTtK57L01y+GHAlFX3
qTL60/gY5a/5DYu97sQb2yaX5f9uMwkzohDMgLizIG9wjqWjSaD4AbcXJjHczdLCVpGpM58mv5Yv
EYWjfOsztWQLAGcrGlYzexZR7mWZiYrdbrjyD+cQsCYOXvgMhzT2m9j5e+bs0DHXLvMXcBNcqlPW
9RTc/N9ikBZdlK0I/hpqcH0qmMohmlucdYRkaVJ8Ygi0misVG9IDZNuJdbD0kxZPj+m89BGedkc3
BxJVq7qbBTQKGpBOi5zGmem0EbAbC4hggPajL5T1TTZ6X5a5LkarIrAwQlNJkb92Wk7lShZzx3fw
2fnH8Q6tBXw6gmHDhRqnPl662tW+DMgz/SlNjp+hPMh0mqMI6aiEk8NvJEyHUgVtTkaM++2OrLMR
BNMQvdM9xInMR7H+GCEuRc6KQA+NyjzUg44zUIhTQHB0dJuV1lQcH0rc2W0EJ5WFA8IBBqJQuPqx
tM0PYWmtxJr8+5FL9c4F+rzZsjkfsGdcnDgmrYQWj1fbLP2LmswT3NPv2un6sVYUQuHu6hen71si
K/eDKz578oVHJVoR1wUNFyh5pQpzPtjVJPzTVH2SVFEXQRYEGVGn+elAgPhoc5a9u8SHHglUTIYR
+53j2+arRcOjKF+r9dLeTh8iopMbF+6ueMPlveDMVcn7kpoMbNZbhiLzlieFOb/FES+LGL9l9iyC
tQk9x53Fe5r0qaYQsou48oHIDE3yNU6ET64tUQb9bIjmEKtYH3/5wXMFd6XoiRe9zKApqTVTkWP+
BvUXyQM+p+IBcG21aofMBQLDpPije5I5r3+kWCBetY+KTrC8zk0uwfc0oxs6W/F10+7JQBudt6Ul
46UqhrMJZfFDIqGn/eWvkUbizKc6/qBOsPoqBXEY4/lgbM3hUsG7nugsSKPTo2/fLipP3/fmRRAV
n84QSDeXgoEL6JVX3ppiQ1zkUXdxT2+LDxDKop8GofxwFhzMsdUbKAJnTTsUFqM6l1M5NZqqOo2Y
yat0jVXi2nHMZ9JYgOud7lJmLSB3U6OnaRGUbfvxWCbzsHr5EB2BgWRqQURK0nr1Lt3R/Xtmjw5/
qbTj3AzGslE7QufDBuYJbg0lgQV9QUxQesSwwbwuLXgxcTXRYhZNbqQHhKwHlZu+RtwrAjfBHxBZ
P6cy8EAPd+g653Gvp7TApqBk0+Xs1v48bWElLqje67qpSKr3ZNIrEjftjrVGddecVGb9d77cGdmg
A/wrxTEPSFa5wWFWJBLaWC2mgYug/+KWcsIAMCSJdZQzxyX9A2eRWBCq4QNAQEJhc7VImskph+HS
1HRIAiqbdgAr4K1EoBLfsFqFthPmTTSRMWBVgP86uEoqBpPCi6TptN1jjUlqzQvgZfsHauxoXPwS
kNFoC7i36yfwBxA2UM6RvyawRyp3yzNZZoAfJP0QWVbQUH64FBCVFapd3Z5SBxT+q9uxFKOt0bea
wrjB1ZtZjAsBqLy1OeEcM67D5/oRGmuF0T61wXS18UiQP60mwL3VJa/HszDd6pSu1kMZbo1FyCYb
KlGOaIjP83X9ykg+43gEVBSiuMW5nNQjqDRjaVeismjZfSAM2VDL15S0wKPm3UZxW4jRnkrc4fO1
t0IViyeXN2FX4LuViFbnZF0Mkro7BP9LJYw3VQ5J6+SPCzIE3ptdTfRF1iGK1u7cQAVyQVKgFTme
6lx9yXkOaZffdu4simMgWeuOXIlfRRTJoucWmjul+YZBLPTfPSasEkSM2MZdAQ8OPBzvmfDmESJk
6yNvYKD1jnmfnJjK/uffe0SuhN9UQ0OSFytGW7i8jCeox4+hANPXXR3wFok+aBZcIKWsWmO8KYZV
p15AfrqDedhYCgQJMxNxjvry73cO8r7pZHPclN93RO20Vrx0sdkdvUgu9eyfxzze47L3YVgdkZ7I
/20cWa2EmSqY3E65lFtbdVAvy1ToGYXJoz/sTC9sF5xlULqzdtgdzjVG5F92CnWZL7zQhYjgQY4r
powaszd/1dImwoM/GMnJ7fsBaOzr7ihBo374kvX/kZRj9On9NWCAuKD3hmGyDuMwwZLyW1IilC8+
qUHfA31jQAixoYoTQcdtoVPL73AQp4TW6Jr4p0RhO9DpyQjyuiywARYPXozrbnDyYiaaCNmDjVNU
7q4u3AqfKIp1M6FNy0zjjeQxZnYXFcTDvSzIEnwaOc9usMHN96Ad7UjxVMKh449claK+Vwi31WKE
nmFze+D5qlStTVGhKqWQcLXAEIlVoyIF8PLpEvDxjr2Mlp5+RYvJ2rWSKPwj1Czjf5ZcPr0CeLpM
rCIMqXbgpeAw518g12i3Yw2y3i/91FEdX+KFy/6ngRL140ngXsRgWq5vBXV3t8GoWa6pYSV59qmx
t4fuQLl2MABfiboMbRV3oeyM+AFF6mximnPStRfUjsSnWf1Thim0QyH5OPuFmyStDvR5BGkVBC/r
82elDv0nHXKHRsHfG/x3p4t6lMFQDRzlJdKFeD+9so2CWmTBUfgEsR/7T20kGEmMccSipq6x4hfG
nZ3x6jZ/OyB5iW1MrYD4QGJsmpG/UJQ/ZpPogRvwPuMytLuRmt/kqGAzPFjzBg7qQB5s7hDqu3VE
keClqcEUaCUn6KsjQjAsp3eIN+RCW7WrABu9fBe2AhySeLISpKaEj4nqDzRTy+eX+IUhaRF2+GoW
TIbwlI0D/aHW6ETNbpfRhwDMgaTJuz8qsgLCWi2cZjfkKpqMyAzM768E3St5SlJDVfn2GOT4O9j9
NHwMrBKK9KSaWnQraz/jVSsFZramwlE+Q3+IMwa4/UW5xZ2ix0J8x942kWIFd4zhndPktFCfI+rI
4Bdsdf5FvL8gqUwC2/zCAXirknkrZYd7F1w+dr/NDALNsxlE/8t6+tK7mk0ESBGlBWs0UI8I1oBh
6GehpTGJAjarTmHhJ2eRBfSOYZ6QYDRvkf4JeqrUdMu5QfLu0z05EksthJpCeICPgnGWRyJs36/z
k76vE86rxDXwexHg+TGMUkl901yxMT17tq8quSLbu/3URx/85/y9D4yRsmkx3loxwvziC8a7I/PE
GP5e5Mx0i32xS9EtVBSgLHEKATgtIybXPzxdGg49yTDGtnGNP42v3BhiF/KeKn+5KHTpW27ABxAF
G67yO/WCUqCU3hki57zX3JV8TeP+KEY7/3Kck4paKOm6+RuGWIb6xyiw4xgiLcBi946EHChBj7DX
raLg/89K6GKD8psOOm6kiMM99qdwjbk5VJ+rxpOkB9f8LFDcwwJadEsFxdxPA/qDH041MnaAgVVE
PJhjByEB//tGNgkZJ09Sq0aQ51h7cK1z8NLMdJWyyS9XsBN1Wnbl+bAgsE3EZMOmcr81RSQnZLvw
pGrwBE+JFnayrM1DnhAgFBQCgV4u7DFWpbwl4cJJSas6LTKg1mB016zKdvd4sDwTjezWJFW5AFZT
7hV+0PGQ8WmPhkKKEnzgeJvDGN3ZAhNbsF1ooGrrVwFHNWm3WPq750GuqmVMhKMT8/ZPLwSDrB3S
wZRGbib4houTA8wrj85LTsONvRNIZsjLuDXtbmmewCxsDhg2i0IoCo6QGYC5F3rQYnoIDbTQe+WJ
mPxEJIgEJZmva0TMNfBOmlgOv1bhSrGGTMIX7FWGImUy1rOqTni9HkAFS17QixQjl4SNtXk4iEh+
3BMW/CGz9sxwfOAYQeKW4MpPwa3ARrC7g1cwsoqfdaB9BXmAxb30Gb7i8terw9vdnKzpGnkknd6u
6k3MjVHo6Hyufhjuz9H0bJgKm7oc+uD/WooWzeExG3kGqzDcnVCtr8orwTgxK1vSws7L4/YHXCsd
lmja8Vc/0d+8O2ZsLkWktnfwiRoNsz48SPyL8J4RWAaHFGeLiDZtGuAE4vFRbEzznpbip64mjjFG
n90P2DN/1rLHeVcLwH1HtfVKUQe60GcfB9GvyGVfzWrvqyI5nFLx33wr0TMFR6QP6cKELLeDL70Z
iO9A6cJOCIzvco76XEr4Bp3ldnbpG4+pTLuf30ZEH9+E88tgAZ2hfrbQbURxj8nlfzNtkPT3drAD
XH1VQQyt16Fak0qy2ULTiKbLm1/OCv9+dNfklQ5q/O1FWFpB/B2l2D6cUBe2YWGrDVSu4+HIjI5y
Ov503nt0rZhLAVs2lTk/lGb9rvM1GUDFGRBO6hboqChw+DWjyfudU5Rws/pvVo1c8cBCj2hckHb8
7kqH9T8fjjxGNCOLGktLpl4tnrpOTgBS/8tWEPJBgNt8LC/b9uN1KL+vkkAtkpNhOyj3JzpRKjcg
S47mCCPP1ubVbhR5IDbBC9V3NRVE74RKaNvsoUnra55bWszc5MNY8LfvYHK6tdS1awo9N59NrpwK
Hrm0eggGoY8PU761w/pmIiN4x69FiX7ccdhhI7lsbY5aa6feEFzXFqYdZBNBQPEhuJEXGTIUY4bC
sQCdLSIzrX4LaDIXcKG6Rdofv4OUn3tpHWZBl2xVJleMv33DgS+PNL4FNYvA0LT2zQoGxk09sBux
UIlkcq/p8kbEPoFwu2RsFXZojDHA76aIvI2b/oaEbsgj6rjIgPjKCznf1hEjitPgVafsy+ZaYp8W
yUWnqcZ/gmq0irylYA99bE10ncOffbsq5vdnh0faclv7ACM3QxPhIZ5iy/CB2s3WtA2Wet+Qow+Z
1A0tpP03/iU7lDDqFq0eCSFnPcoFq35WP6hHKxqUyIu7YLVRAcIb6EtWsLNh36r5srj7YcHtPbHd
rzGuRjW2fNSA5hHqKXfwb70E9qZ+5LKWOrfsmmlhoKQQVT195mA/kYbmA98968XvQnGJ/Pin0PjR
k+Ipq7qRFmr89eXn+Pdb0wtpvy2CSInt/v4GRd+6qKP7A0nlNnsvBsXcP53gEw1HytfhMtS2yWbS
R1XRdPjkiFOJsS69qLRJHiscBFhA8rJmpwJTiOaO1Z3wzwUsjnbLcMHe9edQZ/QIXcRTJM9NmG9h
9fO05RPQ0BK/y4pF0cEXyeCWBn5iNiLrVetfkrygtO+N+Yncf6CUaTtluZjI8+BiVyX9COQ3emcI
tfod6s1mSKbfGI86y73AFYdAqIB5VKCGs/xK3dUB1uAA+HD8En7L8Wbcbh7TPO8f0QSHgoC4cJSI
zPQNUNSNttOB3nd2VkUC8MOqtv3+7U0fVr6t6ESldzCjplDE0xwPZk15SKkWVlX5kFrMeiI7n4hb
lSRWdqoeLJAKMOOYLPbL4jEnjY17ieapdWOoSXfeAHZBULsLrTF7QQDJU/nvjAtYj8INGpXd7l/y
BJdQDwtFUj5tAcJQw5kSdZAi4xvKBJ9ytjEMkhwT18CdaWQE8ixzqRTtHxEw77jjsKT5w4WylHUK
qyThBtJCeDjDLh1Y0PMMb3bQ/Jnxsz8Fsvb3fDNdnjFxGoIY0Qt/1kKOcm0WGx4YNGPvTerxKCZl
UFOXWjYolt2W1E1nbKHtpqBtTgrtz91kBeOgQ7toSA492RxljG8XNttyI/rgGbIVtMd5RMYPUyr4
/fy19ui/Kb9VMEOX/5NjRGupTfb8BdiIIW6lOeAm+fJXwJJYAhALoJWve0EDbeD7HyINlFWkuIpd
k0EARKS0PDnVNw8VarUNaSOfzPE6oJJwmKTVgT18huOALc8K5UWFqibCyXFeYQNh7LAf0CKZGkq2
KELP1thlhzWB2niJEDeiH93va7M5NWUOhr9VMuIAduCk+zCD78Hi/+85/ewc8kqu2srqMXGaUhSg
EtoBbyaIFGf1b4LmcDAUbGjy5b4vzqWXaWNgn3SB5aJLtADIcW7V7MxTF/MmbrRw9gW3YqbcI1bo
PgapEi2CNa3HHXRrPwPKpL7/BogkXm7p26qiyargaRU6r5H7BB9zbYUKZpNUanoBVekfMUCIzQJO
C9x6RVUISZPh703Ct62UAtLOm5XbjzcvXctk2vuP6jfuIA7QQc+5DX99XCpk+bXTfxD2F6qS3nL6
XtGB2tCIUI96AZ46a07TPGsP/6gnI/59MDZG9XMkWTzs7SPzZdNokm5Ro0GJDjDqg8mlsTABpGCn
SdacaB/Rdd78pYA5tGwaLg+ovCRjp+DozXS0+V6gNf9ZKMbK/1KpbN2O70XKnvGmwPKebgrICMxD
zaVdyjsinth3j0OwcIH2mfBlSqVsoSdBdmVmd1FioSp3P5IZV1tAfXzzM6RfTDCcqA60r3T4rKCK
omCKkrUWnGk4XFf/kBMx0I4evmBG5IExPofzNa4TI5W91xb82RKKhNAcSo6sdQhv0zTbc2q2EyON
+9OBwuOgPHdDfm1nEnikFMidKK5YjYpRoIKR4fkZ0Rgg7zDFEA3Jo9t402bXUX7qeTymlBBsOxYk
XWYuf+eWaWXgvNsT9sU9RwfWdAq2qZ6wUAhlEt2W1DZa5mcGpRVZzmKbipjvczaaJmOY+zCj53B/
A5puiio13kGPHp4q3TL8c3L+bDJTnLDHKOFNq5Zhw2/7QiOBdkj9mBUgwBJEXt1iITaJjO+purds
9Js9x2KwbpCr6bDZQAvzNw8/2W17dVSTaj3Av8gqkhSW1ypo2YDUmR5Lp2Q3fG7CZGyMtseO5zH4
ZEwX3CLNbkxnZKxRcpoK/wTeaumQ7JnvtcdbEhH2S5fXDQl864LVnyZBKu/fUSYP9lgsF8EK9Ce1
og+Cb3lj25yP8Bisi2OCwi3rby8X/6yQCPdrK0Us1yoJdMq1JB4PnGQNk/A5/Fb8ea4k3H6OD4xo
tbsf5Bh8SO8drtrfIdcYfKJpGYd0YWBxUAwnq1wXW9+iT34aq6ngDTqcuLXCZaI3ti9toFSHyE6M
mgeXGUWaJ5P+pDgh1q8TA6eBwOtt8FJ9es8IIikfMMl//azQ4NTXbavgNs6REpcI3SzYVPcpGgtf
Co88dsQvML00M+ArvO2WrN8P7gZSTYbF7MJQUkPTTgJC9As3aJzjsephLRqrpi1E/K3t/XhVazyn
NvyxeecWS3FBpETOBbUEu8RfPHQ4zAEzKvBgm/K4IVRjrXeBmvIkWHbhdPZgE0cKw5yn87UG8Czz
gO0CfernuMo4Jjf85UAhTLz7Q2gx65ZWJF/4cIo/j01yoz9+zYmxAMT/8lvXt6S3ln2D0hlvTe3H
iVan+5BCijU++Zj+UR+tPdjVqCNPN/gkSpvBiHorHHUeCmiIbBa93Bohv+BZYc9qq9npv4tXC2ww
eyd2jxyG7Xj5mAfHd2VICX4EYpvh8I/U6J/97eUsTeBMqIYy6Jz3BCxwX/K1uW/uZpfDUR0yxHK3
RKxEYZ3ksiwTFAVGu9Q/xtyXXKiZ0zvNLh/4LdqaHd/5AbKhW2MN/XpCzSZ4IndgjBos5Nq1xLfC
3UkoRNGGs2/3kunFqIaFHlss8sm0X037TMMqKbmqnkuvgJsZ6BUGYyXaZxJBbZQQ3kpK4qRn2sEX
6J2LUniQ9bP0i8xujQIrZ9DKhArjczAYC46CPP5JaxQHq111vKv2HNDnRvuF8psGJlgqEe7Wr0e1
QbCLGvF4I3GQqC5rnaOrFhQszhJWpFUncze6z7vcpzsRXUxZ6uGMJCrN6i1OMRcTEMDYnsnQ+w4P
6tHV/zzyoLhHii7RdHrdFiN0Rx3ZFboXkYguL+3uJeoleH1GGlqn6kkMtew4tNmappICmtUL3v2e
fwPyeN27NJOTDR2WnPqHGRir4XdwwG7vzc2xwt1iSJf+E2WZvvfm1HtySXDaO2YIiAtxqYar/kie
KEvG/6Clv//NQepT5WFupNnZDyChZ/T2gRMGQul6q+dPC1GiNc8Bq3aGiuziok/pR2FUrCMlTai1
liu5CC76vlpJE7qh72GDVvaI2vzXicHN6cFw/eVNNcf2TnXVHLzxnDr9jgx/RKG4YSAc/q56rJgR
VsMEZbXGyWkZDNiRig3dHSqdnxyR5C1eDmteflz/1kedpwe7MyCsQ22iXgLKsZYG5cVLbiPS5eDh
4FLJgNMpqIkw6SZCQB/4tBslg9QKE+ru5acaRJmrJ3rgnQ+dhLRI5VXHUpwfIamFPdM82Pi/0WCN
9A9K65oXGqmReoR54cipI5aiSKtHA7mZj36xF5gUQ8xrPUn/4Ma67TAvgopiZKD64Rm/FvKwnB/c
iBJQj9zL15Q0y18CMH+bLoWEvVWG4xv/uWDLHyFLXmwKgP6xDmjQ3uQtKaY4TPjcfo5oPmqt965N
rwajbGXPknKIOby1DH8DDY6/i0eLdDNzDblXLa01gNjoO1Ph9j3oadMHaWTsMpUxgWz1UQH0QIzb
h13gC7oVwACNC56453WpBpvlhVDdyHXBOLFpyFx3V1mQG0YE5DtZ2n/dliCxSJhtonqXYa/hB2WL
lD0Ve0JDb16ZqhckqC8MrsLNAWHpqf9FFj3OrxjSKPLSYd4V6ey4BnF4i7UmKvjxfmpykzVHmV7f
vv5p7d/I3PKInZwNumZ9zrCxxh85qEG9a1QxqeKzPn5Nfxw+HShXm4Gag2OhImDAK9raqRLAQg6X
KJx526PJsmX3Y7Dg+pUpsyfWZSRmnJJQqGGql8vnDkShKxWSj+LO3Sin+kLmfQVyjYRE02Xq0JU2
CaqwL7XPTrnKs9LKsHDsKSs/PA8HCFzwbsBCfjh6ORVsCTP/lID7U+IIRB7rsAeHs+oukOdt3zjT
3xE+gyivsECH7zNNNZ9DW7LbkdcUL2gVNzVch0LiC4hJAxjrn/KenLjnAKsZjd+0rQgV1Fr9Mpos
ZzD74F2LHKBCSTEmcTcT8xLHHacm8NVDfD5WMs3y6KeU+2XH+iRH2nddtFhxdnDkW190vtxuE/iq
FCpJ4ChpsWGt3MMnMWXQ9Y2y3ylpuSQlzLYy0H5rSYg8aLDeYstTFDFb98nKUmugwDreB0tUV6YE
Jqdf5TOgU/po9K183z3KjKG/O78H+c5BPET9Q0UsHwfLH5OPIBBhtT6E3eZRsb68t1FnE2Tvtq2c
nI2pxRZFZMyqNK2r9Xu/Y7YD23ET9IWFXZElHx1cyfD/S54YHDcZ4UMMYj6dvVpxYW22U4HX447k
ATHp0FDJDwyIWMVDOo5GL2mRGo+nmixyrTouRu6vAd0VBB9wHm2jR99XBAUnZBJcMFWsHgx+/rTK
ZOHJAbHSUW07hb+Vg7JxrctqZXbYqjwju/Nvr50gc5xUdKZ6dg+QKTPgHbWPP/zTnYByDFuLgb15
1YEwc0xAkjgzyEy0Li0fSR6r4mC+NQj1Yqrv0V4ZtjNRys3oPvCxxgyIZ48fSwqnFjz13yQOwLC2
vOQdsR+yPbGKusNB3M161g1kqc6KJdxGU3M9l6LhmybtKu7dFBIpx+zkjXUSrbujsDrrPkp5Qz90
Cod9zDmGA1wyNWH8K95Rmcj5uBFt5qXXW67TFnkJGdVN7LEZlqAOVPN/jHZ34bPm8dNVq67U1xXA
pqSrBUvmau4ZBFtWnRIVl5rDb8PnsnLe3dlSQKrA46ce/BcH5/FxPGte9pnq4eIB9RuJZ/1tW01D
Qom+AQSgY0pBHUKb6k622Oz6rPnxq/zaNSAf+CGZncm3lT52NT7il0QDYK/dpqmg7Pw7ve70Ibje
RJFeqaGXmlhadE/sPM8PyItbgY+duwj6QMEwbTWTdE6pTpWCdagJeDz8fX1eRHGl9r1Ud3p+XCnk
iEgcpx9KjK/dU6CKIgwE58fBxCnZhNZVRlpNDHavQrxcx/MS8gRGj5IFfZJPsnb0r0PeG30wYksz
P+dxrIdtvEAguhKeJchufdBssxqSC4AuRxlWSrWfo3N9Is2iD4U9zkznaILwuNwxyC/935olQsEe
U4EdWCt1X5fMo8LhMhybnvbwGQE/n3SZ0s4lJn8nVIL1zZFIRTMQcDyNO5vj17Hzx4sqVdLbn+s+
Q/NOHXqpp0E94/7QSUwv+POZc1OZh1Gq549KUif76MhypKXuuT/z0p6j/s5FVgmAuGm1I6gKpexQ
CbwJ/WI8m0vBhgAvNE9V/orMsvosLuVkF9pCuujxkO2Ky5sCUHW+f7dgrbdNAVFFxDLXtSh8Ws5q
TmMRA68Hy/G+Fuql32qvDqCieyfGe4GFCVK0J+UJNKYdfTaD8WY8ya7FuZWDeBYdUdhQrOHz2oHj
QkxoM7jD9eeoQEYdgegf3LGJun6pD/68ZpqsSG9XRSXE0WJuiylIEvrikf4XKP7xGp7uDi1ZLq+/
LjqxKTDVbfzbFPKVV+tlocDfJ3FNSShojWZyTTcMrHL8Gu/phXNOcW1+Ez1mNagW/e2Mbqc/5eh1
8pRlxCvtUBMFAyXfm3lh43j10t5VJpJYEBxdWwTRgPVYPTOm+EPXWRzaPu8mDEJ6XFWEzHesz6vy
LDmkEv6WW9aSd6SiauxdQ4dTk8M8QP6gWMKlZCApB2vekf8S92JlmyBszIHgYe8j51uVxSn2Yq8M
B9YtVfVtnJMhM91mUHO9rGUeil4ZYm69mOMKXJDPda7SHm9sGrnlCqDXOH2jJ7hXuqZ9G9qT5mQp
28G41IM5Sm7OrzDpORA1dfljOg2mDzxa0O8FzuNNgkrgrLY7ambqUKCV8nsG7K/6d4JezDUetdd/
BhpXmJ22UyvodkhJu9jcr1gOdBqhuvcNCDXx91T1qo8SODBg5eIVL5cNlB/Ue2+taDrTX76//Rhc
dQFs1QLipHbEplq2gRDp52ZZ/DX7e0Dk1Nr7JbpqDRjgFi7feydT22L/Plc/XU5Xn+VkYH90bS30
G5VkHdPuZ554qGtg5jSzYy/QrJ3Bbm877xU/x+VWhc0ogk6vF5GhsOA50XxVNZeng1OxoJlwz2CT
QriO4UtZc1wbxPewEdHDCU5f5J8BNmo2Ykc9Q3s22KBBKRUCgaBW3AcYJCakW55ZD3vQ+pOb7QAw
ax/3M9uYc2pC6VZNUUFmIdVFOHGMI2G/iUjpiLps0ktIQg12+IA7xKIOT1AlbtaVvoAOBDWBL3ye
MzKunN4rgm53+dzAJ1EbjO02P80EXGkO6rgCsgCxm2N/AxpxTQ2NhGHJRfGvphJfYNc4YUsl1t4o
f11bF6NnhCbLtv86f5LxEaGHk1XpbUIdhZHrpEKpr3T8wNXFaco66lQr9TR9IvzCU+Rz6v/vo2TO
bYxqAtnVPa5+Q7t2I1NBx0NB8+yud5G4GZhfZeSDxqUBpqmO+RlNBYT0qq8t8LcYGTovwhCo26JX
031GuuJXcclPne3UGCvC12FjKXYDEnlsufg5Usn8xaWWrdjtH9jxOV91RfbpvXQoE8EtsmE7sm9a
ZvfKfpUCGyS9r+fnbF4msn3fYTEB1eqfEDArmrb+hkCV+clxkGKZBjbtkEtFYBO7G5qDwuV0xJBM
uNfPXdsLuLIy5hMtCbVXFSwr7uofEjlyZsulzpV0fiQA/MQKPVrrlirHn939CoWCvez353s7BXon
fG22QdF5XdQ5eBQ8keN4Jk2lZ7c7cGKIiGYmCTBGjXoZ/hUwRNQZOudUeh5LzxQLGqTnwpCgIj+5
mzkP3xP/VETazg09g8YSku49rlu2g0byus19AgIQ1MpNQ5qqpcFF4ySc64eeXKiZaeItAkLRaOZw
nPNZMwnEOOjZQq/lrv8jBNq9e+OGNGBPlnZvbJpSG4VGHJsJbAYsub8KMLfYnay1Ij3mV0kqKBcB
WcdIKZ1v9kRmK9EqTqlm3DqrcTd5b67wkhepAvlAHeHg2fApGsgqYAPneBJhXeZkCeC99jGDpLhh
FXmgg28cD2mOX4w1AQjR4Hg6M1xrTvTpi6NHNQhblHyjuezfiLyXsp/D7JN0V91FqT0VzkvH704P
l4MBM4kPV3zPSk3Z3OHpx/aaWFM7CSFSCkewvpLb8NdRQbEks23BSk22dTbdhuLKPyRF+xv0FZgi
4sGL4gR0HZRu9EJsELxCtdQZMyKxSZL5HOZKm4l97zqhAU00l5rEIYsrGK5zxwDbyy8ESNYTQvBt
OAtzaxWFrACMkxdDI39XlJF9OuH3F7Qj9jz181blEIbT3IsjYVnXZgD7sBwRUF4rO791pTBLQgWa
NVc5UbZ9BA6KW7NUIS+wHY573kjS21jj+GyFtgWMGM+14SghyD7k8sKmNNmvbvAB/DaTiebJiWxQ
0cLYn4lO8iVSr0uCCLV+6JOapxfJi8R9+UPsRE/iSs3Cbv1VVQ72cqdOCQ3UUmifBkPBKtIAcP12
zo+qQOfKbWS+73IpdFbvFeN6if37h7oXjGEhFnYg62Xu//tkAfCLiLf+UQ+hG5NvWOPnTTUqFGs0
sL4ADwvZsYzGUwfAKp8bFH8ZkXNdA3VHsn1tXnqa0Oi7A1QC5UrfkyQE22pMOxL0z0SDIYPQm31N
jgGAqNis766gLNXe7bCXtMuXScpJty/wzGlEMlpu1wOozOoT5DuPiSreIsTFZVz/Atz5VWQas0VA
KTTg5bW13ETgwlGAPYCdzO4XGI1gYsTqVIqy/JPUdVpUgqaYOWo7cf0cxnLTfiOtsm0iMIY+a8GH
XPv+I4q7ZgfAi6tkMBnw7G4gkGfTz/dIqhZyrfFA79DOgFHXClpqTDw7Illj6pcQIk5HA+2d6FsV
/t1inrgtw9YDjKicwUeNiT1H8LihBp3cwUL9qlAozVBUpu1byftxsxJjFrN8cIMNGLgXafL8Nr4c
eL8clr0lNA7mC1rbt2Yq1kcL0VRoJ7/EPi1TyEODz3YdZ65FPq/mUOJHPJ+8XUN07UId0vOetpQK
whqJYa9RyRoCIuRNKVBixrlE6wSdR/P34mI+Nqar8INqXR5MamgEkyntUIfY8qUuGzy5d+nbC96F
FHLDNjiBBnzjWdInEjsUNSRvaHL+rXVVTz3DKR53rz368x04EEzsMv1NpG5r/NE9Ibt71C7Is+Kw
0zlVDAFglGoVxnkytMZ2Net8RSA9Dbk0l4GVXToaXoWKFTFmtzY99KLU7gbm8N7Nyi9tfIzmHIf6
OS33LRdHPF021np4O3u9Ak1YpK5fYmEd7RgpqchbDSdyZFS5M/Dk/PYmkFxpPHdYdZ/i9GTByKIv
czCnuZqCJaZwCUHQBmzk2Zk2aH6I+IJo2W+PmsEZx3oxAyGSwS4ZEIeaHeHB/SjG+fDJx3MRNamd
dgi54B+ZcKJNBCqjaoLrDlcKusk8F1TjEx5MRCujZtQCSmUP0kJKSudTGk/WLG9tGfLHBPVJO/jL
hBu0RvIWNjH5svrQ6FnjdF/BP4UdPFFzihBy6BpyweLY/1kTVgkphI4ntXtJoJaamXrMIvg9v+c4
uU7HeXsAuvOlgettWOe77zGN10di3q+FsN4ZmynRmZRM7f6HXZTA6AHFylrtqQazg9deW3F5iUSR
l+W9KkFwCeyFZDSiOjdXgAcH5kWA/DzL8mn7a1D8Sk4AcEgKWKwwojUDVONRkTjov6LFZPhAvr7M
XbPSI6lgAlZGJCQJfex1psdaTEAYQyCdpVrKC9CA+YMu9790x3TZnpQ2HAT/RVhXw8k/YkIiaADZ
hFG8Zsx2ZFRxEJmg7iQ6Xhzyxqfp0GDHpm6S9dngK+z1WIoQdBYyWFizf41XMDEzG60kwyEMxkw1
qj6nKhdRuf/2UFacJQhMaAbti0+59+OPW/vevHCpANMKMEctRuG9bdqJMQaMRvWLzNbdah9BpHHJ
Vz5Kr+6HPLQklGXb43uh3aWkg5d4Sr/oTPRdznRNXNVOCZb7gYgb3LyOLRwnqdCvRZYk7cX3ReM9
plYxcTGQ3MHdJtJtNUwLoEW+77GQ58Ht8qlhRKRJO5bjzpmXx//B1CgWgKVqcy7CT1ZiaERqllwS
3pcZcdA7X/u+gbChg9W51xq5oGx/xjpeoqn0HRiYcchE471Q+o9s67wy2bk/S6CcvmF2EtukxNSC
dVk7kGfuWAx8IX8YKCc+aKoCYxCgxmuOgT/g25Eqii0PlyKGJfDtDd3NRffSPRMRSeI/zrPfbn9T
JKrQwJwq3GyiubiiajndPOz9i0RuU3WGS056UHBN/30mW0CIp1OuaGpXfdMzD+B4o1UGMuJBouUq
vvMa67cNtme5TFAN7ZJbR0uCw+c0joDi2s4HIRR8RXXu4yegJNFjQBSHCgGoFcatZcBJ2dxbAsY5
tJOcbTB9prMvGTMe+WZs9lHi3GHeouXvAOoWJDhZFzwKx1EbdT6tDx91SEuwOqPOCuRn5NpqHSIF
8Gib8g4Wmcnu1zKFUC2Ib4nQWOcjD3xIN0YaiecBRXSt6hxvOox/s1rWJTUkG4UGkRw+xuZUolto
QJx5tYF7Y1dYGCjYpHmq2YDiyROOZvn1jF1xk8oy54IWjWNbEylrqFX2UX6J3hsZOt4I7adYqazA
vyeeTrAks965Okc1pYdCPDOtubGd0TpHTnuzvd4p2xO+3oKr8KN2eTr6uQSiwQmmYZLcboo+0IgZ
jRAHmu0bLHog8nTnY3utXvqXd8x5YlxUayXG2/q9hgk5VSYDxrcvDWHj3L8My1k8VQJ4r9BHbnA5
R9PaiUQZ7quZdQg7hQcJ9M+YIlxPKOI1r/CuKrFoB5YWbDZwj/TjUn2IMRPVA3atd0MW2A/26upp
iHrgJBAMNdXlRST0L5rzjMhi0OH0wpJaKvk70t5wgYiezag+mv2qQZ7Z0RDIU/O0wJm6fd/Cv+Q+
DXYQ+ofkMcXPcFIso7IhqCVOriCFcWANn5TP+nJWMtpbfjzccRqLEkCtOfok+YfSADpMEKHNNLP3
iE3TEPnr+KvEjJZKt6ZMuwYKqfbScgiUxgRiWzxxwNX1iTDJUjA/6yytpsBjqFyleRHgL3YVMpHo
jmQuCCEOwOS1+nLzYgw/0vLxqAHBbJ1T8StaIquI+e5AeHdk7LnvPPowMpjm+2Qz8VO7MRmfeQ4+
8QTHs1l9S/TJx39JkUirb0zdufW5mRqBF8SzhQ1CFhARuBuB/RJlA/abxiExfsnPVXOAtZJxlzNO
j9WJgWVYAah9QQJdiBsD8V59NpPf4BH3QrG6ipEyw5YXyfYGQPFYtaQsEPLap7D69o6HXacMrz6U
YEUQPiH34b80KMCdEDiGU2BKevAumuXQNg9W1lH2xeI71tbKLVg6re5p5iRgiEORttKOYxkJzp/i
CfhPgbPE4DgnTFaV4fanPlcViACqmak7zlyMXIQpncC1ay8dZCxfCgwoj4/eqa/7z3UsHcxsNkND
jTCzDu443dD0mdzBw+wsxDM92kOc0yWJaH9FOJ/g705FRExF/U6igQ/2ZdH0VXXGAz1LZpAKMORk
JCgf4FKQUfKV1t+GbGtzpxbloxtoL98qVMXJqnNf5EdFPZqSJpGY5r1pcPmix0ID1yh3Ymd8mGRH
ySQOVbvjErRn6Gx0q+vC0OEA6JlJ1kZyQg4ZZrzvvyae6LKDt5iHR3KmW+JnDX7m0oVBDC6N/x4s
T8ZJnTdGRZ2XkvGz/zMWq54heEX/4fr5zoy0UoGYVN6gQ5ijuqNgLhyZRXXFwllESsCQ8egO6VQQ
qhkZrRC6hs3M9Qqowu8wGQxgpf0fHHB36pbomBicHcrRCNblgCm+/yNXMGYKn8vXiSFk73Pqx6jA
EGpluy9uHdBUHXHj1OrjR+8CJecbua6HIUcOZ1N1sD2fLK8MOMSX1oA8PJBAoEA6iYBgWK56xBFy
BUu2o5QN93EtGtxuB57f6cy4fd//4fheeZPBeTGNsCnkE++nZBfWnYGUZBIx0R3LOcjJNOwr0sED
F4gxLrTE/lNem7O97rLK7EYH5pPS4UZzSISZ/6cINv1gUS1k+b9QFAN5xPN1MrEyvKB0HM1orGWu
JV359nPGFStFk77lFBZ6nrHfH0fu6uY4y5CecWBERhn0Vexd3/uOBcMORGXuR5lrKT4CwhCRnEr5
fw/Ggk2yfTzQg4eZ2NkjFesYvdxMHQnLfWvGZTlQS5iHeV/NLKo1AEApYIEh4O5zaXSNOsmjKbs/
rHDgNL7J3QeBlLF8blwYHVwBj24QqLiQjOt/byhpKiaGd7gpEyR4a3cgiUNDdAwCGwVKbDNvGAb1
3D4h3r9LTfGE+OQnRvvXQZtJfBCYuHkG0w4KEf1DI+ygG9niwhiSLM17FqIMZIi75v6S75lvHyHk
3rvBSKMDRXo9bu+TcukUegoUXgX5q//j/81Jn48MKXqVr443WEHvjUfnyuyOGir33RQY9zFmhXaa
4BtOgtESDyf9ZyAYnQdoLdwWnz0BBqnE0eS0IwtxNuZ2Q9Mks0BlnklOd37pKLv8Bptf7D0xA7Ut
8XV0mt9IdmMhkCk8XEK3VQNRfEOfsnlcmzK5Bu6+kw8e1CKaFMDlAsiJzWYFfNGhTVYq77TqFSFB
j8kWiGMLf1r+hhqS47Vo6aaqkDBqwtdm1r+t1GJAaoJWGTtTHsXDl6xSJhQnlIExQuAbvMoh1UQ2
5kc28l62KkERddpvqxBAMCi2VxTv3Gv15PUvgxQbUyc+3TbQJOI1adQQXcIABTUDkeEXAxy/51AZ
LDp/iftr1tC/rRybGVwG4IXpcFr3HjfcFVPDgi8PFAypJ28zRag/mb/iidYhw9xIGtY39ZQhg/pJ
xujWaao0fi+cSNO07iq7DVr7aEJs7MFQpPI7lDnbj/wn/ZZvYtrS/1ThB8M6jIXIJDrxjPWLaZP9
M8p6rRLffHuwytphOsRZsuDg/0D5hOZpFKyKRQ1ymZQoqga33XT2BkxaDUuBg9064/yFyIJykyhD
cN+onhnLdp1JAMSx1YQldrrr8BX+myole3ay07mOZ/PdDYoRMycfXloc9KgtR8PBn/XBtCUWuLjL
un6sFdTf0SMo8/jjrUSZa++7p6beYCjVuTghZ7Hka99adfx08LxW4W+IDNdHKuxrYvHyC5VcCyd4
HAne4pv1GKBj5tdBmvSszsa2nAf0MEaW01ySfl5MJEHLUN0r6id8eom3gsi6bjz6R2PEUOrwX3Oj
X6xFDl2z26yQs4bhA7w6qv2CHq/iEb2dDuGut3XoLIv6KYaxZjkkolB40v96n4ijqiMHm33VgTVf
cJfKag6OHza3sEqPuWfU856kAim8DAcODRuv1rCU7Qvw2dSAhJJcsFLaBTunVTK7Bb6a6fTeh+Fx
+VGCBDpkD+fIwnSiZ8Y6g64IYgPraMNV3A8NUId3PyHmnnKTNVXRsv8SQyIukD6iNJxrTLqON2aq
hepMBWmueD3BuwI0Bx+Adsthif0SAGtKXwUVC4yg6mt5XSNExNHkkeytjO1+gZNZ11FAfZLuB7NC
OJngMwjPzZdIUei6t4NF++6xKD6Qvc2ar+6naLScHUZkXqiba5vMXYmLzXES2tkEcbbxZRGUix9x
HKySCBxTLpprSjRposRws9RbG3qP2IHd/6Sh2Wa1is7HUUBYujjrUoDyYda7t2gA6m8ji6lfhyJH
ci0UGvVQcYpe0XdonBXFy6lAgqB1iq+q6H1ZUlQw9wrXWVkj7kjNRkZbpbxXeujlL0o42ClzAm7F
mZ6HHPtM7uoVcBFp+NzxOCE75n6OJl2EQxyLRwSjzpK1FnRpjFsiiar70PtKWUMrhfG85CAi/cnx
GkIHsximhNgs4a8IoYQ6NClObHkEqI+p4Llr9cpfoq0rYP9Tn90I6Xu9d66SC3ZgVEbmadO4tBgl
azyZXRA+/Ytn28gjUibNB4wIs/sOdRDbs7ELW4GtISCav0fpm9DKF3hLVHI0pdTVyNL/fhn9WHm2
RHHadVXLUGbjXrPjAFZ5gSVa2DEAfHS3eE9j/cPDwjzm1lElk/bcRiBjJ5/93Nul41WPvSHfMYUJ
8OGTVVRDk3EpXGVRHJb0+g0+krz4NtFAxAaPbA/R2boGbCHSOG8+ZC3vPS8ua1SKvvrPLVVs4Trl
HGB1Sz6yLJ5v/au65eEvyb6s1pk0HGPU3L4iDB+CkzRHjfVHbwVs+/PznpomJUT3TdOENwT7FBgn
xwQOowUgrm2PFD2GsJUL80mB8etDWuksJVZMFamyt7hy8U8+W/Z539ExooBQ/Xc/uAW+yJuQRGoe
a1bP1IwhDt4OctvQtrWkFjR0TKZhAkf7MYvJ9wEiXXueu9AeGbbd+c+UGeiMFzcGplzkkouVUMFh
O4xfSywEM1VafIi2mG6G+2T1XymcUN+huezt+aF5wtaeDuPwJN/5yJIdNk8IIlo69dxKgyxTF+Hd
nGaa5s/YvsqXnsJEdjXPeNL8tB2rlv8ToO6Mu3KaA4E0XiUVMba6TB1ZyQRK9XDtR1tGTbd/oPAv
S9gMCwdNEgInT4PNcWwphCe2OylYgexNxFPqfa5mXclTM+TQAVgNSle2s/tcF6z/MgtUqkvkZ0Q5
uofJxurqdht0IEps+lMd3fGew8U7Tx1AHB+HmOzB25p+U7UYkujmiGdnEsvIBS6ucsFPttiwnsO7
P3q9rvRxD/zvheTK4WfOVEWrULiSBE3RXZ2giinkUNcNwfTAVkuP+0E9fFCS4FM6cSwOn278aOV/
sQEY6B8RlxyAB9m7lpr7ldD67w0oQ4r1ej2tMXFHXDnB3HhlU/zPMFrja6It4RLvM5jDxgey6PSX
Oe4fpD5MTBOignD79kjLnEkHoY1DqO9wFieiBLLU3tmEZ2f6FDikJz+RV8Xj4KwO3+M8fCfSA5E6
Q5omVNHitaxiBtcB/Ky7sREq8xsWiRzcaKClMNNv80x2LmP5+I9XIc+49cmPT9fWyguyUfdmBWMx
DtES+R0yH3sezvJSApDy9F/4MPuZFwY4c3s2nQyS8FNdhmRDtkeiIHEYI95D0iaAewKjX3cA/S2G
IvwD7uAz1KyNz+TN8U5brh+LHY5hP6hk7ZKY0PJIaZQypz4JhC6m8GZWxMhwwfs+FRzqttOKzWf7
+92D7aLc+0cyFNTn9MSDSgl3KTw6HEfmwN9x3ocYy+9v0djYhO9Si7lUiYDFr1TasusxcaYg3X/K
wcXVdhDZ0T9eD/EBfq/hE/w7OJ0ONrNRp2xblFYsOBf8AoMrTetTNRtdz5QqA8tLqxqnh7hP1htU
/LtpxRqlhas3CRTxcg3GYyeG2xGQddm1t4R0fpFI3EgbB05pg6Zul1msLSZmXO9MlAvqoLEjYjWJ
TCF2vUNeI5KtT2Ce6FM+Iy2oLvv9FLyrEvhGTpNO6eM+cW8Z3c0pIF4oNJFIA22mWUrdzfrjtNAr
4sVjmJUlTd+LZ2Kt2NpfvG0gnRGHxJwsOvcenLdg02pQ5B/FHAcW2Hgazt4e0aIFNA2gTW6oylLh
LnRD1b0CPIGjOzXgJHmIPvh3K1dox6DhypMNSIEVU/lcE9HgOzz0dwFtWvEA4H5pT55F/Pko8J7R
v2POa5iAw95xQktMugb0ElW8B8KeVoysPWfTCvBcV2YW7Wkh1EUvmRUEpBNTC89COvW7H2Qtdd7t
aclokvdVROUcFG/m5IBImWIfH8/se2KCndC1KhbPPX2v64i1aNVioHCTXARpW92WK4z9RAmKm4yZ
uL8vIqNFIWmmp9WxEyYW+Q/jt420poTSpcrxPx1CniPkeCEKjJo/mpgWfH+sni53tHTmFmsPEAdH
8HViRafVWFWZjk1EyWkLf+Qb6Tc4ScXABECwpS8Kmrz69simmZ2am0N4mN8oLKa442HymuBwdjrm
ChgH0mqLUNfurYUTiKHFWA7wSzFpPwYhe76WDS3GoahCxc5eZaEyL5hSoWLxsDQq8YZt6ND25FPW
Q8J+hgkjmVcYjoakQC3szwFkoUoC95qs5tBRkhfijxJqNWv7r4rMc/yigDWHo4wo+91n1OTwpOpM
wHLN47kTfdki4BCv4pXses8IXlzcqMDxmwJpFWtE8sBOZuCJcE1nJBOM0YDCUCAoaOoTFGqjysKt
35LSOE+nL6lHoe2tQIwolJGZTDSwiweLilptVlWXrgW2+wfJRAZb2KYkxSqOfy+E8f9bR29SHLLc
Zib/NXNXrZ1hKOSFEKIr0uPVk0TyI18sTbZ6pemPhH2Z92+x0vjaoJvBTzEcAjElWytyzlL+9Y8R
W0k2h/C3bNWpMOUrQNI8k82d3Hm1YI/rI3qVG+fVzG7qkLlvHTNQ0OcJzA95azdzXPz+BQyfcW5o
GAqfXCeVMR5dYH+3X67mst+YjqdgpPdXVTkqq7lKxeqxD6lVyCJhCQeN1ABB6SwaUbEnMXlZ1svh
s6XZw1us88+QKaDZs2xy62maA2F5MqCtYCGmAQTxBW8dh8rOuVOpE9nqwNXH6A2Xa8GBKkYTIW3K
l5yNoIEP3Yy9X9n+rv3yiCWkqZ7eC8lFpwCtlGVqt2Wid1dbDPZOefBAinkSw05GkCe0EFba2i84
CzpFimGQYEVkfqSryG61KtbwB1ze8B6aDSB7Uf2bcNUBItyBk4g3xnJBanURxbKhCsEb7ZpRiMb1
ZYDSpzjRFw2aLzLjBlyllMr8JStZsHuCPaeEWdoUA2LK9iposvWXte7lnmtSlp4MOl5xYrKemNuT
Qudqcvm9+6snJM2+fgX9XfVh8aOgc2e8DTNDPBjrMAEjLCq8dPVMrGaZXGJI/09+0KpRRxWDeXsB
99aNypX/jYy9ASBlrOlArzzOatiH8GmRvyN1ehvcEGGv1naRyT+UFwV3sPiddFKDfBVhnbb6YO9b
OQxZVz+Cz5BOMN5r9pUcGthqmZtgyrx3uIedYrJzRKn9bJIZPeTxRMJrSlLDDDT/eZJ2KAWLMZHf
zjTH4xYBU6UfbzsGPIEiw9Q1qa8vCyWgNBdwBUvbYC/dVKu40Qgdam58cS1ThWvq2vDDBAzoorDR
8hunhAWwGONjTbTKTWAYY5MpHTNBL4yfFMDcl7vrIXvJrNOnUn0TQw03L9ezIav+nfiA1hD0v6Ud
Bdxy+cBTPjJlRSMTPwtn7ShpVf+ahPo2CcaB+IlwtUbQZYFvpdyxBzjdo1SBVEL5o+qd0e9ADdLf
udUbI/oLu230/L2ZHaC2XLl/QwoP7E4a+V5JkEodtGeAqi+f7Ybdy07irBmKKas4QEv38bre+R11
2VbFWRwtiAayID67XyXWLvaky78TR40qVtEt3wJniHlehHROivGaAYr+r04vijBnWdLmvL7uqHh7
vjwCw4l2W5eJ/d+cdE8HVCb0irgnlL1Qyov28hYX5fecobLMl9o+4BCD2BC/M6MJxeBkdut4gmoL
Doik+0A3LISABa0mSmAQoLBm7cCbiAz2YmgwVDWieqj/srY58XLgZUCGAM6Oi7SCuybooTRavWwJ
ODjnjru4/DlGi4wdVdUVKovpun7AusUMlvCfE01g5rYj4vrI6cN3lpfUfm/LsIkpiMFaxH45R00J
ky68VV3qLuQKmn26swWXpK9tXIvMpbB1+rQTHk4eyjym2sYGshMX0l2RCEJMWAAYbTQUinPahlh0
L/jSCIx/1cLUcFS+Ysix15ld3eJuTjR1d7sLx3JNPikBPMiMCYoQiOHDv66+Ne4rl8CebGLPnCjl
JtDFW82tbGsvfx7WDD6HZ4YVdEuYNPyG9+mmwStju5NuOZHVklOTfbMQgK972Gzz55XEz7XM9aXG
2CH905OWLKItSt1bwOXviAuVI+8gdLDumyvZAQfyapv8qFl/QiYukl0Mznlwm5wl0U4koD/lkFm7
B6CMdbZgs6ZvZz1M2OHzKcwo48iFl5y+ms2BtuH4+atpR8NDOneQlOxE9qYBwvBbE+jraVJ1lBbq
XwNac3bMFhrRlUvA5SkpYM0c4zS4KoT7XKVcfc0Gu6xUmYq6+ZZ3O4fiNDCCDKqHJbHFPSgQlRMV
Pdu/70HBLRQNrvm8vsgCGu+Z3Zz75aZhIFyacyCb70VNLo8FJQMzxMmWMzXl2aCO/dZI1ynJQFMJ
Uv4QRaHPpV3xjYPj6jqR78Uef4yARmgta+MG2qqrBYo1h853BZJ7GM5UroAW5NANQKMakhCl1Uzn
6zeVxiBpfCOOF7qYHpnqN+D/a5xelI504dwDRUp0SgQ9o+uZyETalg11zBD4JvCxgfCokaKHpoZB
u4x6LTqEI7luqU7WGqx5TOxiRytc3OXu1Dt2/9Ex4O71bxZMDaGrPoDv98ukFwcNUVr4SZn0GnmU
Whfkhqc/tz4hbh2xpFK6EdanTj78K/M7V/pr1G63wIi+0yvC15sS74UIbramjGqSJZHAqNctOc0g
TNs8yV5aWuEnMwN1FMYOnJNN36cQ83MeZirzfwNvjmT52wtGmC2SelW8aDPRbamxW092/QP6S4QT
GMINMDqEymQMmpRLhVmdSbd9zQd3Yzlf95S1nS1bHnBrOSOIB5Mw1VUETE0qv0MnEMjS0okAGEUQ
HWt5y3vl91juG3XKs0WyaTd7nLTXu6L73IDzvWF2Krwu5ZNaXTCfGb+SAedOU6H99k2/A/mP9Vfg
H6/XLY+ExnlqMrPCZ+FRob5JTXaafZn9d4j7wzNMMTjUZHzDwu/eji8JBqTowDj/6IPvd2ds7Stw
F72O9bX/sE1kwMlzb3t8y9IIu9N63TiaFMHm09pz4aVA+i/RHK0IAo7G6wq32AE07m3vrMcmgBvv
rcTqXBqr/VrFxUeanRA0GIJsMI2XxG6vo7wuiILosJkTPpNaCj1dHyOXsoDm2mkGbap97lehPqvV
pp44KIQQ1tqGm43LBEQ6iTDDZjLFormGCSfYRJ2Udgsqp+GACjDWoshjjS8tCUBUOccEsT7DL1T7
NQjDeNWY7CaaOLt/rjHdyohyBnKh56Oa1RqEUte6VROWGtQIfuQeKG+3Lv9UQyebyYto3Q0EvfVg
JYcgrYY7eLaEP7AUIHQZFa223YnxZ++rFaK/UA+N0jm4y2WVpMmeiKO3N0q0KEiosrM/2gLTYjCe
VK755XV/iIkjxg7mCqONXEMAnNphdWUAyzg75X3Alg+M851ZaKukwas8dW7RMibAm3ItZhFLZrhc
E/BcTnJ2jLeA841B2+5R5lw/Bf2sGFOKhyAdBuYXn6vmEtultuVoz/hQ255WAZ2wgFL6qjw7JY9U
2jvh3qZYuD4YrOc8IdFZMLNyRNd9c9dkf5DZkf82kqdNrqLQ3Ax7WPGXYWgzc10UmnTwPlwsSDY7
Puibd6JImxDOTD2srpAbKPPpJIAopVe7Or67gL/4u/j/XRQ5SxAZY5U7GL0m3g2hzxnxwBd4jOGD
nRY9fn7QItFdEG8onnzMUGhNP/EGreR+LWm8dxjM7dxSq4R77cGCLk2JSzWET4RgVVq+qRZ3V3Gw
xGH4GJS/m7WEX8V2fYfQHucQl60N/nR88xNd2Eky/Em18sVPXS7fVlt2AoJ5+cT8Yy9gnskgDlj7
gMfEweBtPNtVuLHjsiKjjjWb8CcyREQhExd6lWmFWzA8uqu2q8+6Vsqaruh67SkwUe7d3lItKf+4
OeInxrI8E42r2WJi0qptSlVIaHRCRwagJsbV9j3Gpd5iL6NnZ468Bjc8e3SP5kQkT3EGdiFaNef+
BLAAR112UN/rcDok8Fwm8rY6JehnDpPiM4vcMLeFyZo5O1TwO7D5EqKS8SF+PeICjoyH9kniMKdg
ZJ3+dX/5P7wKtGVPDL1rahKzKbGDEIl0iTX+SEBNflCIJ/vLPmPd9X1gphZR3z0aHXVwj21/7IM0
PC+EzeABUCZ8wFk+hTPZjTlpYNrSAjCxfiJLhLgi99HL0IfKe41FytBd//DDt59jywXMhTVQztOT
Ov3pXY2QlKkU2z/62hiHVZrbdB/13pVo0CaB8sZXrbGbqYimvNlbfrOqP+A1xWNtW1GXngM9KAJk
scYfhdOHyDfaQPzXCJee6/capgqn+rH7vCV7ckKtO/2F9rRN0m4EZmbevadVFgxtwntrJCw2epnE
/pPs2vf/IB5nLj7+pcBTHlDjjFN9pKS0xry+glO3N6MMdnXNgdvZQs/76gpUtOEQV127qHnpgccB
MEoQVVZ5zXbePYOwBSwUs1LtO4hmVB4Bqbz5+A0zwKoY3ZsWqTRGk+5WI+qhNdsJGKK/oJMTpXkU
aIOsGSyOvjh6d2gTcdCeCEz5TOGfbD0R0WeFxyTqOiVDS4lOFEoS92UOYIL03Oaumnpfq5rA1HNN
VnZd1Rc+DUSC23DfPv2+RwlXZBZK7ZDMghMULO6INu1ofi/nNP8Ypb0PrGZFSnDMb70AwmShm+d6
9vdgtAtjX6T/Vjyc0GSbPz9dTOas6IUp3BwQEC0COKmweccLIIEJ8dn4Bs1/bEuai0iww3e8+xbE
n4fM9dWsj6j09MMAKmISo9uNAwa06Rv7V7JKUjpnQQKsJJqOEJrnPVbND7JFwXZDDxpxKvwDW9/y
GA0UssouZcme5tTyU1QHr1KDrQfN0o7q2ce3CrkP1Ffx14olkb/fZ4IxK6xDxFpC+CwufN4H51QE
PryLYRVfN8Jgymd15TnJzEzYPjPRliltv4Awo7bwwYD9jsfGctCHVaNBSDja9PIVQsWoC7TEZ/7U
YuhhfdGtcAjgJ70eU6f+NsiNtP2Vd+AucfhravWZWr8bijlP/hDQgZIn8yiRAZvgCxQgdnlHxeds
P+mKMep6OoyVHdvHVkuQfpZDxziqrg3/VUupB/ioBEW2O0ZWpqDFbOIvlh4G/w5iEqtMXplgy78G
EMpUOCaDz5GrbWrWUDEGjxM1BZVkJX40JTFySato2mfmoFm4j3I5fc5cQj7t99vyWebniR2/7URG
9nDKzWiKJykpoSwBHYhmsVraT7yyQJU956/PE6qUeQgVj4HdKWH6RQ8bqwUehvkd9LqfWG5RoygM
98g/nPlvQE3Nxl7DiQOOq5Dgqrkm3AerxYSoXb5eBbH8MXG27uuYgpC4j1EDDq7bv0DVzxueVJ/T
KZv6zMoyvNuPHDsP/1rj5wNXU1UeE/dYrMzNv4njVucZZTjfuKdTh7zNOqBLyN8r2F1fSXVf3oQ6
9+6SBWTEYKZ3w5D7fNISCjhStmuv8xAeOaYGegZI77gxs9j19rF7Pq+DgCzES8kPWIB4tC+3cRWN
mCb3JgWpr7TQZ+PaRcMV/QNPKlhz3Xv1Ujylk1WyTbV4zGIDMeA7/kQSsidI/IUncIDqmjFvvrCP
RMwASzvlmgF2SSMg3sadpw/lirr5GzjYKDGZY2j+GUZZgOL7AMhE5BHY7/9x3Oa+myxGxrMoqBI+
c4Ta0ztE4DR7gVLLHE2qOh/JOH3Lpw2QsgGJl0gvquhRd2KjvZNmCqRTSvKsexv8jgZ26IzaCZ5o
WrZNLLjTFbke5qAfqgtO5aQ3xl5XZeIAiU2zp0w5FQYfuD55HllyNZQCszfpYtupbaQrATo/ykNQ
oWdhlbVJHoRpEpKkAxZNl3U6TtbkPscyZvKlerhNtK7hvJwqOOcQicrwr5kOsJdwUwwEYKP7Qtqg
AtFsJD7TjL+0zpSX7MZs638lDViDVCpzmOtvjzXihtFmVVkYIwr+L1C6Geu79RGbVtX8qfajHMVg
YG5iHKwV3mfDY6gWhvPI3/K7RDra+bKSu8o2t4XH0GxGcJHRnovnKx2ILNQs0RZdlRVDfxnaLNER
9tazXVJU+CypWj2qBHNKLc0ZSGDv/FLCDnEYnaqAP6OKPE/ZRR9nSyukVq9+YVIAkDXR/LEm0dqg
SfmStjaimivc/cT96z0CpsF8xBJcLq5JhSXq12X8NbJEjxlzLOqQ1S0uhvMUKsAM2d7UnAky98wz
VMBfxMzIPsmsQkhJGM0Y0Sz6OYZIIE/6rrOcGB0ONHI0ZX/imvJsoqPgcEQikUTk1rtrWyUn4aj/
oUn/Rz3UKzx1iBc6KK/LS5Q5k9g+7Q5t+DJ0L7y3MpbpHAazIW1t48VrYQGPDtfaayOd7kmtEEIq
fKa0M95OObFDC09VVZQ4cmiE6kwqSekpfrS9/4FwNGWDdSJo0lGYHfPgLG1M57T/eEyZAHDG8D8Z
y4g0SjPgYNw19Fz9OzWURbOmoMNZOEyXNF4izLv7bW+MJU7/4GhH6nvdCk3xDgRI7NHKn3ZGcngl
9bBETnaAzvm5LZw7T5wyM7wLZNsFV19awLtc93XHtx5TOcDoXoU+Gtw2XdP4z+XnL6HsIg+xMyGv
PEW9tVk2HWdLt4Zue/OXbeoIp7YVIL0ugidTXXP8NVQSJ/G8Nk+e6Ynahe436Ega+4ErHMj0LUjb
zJ4aSqdKfSfl6FG1qEyY2aspyCyF5QxW6wQlsi1XCGYX954K0A4Ud4dyMWrBxODaCoJ764Eyd+Nz
gVISu5naft8/JGSZ/bIfivUna5g/dvTaFIIOgjUwwLMp6zr4SwXrlR0RNJjuqg4TjcbzqMVcCmpD
XF4TpTSM89UTWSzAbhxsNeOWULnCkbsViM/EB6zx/ezoncNi+FfiG4cRePBTH1MJNiXQkKCiS0xU
1QXX/ISFXeeaT/ZXIE2D5DEx4UldcioRIxN9ok5Qug+rRYGhrnFtYShtrXob2x6hGYkVpGCz4ybO
Jgg3uElIUhE6MX+YAcUXuB/5of9j/ECkJawR05weSaJW2cZju1o8Cj2Q2pHVrCJ5SCzCI5nJhLY8
pNnHjdBPGmP5Uf7qUIz8FNpdUTnGDwwbTpzXw3buYRqHSsnhZGGenVkfdi7ke57RvAwb4fC6nToN
1egIpdkGbfKMofuK2M/oS8v2Mr6jDUkNlzg+p5dK4Xb5LbFO9VjEbAh8iGTJ9emOMh5ihSE9vPUm
keDXF68vhgilE3hLK63ZhTx+7zZwVY77Xb1NG1HeLku01pzBf9W5NIApt4PtRQeEafoaonyHKZox
hKjMAPIpWfXaq8PH09DZL1jZKAJ6t9LyXhpVFhgDuwaGcUbI+6TsPCd+cEQlaqPVR4SzZUWbFqKa
BX8HqYEQ5Lidk1jAlti6PbaSU9cpyTxpCpbPVHjblFSwlaAXVw1ucH9WGKjjtemSogoydVcGFSC9
xEaa6kz0bNUH/C9bkFlDkTb140YTBNR3u7KwC2MQyDkdZm/CUOZshGZix1X4FRAWfpNbZvm62pxI
Dm0tTWRv0AZwd+oPVbenWOUDYjuekIgSxo1BcpgdwgYGDbthnUApL9QMSmGZVuM1GgYqUYO2n/iI
OqLtX/56fgacR97s2+0ipFI+riJz1+1eMwQawkUhb9Cy+hxEO1NTD4cMp+8SDNOMXGM5ZSXTa+FG
DO0xEbHC5e17akq7SkTjLrrYPqMwWryuvp8X21yxFn4ap8AWQOa+tRNB8Nu0Wi9UgKQ79c4VfolL
v+KvX1iLfsOAXi14e7Nc+f+q931qRpMopfM6PbGK6OOCHDnAoPtewAYuvvllNm5HY1styH/bJiZt
7Krh8d9q2KV0IaI58lAZrFNdeb4BShiKm8sA3+8iPGrfZfajvz0f9S3oD+vxpRlIWfNeatZf+BKP
ZVHLBxCwtPULrA7dGTVjO5xl6wup3BD92Y+6epshuqC0XcDIhKRu6QqFwmky0+bD9veaP+JmIxS4
YDi0CQ0pJx3t1v8+fsCAH+WPu8SFAB9NkfIXx6Fk9u236VKAa4RK9Cp2TQdU+7KU5MecUfONkqS6
Wndi3t8JlxSB88BMu4iw8K+9alJcCAEnzJELftaFZoh3ZsoL8YjCXhEuKNrRvijfduZPoWMDtDao
S3LHIhRV5ZgUj+U+Xae6PJ9BAY6ZSItuPg6EUMPcGR2yP2kh199MzdfzPuEcHAKDpm//OcbPTtfa
Kme5NVtDfxsXH7FZ1VnbhDbfbkzu0EcY+KUSeH0LY6n2ol2ivB8A4ueiXoGW7BSLb5P9Jw2zgmWY
1QafJX5pgT4hROhoF7BJX/anta4bcPUbsl1dUV9mn8MObhwt3sbg6m+ycuxcg+NBmPlIrnxI4uOL
QPxL2kRk85fd94qIZdCV+j0b/V/acQHGgijC8TiRdKLOPglmqi02mOLp/enLtJTIOhPEg/ApP+VZ
Ftu3eVEnDmriYOi1PGcpVrxwi+qx7TSpP5NAomfQqR5NHxmotuHguHK9kGYFN7DKlOdiVGdSfKCb
KQiJzFXx66FHZQCBmSUjhvRfDKrMz2iH9QcYu/t6S5LmnEn50vw6h/cQEKWtJ9mqWN+trjTxvybe
X3ODAEJttgtvGrspo+FbFGD3FfRf7sdBuKlRUjNHCEwulO7g11dz3DXZ93dGLGVu3Pszbolh7tkA
IYI0utvWGQBGXikOHDCoc6/QHCnqgU56nQjkaTDXLs0yFushDxvidV2ojNn12ZFr+uOaSvIDjKFL
kgGK7wpIzFqx3CCEsPM8Do90YAhvdr/uJY8lXkyVhe0TCDOCSsNfe9XqLlMJPQjboptCM5ihgvjK
fCz0pW7XQe7kmr3Lowsor3Mda/LeIjMDJBc3tR9qVrYnju5QzygjHm8fZv1JmvhUiyH6zHXvORn+
u9tVOPev+7f9uwV/KD+nL19UHRPwQ/TvxrDqNAjeNptrINDZy6HIzQTRKsPPhdM7YGm99/foIja7
dhA0xqUqsSGlJes9M6KkJXquBZeoHq8Ez464HC9AJJaHuv7yz+/hDSxWMx0JsTTFk+ezzUZyx6TS
yUoFyFuiDdDqybgEG28prIusV+FD6gOVVmVtIYQpVEbzdFIxRvhKDlQkXNEe/pzL+jxpVD+joUCo
OY52pVQvUBuidwBkizvNWpBsF7LitWZ8vroBYunghSm0zjax5BeAY1AvgsO8yUCrL8PIQ5xU8jb/
CnZYUE3zVvUw0R5JTLrLoDqw4BrSxzzUgHtGakpF6hJ8QguZtBrPlAweYrP4ShMj4Sq9H9AaU92M
NvsmT8a1lc0B3fK7ioyVq+RP6c78Ag3xg39Te2ybej65PmSK+L2Nde2UR9/xgBy348tf6ROAnW0G
A9n4Toe62VeTvuIBDc/2Qw6ySWcm1QdbyuSWgtC2CQw5YgzgkdlAuAqZctLlM3LTM5K0YRGNof/b
g4pr11vfGvAsXh09uziXLMBn21VZCrV9T/Tck+IMqfiHXCA1uPunb6l+DBgUXlrW2BmOk2VbE8Wf
WeqdGMw2/9IMR6tllH2asgt1/Q0wGk0Q1VNBmLgydsBhjOwGuoTWY7qEobSH+6rpOK9e5xcR0ehj
MqoVoQ023z/STSBLe26Jiv01o6XbastEztNbMhoLumZb11OiPzywV2kHxpOr/A2jMu14un9VgpU6
sDpaS8pKwDKsFaNJsEfQhve+Go60owRCqXl8duCSvTgZwrQPD/WvYp89QkBry4+hxVcox1vMB1U1
6m1UPjt7ez6+8FXMVNfmW5pGxZfIIPwMtorRaPvEBKQlcyFcpXefLEVfS4JcKKLVf32jhPjYdgMz
jGi4+PJPU2vXekpD+tbel0/rveF+m0gmZc6xPZbU2dBkoU3wgU7Lnd2rAmNw3X1X7oqJ2SEy+aJL
uZ3Lwo4ZlxG3HSAs2/9xS4DNBcsSFhQXAfoyagpkKObr3ums43/vdnBwGi6QYxGP7xH843yZZZ+F
56a5TLv6QUXWHl40xY3O4K9LuxJeKvXlXblg/OKxqKmUzlsc5v6PF10C0+K5+hcIu1Zuk0r2RxrO
lRKd7SBNc6sLmDQxXAy9gfee6f362et+3Mr+4fkaK+FuMyyDzxYcBVIfDaSv+jKyRdFhnxM6Go62
OHz+rfGFbYuwymj9vYwuu01J+SLQO2abrUhH4INOCWPDNY34+ZXQ3SbmZ0xJI/9n6/tFE7uVDRVj
+bYVT+YVMEFo4VMDqEBANIH4cCIXjwcH7XFxn8lA8fSOTvl517CV2zmHemCdq8ZE6y2pcsrtultW
VV7KVh/WslAF5PpJ3jGcTIthpJ+VvKRhUOAoDZUcpsaOHVd4mWTSrP/HYo6WSx85rTi0YrHAkz5+
4zi+wQW/b5KPQHNRyKvaxibz1fgkoKZjU9mpjEM8UhC/H6TzJU9WuDpWqyTmgo+ACXXgSJD4j+MN
OnGBhJu2EHBtgINajWRsw6j02Du09KECoQPGpxIVjiqMmtfu1oFS37U5ADSa2/5Czpu4Aciv4E6X
NrLspDgkc7lsB7tQ6ps402P6KGdRsMmcr4mupZ4YTFWyTm2V1ZXMltDCqhFV4m1SajwYTmZjXJpp
2tcV+dsQtVGim16H0DPpZkD4geT2ennCT4iYAtsFurglhFNILs7kyS4fHxP9f7mhlHLCDwAV/dt9
n2jqHxFayEc2z7YRWd7abbMbrJwITa7uKjYch1rx5aipkV6s1Lif0sINrzezYyicnqFetbCplh8O
00vMRFtGut5CPZyM9cWKa6re/U6Aq79q2G+1WVOZB1538Um31h1ZYcWz42X1lPd3phZTGFwoOWFg
FsvR6MKN44ISG8r2f/k17mLb/ZLjBteBP4YCodquBxERvRJrkckKXw0ODZ7lCN7wgF0sNyFsOmkn
wqVSpGXj4+Is5yoCb/aYwnsXTua+lbymRSCRjNiU+DJMqH6/8ln2FkOtR3G6C4pKRcuR9XbMluy7
iE/ft0gnBcjE4v7rqm07qcYJ9ZsmEMnE8s4TX/a+vgxgiHGfGXg1V05j7ABndHnbzROMPbvXuPjN
maqcJ8QnfBT3FaQALkR8SlbawnbeKnSPSMPuzmhKfn9+aXhhqMIf1es21789wDA1NlN/c2cMpoP+
l5vycOkD6bLKkmb7jbk6KH+9ohIKeSOQJDn5+b4ClnuyfB0d4ceoQ2HA2golk3PG5+1qxCZUwgp5
hF/CVx1mYyJJuaDN3/1/RVzdOKHB5NlNAtOBlTSy52o+yVmQNSLbYqFo75CgSpeUyUklg0/LRc6d
JtpQsPDfGzgC85U07cmaVq01gmyoUbMxeum46apmRVxWmvhA8Q3YuOpzrgRTDROpVRrRARwqqDQj
CPa7zR+bQsOFL5o+3XrPEAUJKOZRlvrZwdKWLus4CmtXHe/rLA+FIDjekx9SYzgLF0XQcBdYhdOf
O9W1ldgSrvW2Ts5ct/ejfsnWeQC2JtARcPi0b0KfQ+IXIYVW5QG0pByIKfqSwsA/+DTFR9NrMnFx
ngl6v7pup4GP3iLO8WqZBIzQclPMp6bShprOBg/qwsLj/TATpvmT/j95fpF9nnT6MHt/8NdYndIY
T0rKu7Q7642o/rNZEJsZ0gFthLaubWIZtejw+k2cGAspCa5U/TJJe72jv3Z301a1W07ve440UJlQ
koOT2Er1HoJ5b82dBp5uM4+wvkxBdvX6srLfAWqZSaQ8o93kyPCMRo42raKybO3ON8obZJLu6wN0
83RAWa5JrScILCX4XLnL1LV6uMCMOqGh2jXv/P9h7tZ0HHW7+p6wpQdeLo2mSCZE2ZaqVWRq/Ntu
8CV0r32WO/jXEMAr1UZGc3u0ixVF1z1QcMWvstuxwQ6MmLkaSlHTWeMXSQRHBzCbh5Vs6lJdrJdj
hwbCN9mKnkwoVJ2iV9fsjWsKYmQY4aJOf7Tk/rSXy77j1975Xh9m+frwAMwbwvXnoDg7xwdlgHM4
FZmYKEcgho6K8xzhdDlptJ4oT9SVML/S6vfScKlPqQXgXvlL+raDmbAAL+gscOrGeDp9onD4QUmC
Tc2ZgVZt3pjNf3v8+SapCyiwWKRpGHZ7G26j+7k26reNWjXzkYhmh3EdS2V96pTFwxJ91lOZPpD1
7CnQBAPMNie6ScxW808WxQdxk2SZwv7QtOCTmzeE5hkJB0bwWiUC1Mu/KtWaRLIrGQpeu7J4J1JK
J9eVZ13gJPMFL6QiIwdClbJ4W3IwpW9E5p9LzUvZSfOnRNkFE1GsxHOn8kye90Uga7UwiCWFdeHC
Atysaf9S7gQ3gKIXLHjoy8GkysEXH5d4TJ7NBOOPTtndp3zwkcUR4Lz58tftZW/L31eE8zEp7NQ6
+zg3M4mnAKb0Fu7sU4qffDQOWixh9cbOR1CX8/PWEWKQbxzlRGkA4um/+rjyu4sSxeFQX96zY7ws
N/Focue5PvI2BIX8fRMtMZAxHHUwtnAsz8NTeEaJz3abIMon81Eqw1u9iJPg3+ho2b9/BZDcbgkj
Zi93ZgxK2DMaRag/TrAdodSOA9Rq4Yw6Vh2xY0lJFF+F25Sh5BLIzRzdHRmm4njxmDplo4+pzy3I
12KO+mEwcGEQJPIlZ+9zPQezpqTVKRNeZF2s1Te88ysb0K7xAV7VXKcsTD3VHkAbLvIzkL84LoQH
sfrV2IE3hrYzHukdks1FOi1W34MS/dOZa19Xfj1thDNc1lSbN7ygDx9gOFFmj+Jbqb2PnMG21i+s
ANNngH12BYZv+2eVISI/icwO8eNCTAleYZshirx/bb4P/qhrcld2+1GVT2Ys2d+qW3iuBjSPrbvp
xjBXdjJ2LLC0KFvIW7IHG8dz3LGbwJId4gZ2Y0Fy/yVVwLiI9hZaGs3PWKvnqq21UBWzvHpDg64E
awwK/4CCzurEz6qD1WCM7cGeJZFmUsc7ZHegxsTFCQObQ18TZo7Sv75t9MncOotckPp2ruJYB3eX
WdfJXndAIa07AUEC4GmpXUoITonPHpMbpoAQfueNE/U5SqSnrgvUIGTPE5TLD3FSAawUiLZZS7/K
3kHLRcnMyMJ5Wrvbq5rSao1EvNk0erEbOjjOO0YITEox/eAlV6Y+EPEq5iOODDmPxwya2vadxDhf
mFfVqdKKyjqlYll8am2fsfLkpZooRgY9aI+KoaOIuIt0OYa7IwXEfonGo1lmn3jUPADz1+TRLcia
tP255EfcV4wDDOVtFfHPe8u9CURtkUEkNTrJZltLNxB428/1hRzY+Gu3cNS2LiiixiCcva5sOjuW
3dxsiRYzuuuUgSa/DN64DnOuiK278dNzzJRFrkvPxi2P3b+YKcdQ6X50f/qZmdCDCdpFQZR36IRm
tTIvFiJcQq60jb1D4YzdYPoQdJqPBPEWJ5vlmlStWCG3YY94nbKwebEwu4/MXtiWDug4+y7GQHEe
6y65f7dR044PDw6dEc7vRRySBohsFVvbx5WT8Z8K+eAajRbugMD+7TO6h/8vSsFW9AhKbMBy0Fuf
Vu3l/B8HJnxw8qIUtGF2CM3XNyLMc8kTDF0inCvQaIRSsljZz/2C3JbYtFDrer9HoMEnbmaZRucl
6o2YB9YVZhWK1NEZW+3dqIkb5xEvFKLDcIgsked7Hpqj1bsL9i1yiaWRWdtS/De7Vu8ZL+luld9o
1TaP82pXGeJxaACNUERDOSBrgZHSfiWkZ+K5Mi9Nwfm9vZ7LytDXodcJ6pzk1give/6NDnT6V4T3
H7J4oG91U7zPpX3ZjnT0Tdlyq7OrrtX2f+etsjOVoj+xkItrM2A8ysKvEM4rJO/dR711t8Yx5A55
5ve8/VykdQM4OzBOHqjUTgNFScMSnnCXiEFdjnMGt/mmNyyiD+rELwRPv9TtycfeznvhUOOHIJpV
WP3yY0/EKOPiOPjmL7MG37+OhjnneOiVJ+UMIy8W/MNDdyG5HlsAxDCMWgFlpcuB/nFfLkyDiDDL
TcLiHbnEAfOXiFbwIYWITXEgw64atWCxqLW8x5lDJP9siXO9gYXEbiw90hoWj1N0tTGxyOExVwiH
vmZH+djozwnA5aHykf7AxLIXUOT7MH3ZWBRPxkQonFvAhUdKQHJlUotZfKZQ+9PkD690EgQ9VA1q
+iUE4xh3YAqOWMfoc9jdRuuhxbbRclK+2P7ZRo9DGxpUcs4/NTIl5EwElw1FaeXdvpAs/nlqSPus
KBhvIeFlu0O8y4f5K4eGT2GCBrkh8jve1Wuy8Viz1FYZtxYK25+nsDJjyXpp61aqFyUGslgkE6gC
yHix57qPZTDrxcvr1H2LHArrfpeuPq1wpLWUx5aztDuhBKieS4TjnVm900PPTV3BQdlMdbxFKnLL
00TDIQ6Ii2fp+rLreaFAbBsFvUHuGKzk+jUmfRyyvq2fLzy55nbglPeuWYhZym3R5lX+otisA1kk
ZCI7HvPxn+9GhStqwqgP/TC6h5L/MDV/wxVtAlgeOO/8w/ziBnVfDmJw/8z5mkSI9MwLFow/VNTc
YoI32jPWAt8V6KGoKTfi061fkLiA65E2dSA6bLUmeZkB4P1ypdwyBFbADbrkghwNyLxGugaNG/hM
62gqTYo28bsjqpS1BkBAsyxtkN4Hs/TtrYdry2lxnj2hxowJ+/ctSZTveg6F6TeIT48f8EFGI6L8
t/QtNTExOhO0aJdO5qK3xo37MfgB4Ytx8bq6Ug3hvlF3cqCHj7YsGL3d5CKNjIZ/E8GSYW5K9yzm
QwnQjhCClZCyFaQLU0cHFUQsaTN3fGotLvBnPE86V6GnOBpPfki/jizVgmfSTQ2DCLoolBolrigJ
o88SJi1m3juJUIF8IwIOEDnZkDdUgaqLuc4lNPDkhVS9mjPmFaRVkDvi6z7AzglaSjU4WSyynmrt
wQNDeFol2HvnTpeOK21ApPFnVS6joZdIXnh64uyR1LahUNyAYOzl8cj3NqLk43a01V0kU27bHw5b
/hf1SjnRyrV0onQQKCqZMFf0ByW8KMSZCQ4Fmqeoji7onmOLpluU5IFKAw3IQpIj9iUf24zHURgs
65gGvlgPfqK6kPn5tMRw4f5XwJwHYhonWa45K8TFq3/d+h9C8QadmwD/n6nItII/H6bsxJatogmD
/Do8QLcxvAbV3jPX4ugD88K6h3NYmOQZAIYj/h3hsf/Zyyivp4dIix1fiP6om5nBLx+RszIAm59/
OaXZdBMGkhSNIynYVfkiOH2vWvJGOonUabjcrYQsm51wkPmuLPhAQkGFevXfvYjY2esWos4MAsBj
MEO6HfLz1e0oIYn8PUTEiopLgxCoQ7JXWzH9pmEvfrxlWGRT+nltL34T6gC+qv3Z352q6kL1E2Q0
tMGcoSlEGqvyXJHIWfSe2W0iRrw+y8zhBnT8YqajwmdXrlf0sevX521xIcVx/5isS60oIFjdhPKA
Y73a9uuT3OYTAcWu8csrkO0T+sq2Or+u+7ajLxj3Lgfg4yPyn+HtZXJaFrxWvqPePFsJu1kRYBaO
VhUFZFPpCpmVR9ml3vM6bwt4zJRKjHWxVC38XJtC7ZquZKzjfD++TsBGDT+tYKFTIo2zj+iiG3uj
q3Fc1LA/+j43thnWBaaba7lKsbkjekZWx7iriKvqX1ecdN7j4Hufdk7tJFcmKGzMFfpfFb4MIf/f
zDspPrjIcYKqbpyeWDnZoAw9f6slYMXL9fZcth185ZwTwRotLBPj4aloF/8Y5vipkY2/jK5KMKyE
wch5xTofRE86Qym4WnHbU/lERuyJYSQuoYJFGEGBvVfUaLpfLNxYJYAXI1eMTyAJIimE0ipAqX9X
HbwhOSsxNfmtk5YIvEpaEqfN1cJ2lVy8hyzb/Kb1b9tTiHebugLvqMl+4vLCQfd/Udmz3PvxdKDL
tDrWZZeCFL9avQCwwhryB6aOMIysDwtSOR7eVJ0nPYuxTL2/etxw/eX513Ex34xpL+GwSWL3WgUz
tqc1STr9pdfEpCIcmkPLI2Nren4Dkm7aWqmjaZUfNxVWitMHx22G60kvbfbYzFD9LpWiw9qyHIti
bwjXt9SwnKKrO/5I+HE70ECho9tT9hR8BcrR5R1Xh8kt9Ho/UlzYsH6ljej4/r9HvmkXA3qtniTa
Up1A4jsE0GgvYSoTJQgxZSFM0DWSsLjlJ9Zl1YKzAjurJahw8KdBuCKYsXZV1dOfVc5ZJn1l61xc
gw6ZtPX4Rb+znY0N5po/H64qLSoAszJ1WUqUMcu/m6odGjLhC/e/4djsJCZh8ENC1vNNTTNxurm0
g+47ZUdViAymvd9nkUAlJWXjhfbF7h41LnILZ0zT3x/LyJqWFBjjE6fD0hMC57BAmqB2AhYKiojx
UpJXBGRE/93mWf411uFunUEHOFl4WqOudWYO85dILtHhJJw02LLKCYruVuS7RWYJ6N3U/SrWP039
iiiELvcnml83MUYAeTN9aTvpkzC2VWZEyR8qp+bK/oE13NDxWFlIQMvVSnf7gHhpHa9w/bAKuRoZ
i5JxJiKUfty0Gay0dKnBW9nfPwMrBeI7mdXNkI95f6B9lysyyMbME2Q8i1HyF9jVtyi5geWIpRAu
OhWU3L4HRyxNPHQWvQVIF63Azd+hCBXnjovvHCX+iwqiVf77bziutHW075PcDsqfvw6oR9kECkfn
wu4rti8k8yRbd3Cz3FseeZXUJhBE5TLDgMcX/9Lqb5jrcZEt/wByG3bEGRxe/eMX/W/ZpjLACz3A
0DXTj6z0Ex23rzjVJOtNnGQnYmlA5GRRjp/03Qb4hHy1uYsXU9jp1hNZvFGbJdcP1zcdAleb2CuN
OWb4bpOJ7QS3WQLUGab5Qasq1atL/cdMoXNn/grfkSnNt9JtYOnLsMiGEJxq0wVIKlUz91v2cv0P
nspbFixTSeQHEx/rS01EDEeuR7b8YEXHiZ9AWBHLxgNTMPA7JCrc2j0IZT4tSZu83kk2eBerxBV0
1ClfqxeltwphPf6tubaAb3F1TJR5pd6HqhCYUnlO5oK8i+cVDznV85dGpDxZX5rWO0IRIndgP/WQ
1Ejbc+TEfZGGw7JD1s7yPPRfr+OAmUXrIBJmWQI4pyVbbQEIafje8s/H89cY2ly0LvNyxsLK2d90
Jsain6RnV8TG9hm1OaUnP29X+OTnwfdu6deo+gjgQf6OSF3akYyVdLeU0LdBQ5jcm5P0U/gulrOk
+bJoh/ejI7gPRyPmEyBseuhr0YL312/iIOW7s0WLTjIyWdi1zabC7ljoZtEVe/kzShsebw8ATebj
RwCld9WQRlJFZrKfgyq6SVPXM87fCdY9ePin6JRz3ijeAKtFQUKWshLnBX4Uirovjl7AWdNDMBoc
YSMB8YfwIMzKAauN1ZZTSjoZAcJMpNy9Qt+5cL/Wn33k7A9p2Irc9TqIi/AaYJ5b1PZ68uowm007
aRxiU+UQ902PdtJwpyQTVWOHwZabkoYZs6jPxnd2TQeLxEkBxPG9F2yL+/2W4SUSU9EgeIptRX12
SHgB8DhvetAqKHToyGJbsccbf/1MrIQ5IpBY6JeBpzqUiFX6h4/3Bg3OKaAGVh6yGhpQsN+mmAUs
sZOF8BCY1SI1Lc1a4neyfpB1X9z8hsZufKjxKl/nrNdW2k38NIuFS8WcKdTFG8kKSF/mMtqb16E+
jGWo3IShJpSb/XqXYsq3Gc5LMCaPrHQEpCxhD6ka8fRs5vDUNhy4kU24C3APNGW8PIEXM3vlxGsk
6y+wNRgGaRTjinGQdep1iipOy0Sxo6gTBKZe4wjhJGMchN5xF+hAO98cQX9feFP8vT+YYOWJ5VP/
YFGP8Psaopv6E2q1gxq7hX+Y0+SANDpITV6engLf00Sswx5xX9Gb1erxX9GuSyxVJZKy+Yh+ewuO
uHm4E/UtAJBxpgQPtU7qdNaplhmKT6Blx3ckchQoFOEtwm0v5XUOReUNfJu+faFG3JgXKB+//Sk3
9pSJHO9SwV0bJXIrE39IwNZJoK9Rwtm6Eb2PZgntdZ0GhNuPFXSb8ngOwKv+GMnoM40JBpgfIzks
LC6Y8JCvO6et3ohcKBPjvJHNyLqbsVrVGRxG3cG5pYtWHqZc5sJEwcs0NouNmRjrEN/pNGaAcpuf
S15+Dfpr04LJBkLEiqQRwuDvP/pBHmv8cY+fEEC4iHJrMdb7qBIMYJOxPwTeutE/X7COv93vZ8F8
jUZqAM1p5hLb9DulTToSe/WvyRP6THiCwxRtr1bHh0gJborkHDD86NwzeEeO9gVI2kmH0Q2bB0SR
hit2cc6OiBIP07dyvHRe57qymvjWPZKKPf4PHjWH0C+vbks3T9Ecj/gpWItMP7ptqmHqeVcZcqtf
2u2CsKbjGQPlODVjaw7q5qs6iF+8Sb9psv3KANuUXJn2n2vLaGfQo0RR+2jcw92LiBWWDlEwSCYh
R/KToLVRfcehNRyFXIowcnprEsSY4zFz9MQNifk4wO/WWDmfcvQ3WMW+OE56c6J5rsLAlupNd+Vf
RjimkSdICFFhXk8U/J1QlNWbqyt+eFzwAHRbhR2RkV/svRqxhQknkqBtIJLTiVz3H/Q+IcUps6Pt
q700wGzoL/h/tLn2/qBXQ2GAyT5mQCvXJzJTVsybUrjhGTSPauHvP5iB7DZzxoYLk64JA9gmwrLz
aHT6/j6V876vGqJOeuVNwknJn4b3AvEuteKFRHV+uu3BWENcy/3tN32g7QzgkVN7YzSn8b00UVEZ
Ouqnpq0xiRu4jaUAWGnBtb29aQnceF1CFBpXlocc5HizpaEwnpPfhaGK20qrp7M7ihP6CsPSXSsX
rXdPX1vsXdAeogbd50vy6uekqrpl3VSPszYOgTlvrMeKGszzRyxUx7JrZkKiZ9E5iZfe2lTTq0I6
TLSBH/rJxxWvaVMttq4sUQXCQFD/1BD2zh94fok3RthFMkYcTa/yTEZwB9Vu5ckovlifk2/6zgrN
i2Fsbo5p4D5LR/Vh7ZaMNyPvxMRbBpDDBQYDqqG/5Bq/mlaplZBsJnVSFIS010STfn9E/Q4DWp/8
Q5RaKH/47CpV6C6Tqp82HKcPhQD73oselKM2WRW+EXIpCM//RFJciEC7/2Uq3CMVNWCnBTAYC4OG
h1HA5VxdW4795mP3Z5GKuPE4OZ9vHG3pN5EHaTGOjArRV6H8JqZAQJwDK9/4BZDtSfIBY6hKKDKG
cMGfrfXZ36caSGEAaeCUnEkkTdhN8rnadYbW+1fbE1uUD5DXH1gKyaelAHXKpqc58l/e2tw0x+E3
2JKqs//Fbe6DkVciVR+NEdzAHYRXtelQyqdHw2Rdwrdctiiuu4/xrQcnJG3HzZs63OmCaxL+SHnu
mnJ1BiLPLXSaXNjmNh2uuviXOXRaG2VtwHFkH2UyNwuRhvaz7coAAYt4oGNK7XIzj+tgvUKepGIE
dqzyPrWNTqnqe5bVzz6JmGJFKs+x2ZTntnmG5vcFtWeyMw32bxeoRqRlxauDE7AkrikOLQUis7X7
USDaxIkInjAKR8aXCtlj0NALE1L839y5qxG/76IZqWhlIl1XXoMP4h+ZBuLtH0rNgHUIxUkdHGqq
p+7l2NGKLsZdSwxMbWf3fu/nFCVR36dVhVra6KH7d+xHGTKzvoWdUqOboeSmfphGLQRMYgBXtqjL
w+vn03DViiABt7k7Yi6OTc6ErgptaSxFZZ8z6wssXYA9A0UTQGKycKka/UJ2srXhbmXXP115LvVQ
n2dVoY3xdt4IT6Q/odYY2TywGZsHOXupnszX6lEp6mu3Empx4PCPzabdGrcB6P8FzXwpo4mdVCkf
qBOwThJ2pSyhJG6w9kep6Ufq/E52nj66YAlLjA04dDSKQVG0+q5BlD+0fhK9N/BGbt+vivEEpIV1
7CEXBHB0XWIKu6PdBTD5Rinck/Q1O75mfj/s16IG5qdZd13fz8t9YoStR74b3i/JXbuTtQgwKaeg
bsPVc4+pDySgAIYnOiJG5A//ZibhkietIwvlk3im81A/LWl8IUtNhBwdtWAbH9sTwsNwzDJGftdX
407Sv9NjqtNs1/i67jXgx6IZttiegQj+nh4LeKcKBEXHTz8HsZHOh/4MyG1GcpAkaYwlg4N06L6H
qYPd1swLVlk/50TDqG5/uqtrqAMYNNsAuSPJ7GsLgU3xh/p9BJqMhzWFtzit/FzrQWeczJeg7+tW
bXBZFTBOIlQ3ZZCeU5/rXljjt8HRf53FBwzouZQXcpEGtYlNLo6DRramnxkZzN7Oq39k7dLutJbQ
/2X7JXiM5lvguyc6wZOMtBXgRe0JIcCQKoA/HTwMkAff1qBShPAxEnq524qh3zl7i6hgZa9FFtiD
WM2Cm7pJBLEDKEK7L5GN1tLxwl+eg+pWyoAF7n2AfVTulAXU6rbMeM0JuE8Ikk6sXn9sxuC9TdJz
6XlxRMbn4+US21YaMMyENNvParVdpC60iWe/cpaGWPZVZXwfh9ULl/aa5bwZWYRkBpEzNZ62kTay
MUjDBbQzI7pAnkkEogqdOGW5CIu8rtmLHycWwuygL5808GDStMBRcN/Nb0030h0w/qYGM4O0Hcpp
J//GiUzFzFMrpCa5SGtUJs5JI3706v8LaC1dB7WY3oCjRlFJcFADMj5KYQVGboBtK5RwyqkqeyoQ
cPZ0vip5E1JzMRlG4UmE6ADdgruWZZeOAL3b7OeLyKnMFUXSTy0hPzsH9s8Pxzl9wF1eOyX+nhPo
/vopvM0gP3jmkxtXsZh85wibCNyG8kT8oXl5tNiSIS5UThJCAypiH+6tgXGYqvA/LT/Cu2XQWXE2
i1PwOMbvl7zEpetnuVju1SoydN402vPHbYl86bijKTOdsLiCsyr482mgpf1OjreKZSiEhA5cQ46E
JmNNI4nRIjwxGMvU+I+daJ41xNtb8utFJbva/ZZtyvhPh3kZr2BuKwdFwfbZsmmlUVXKLF8l9hcR
4GQeW1Bn8SVnlkhcs/zhitVFQoqMcK62dtXKXOHXdN2ZmX9Qjy2Rj6RTaD2u7GOP5tqWXLo1nwMn
20q8k9ahR0uCQLdJVzu0OUvWMBwH869ZgOux0yW3ZbNIuu38ndsyUVyJNsZge+brfPpjLyufZ9Sa
yOBQECU9h9t5LK2lTvsVAhturHdds/zkkZAh0LGY0tU8uJ9PsOtzKXvyoPYk7jaoLEwHeDugshPG
ecHaZNt9sknwicI5IMTeCK2RDckNrTpSZUHIllddRa+HIYJ6kgyZZwNPr3CkRtIDTbjQQ11Dwlyh
6EB3fDRVXHYXo3So0ejsOIfZ8MFqy95Te7U5R9uCFWcSf/dmK75khPa2CP0YfKcclpWBq2RuRK92
U3AZonzhD9H/r5rL6LMa+uX/boBXCTyvizlCpRT6L9jpnBSN6Hk+RJCzyZfhSiwA3Wf7ebkpK1fV
GKW6yakTvAqUuIvCDX7+yQNXirqeh9oIgS+0ypNdlIxjHlTgC2hrDuZonhzQmSsXG/KgnVsOl2Mz
Nl0/FD5vvSSatR3BlH82DYxfuf3vQFNNzagRcGjd76jaEgl/JZiMqOuFrpVygUh91M+EDxEGoB4o
hxFoDcNBKTtMWGtaPUOgk5Tk4rLy+pbD6NO1hUXbFis1zWB2NzDSv2+65wRG1vPYBJV8Q/q5tlGv
tEpRSMzK9xGGOpLm0A/tis98yod9MF+IySAMtMBSUlXGgAtBoL4QHMeEwIjHfY2j4i0LoSMEV9+n
7rfji/ffh2u/SWzM3TenSS/5I4jsWgXhzhr9nngllpfvb5DZQJWY4M1YbMfIgqhKjlzHxFayEmPz
w7tL/QQPySKcfGAw6Cj8ct4pbi5iuKVjUJLpAIaT7gzgYO07GQ5SZaqTOW7tVuxe6E5eBpgSuywG
cdko/V/vekYOsdsQn/BDd/zWRibH9zsHwctrKLADiAB4ZmlL9AruzZg/SN3I4SJK3Bd+meqXfgMU
+NkR94YHhPORahyzLggf4Y3EBdvmPUz8sJKhY/KU0RLeImXN+OfEGiQYN4M4o/rUk5xHKdq2zU2s
AaBxxKeZ5ViIgSDkF2eM5SKcqU+S5OV92yxUGlJQGlL2AloI2OXRl63512qA++BldTnR55toj1Bh
/j6BOhLT3ng+nFqfZhveChgO8iOzhb2qlKvKoOt5+O1eqotsWuTMoVQlReUk2no3yGwatTr0Oj7H
H+KiQnyqaFHr0B4odM1bFjZDlSLdGR8ngNO/foRgXdEd2NYy9jJjWgJejqZXX2fPmRrjQJoFCO0P
upsBKm4w9gQcZXsy/JpFfDs/rpK2wHlTlXiorEJy3UujDU8jdSXzhPXksHyStJzj/H5wywlp4Am8
Wmsy0vAGpqu0oAGntJBumg4VFkOGekX0+p+/wp6mnFdno0d3m7Jzz6hs2EZYg60cl51yU2v4Njml
mN4AWxk5Ci5OwMDviqbjKhsa6lu15QHp6GzDqnHgKc80yZnmQphqHeakR41DxABhCyJceZxJOHgh
1VI7PvNjPB5MWRZ8nAuNiEDNbalWQiTXy1B+cK0NAi5YYUYum69mQfk0ylNx03nsdI+LUf/A9JFJ
fLUPK3gXJXap2L8Ac0V49/cpbRIzoDbe3R2VPJLgr9HxAT81qFnBb5KyXMIpw8fu+slkYFpsHosb
YyzyfgVJ+1U65glnL+bLryx/GeJxD/vEG2MjAtoH8d8nbJqjKfrcu2YPRP5MdC8W/1GuGv9uMnoM
uB1iRFQ8BD3EaIxTLsKzH9/f1ZcYtfujXqvbzYnWSgWjwWURnvxBj1mgfziR31aubIyFkgJXkEp1
zN7TPgpJIRcDKDmYjfApK9a+xpq447NXGUuyLsZgMB2hyiih4y9j4aFfkhW1idCQkfnjm+v/98g1
ULgz+c8VFXaJHGKHcgE6+2dzRUqh6u0oQ0C0rE+u38kfJzxlDoUfONrxXCMoPo6G+4nXU603bNZn
vKzE9fPMeAgMPaTkpiECEaGlS44mDgg/LMl1qkjs1ZrZxkOhRloy0Cnxt6YsSnk53+oCN4j+Gn3G
j7luGnIXlpVFzzetq2Yv33joVOkFHPmS8xkGcKEhGd4WvaHwbVDngLhHDbuXQ4dEOQLAhTGCJoBo
/JwUGXS0sExnrOv7dxMKbdQQZerGWNv4lbvb6zqcH7wBmz1Po2cUpBFGnK/Q1LDwjrJ0t1PKLcOz
Tx+kdyCX82p/Ufc5W4Dihol+KKVE5CEraORZUMAeseMC0iTwPpcJvOULYh5w3hyeDoc9nW+t3f9V
OloleOGRxOx99cHmImFSWZiGtAL2K3Xy49brrjKVZwYUZPmOlE89MnM7RiU3NbeGQ8vuB+9fySpL
T3SkWFkaQ2lTAz/aAE0W4Jm7ZOffLCWDBkDFJAsFnGSH9vLasR38c/34FkELgi5YOyo9vWMzgk3L
TkoGZvHISJJTanaGS87LFGCa0N9nPUs9CVaCti/8N22tjvAVdVg+MCPanE1C4OK+1gPkNqKER4Y7
jP0C9dqLJ03xt7pRhyKBGLY3HU5ussbg4BQfm/tea7aSbLIti5m0Kb6xZOnPu+tsB1J9ypWd6EUe
wrj0bp4/u+oBdo5LCabcK4Jay09IRdiGW6YwSieJgdYYFGf/1IbdywxkYu8aE7x7JaAT01KjnTRY
GcOKX7qrChISDw6UN9qyiMUjmgaW0asPnicamb8gGgth1HLof1zwewTABBKQ3L4gBlIfmfGiX5+3
Hn8FdxyXB6SDfCU+bcGu5Vyo+Ty1Jf2l10CbK+dy8tulU0Gm34+9joRVDNzd0vZ5Ez1FEILI2IPF
cfy5mHh3O8n0M1eMJeHsZkSQuNFlnX9o+JeiUC+pn/XG2rw+GL73HaelbdlrDsELswZpjo1ybJWF
2/Ea1ashPzxyZ7+Xp9yNXug6MYVFdCQNWhTHiB6KtFvlMFbCdGE9QKE45h5HjPpOLWtCJOqRRoxE
9dLHP/WvRwgVPR3+CfYzElBGsGKdeO0XaGiVmOKNyskft0Skmq0jRufncITFzSu1T5MXTZz/ftxE
3QPQkuqqyc20SjdIq/k05gDpA9teQ4rxc0e0973ntGabEX0K8Jiy3BGUgRrYgs40mB2ItZvLIUn/
bJ06URwgwix6TlbI/7C9cPrPLK6p+ZN5s4osTG2KK1nIoFNMxasPqIYEZvTy4yUeCA20sc+lmxEi
xs6v2m5GruTjAvEy11yvFHgvt2xRi6t+ISNTvesswk6mNy5SwVvoi9lbz6Mhm5ffjLuCEbzxVWyb
YmzYEvUSX5x+EG4pmXbW+HWPC0A0fZJUpIlHoLN+F3iSQdLS0jM/JtYc11KsXkTVu3kmPOlECMHB
023lgiAoAPfFeOG3xBp0zYmm3aAWwAslxGgY0BfCuMRiWhOVzb7DbbGbWh+TgvuSgCPoSCoT9ndS
X+WsnG8qw5BBcuWoBSudakpl7O8ATDVLLhIAr5zQ/R79P6dwWOAubMuh+O0W4Ul+jFbviIEJCrb6
TlXmExzwcwOuF/8qjgQIvwCgMSV/iJyw2b9hujlJ7K40Gx4NaiivO7LpNY/Jkp9xcf4nqmNNo52R
fKkBpsFNDWk7XXpF5NlonzWg09H7tYRRXsGuZCxaeHJEqxrjSpOsGfmIfZuHEplgQN/k8BctGEE8
5qHBY0Uu9H4ccyhCOJDmiat0Da3k4964+v+qpPsBZfg8u3FJO3/VCKnCwGinPWy0t3J5Nikggl/p
0mexpAZpaiqz6gohWHZVC/oz6WaPCEdZBOysIMoxy6qO0f5Xljvd+SF4Ym8FXVrC8HnPjfzsA2B7
Eiju0mLJrM30O/RkCp5rRr/0x0LKFzerDTtaSnFrVXYi4z1W6pT8/p4iznidTiSC2pb1cyPxITZ/
zZ8vDcgS3z+XZYaVjFs5oKCNXR51dYRM9feTV7WrqI7/6X2O5dD4ZUYfPZt57epm0k+wBEdCoNku
TgxFdTiotgGZkvtV0C4wf2dYad93TLSkm7lzBUbCRhpnKPJgWMhncpDQqcu2Yvds4/SxIUQnWI5Q
OEHLbl9n2OoUxPObpvCeK0sKsPggU8phATMynZuhqUoKMvRuz8o8BXzAwcsGi+svj30rhv9RKSqx
cF/0Ktemz04WmGrw4FecesWeZDWhGjtOy0O/SqwQ5LsmKcsfcZlvhiut91gP8x08g4Yr5Gh4wMLS
ILPcVEYue3gOu+0DWFq6Q4Re49WeqDAticgW+aS1fOTbiQPMFU2L1Pfw9nZJWjKAGdFxLwu8O3r0
buUWOOTFJV9ei6UOtE6wPooZeB3Av3v//4WL4ee6bfJW6ZU8RobWpdHaMeWwdhS5Jytty+Ua7o/y
5VvsCxQxiIJvom0AgOgqLOyKSD21tlJtwms+EDInwHiXQUEuloG/K+hGeLyFtqX24NRgTjAqWSDY
xgyKXpm8Ga6QWxcs1vJAJoOZ8UJsRfwA8AIosd1yuZ6Fz6nT6IfhtiIUUFTe3gVvQ3/ti6AJEm6J
x4I6EBF/lMlpdL1mHIDGe+CagjKKRfnEFTaBxFHUPRVpi3i8kmFGkJmyOQysGNtidtJkup30FIj7
EyZqqx0zRhH8P0dgxWY+v4MAZkv7rV6mbGLnu3MDq7EYJ327uhbxzW9G/xJ5wLiLo1hKh8AE+dtj
IxbSZjHHs4TnTPCudKqA8qwJKN/mUWnSQC/KeDC5L5/IxZIBb0V7m+03hbq+Mmel+04VI7Orp+rk
Nt79TL1T8j5mibO8h2eJpcBHhjQpjrJcGqYg7mVwZ55n9w1VEys2n5z7keMFBsR76zP/JqKMGeUv
dtG686duEy5heseE/i7XbbaXE2EANAnGnAW5WtoHj/ysKB7gVoSXxlPdklT4Lq9ktZMDxmsfuMCc
paFROWgwdSnARkMo1S7MCIaw98UnJabV7MXQfyeJNJgPqb5nV9BhGrEMnWRWI1zt/79wHfUzw2m2
ikIxErdQgt5voOmOK31vTCHLV1qXOkrdyfuhcEQs7xQNT5Ig7LgiTuXYNXQIhBkVCIGWyCYq+5ws
UnYjVdJx1oHL4H9nX2XafvAE4aKs8doGmgl/jUqId8zHRy5Wjl2WFq72lSkwUgKfPFRiHFqIBg6Q
fxfSsQnPY4fS/Dl1Uo4uAyfpgD2p2tGp+8jTQsUFkXAuYABpVwUMqk0wLyYUQL7qrd/XHrgeo5Oh
Kdc1hUd5Y+KG89sFFLWB0B+ggPIcHqY5tgM6gAH2VuIsGWShkYIYaalKVzsEeBE9AERD89BLmQdn
MYTl+jjSjqeNQpeRmabPQX+z1WSzRz1+oXYCenUAwEsU0T+jDmlPq8hYhhbSVWVc6CsVfwRrV6Qv
nHejdiEmJxdCOAkz1Rgtb3DelO/aneOi9a1Q8BSJgviPL6R5FNLIUYg2LsZgbu9+rf+9jWDxucIr
v0JI0+O9KONPvVuMhydK4GhtLxDFvVFwmABSIKLrMFn2uR+vhnnDdjlhWmlHXa+iXlOss8HOQ1ww
I9nBgLrhX17DmZS7lJgyy+ihx170VDJE3f43N4wmI6Q7QhqtJr23RcPr+C94Z7anerIBjHu82dvR
MbwdEccDFaXFlq4SNwCNfk/4RB4nr9eXsnFG46zYOOkjb7OhOYv6LqZim8WzMfPvNTaAGJ8hD2zr
AE+o/IZTkcghRQczlmMDNtQS4WrfLfg5Xp8ya9hN5bAidr3sEeKfsdH9uuIsOLdfzrGVUm8iZZPp
Cwse7uBJGx0NDIrdGg5RS3sWQWcHe3xzQZjeXF015nf2kQQ1i0ZcygLfzWSO8SmcKHBaa2SDGvEm
p5NhR6k3kdt0fOCzfzQPka4OxvA+4DcyBalLf1hnvM+kKY2H4cXRCcMJ1oHO5qHTdMHyCTznEaa8
Bs1Exkls0qoBsYjzAwZ9DIDhqZE0JizgCMOPA6ch++B8Ctl8ktlDr0SM+B5ltiPnCj3xFVQdpApD
Ubx3tziyjUuFkyjFb13pmecKdeTIK1oZK4WEWbgddLd06+WN5QZOVbiYf+xc2VaQ7u5jLAQ0G4E1
+iN3Qk5VXvhukWHd460jZvn/rwz1tUvmR7snLkuXUqXwdk+3cuAaarQfAMnvVFaZdsR2xcRG68fi
mUf1k3cj+HFsaMZnsmxn0RPiehTj1YC4TLRaQTPy3hDNbVudGoTF/NfNNbr0u/Z+AHk7drvwKq2r
wexSRZ73apm685h7mukvP9Hv5pa8iqXhMxFIyljsx/zwN4cuOCKPZ53T24c7envcmgzZ0XRsriox
p/L2Vj4FoCEgKQW1hcqbp/LemuwCRUlPoK2kWexFytohDbXYH4B+GZqYHhPPCGaPkreRHRAEWb5n
+tQhmR3GFfnCEp77MIaSbC2iD82IPg8ad/hVm1bhwjPviwHvoxSqdd/5imkr9vIkdjawl9ujoAE+
xOMqvMXl7weqS7kvC7wtQP7d5Y7D2OZ2HZys5H2e4WqWZqUtj41XXJB4GOYciVbbe+OT16lRCcnp
qg4oOP7In/RZR6mnWTq4ddvJ2kQpHziR0awUujBxeb4MaENj4tmBTcXLIaPsA2uyzT8Dpv2ctHoA
hnin4XpcixN3r8Hd9DuB5zmrKKhfVkWpz+J7K0cHBAsS1s5DyFAYX+cG67aMCKEit6bnfJ8sY0X6
M5W3AkiofcKPdN9gR+HVPDAorF8dWim06U7nzL7O7GrgFCZyYXyNeJeMy9oAk8o9pf6y+DQIf99S
lfnQ4JUwDqTxaGlSTs+wjT/NCrZSuv3FmnomDACPp7fnhwK4TM8e/HF2oviambiUlrXd2HIT/N+O
i9+CxqNjLGXMu6+OWeRsIuhVobDta54pMV6wwS8D3OpdNVUNpL0qonAEab8Anvf9X4i7WR63EOiy
s05x4WCHtMgGQKy7LvR7k47xdQd6Mks1PQopSZ3hqkF7zS2g5x9DHNhgOoxNAhJ2TmHMzCvOtFkP
0YZjVnP1ggGCcOsn0CFKMetLzmPSpBSIqyRb6qrOu15S7Nxddf8lN/u9GREGxCCecPBKm8f6mQ11
CR4IDYSLimRghudC0Ply5HjpRBrtsp+IUazIroQJFPqCcW9cAFdze0dIEeoGd65q5UM7tH+C2+k+
pBC9OU9OWqqPg+6Z7V9yIodX4GDHCtcCCHKhONzYo/eT9Vj55OFODfrhZFMMMJvI/uShEQFhWKz2
BBkncoGwo53cpqWycIuFw5G7WsMi/RDO8JHxBh72t6E9NRHBS2I57SR+k62ySJGKeQOyhIrodNQG
LDTcebpslGylra0AY9Ul3W1V1XtRwWNnU5ocfBJEKJctto279OsEWrqNZyi+Mp4hqlj+X6UVg+gD
e17tQdL+ZUkgI0+tyv8ebecxQl30pQM+ija6fsGsT6X/iVuBZGHCJQb5F0144hbl0bD9tnBzvDTG
6mLdcVbCl4K/z9E1IWjHXLWsGG3QHyzVJwLRpPQwiRDeqPqXj0ZxgkMX4VJniqny6KNCBefunqOU
WoBlwWkHiEyrpHLhRS3SR3dpo5gL0Mgj/Bg9yzO2wgCtocHhEAIP1pn8+v1gROD92OazBTmh8HdI
bFTujWBy5esTRUOZlPjAssbQu26g5KljOkVCNTDVx0iu+4o4Aj+ddw/ovBp+P0WgrZKJ1ZesywEs
+LcK4ZbeH2bERwIBgqTBIKmLHvgMNHHp8ePbEfXTax0ioI2G470BRZxbR8o6VWR7yovve8A3JypF
dVpuytq3JtLTP5wa3KzDms5OwXiDN2e95PUkQhvMJY64kTJy63PhWbw+LonxbjDWIAHRC/kmjZqe
7ydGf5n9vvkxLQNSy0kqDYiDTB1WmQMjxa4AZxc9/Qe130/erJ5FQ1ZNag7GJEljLckfphXn5RFB
fkc+HgFQZ/c2prQ3Ek7WGa7bEIarFJJOGodhbE7/BTxuMtjcbhzosZLyVCtQ9ah+N8c/ANKI8n4X
cIdcb3sGeMw+MO6g6YUfFqhlCSDRlFHFqyub/5j2CBGVEut91JhqYq+M5K2+7g/KcnIkAfUYkbLH
mI83F8N9C1zSYlMeKwAgzHCIRroRV5RQtKO5ucH5gMKjJMwwiztPVT2iQu+mbox8QzThIa10Gh/8
yJbIq5P0Y+G/SgYXTEjlHfsMsmPKY6HTRKOZAGx7ma+RSrhwg3SXLZxJYb8LkgeD2t45sA5fbjk9
MUmEixOSJK54ED3n4jqs5UbaZ2AHCA7LI9xSzVqzCoqMMF1NSfq/XdLkKZBrOD8X4VEuxUtMecwY
qSrJ01Lw+EPwelWx7K+X8k4Nezu6hu6m4AG+3q08EEqgioZXMFIUTfrU0Ta61T0HJihKs0FE5+PH
VL5mDcW5e6wBa8Gk7j/YzXc+suB+DA8wzT+/I9n7LosI+w9u4AtlnJ6YgzLYXViHmEZ6bNLGczkO
iRR71MO7lLHwuSBB4GoWE434M4z9vgQtVEqGDcpJGdOUnYjRrukx7cyhGHG3IAcjhzoH82vXRWCF
rY5QMMFgrVhTWb249tA6konFDdvobzbobEPL1KzQGKCajg372nXDtJuY/Baq7aeJtwXmrYm9avJ7
xGDVA/RLHXpy0eiv1GEjO1AhuNXNgY0yv4BvREZ1HIK0FjrsK3nBWKrx2colkLtFWLFDIubS340r
l3TwSPcs+H03OZleImOn3j5VyWv0zuQg6qo2YlQS72ZrBZmNk5YV96+HXscQo1g2PRLs+WpRdu9F
feC//dccv2nVM2hDhbWQk+ig/QAcSkUUzZEXppQtK+Tf1fLzcM44oP83sOBlwuw/jkfAicn3fuB8
VrIOhT+7+M9meiA6jw6C4gNUCO8t0R6BlmBJgslrMsxwsR7ogOAx5nJwjT0o0EHsgykvV4mzO+jJ
UPikUsyZg4QY9m7FDAB5lD0EznQxP9L8636HvsO83AiPiFNyuTSgq59SYGVt7UHkl3SsVKJ7y1R0
jnmgtZXvzSLZM1DpOz2CqickLk+xk+6n8qp1PUIav80W3rhc8Pafun39yxXqhlRnc80sve37W+J9
oZ1NBbjzx18kHkRVmU/L4n57L+CYxdVwi+homnpV0cIy47goCUd0GnYzh+FASqELmDNQiErlBVA1
+mTGnl0+I7vm9yk3bwqLVVvpe5FACtR0z5PWf11f+iGf3XCEWam8efxycent7EEbIxfOliHQfoys
yp5m280gFMw+N4SzojndlBGGmvR0BYAY1BvJjVEKpWbyvNgyHdYc6qHEPuKnwv2ogpVoYvQ2BfUu
BgxT02wB7lvnbWPkgYJh6ugGzbpuY+M3tO/b1l4A0L23T4RzARk0A4Owjj+Ub475c+m9OOJ0qgHg
f/na/wALrYYGUV19RFepH/bqNyhDmT056yWMa/WAq/YLiZUWTs8E0XZranbpnEavZV9bXUR1zJPs
42bdrV6Ua7h4L+wIWZ04wHhMXFyDb9ZsIsSk69n4+s8LtS0zpIvqznhfgkD9Nl8tLxj/Rd7DHl6g
J5Cw/RSqayZoylr2zWy9bxnD3OtzAxwnyxuW/a4r9UxhmqapmVHC/j8UVKc1Va6MshdHxa975qEd
81rNvwAx/fi2NJ8YyXLTIAaUfWKUeqGNtypV+mvB0IlSHb66G14uUoeOxd9w1QtADuHpJWDdLF9U
XBs+kkOFeCOVee41By5LOfmU1X1rY3ezTGINNxv+naqk4pcob2oIu/SLYCG+11iPn6DS+wf++/9g
hwoMYy6fdq5NITxcpt/c61/Ip/7SMT0FNTZLP2KqLt8tx6Inb+lQm9/rEL1WkPogOcKh5AZZsBlM
g5BWNH49HaNrqEoCMe0DeU1cbf1YiPbq0lKGISdVIt0UGj486BFoQ0gw+8JE68PyH1Ol0zcEYotf
UeSP6JE8157mWZO2Wdh270d/b9hhLqLmS3+ihMOnle2PxYw7jREoIwOSlrLVAN9nrc0Z+fCgMfQr
Ruj+0IItXmW8mXnsE773Lpw+Em4Ag8CDnt46K7/myhO3mlU5nKeerCdZpgdMt7q6phBkTF/WaAE4
krbzcOd9A6ZK5IRjCagKHm4kJUVCKmvUS2COxmun5ndO2gdHhHvk7qBnYZtdrnFP36vfbR0MLm3E
2eCkKT4nJ9vvpIUCworB1ioNAZT6fAAdzuCWx888kgVRhu0f+Yf303E4s5/yACobpGSktWDnaPjZ
AqNEHVe2h34Opb0cHSYvU+P8k04QXLQxVw7xclo1GwH/hO7EJdb0Sa4a/6LbGFA+TlwJC6Q8AyXL
B+gnDuXA99c7ZUtkLFLCU/aiu7TW4iK3BGbIyh5k5FhAlaPk6F8at4QjKwWBGbllOWbeTDymEpi+
FZBjmW5SiAXV4+1udaoPU88S1s86FElOMvFaLgzmDgi6dEl0LRtTiDN6LctEArcAh/A/B0s7ZXHx
OgBU0UKEMyUOcdDq3aWOtlcixXkzMoclGjLi6qiqQikJuzRX3hwjY5UYCk9TTTRum+a/2sHoVnRv
NSy96/uhH71t99/81AOSmqOcrUz5LA4G0cssz16m/J4v1whRDgpaFEfpMsMiBWivqsnQ03NKM0nw
ki22xubkXV6vhwmGEQqe9Y9oafKU8oireIkKbglyOP6e9kDAKnvsrXPQWa+6LSycY9RJJzApv/dn
xSBWVe2csAVnFYvDPIQKpiWCvmO3EXWArVeJml8FOql3ymW/SiUCqdeebmanLTczo8Jx5JczFX0y
krVXCyyNLOTP6do/2HDKoX4LAJoFaYcnlzj6Np+MyLJieI7WuIkK6BJEB276zplKBMXiLnpBQUhz
E6R456Pj28z98m6BuFK49M4X+YwhUlO2U3cBiXh0avPO+Lie1hDQgMaLdpi1fhstfRDdPybHAw46
emJFOGjQE9CGqOO0WSHhzFIqP/yVz/A2QLJM1gpk+yAPUC96AzdtibsdOQM6M5RT/PMtemRe9n5L
40tZUadMObWWZVddypsasavzv6KicGrgELX1XtF/4V5rKpETZCBmx8ooyAq+I0wDcGH+igBzrEbj
oyfin68FUVf7A/OM2mPVJig7AdRP0Z2FcwDOFUmjwxtv5cHEyWrRup0tQ7OIpluExH89wiYkOlwf
EU7DxnqLfWEGQWaatJLhHJ+lel/+ahEnn5T/J8JxAvTZEyKuBV4tLlOEmQrORRGxAsUTxs5GLPdc
jySiAeCrHZSZLkSnj5KbDdR6vPC5t8fJvRRCNWygS5rDoakoJOmldcvsbgOvXa2yANMrIJAZiaxz
1tCZOCE9/E+QFjISJnyS+XaMu69gJfTPZnQQUcUBkkeXTOOwer6a/PY40UUQ0+2UBXBHeQILe1Ka
ems2H/Sm1kYFWGs0RNZWqWVWVRT5cTmL6tPHL2Mkud0iiFqhw3y6EdhJqaTu4TMwk659OjpRD3oK
UFpPcvqCSkrZdKm61hUeHtRrKdUzV3CHF0LINxZwjR0zUKyeC6/z44UJX4UlPcbeMflopodCnaY7
GZZM4r2fOz7atUR7wBtUyt38LDnACMdq3/3Ds/G1XX0w3KzjTF/iz7WpA6jGwlpOvjIlADbTkSNa
GpHWXyL5D3mZ1/eYdVWcvtCrH2OBR3x8JlPrMuuTEjri7k+Rh5Q8uuWtdDTEts7eN9XcW9X4El8J
utbHWyRNr7Bv7Vj2zoKjZUsXreQLukya1plKJnXJsSfZFq6zYSTMybB7Xe9+VT+JpTjdRz6Cd+LL
i+npfNQ0rdCWUJe+r93n95EUrxcytUZEG3AEUK6lD6+AxTceD5LYLLovpEvTPw0IIX7I3YCBnane
m+jex+hAfIX5D/XL6RVLarCIoGXULWlReX1PR83LsX8TC5es+Vt97J9eHXvOvQTchI7fwF+o9cse
4biouvwzvjehFGXNxNX94RKiwu9kgzTq9dhvsQIBBEhg3qr2aIIsebKLIMsSBANdOhw59t65r97H
kFDafU6msEXPzlAWoh1TcXLe/dE+sCh2E0G4BntDi8jjlaj+kEolVOeecmeNCi87++LTM+jK+w/1
gpwhrC8xmuM05mImzuu5A6K413MsGScVfpeaMzYef/hHopqAjJXOft9eC8xHip7cYyECh5JUnZGb
5zQlyVM2sW4C9w1lBZ08wYqNCpy2xpts/Z+SCoZRNtZ5w3X+rZoaFobaTptshxqxKhQvkkNbwYa/
kYBOF+Pbd9HgyqrtGraNKkcMOuSM/hqQHWBusQSX2J+S4hcrevLjyRfBI4mJQv30o3V6XmQiWmp1
CUZH/AALIUpuuydbQIv+A6UH5TMujquNp47TjYio/IVFviwapKeHourMTfmOBI0qqHsQO2yQ/fXy
ErTtrPhSayfQOmgPbGlNHKxDQ8Fs6xDn0FpFQILYsp+yT1upXY5eMhDD4KjXfJ19WT3HFszBd836
Ku01IDlSaqMdgtbZsjo0g1i4rtPwJLQX0NAHb9N2LyM/3A0Sl/64H03uZX2b9taH+sRtdmoK8p0J
p1gRcxASUQIzLcdGREK35HGC6Z/5pluMsk1mJE3BhLcFzteBjhAayfQL9/HlfUDcocHbEkmn1/bI
uS2GBPaTfBPgtLlKKrju9M/iZCRSLFdNlQ+MCx6zkAip2Ioy1VLJ+IUY43s+N8vA295jxlB+L40P
3VqUNNy+jGgVhh7Rz8jFDK27cja5NEDEYPYMM8+N64Rr9Mrj0/yq0tJv3BdBmyyb2bT7iOBSHPOb
rGYUxVqoT3cNmnxTecH/n/EtvmMCZKL16xzmtFMLYpi9nAc+qpCDsBJwl31jeDFYuGkgBmomvI2x
7QCF0MXUbqMXobRIXGA8CddPoJY3XBqoRNc8+Wm+ROagEikcK34Au4xEXeDwLq2wgdOIu3315qOW
8+qer00HinJf+ZQpfL+dUmf2PBJimuwhEe4bld1677NeCPDhX0eMb1fQX5ufPaI1Rf1dq4cK5ltQ
QcOHGfYw2+lNHwtnxfNdvsQniO5eVM7S4q1H0TQ932d/tTxVJt102heNQP9zcm0Lfz9gGnhcOJQT
9CKKD68+RC9dl6jMkpnVV9P2Zii112qpvCk32aPC94xNgJkIPbHCInTF94LHSfsjL99tmWWo2Gjx
ec8AlUNeYKt3CBPonsupxUZk0swF3xsn/ca/vPz/PQLPd0kD1p8FbS6b6dfqikJfGnnFsEPUwWUc
HHPnfbEJkN3GYcfL5n4E8Ki++vP0ZxFCnOFGauQsSM25EFkGDGM8OilZYoJ9im8yF9TvHkY0Mufv
MHrFRUdVUL8Hjrxgzi++o54zeD6PjkXhwlXluJyx5TVgv3y6OyFkY+8PE1kwbxZG2zc3BbZnKK0V
Yxl18RgqlyG362+dj5VQ1CUIrvglUUTrTpuaAVHUFMAWEfhpyvAzkSl83CUbWtv/krOn/0wc8bCW
LuV7uuxHEigRJq6RckUEgIQu6UlPTPeUs40R64GvtYy8eOFfaqYiT2WoLMRuReKBh8f33Ag4tCqt
bcw9iqHBM0JoizExpk6v/t7iEXFiJFDXg/lLMDWWEZ2LKJNf4yuq6Ji8YnNBiV5NwNHEG9UqQc6c
vvt2EQzIZanQFu3KIkY2y6D9hNfy7NZDyS6HtptG2FuaweJerzutizo+oW1Rdd9CMFFifE618RZH
JQf2fuoeZGjG7248Yj7MG4OEkhMwxtwMf9UczldqQ5eHc46vDfatWqP2AKTi2oA5vXKr906SBVFf
vNAyFapDjbIziJTHZrpKKb9SBSfEh5Q/eREyaanUhy9+JzntRpQd4USOY70bahia+V0FNfzNPqdf
OHnIwhZd5gVDvIx00efB2fOuKVTES4ozOfCOk6BzinO3iW4NkxkcljL/ZRezLyHGzj41YY8D6JcA
rMt68ZCrtSuK09brjDgwjv2V4WD7tHZCixTEHJCjlOUTumVULSmj8UgudCHWI6TpdSkhl2iLaVHX
de6dleTW/Cx4XKPJZiOr8j2QnElgrQSNWQP/jtzpeDO9xNNF4jKyabZZfg4sEQL8FqrEqvoNteWQ
7U4Nm37fLyl9C3CID3AemV22ZLDGSfUGmw4QDciGLrnhMJId95YZXcCa+aQWpeF1pgSKACv9qId9
y6PZhV7mvp9WCPS1QjdWk1e8zJi7ccLK6zywLx/eeBg9y0A/DRi+uD7/Ma7FLr+W0PTpzbwR4Z0J
s7ylglnBjN7P6elMDxd5nek3rvxeJsW59z/KUuYG/t2EtTL0ApFWwbwEFswNxA8vHaNzh1BrM9Z2
gQM27uh+w164GpFQfZ76MCO/8Byqz00BqqNnQGjX7V63NcbYiulAU1jw/Gl6XrfPlTGhOKUp67LL
UvWhb6Sn+I2Jf31t7gv6e2iRJJUcm82XoqB2GaMQZkMKm5elF6FzAncRz/5BV3DXsaLFFz2ff27e
8RIRHkDKRmMIuWs4+yHQVr7qbl6/1P8KUmfv1tWJh9x1WuFrY3WmTWILiUv3giDCjahThdailZXo
ZRegJTpYMuHzDpqH+pgV8S2FP4oEgNbd5XtpGwz1058Le2NYyfWHHNakEHAbCAEGj6MhaHbaYaPK
2cmH3alLlBbPLq7qw4662AikxiduQQWicR3wz0TgayT9vxGgqdTHieR8YajHi9wmYIzTHiPn4A+j
lMBRpER808kFQMfDjvLOt1DogAp2vy5vGeqrlNY05oJ0GRXqean9m9TDqevvkcuEV+Kd7NlM21XR
Mrh+vjC7t/JoC7FFxC7BbKAW29Bt+zaJSUggF1WzKF4Iqlz6Cf6MpCpiJB93/UGBbnNKG7kw+Tuh
YDkAZSuPOf6cl0HMDb9QmhgABX32SZ7qS1WcvvMbuGfsVe2/CJDrPFxjASY1sMeRa1+R0p8mU5wk
i2PBKApcloWB2EYHz0XpfUvn6oKiR0zh0zjBKfF/g/qPbNVKvnaH6jA8P52lgE+S79QezxOtGosn
TQuCkMbOiIU5G5aqsnLs3Dc+Z7HTaERnMajrPxk2l9h3GKQyjadbwMxoxkT9v/Utmtn0wV2Qc3bh
tap7mYQxuk6VOdW36BQCGar3J1bL8T96eM0O9uMbg3RDbG4hmq855rXzNpZIp4iojLMiVlV65TKk
31pFkZs54/0v/6ZJsK6vr/UkbFDErJzqp8E39kX+YY9+heLt0xvBpxFHhCGPuNyhWkpRMJqc7+cB
uS6JLC30RbUscHdPtO1VsDgPnG5HMNybpTZXmLVgk5ngIZHXBtTDMNZgD9g3qKI8LYcC8hrOt2/j
FyxnOX8B+Lc7VJv8plhl+nf31IknWVLaSv86fEfdzKwFXmVgk23qoDlKPtgeWxfiwlVzR3t45Noo
EoFX1y9Y4kAOXxY9CM26Pii3VM2Gm38e+8AGQaWqZOd44GvM/4tXflg1tajWLNCTC3rO7qFnNMBg
s8HlWJf3OiNqexds3fQCp9pE+rjzXFtj38mpsa6BPrJ57HAwq01RrdO1tC1i4aRIbZVNadJ/BtRS
V0ieGGbkUBmCXySJGjCWI35G467ugC0Jy6wUjXX9MalnlklNAKn4do73LeJYxrg1rwrNiwJ6qtjX
xNtuol3vWN9/61QOWm3QpVGVAUfF3X3Q6PxA/7X38XB0A4anyPP2mMk5xqlcfPR0b7ZqQwhHYEsx
2MLZYqvylQDk/+oe6GsIJxjRNrhpGZzbTH7PiBbPbkzrOiKYVRCK/k27ZgrvfL52kpVqxy/KtKDh
9iIY03Ie0QJajv9aZPuyRwKTV1+ePhC35ZpUNbLrcO88vC744sDBH4YguXdKBtkZf32woAdpj+mV
WxFedWUSpqRmjO7RiFzXernTsC2YbC9SDueo1GHCZH2FCtjn/a5JkTXdHAZsjzvMmj0Xz1Gwedjj
Mgb/e2upnGF777U8ZZ1ok3JkQrdSSkJCcv8hCewepQLnVNBWxhHuh09xVoMBf2RHpmceQ4ObAnti
2ao2La2GXz0lov1MvYcPWMZFjqh6dVV2gA7Ahd6K3Zn/pdmV/0TGT6u1HOpPEhjwUoU0LyUM18QZ
XAqHJ1jXkWhF7L6D+JbJBPKNyvzDKii3A1zu+lRTke8yk15lIr21uoAy5VoHVHT3axi6VNI/GLHc
eAD5qKfKLE8LVzzd+/0F4X9EM9EHAQNZcRWdY0vtyMw5FaLvuus9SMlcCa6xUrR+/xz8nuFYWu65
Rag/lFhxNEetaxughShjfWrrIi/PyS+EW+XdsuR3uAqoydFAUWoFnO+WzU0Oc621ukzaSkRMEqY4
6sIvRnySfhYBIk+8YedSxys/gmxIMxJaYvewSke1OEtIvDKk8xrVZAT60bm9UFw6VyZ2QUzOHVNp
tJSbC2eiVXwclEaFNr60YI8pmoOA/pLyocWCdGJeGDb9RkcLsqDVWtk75T+OQW3bBoJhBa/3/dHM
QY1Xpcas/mp0wiPRHh691thDJVndqhsnfAKT4c5T8fG71p1SGbJ+/BhKDGqceazWSLXKaToJAj5E
x0VnAaQnwu3QB+hgrgUvKTew5i++Jx9sRXoLSDFqZyDMHuTJMfnfNn5yyiaD6BOPlTherev84wXH
G5w7d8AduQfDXhDPiDcGBkBXMg8Fr9V3IWKtAMNw9k00qSWzFA3iLWorALeMqwtvKZrTAWs7dA6R
nQ31GXq587SahgscubIAFqoP6zCLNwlE8OerbMLjwZqN7FNUA3lJyxEAoJNCLHEIKqasOuwq7pEG
3xhRhfsX+94IkN67VZu8KVQVrB+s0QP/61Z15ESZPysG9b0mMtM4a/ir1OTsqdB8tjWj9pQNBW5Z
LV6gXMbk3eWkV86t+voDNCz7ohn4Aee2MvcuTO2ZeQTdfI0zniae/mbn1zTZwEP97jYPm7R8U3R8
8ON7FYk4m8dp6oS4K3QSMC8KMmKUcc7EgoIbjIa1qTH+aLMWvkAA4UlgC/d7tsx6ydrC04liaCtJ
tbv6gHDP9ZoDHeGrT7VapJXfkFWaH/3d4i+EVA43DS4s5Q65fWvtmW5KkvYb543x0TvCTjZtGg1L
guSL2H24E7omCE7pR0lsYtJRydQw3iKQIfqjfh6lJLglc/Ro4EHmwWZ+4Po1gZD0vuUuAALir2rx
pqEe7Y7arLTuqGSeMf22yXQu0ELkrFb5l0nRI52gdAK5dVVN23Xt5EO/jd2ZmUmbrxJ6jFbI5BDS
v+iVBG3mFOF+EqTZva54zvyy2j9TwQ7Vkl9nONp4qsbT3X7JmsQpea8KxknIAnDyPZFpMU80jD3q
GT4G7Kmk9pQPj8crSZoQWFLVnCM8RDe/1uS7gaH4az+rmWvJSy+2ocn0Kx/aBd4M+0pCpj/Ns0O5
DReLwUPgEeWGgNVzEZwFtYk+FaY3tuxtrWKk1LDHZLZ+7sXviLx49Mus7Gh1Zan6ywtMb/DSMiiJ
2dh0zXmrbZ23iiXsEVN2XnE3h8fNZfdE5u0jOmJTCMcZkzdlltsXyUmPFmCNrNeJLxOVIIhSToQs
v47VdwKbjPuGFDmt3Ql/2eNEfbXSMQKLgibFp6Ak70qJehlmIr4sWCUWCaC1qH8QgP8yPYRLYIJc
YHrJRjeOZp12ndeWsxleN7W0lqjTOBt73NObegAp2cw7Epb/sNN9c6HvN/WAdP0dAR5ClEpqcXFv
PVx7O6Vp+Jii0IZWY9L734eMIiRcw5N9T3ezKMWaG+2BZVp5vx6G7dxEabc5Rb+ryl+ZBYqI8Pdh
sZ7gs6ymmvsaFECaCP3sqVoMOxBX21J/MB7aD1hla8dNGZYd3JPjiRuUdzW9bEVojEm0rV5u023m
msMOK4LaNp5rW4lOa+lH+NceNZ5CqezvZqYLMH15yyDk54vVaQXK5ricpq44bNRW92KhDaa5eA63
7E2LaA24efvyUSC4NDbWO0In2Z21d2idcmKAkHje/HqhWzdhzyarvcH1bqtINgtTIEjdcM6eSKvg
DcaDzPQTXcqMm9i+s7fd1CQxHMh73OLDK3iC3/jaRs8xcV2WGP88HY+DR1tU1Rz3bZdI6duW4VhJ
fmDEiFP6jM5RQxB27v1m/mO/Tvvw/NEnPQRd9/7brHGjx7TlUQjlA6QBi8oDDjesmaHBOg8VJLK1
g8oCRv8GbKZxL7MNwpJ3wNSG9byCMZApnucgTQYoPP6YNMjrH/jMvKm/DWZtEhhRQx1VzSmj3NFd
PVCzKFHbiPVxbdRq3VzaoWcHMYy50VTuyLjqon950Ow4KQk9+X2gWX4fZnr1z/Wjkn73lZEjSmgz
4Th2LW4US/tuJmEmCemUxH9sAqBkU3t1qx+2rhUi7m8GPPWxHCmp602zMc8lCLU5WiSDJR5fQJnv
ju6V31htwSKrrer5iI0murth7VUOTBdfIBuQ/TmumztlBGqzEbjChUfon48WGDjU1RsQYpJMKA6C
vsnm/Cx+dagU7UxZQo7jBeWO4LgxnDQINk24BzW5KDtfa5WF4n//8RIYj0PSWlY49CJJ8u0wUeBL
3SHN13wYDR1DvKmDWbj5JET2JN4vH1kgPv96bxLYEjNaTgV1OXD1+gToGFo4vwrvqNZduCmL1+5W
IKFmDkx+u2YHDSFXqb1ITUHuzM56DpnPP+l+fOG+Ena3IvlYyBXulxES5BVughv1WvzLvxlzbC5l
DG/L+g3oULrwFg6ko4iedoAAbOFi4nySUEB1iIVP5ZK4pU/XKn8GuclYbJXD9N1rl1iy8Q4CreDs
n4Q+R82oOaRBbjlPJ0UbGNPI778+vHJ3dmECQ3QgygFRGQr/VpQZUpvcP3yv6X9WzcLVaXlBjryJ
eEzcteQ7wenJUEdmLH9V07KrpMOEIjxdt7RSs3g2QOYStxzl/Moo8+vfqMzorcAm8Pcd6JnUh/J/
llb6/rJ5JfP22OLFbufJ2Ms6biTnyoa6zVxc2ztimvtEne7PwRg7tQI9vZvWC41/qh001yGEUg1a
affS8UaCp8+QcGPIwgX7sCZVs5ZEuNQ10oxXUKCZ0GpW19HG4Gdvd5H4/U0Z+JwuULzRUIseXQl5
/C3e8XZSwQH5qqxT7h0omJm3jNj2lvkgWckMoLrVOJ3kGtTOEvwpRmkyKedD3wZYzhAbpLF25+h3
QcGHfkSc8Liq/UelRwZoUGx7d/z42QdBYP1sGG675eTIKF6NFlZRwQhaUQUkf19N5CbvLRwfv4hE
ZCQzQqX6pReYXGGGffSkcIKUJuYuwoY/pCoBxvPxMyVnVY+WGuF43lJYX9SABIrbyRynsG2XTEmt
wddZnzVvZ+7K6CQmVMn5ZnbX/xk/qmqq7XHolSQFAoo9qX5Dr12hMm6K+OB1ZbG6r4kZd1aE5Cqx
vT9nDI6dZeiiUW5DSdXaM8e8WxUY8C4exu9RkiWJoBDLeiPuo2SKWykdRBu46TayQmpRGsv0p+1+
I22CKoRF6HmDwxdRDddUOpUw6LLC3TpydHFBBFNov/Z7Vs7GTlqTiJD3LW0GTPr7BgAxin6PtNuZ
yg+EsWEAcrCFJbvWEkG38mqa/JZvSCoJ2reGP0BXQJ2YUKKywFKcUMNesNS1OxQsbaNy5vSK/uKJ
9/k7OG9VXi4To3c6fZWUEfR5NnCl+2Jv8V+jbiAHUNHlkHb/wiS9dr9TcV5TcVTwV5aGkd/Uxml9
isJ7xINoriPij6tSGl3AdpQ/IDNjT+RIPnh8ph74imgueL5q19m9Opqc7nHNA4RWjpeywE60hqfw
o8I4UcZr9Kax1hVENr3cgYYasviKIzK+exROgpREvQqt9w46AXt4p6ZeR7qEGLnLAVikVw605iu/
ODRZufi4ApEjozovwUmdjtNDdzxk5+L8h73mcggFl8bfB2rwA3PC0LvjZ/yS5LWAkjrU4AF6GqcR
U35qS5lSC7dBeHeUFYDioRu/k5bp1gQvyTjtSmuuJ0p+y/F5grhvLFIalAhl/gxXA20PyGvJUmFG
eruTs35Uijs8IHifJ1g+3Mf6zBkoLzbdoCKVndWDrv8rAvdx9a+p4G4tb6Us3RgV5ogKj/Ct2Tma
mQRhxxyO91K4/RUI1R+JlkXWFxVFc/dcVh6Wl9O3QxXwWlqEdJni9JOE2fKoQDYOMYJMzW5s2X0U
jaWKgtVNicjTHFlyjXccaG07HDWIjlCLjHMU5d3uPAy/9u94Z9mIXZKKNshNui7oMv3ZPLnVYQXF
Jm+UVKK2JLjGIki7R8IhLe9IqG4HTGZB4G9GVN3HJk5eoejr95yAfDUfaA7E2/SXUHLcqnFzJTcX
jWV4JLbDKrKCWBw0BLDHQPx0cG7vSx9DrrqL+4Zv65ib9AwSNQYmbewQbSiGB0T6vdirvD6WcL4h
ucRiADRZ6AI1AhtAZUlXwvtUKKYofTgrxyI17UmPdEPlKwKMzzI3qUyBpKrOD0kaua+MqfCwE14T
vI+1+zY1knveI1ViZXcM9+gaQz5yH2DxtQOhjsxVOSWw0GTaZk4ewyMElxkKW1TVk6ZhBjEPxtzw
PjUcNXLPHWt5+h2lsyzycyn69hzm+S44SzuCNJQZvr46RnbGnp3wmPkErXkA0J3bQtEQqORJduXL
aIFTs3EvKvMkNiNrV47PJu+VvkwBl5hHfh9JCs3Rf5Zul/es5vIE/3sxX92UjmNbHRqkcRvi0w7d
Ohgn/oVWWkn92lkKXUGOCFn4XBvwOu6/4bF9OPMYNYW9V5A1Hz0lRVwJxe1k9uUbEkZ8r3E3OWrk
OI3//3d0pHoByDBKkUy028Mbc7YCZ/58lzdVLfS2uihd2TRZpgnDhfgMTxF7kvacpIXi65nmftt0
EyciaefWMhgPpsLUWlPJ6/AWbpclBXvzX9tWaX7syemp4HfQsYKvwACF8O5jLCUZyVrfaLh0NMao
ulPvPoQDIzCtZ1+TYNSWanEc+bkwC24ewMR7DEc6193O3D/VexIkeo5QFR7zNH967zVe/jBVfrZf
2jJqA1+j6LB/5eOZsSN28twCbwDixb9s7hAUjpWKd87ORE8k3ESEVhUQ7kfR1S/fQs6A4UwmReGz
UAQQx9gRLSLOvfBDeuAq8WAKKDMd0Par0JRDBl0tnRG+kvBMZ4MXVfpLulk7khVgDvpU91ZTYO/m
plIXtrmyHpOgVINYf3HD8U8sr3sWTTUGqOssKnncwxsWqeaHZpZJcFjdcAddH1TMIyAgeKWBMvUY
J1xC+DY19y3FI4YJlDHntyfG4VFxF8Zy8ugxbmS/6wTv8t+PZITh36H666IHBnPl7miXJEvakGJe
vX81yUDtDy5WUSG6iMIVdLNzxzZMKVq5f5iRuXp0TbkNKnMFLiycsaJs2Owj82zEygWCx+MeT7Zo
WKLodsSCEp+zjl1Q9JvRmwIlhKeDdpN5s51PPAPJqAvWsVvx9IotfEwlZ9hct/oiRRSULh4OhVZy
AOt7i29cmQTi8Z1FN+sjMJrnpIKBCjgqmwaPTfkPSLGkDEYq/8lbAfeUQi3ejto0626LNoo8tF8S
txBvmsLq5Mt5Dydt9L7Y96JRbnPcYy0Mkuamtaz7oyJEygGskZHHRe6TDfkCZXqDDXhFY7G5SmNv
RNbRudN6LFe7mTPEZH2JwgnlSRchlla1GB+6gEEPt8K7hMa0c3tXwmM6joURtAhby/D1elJZZLcs
CIt4K29Zg/F/D1RkYZf2VjxXJ50fI9qiOlzwnweofbk7t/n/P/wvvl2I9LuFxMmsv7pqY4XKJl7m
B+qku3WEUNaDtKOYesFwNThl2LYou5KSulcGvmL5AnKwZLmqj7s150AeUZj+tZt1XRz6OYS+fhw8
Y7w7ywxrorHRlxBXZeoYr3L3eCY9ZwptdDAyWAO8q/dNAk56CHWzrMicoASl3x6pSd/VOXmWt346
DZXxxFd6SFLPZAqItm2B2KMElINjgQCz+yA/AP+uJJt+94BSCMiXSNk03akyRQJYWI8+XcFld1cr
sZwwiqifWdHjUJo3qYuFJEAxjgVNtPiFyBLS1h3LmNauJwYq7fGy+DzBAyJuxH5vVDcAovBvImIV
p177oADFP9F1rEa509v5de9j/3H7qvi05NoCYeRIEUplN+4KzY1M0f4zXQ7B3bRO4405GOHdaNjL
CfTlz5vJHg4IGGV3GzUeOIXdkmeDc0I6gkB+uOllZFQRfEyDi2y1D2clQRtm1hWBce9/nM/HwcqS
pfAF6hJM7wxxz3z3rxt8v4TW9kBdcqZLi9lavpacAbxXqKCnNhPVKB8+mlMbjD9gTxhBxsLkcLvy
4wl/BLOLYnPEz0VpZCowdfSWcgHKoyWr7F7VdZDAvQ/6bgIzYKVVp5/vNLQdrhUOVtmisZIM11Ha
HLhNDAAbgFnLhzY8OUnVpPX0Nwgh6sG8JGwuR0RPcQvXa5yUKNvoUgaNwqXcVLj+9vmYjo94D9UH
aLmY1nWeMOA5jv47vVgDDdaLlH6EKDymBBBjWrxOiFfaT2Lkr5l2251nGeXhB6zTPTW6M083Nt7M
NbfmuTHUO3sTgmvrnaXBwwyycZYiAtGtaYJ8n+BfBndpsGeqLuwxSUx4JjIE8+f4rhWIElN/5MDI
7xqskGYQjAqFeZ08xeQmA1LzdkyiBSXrIJ+F3gPWWQKWNVQFdF7UfUA261fO0p1lAHyhUn3au7Cl
MlpFmjgG5G/TBo6qvmYOQi9FsNsrAFvFIXOJHnPSD8uE905zx5hbEX8eu68piFXAtAi0/eZ+Q1LD
lOI9QeGlgONIbkor8JxLFqaOWXz4x0Kfkp7vj0wjPUZRb/rEHfYznusPQ9oaA4jvsyRgRbV4qNnE
hhOT2wH47gd1bxl+JlXh9aI5IowIXGuSJuJQ7Gl5mg3sCxzQncdum/1Cb8NgpBlD38OffcJ2bk9i
kFxDU6Bw0f7FNFLv4mQ7NtWu9w8z8G/xKDcz0ykxXwmMOioyws4jE7xhNZUQaf5zwwWE74HJhOTT
hfcALZgkcMWBE961LcP6WZq4geLA3o1wTiv5LBbfWxkZtQz54Q5Ni304es6Itn6qzgrhlD0nVq9b
emUbpujWElamYGBMvRptlbTlbfgLWm7mY6cHYBSEblU0Bx1d2gSrb5lvwZM4R9P2qCmaNeJDNGQr
vGa3U9FFMNTgF7EbAeT+ksrcnOgucShr01MXd2dAvObVrow4Z30JmJ59tNSatqHfHGqb4k7WRj+X
v+2Uqisc7nIRf4VrutZBq48Aa/71AWwIbXKH3kyYMXUkFiiFBmabs9GZ4L4a5VvBzcgXvMUF/n1a
W5ZZ1Dl4wi2EJQ5wIps66ZhDx/xqMNomcH1ZXpw3EtJg7MGZapJzf30Q8JH3vJ9yZJxt6a/aUEsB
pbz2rJfvGlWtKtvpLBm+16bUoIWZ5kCWX/XzKa1huU919YXdFHxAqSwBV0pF8TvNsq7AZy47cyZJ
hAo0cfZuqftuV7doupnT/HyuZ1s6ndd1+2Bx1yMftZwPNsfAn9u/LSXH26l7SfZjG0ioxVF8C3BG
HwSKE8l2jegnhCoFLmL76pWopg+q87m8+jw9O/n8OhHrXzoD8Ot8buS1uVPlo7NLm1EDS/LZzGfH
V2vcFBcR196jVPlyHkGPkDlPZwn0F1jMhHbUHN1oULKtt7e7IogByROpTdzw1bp0+53OY8Xcgi3L
3e9LiCYDQS/jQs+8rcxOzNOgNjOMuhyv4WhdCkT8sdtF6uI8FmeMHXCyyyBOVEufTLX6n3h5kwTP
NjkJNxEcMEGIVr1ZKGFWNTc0qDCMhWG7WxnRCiQDqqzUlEupik5QFRlSN2sb5lN3fqfDbOca3bOK
uHdABMfq5spw5s5AaY8si63UQuAc4ZdHOs/qDf9uF3WAOZszKpy+y6b62XH75IJ+Qonbw4tnUF18
jrLtsPDT1XlRszNcgVZEjmQhoUwg63ld84ZgL+b6wqNBcDOL+4kLfXpo/H3JXE6rcquPe79JVzYr
J0GjHMojAuxV0cgbkOdttZOSPjyLiKSqu2f9sESlmtXg0vUPm9Us2lOCNEVNAhSS+7Hubwa6GTdK
KW3mq0Ve55twDVmyuMkl2p2qyBca03+TP3XgitpLpUh6SBjfa+Z32tImJDvyzWW3p8EpvRkUyeYj
wYdhFuz5vzgjEohZeOhQeudXda94+hcv5kJMbsnkK87te5fVaM3IwoV/3If7ZWupKGx9I8dZV3qx
uDEewGTV8ukaR32cppX7VK5NjwlatkExjjLQFoG5jc3m3eUqhRTotl1xMOtvvIZiMGvco7gKdkil
Xp14cbJpYzDRwoBDCQXCzVPQrEjC2GMYYHTBuVGZI40hZHQXsWynW9InV6/7fdEHQbd0Kzo+1kE6
25OO4cMcyH04cNLKkde+peB5g4klK/X009RWqXGO0/jziPcqVBbz2mLy/ljsnHbVeea0Xu2CsH9l
aUUy5KNe1s24RTKu2olJleB2iaTxyBwgcFVWPdtfKn8bTu+DmGl9PQ/F3jljGIIm4bxB8MXz9vdo
JF7olPxm+xBT5EIEYxf3dm1MEDnIYuunWiGfQZqYaYyYd6QlQZGqQ55O67t1Wp1ZKmeDNKvwcOfQ
maFJGddbMts0heRK4D+8IKalUdH+VAUtEig8m8NmBab+BlXSF7yE1DBGXtYPscspWUQEu2BwflpY
IWRJJyn7DIFLSqGHz33cGdWZr45ccokCIUVn6P6WcUECfyQIcj5kPrh1W+ycC6VKN1HbazTSXJ2M
wMPYJxRBsxAtpV8tjMWNXzZcKdkk99eBLUk2Ycu/wQgB7vFoWdFj9dAsBN1+6MR6dt66ohCw2kEw
mibvwPgw1ky7gmgUSz5xAIiqc3s+ng/Yzb2gVvpNGp/o77p+ioWY9/Tb9frLvqhFH/1dyIxRvIG1
KOSipf5V3kumkFJ4ZiXA+DQPdEOfRtXDdWNmGed2mXStsNFOKbCv042M0qfMIi4YranmmpYRTJhc
gxq7kxNU5DqoOwpw3xEpT4uDTafAKFnpT15p/CZ7UADyPznMtL+L5OEGoq/ISX7NL+wpbkarEqfN
SezcONm03p+Knp5iTocE4LcXtbT7Hkt3uZ9Ky7bLjvavwiVFeMhVH8vs+7GPqU3EcSS4CS0qPn5g
17bZgXq+it2xl27f7Qupu7riNWDtTt84gqUmDwPoGh76IPki+slQv4IpRLRbHKU6YY2K/b/ZLzh3
kDEZnLolSKfzQ0pprmM8G4wixkECkJiR8yfiWuyUS7/7grx4Da+3gT73wPFmmKoH1oavB7MH83G9
HbjdjDVJQjDJdRYao/nKzHhzslWosCkVy9N2/m1QV1omik/m/HYl2sQbEb0T0T/krnZz4/pt9SyP
OEEEZtrGjN4/rf/k2J/snIFOOwLoQ7hp8PBQrUPJU4IKxwWfDejkVF28Cyo7zLLpaLCWi5zjcQ69
UO9/Waj17bdD3Llc6evdjmq2MQtmCNz3rVFlFlUCxyzSt6fWwy1cOVzy4n20P+KHng5pXXL+fI38
0YVvM+iBmK8AQC/M52shis4vU6SGd7U/A8GAW+xigXATXasWkcredCCUww1EQxTbDFPKuROaDJiN
xnXbb5i1fE0m4huc5gAQ17I/vgq8Pk27l+1MDPIwR1L7AYjdXYd3siV9pC58TlDMOFZmdNQqveq+
ubtUJgo3fwSO6t4aEVY8JKeG52Azl4yWjnV+urgksqHHfDflHvsG3UDqJuBmK8n+dHvuktpW0ccC
REZ1jPcQxMGFaMgSwOHD6v1DEfW0ChoReDT9p/iLZKnNUZ0lP6XqICivc7iHQZw7ecRbYPo5zS+L
Pg4m7egIuPLLlR7aK8SMm604+uHd0kb3IBbZRHbW/i9K1dZXR/mkxnW62SUjHA7B65ymLn1iS4Yj
Po1bjEp19FqJgRKONtW81yyb1mUugf8FeIxAeA+BSRNcp7IOI3cT1ZHkOQZqnmJL4h1En7uQONy7
YisJb45kFFOd8Tdmrjt654hH3I4kqhlcF7lkrmKRusns3Ayi+Ru4xYRY8My7HH1ox71dfuidqsqe
4cj964V0hxertzCrN6imCwiQZ/sYXrMc88I2rnbLtnfgstKSgGeRjUFYB8FChblGSig68nTQhCOO
aJJxpgob3u24NNjinOA1mNI4fo/XEeG0JKJ+eBGIIcblNuWMyTCDRt4iVAPj+AnWu6yAkfJhWpGd
usy3DJZqse/ET1K5e3Fy28xdtAPo/X4ecl3FFy2cFDJR0gVesD/x8tT4xKOirYSC4FNp2NXcChj0
s7bJIjmuIy3Kh3PEVCEcJlF4+mLB6ej4eX4HwHpYKuSnY8hoNIv0zzFRc5qE1LJQJMM0qPRJkuFD
7qx/4BKta+WLQob+tvaR+NT750XydP5UGLIdMmedgDC5ekXEN9KDMdl4IFKRwy2SXtbqsWkXjT/V
EYSEv75DzCnszJ/CfdmkAQw5ckIfdW5rX3U11iuCAXvzNDzGUQ2GDI3mB278/iquYGkENIkQrlRH
jQPwzDLw8l+toPf07ac/GOxCHDk43TSsuEsymjOcPQ0bioDiyabOeUATcHDAVjDx4+bVvthr0L5t
l3T3s+RT+0W/Lgx4bbMSHYitk8rPS2mJgGvS2kU/8oFp9t5ki7Kgy2M96WaZpp4L1DevQzpoQ6jL
ecNwaUvURPgJn9h4VHytOukPo2TJOFMEBsj7+GHhnLgECkotH17ihNuET2lrq2du/0wuW45Pv4Er
N/LpCZcN1pjOABw08nmqQEk8+/aCE9d4lx73TDC5C/K8fZarUWg3GJO0aMTCRAmdZYF7ix8H148y
BsiIllYge19Bcg52Y2pFYY98hBAQudLISL7VUodB7f5umR+Yz2aNpC833TOwWxOhKlZPbPNdv0gC
XbYjaEkiqYQEeODvFj7wIubzq1g/PAeTK7aff4j9sr/LBkz5g/yGNYtcEwKSwAfOyKAMxAs9kz1G
hAhx/avGNAANGun/UTiKRVceEuPXudhTJqoqaBmbKjVg44lWlxfZ2u7wFwrMcNi4fn8n1z1CEPr1
BfM2Y1+7MM5gE7Y+49RwfBWty4px57NIvvnp7hGOKGI4B1XnJv7fDva98v1YM4+f9TaOcHq6o4VL
ndVShd0KKFJNvnv3M36M0+drbnUSz/BSezNInlcli8cpf5iydwZsBAY6kcx7TmH+cdFN9wLT1yC6
7UyXsGMamJK77LSE2+Gv0eY9MQ38N0J/8HiE4BAZp+MywV9mTZx3vwhmDjw7CurEnXFKD5VtrgPz
NfJgwFfrSgZWWqBNaceMFJPyJjGDAJCscdf5lG/ykzzA3GtC0rtyXa6hEUv8+3FU+H39SbXgro81
/YdkqiCcfbHNxl05K5toPTvk9n/yDHlndc9mrPpzntJysjftZmTLQtBXaHHfPQPZ7KTjQ2xwjvsF
H4kteKJR+Khh3XZjfhcZJcPo0LFEX0e6TJS+VJsgi7dsl9Dc3W9Mzyu3zLaWKHBORgUluvFHNLhX
Ykm18BeYQDd9D9jgg7oveWHoKW6F5iemh8jf2T1HyuXHerno2/jZJu8dUjHESabA5k8yry1Gv4oh
I3MHTFY2dRsR/Jai7VlXcXPr8yne6PM4Hw7IHiDAVvFIKX3qg+0sT/1WDWYI9nNazKtFdXZBnQpj
NN4TVftRW4KmwfFYnOhevjKj8Ki6AdwSosupHQIPpdWLdlDctsa90SURu47s2VtOjnq1Jc2loTOt
6pTG2KX9Epe/Ym0uLuljONtAjbdaZaH94GBW7kDbUDvsbD3DqWIC6qNSoxgVrTPHwrdms9jnzDbc
R5c2SB+9BrpaMBBdCKfPbxfPRp64hT0cCnwahI2V6bUJrytnKh/Z+w1KizDp8Ky4TgSZCx7CB4ZD
wzR4Ov7frVtgUfH95ICd37OYlgznhA41ZMASvZQU8QPiZlFXf+vMeC06wtymnvsGQHj9ECFKVIAq
GsgxVwpXwXqyDB6wpvTIDfbP+7dQsi7s237mT6XN8eMnzx8GEiunct1KA9b8GHCTYc53hCikJFV2
HuvmOSEz7thdElaKNY6a3R/wmaaOcd0T3bVyczFQG9sgdTBXRzkxWomlrhIb4QbXnqEywluHaD0h
qdz7OApPx+dW5KYh0FDfvSUqZcnSlJPlxgBQXQnLl2nSXZWbDRmUhD/nqDQ/I/2EnB2uuaeAb/yu
dKSv0QSzByAH2sebGqCxvBTL4X8GP4Z6KVIrzpp+RDGJ1Y80RJD2L1Gch8JPu3c1WKwGM1Hfa1Cc
kBe0356E7Th0LA0bEbwttuWrbLTMlQbbhyEY5Fyfocp9Hot+ti1RyjI+tKzvLhZOI+faM+K0TBnj
pyPkI3bJ+t+S9Auv6NxFkdoT+G66NT4AWLqx+Ssh0JGuXJ4aLh0lva272dAfnnRvtiyooso7wdON
p4/VG4dT5R5GUbbu8GAur3K2hYtaM9PD2+NoVclx0yz2KHqB5m74lkHeZEBPG0+IRpGx8Kzdbq/V
jpnz98jfJPRNqQAyhD+xBkjgsq5Pr2rVS+OhLhf7iHU3GlNTZ2EyC2pCnu4IEb2GqijWTEuJoR1E
JS0452XmB5uLg54CwEkKWDc0Pswc0d0k0I9/TrQlxasHWRJfaVTft7J6O/HLs4T8tAQW8wYU4AfV
QhW9r0ACLCUXzz56dNWuE0PHMJ1ZpTvP9Ge8rPdZci72yhjEd6nCGxj5nGqGtwrY8Y5mKFmfUJE1
waz3fglHXkAjD0DpZiRcsOlf5jfMperTXKhPQcKAAbT+EiJWvYOBTXac2xyqHYj6KaXdokpStg5l
qNgsSc6tNWM1KptEyEgwDoRMhCN+Il+fDcuDNLkltgokY+aubzFRH6+qiemw9S3ciDExUOB2IcoY
mxIn8xGIvctAUrd49lbblMuQVlJ1LhGbgQ3rKEd8B0aLZFvePC7r0Kkq9cPSNly4ysSQHTMqwKbk
vls3iInvsuVrawOGxn6hfpd5SsXMBgQsvsfZeCl0Zc+AUXATJ+h9R8hq+hFPBKjvtz/FwupS4NN+
Z006WJ6bykfr9kOaPHnlfr7EHphJWW2FrmUTpcepg4ffuT/l2BlNAEgmdgt1suHF8mEFikegMRvv
4lL+TBZIiexUtYZyCpLx1ojqCKSb4exOiktrkjkhp5WFhJwqE6+2IXTPrFJKc7ipUAxhA6Xwme6Z
l0+2GfiXRg4bkDNGFl7tktcgnmpxuqh+XDEepJczb6fRYG1fqcgb6nschyM90FrrEzT+fynJnVv8
+lXgi43mjFuHTAkUHL624+LHJHwbRydCPDR1tXevo4vFzWslrvqYyYLQbOrr2vEOGBCjLG4kh1yc
PtKVqttJQPWdrk4VcHSPkJb4m3dWh/JTqyGskVNm25JbnwvCsFkytetvwIQUiPIMlRl/pJF23JT7
DOWojSkJ8+ZkDLSUbxp8wrBOVWsf1GN7PjuuD4asSZmqXz9aOTHqpX2ftfQCpZWcY5I1unTY668H
RIXsU88SWwKvJwmggu4Ud7WABV5rArZ7A0UcI0lsupXxjbSUPjCAa6J6PC5Awsj8tf2nahei5R0N
3XuVY+2YvU4OOnrH//FK2Vkhok/i3wvhTPPMiSqdE5siHIV9SPCcrhvAhBDWRotCcHE9ksjC7qF1
Yh51hQjOOgEKwvFrh+DWZjLmtzoDvZGuFMxpPshreNd1NB/mWRHXMYRHMzskPf4Bn1gFAAakyqeO
pmZ7DQhi/+NtMwHSHZCnDGIoDspOTkNj5aiHlP4b2r8+Jyj/qV9ibrQTzeQVjvhxRx9nfr2erhHf
TfuUW+2TrWYJ5hO3Wp4dyFFeD96VcYF0Cxm5130anrJC08pCY9OaEBlVx5L729yr9bWeHzXYEa8v
SFCk0fzq6Jwbrhut+CbPCH3Y8+UFrDqrl6JXAWJDT1IeAlPFQX0MPc/ReCgiUE5AOrB85F6U332b
TBc7xlb50q6Qv6CqAT34/LnYmWM4zRfQro78IXkBwRaGHxMuSyuplu16MWSXJclOo2ou4N6pW00W
5NiKTDNp7P+uGM8EXi47aKDNCiCazxBvbTMloRlPEDDQ6bV4PHnlnjcH1r5HcCv42VYE4R7qJpjI
33/YtgvgevvsODV+CRtgSN1mNDowqv5iku75NISW1iQDbvkJVcBeSvCYdUkGY/rYy+fdI8RVsoU4
zjlPucR8DHyx1/X8ndFaBc8sysRmA+n6o94NqPzlPtompe7LW8ah8ODp5upnOWyimbzXceCaK1Cr
0ixlj+3vmUlOkeDd/rpKRJ1fj0INdlnfahN1HGF9X+UY0sJmmrdGxezag1Wu4XqX9wZ6z2g7GUnV
RfoNSDEtZjKpWAexZEN89YpXBM1DdRfRA5uLFQnicZAhaF5XUFyDC39ZTCUaYpWwrcO/5ZjhidJF
bFOMAaJPVsXIBU1rlfri0vCkswLxE++51Hami1UqQwdfJC1oSaX6kRrI/mH9D4Ginj7u9jCc5nDZ
zeLk5Ww/lXaOYtp6KGgsDcjq4pXlRhuCj4OsV5pFu/O5Fxqv4uPlsBO/VWTRZlW07L90nk+KSToF
a6jfhZLkrDFkKTvzb3/UWhQaMPxCaedwDRRDgqqddsyhcH2dwP8XMfYCkC5T0YIJid/dohs6E9Zp
Xe/8HHu4pusPTJnOB6QqGfUjdzV2LN7jjaRqW4Menq2EcjMJrHScSFa+iKsEFJiNLuMh/P4sSeYP
3iVPAkzBKLl2iiL6BRJVjGbHUG8knPwvFQQBcG0+J9d/N4zeIGQvWJfldW34qfnvsv/A1k/rY5RR
pc4kX1WLuEKuMmWhMIsTE0LuTE8BAEPp4BB9FLL6MdmldPGvUmjn3OXy42hVM1XmJ72OOy+u0PGz
NX539OGDUte4tXnFWPWUtDmVibDp5X17WeVlod7tOmz3Gg7TMOW/l5EZ/MzSubiM6IxRietzD9Lz
ktXkD0ETxAkw0An2dCbP8F+MBKqEgU111LOQpl9k8m3wteUEu7isykgwmngrWl6+dFKcd+zP9RA/
SBw7OabXDH3gfB9QZwpL2iMVm+9bpJE+1px/a5wYQLcyD7YkJgDSqs+lPaRvsoGRBx2X4cZelzFu
Pr4GYkWDsOco/LQrrWIQojXqHTUROtu54YpSfSeqD9GLRlHWZ1R5TJa/M8MSdphVNg6wRlRfi/ix
BI2UjDqfDKkoAcKEWgvx10LqUf9632bCH0biURfwHX0DthA6zkZDGTJKHJdH6XCvQXTP9t2Jzhdc
fBJd2g15siAaeRpfidvvyn1To9lehtOLZNVMtwhHxGLJ9dMLiSoVh5YyMHMlv6/JeHroncQ2K9MO
UoDNRQtar6Trbs5gtSEovuwEq6BrpoxwWv0KLR8v5qAcuWDhO/5qJWre+L5WbpYt4ZTs3+nfbFWs
vM7DKA75l1Ow36q6usRqHalXb3f+tpdbw0pMe6xjYfYG9K31uJLiHLs2L97ZF0itLILd2bG++2jK
WKZ6WMHVNW80yZ5faAr8t+q3H4+q5YthL1XkeX1h6w6+s9Zqd0BpS1wvN3L4mzXPe4yYAR/feW4V
jsTFi+9puvSRPzieIbIoie2lHpAzr9itxuBOYr9ne/Q4fCk9UpBxJHHKLFM/IBtMQYJWQsDD144+
y9aLL2ICf6lzdxukDat67wctzlyxS5XGX6W++q4DBZiWy644Ac4fSTAYvrXS2EAJAabYWM1OgiUO
g0JxsrFfK13vGcc+RWyTPSxn4HefaqvBhO8n/9Ux9ol+jw8yxXPO1sbM2ceI1d1ttiOL+S9JOVI6
ynzwly6lWL+mIeO6TvPEFnby9fpwsnkHkC5XRWzwqzaXvUjzvvCU3gm95eHDCcNojFXaAGePYp+e
cxgDfvi2Ayho4zdN3rs+zCjQ0yJUVMSRiGMSfPeW42I1fyzKP1N6lcElLYd4ErFXc6gTjzdtMOzw
5wGykuPka05hjnWDl26yCc2TCfl678EnHm8ycUpnQHwRxGxlgAB+ANTplCzFS/aeRGQrKjrExDRn
IsrJ7cxVetdNlTq46zIz5r6bxmYkQ6nxbMjj4H4sskjy6GIPqrjH8XfaeLCENTgkmAwFm4LRgkf0
W4AdmHbpXNrixgUCdKbcvRP6Yt3nJJHhCZSwlaDaOGE9AjNWLDWG3U3tyoFA2boXdASBhQx6yS35
/YNUoBZcCiA+wV85bQuQoZO+DGuxI6tt+OJZYd10tO3ctscgcXnL7qkdb7v6Mc0XD/euD8QhcWMa
G0nMt5meNvm/9yVrsHpSc2tRiUywS7t14J0hKL3YwAXPBPzp2Lza/qHtLjx9Isdd4srjtKZ+RAEy
COdFD7c6FSIVVCZlg31wDCioKK3UVifzcL4/sf22a5W+BlqmHQXLo6AYIcmQJS6C1If/tqdFdA4G
LdB6kTfE9ipQBMk7i3L2EYNjBF5xrTOBfQ8TgCe8mSS3LzH7NNSOWZqKY6WNquzO9i3RD6kc1Bjt
Y3UsByaKNP65loPLSS/AoynB1OKiBOR3hWdTMCp+O9Va8k1RLsoj5qK0XtU1ayabQa7q89we5ajm
YB/jsEhhzjbByUXe4jWjYfrs8nLJxiZTr2fPD6Jgp7k7Yj0GrJTl0655Z+CCn7nG4q5k9pfEZUNA
F0X791myP11GYW78P4dUQQUyBW79m95sKnH7pa7zuAAT4+ztRCYFa90qvd/0WHRKx+/JMK+tQIJH
v+MgKvIdEiY0HagUjRgkR1fcApkkIQsLvJW4zKt6QaNMR4yBBGu+GiXzOwHoMTovQvbnNAgRZFCK
ogXYRwGsu/Rm3J16AsQEGZSzVoboRaLeSWkQXvqzjRpaDyG70Kq76byaeM1PPBklOeie91DPla7F
imgV/oARueCaAPx1bZoX7TQy3AhOV9tOVam3Oarw7303Xu66Dr11L5neBUChgaKQte+eNS5V3s1Z
eosFcDnHGynL/yWrNXACCmyB9VkXgSwh+S/w0VutzNhHe6KwAGCCu+jLF1doFnypPi702OM6h9L3
Xeg43uq2m6J7G2SVeH0lOtI0iItxAMgT+VNwKB68uTvtksh4cOU8c5jyGQ7P5Pw2Ul80QZLCcyRK
Fug839FAB3yh+d4aTo+5ErpPPqC1LJLBIp24B0lv8F/IrclqNHgPTd2yRJZoUZTT0iRoGEYQcAxZ
P2BjB+0r2b5BIcvTCdeBQxpQKMZOIMLRXc8XbvueXOsf1PzLsuvS8t7fmm5ABjvSQkzy5wJ4AHrw
SgL/ir6oxaQAObenx9a2pD1AOhA4LgnW7qe9W6SJgXNCDzO3QdPIt0BZWgDPaMiLzXepn6oda76q
T7dlUDBTovq2GvYDl9kEpnSjqw5DY4md5GS+n6IxqMwgQ5dnGrIXzWMILKpEiSGl1eJiWzaeTmHw
aluZ3n19ZylStDSZO1Y8lll7JYvZUDNkDwy8d355IRv6NxXm0+2Vy+kwHQUu5f91pi/clpVp4uGk
p+4frzM1Ct5Gyj5vj2GAyVdG+TahuOH4+CLwJZFf35p+jHWTE8tvFCl8F3UUSqbJ7RgvpI/T+yyw
Drcv3bvt2s2X7k9kCkplhKZ1nVKq1oZicDQL9hP5Ez3QlBqK0VWgo9V92xmdMHCaHR9DvpTU8e/j
ZbtEeBK9dsOIa1g/XJfZkqV6CsPA5xDIYwKZvE/Rav6a68w9VXKQz2E2yqzs5jPfspKnEBJH7ZJ+
WSX2KZVVm48BcpNunTCKCwR4JqlTOa/Zy37YivYTONr7zbqVsDo1On4RRrbr/NoiSYtoz4rzrHpC
bHYtladN2e7dhd2r274yvmDbo8NomPzg6Ak59owbz/DtgxXDHhhEN9jdjh1ffmzFBmU4zVgVn6zk
FvRi5AKRK0LnUKmdgUROa9OG3944kL9jT25ule6ARQnHaFqEF+z1F7cQGK5CPgY9OCXqwyDQZ0Zj
zMT+WyqYcrigTRlZol++ZnA1r9kPy4obWI/mZmK38Vh4zVB2avh0h5+UJAxnuBNFREHgwHkZfFjn
pJvuGbTttpMHn0QnFgT78JCNG06zqDO534O+YiDYSQrNmL2yI2RvBmWxUiP8Kpe91FzOH3lwmEac
SWXthPD9SbK8SqKos82LUDZtiview2PGhoqiaZmBCUsE7+evBvpr7MYuDeBUQ3bvUZDBh/JC7uYT
I6BawPqxQ2Ak5X/retpzUkYIbnDu3/hf0WqanlYU7oEBrwYrSwMTQhcz9GVx9A8KVWoxYaYpBpVz
6043NHDRMZPnBw5QQrec9A07V2Ye0CKKSowBVqT0ktI5mOy/pHNb0yzCLOja2+lMI/6km7eb3bHp
txnCQwpZmeS2FPmFNHL6M1prbDnPm9h5Ax+sTTtV+ZxEaRXsDI11p+fLUxLWZVeWpMXDHtf6cuXm
KXcaKJ6O2co3urUdeS7AVg58fykbxL71a6u6j9YDpbIcVt1PL0m7PqznIn33ftUwh7473C9a7k6l
OIVNv7htz+YIj9iusps1ViG1NcFzXv4VawiFvzUCsm6efHxtx9Cn55Q+HVEtIZepFi11umQ7TmCT
k5OG16FBo37Lns6UrvEsj6M5wZXL6S7j0S4w7O96XraZ1Ief6fQCEoRjptPts98hVcR24QYCLkpk
mpNN2spCJPBbwvlFOtyyGnFwdBu72Z1h5sVF3BMrsV7vLzM/O18Tdagf0U7OJjfkkYMGgajqQw56
pnLlRw1ub4EzZFVMzXeobh4UWg6QjoBL35KA9fVGT4x2CBzr85YWkv23U3BadXvuQD4Dv8eQW8Af
gPEr3p+ug59LPZlbNk07NrdolteRNWN8GnCUB+l/abu87xkJWGKxI8naY1aaqQPVPilyFId1s2VH
CH7vlGjJtih1EIPBzLIW598bJZLCqrxsEcS0Z5iI7Kn6ffSxasYnYSptUGzbOUu62JN1/WOmIXJC
iq8kXcAj41pkayhv5HgCZwGybBL2Y86d07WauZ/oY9FcAyJkm/4a63bkUv8HUZBmdl3hvquZUSgd
eoxx00yk3jszPwpKjT8nSCpC16TSafkWxysEAQp7VzDLb6lV7oHbl2uBv9ME0HYZkWUIx60e26z1
o9VtBQ9+NqIiu0Zzh9gvjUHH/gGq3eU5x5qcXwGi//PDfwibfUIQgcASuFjQNuAnJNd/B82Z3dDc
1/XS0xlARrvGw3RRiJwwmAyZXw6wpa2rEwv+44hdLOp9p0gHNXh6ie5jBUHcZcVrXuomFbJTCZSO
pL+lcYyT/ShAOmfiT5Gdn8uBj9tnFwTPgE2NrkZ0z5sxTGUQiRuEuBXofR2bc5y/FAOTZ/olUlf/
pRjMr/d8drYSO7z9cI8y1OMCCdq0vJ5Iy0Dok+7wFTsnnjDc+KhGLK7fUcdjuN2fxnT+yZaIF9lL
ygbrfhkrcJqQxrjsG9dbfzFXcC4xV2Nrn0XJnj7xx1g2ijSZNuUZ0ZtlTMA6oyyBRPySMtaanP18
0o3CniOd8I/5f9NGUI0hNN9OGao7sGRNdpqXLwqTgTABhNXHn1AP7ZGfh0HtLNWqy2VX51iOHZKn
bEJPqq6RERFBkWqpODb5krMbePacwcHy53s05PWoiFejvqcLKvqSQ2pbWAQViGDSy1rbMto5TrPw
L00MrRFyakK+n4T5xXVtDqBbMtSZKYa5H61CqchAfxrdhVfPcQoae9Jd6AsH6TCzh1SF6WnD2iSv
/mWO4lYCpGMV4PtmW/BY53eORww0WRBAhqoMXxcU2wWHkZDYjzskkhTptXO9jmn8NkbLD8t2Mqjn
XKhUtHBRDhaL5IRInycN3M/cFOE3tOqKvog1WjvcQXMQQViUKUU3YyAKxadzm+/fCPQ0NAbIIcmv
WLggLAJmlJOOnQ5DNqno494oIOumOgZrB7L05yUhV6+lu8uNSxm38I9P9xkAh4BH4CVZElMDGHPe
8f8u6QPwoYp2cXSY9pwb9mDzFquQnmPrhYVR5WvZGnUUinVfVm9lYMcSWJYM+2n7pXH28NXYw6kr
VWL4b2cdm8ptH1cRotHrOBYe5yKDus0WTPvEOwKDimVWjmR9jr4aGp5hd6uJuZuvCrI67+Us1Hro
N2emYZOV0N0Vi84vM5bsrbPh4RoIMq/38Op84ohXf17x2p6NFDhHQZ7+XhaYFKRuFbzJ53Ux7eDD
5of40Drwzdv32V8oWouhUTYWBiv5lgk793uhy399/UxjwCOif9RJ1jjV2X2koCAB/QxCNdl92rL5
1egnPLDVkmvqdSJ+rQWahauz7YenvtSORjWb5sH8nyiBKf55rA1glGVASHkRPKEMQF9X9N558zWZ
oS5GrxWbLukK+PQ08Sz2SKKqD+DX8dzC3nEbsRneSDMnJVmI3/RxRaegIDIncV8H5q+70z7xTQpJ
bIXg7WdYl2TIGmhf2TNewBkdMZJSr4I1/MsA8q5C+6hXaEWmIG20WoDNaDcXZy476Gs2bQZAVtqt
MKS+cV2BsMyKH8X706834litwoOUxR7lS4k2x1ClB7X+es8M82chrXIHo97mTqQN2M5JRntSDXWw
8kcgELkawovYMRjQoVR896MXkiMXhZNqG3bAQRDv0uF3Al+IonUmFyyQ6OxB0UTL/lp6W1OG5UYZ
PoVsxGjy63OJD4oKurTAB6UWBTWYvOsCIzTHRnUy3GdJuprTHY7mt/iq5YaDcTBmC5VGWtyvJqja
gnOv/7y6SaNfRMrzlDZOze8M9pfIaz6AIGeMoAEG+sISC9OFWXPqxLEFL3d8x+AbKbawl0NhdqQ4
IDpKcQrOPleUnrxrREeuiCyR7PXVvrNVaNxZoLdQNf480v7Mpsibt7XxGZuFAZZfPQ4p5XiiIJKa
U0m9ghVB9ygEv6ysZb/Q5RR6u2F+55dlZRY8neR4aAUlhrUOiUT0VAvA9HsrzyPXF3JvFUUXGztr
ohG0lQVAmdOjESIwnRaEl9E7e+Am6ioV7fdV2rYBHgkQFdo0mrzu/XLKJ290zzwQMUlsOUMLiPg7
oOhhj0Y76SwRQbjNpUvOaAfpxqbw4aWb5ST0ZQLxOB6zPl2F/ZRkPkB7rD1mPrwZJl99woqDSTLR
vzH0tALQ8cP8J67SECriA9i7nPb4Bx50FebuYd2Mj/rXGyKeg4JsjuyyjK/sps9zFB1sPTXl8hcD
SuPNSBi2aO66DknYuN9rWevrNar/a9mUDm3t4ItxSQ8d324h+PyPlC49Knhbm60M18XdEDUNKoZ7
ocdw7r6wkfDZ6XiX5gdmjGpOqMS6m90kqVQtORqSV2bnCPxs4PRZu8U4K88+sgwAcIXqY9qHIULp
rP2UpCb2Kn4DHKDrqPOJvm1LAsFXRCve542+VQ83EmwJ0ziTeGYlEB5jQjSjF/RP5dEn2dgbmuML
zuUg/u13qGbNZqWqPCP9TFNwD6fmbF07FNrs59k+lL24bDPaytWbq8zL+S+2H+L/dFdLE1VL/JSn
z9eqS8Rkt2jB8mrrMk/LrhOI9Lgw2tdIQsUCzNjnT4+btHhoQQY7ws7Ueh4KkSjTrxTk75Mii5/P
V6H1xFaVMK4cJZPMkvwBrcs3ObFBdHa5G4HutxNFXx7GaTCoET8OTMV0UuV9vMuXMxA5rqU+TUw5
XLdFEIvt/L+MKTMJND7acaFNXJV7z8TsNH8LNJQZlK45cMscnvZRKQjegm/ESfRhMPfv4tSdqWeC
3LKqOIApJYEgbKfvVAQNrxQs/7BgHhMjD1HWbBcPwnEqS1ZWUQv4LDQvOzLJDdo1dFvj8dkrwzHQ
FCHvPOIy5pGu567sdW8OWuCmwgNmY4jI8Vb6A1ntxJp9lmg8lF5xazfP5vlkX36Blztr4Kx5i2Ty
O2rQs6UT8ALaXhKqBypzA4/3AZnb1keT3abnqXWIUktAEVu3yeWE5seywOvgAgB/P81S5DynWQ7w
p4ngCxF2WOGdLEAKYkGfiW7O3GwRxm9lfA87Xwo4rOY3TcQV9HHkq2FFEoFJFiya3tjvGj3OrVBA
5jzy/D4jBncfgg2N0oXVZesIv9HL7lcPSPRvnEgIs0vZgH9sRlivLgqvUZVMaIKJwMqswiw7z59b
Lliz+eaxeS2DTzg0HaW+gfb+mLPem+1UKto46glza4rvZ9xHeigwCwX18W43tU/vfxz6Nn3mSFey
h+xaBFyGhxEwAyIB7VgIJxTXcVI//3hwp0h/+vuiqi4IEO1RmDa7DlCyk0GAxttQFWUv9mAJEJc+
dDjuN4g8vWfezKtXrHDZUWEKRhBTNmcMrO2WPkfafRcOuwVCGaJNxbRckRp//5UXu4/C88+SVJr4
9Mt05Ag4kbXgYEVFeoHIhOYkpKo4oULWfHEG9bCQ2S1Bo8somunVjB7qzq5uYkjW3SsaqeOZ50Jh
WtjnDghGgd7BVbVMuTBLSXc2FKdvbXMQAe8v9XTdu4CKdCv0BFAa0OqvRMQD7IxSSa1pynw9Lj+Q
wCt9GFUrRphqTLgAd8xkOGlSlHjLCMGTsD7PQpWVBulnAVELOxo38W4n4rk6Y+M9sKQ21D29aaoM
SS1zT3hL5dzoaBxWYGVjqhYS+6X1viJf2ggFEZFAosD23J1S7+VOjIlXRvzLNy+jp4AyvEi59s1e
ESgFmG7iRHq3x5mr7PgOqlZnXlh7JxTR4CC1geSkXvtz762G/I4Uxb4+9ydBt0Y+aCIfYf4npvgw
8IWw9a9bJv54TsQ6U7X3ofEeoKG8yW9beQsRiAWO9ZXJyz1jeQeExvNH1ixarA1tEGlt9kxzWClA
FcMH1eIbsjih/DLtP4+72WQVwzbCGnYBkxv2kq3sbpCcJeiajqtG8+s8saj0ZFxs7EiEVF5n9R2B
kzLG5f7KdBAgZC0ou3+Sq+DT9x4FzGHWy3JmCqTSNFb4/uiJbyiA9k4eHtOBu0PYop9oJ5KgUinE
f4xG1UyWAHnX/vBKz/hSoI6D+2ERDkdiw2bYKjmwKMnTRlX13pDwNynwiav9EuVeYI5JJYz6PyMv
7vQuRESHQJKOpXG2r6Nr7SF0KwAFTg5Ukbx1rXMoqAMLYVw5dLRiiL2OXg2u+RJX/L/EjpX1TFP0
2wG4sUVVCAekRcX41ccqa+NyduMjl+prjoR15sGCa+9PnW4m2FpCmTu9ZgUCp5M/00UTRynj4mAq
7VmW3gjhhh3HBk8N9177CKC5Weqb58X7Csro9ylRUvBsXpjg7WktwCFVyjLG+OhytDnh1dFqFq4C
35L6hX0EEBnLOtKTqwd/C39heP8n+x0ibewfOP5xdJlLDyQpwqiWUGJHph8ZjNp5qeUQITKQitsy
asjWBxHuUJ6gu/slXipiZomEh2VodZNldQCDl21ssRe9UrmopqClatH9YbRWNrCLQdLdtK5Fi9g7
rRcWbUFXlRoo0m96zGOkxoj31CzVOZaDGc+xeXBpwWGcsmwMvowe3QXO5g0NjRMKWGlYD3niMbo/
EbsOOBzp+Hvs3XUADxdZEHrcnRt1nGifEcFnGRz7UQPelzardCB+3l2Oi+I9AC0xywHsIX6S1uWz
Z4X7I4EDOpKEkxbRb+FVIjm+r44svxVLNHk6o3VThZo81Pw4DojkiIYeYN39BupY5V4EW294SDJz
usVs1Cm6x80y/Onhbbp1Q4PRAkUnQ/9gAK5AYso+TYyuN/n2Ac2ysVm+e0ZCYvEAxdFj1KdY1hcg
oyS5hTdo0oZMuCTymSLSv8X7YTPwirqffpQj4fQBEUaI1O6iDQJqB0BElZXYA6t7gjHDNO4Wb+LY
hMQJ6zjC0S4U2uTRTrSjtgjdKDWGtZu92D4eC5adY8UreOchTbSRvzFxVytHcS/PItbWRxRxLv2f
H7rGfmgeXLG/7mlCEWDMWEtkRyI9JYtmXx7D4ZXYNS37CArglDoU3DgMt8heiTwZRT8b6XMCdImV
NjFoX/vIoIl4OzSCTDt92qv+ZVTltxTt4v+XPXPnv9/h7KRjogVr+S35MNCtu3EFbM0qWGBbHJYL
Cbpvw7xGWYq839FmoJDoQPsrtnTYMfU7l3Lz6Yn5bgKOORhvOZqwAW7dnm1EMTnJMfJAXdlaMqAq
hJO3PT0olYZWroyEn7BhN6/MqGLneHcHN590/fR5Y4wbTHVPtbdYbjEJPYzsKm/8dW7dLeuMe2ej
W5Q6CI5iaNHwzZ7h39owEdkduoCSHqaUaeeHmHxhRrcC6Y5BdO06n4b/KogWIjXr0rSKpNtY/pgO
3x9xQDz12lbFjHZxYVDZl45J6nD5fBcPB6v++L54rt2/E5LE9XXJ6Yoj2NsRDJ2pGmNLuuVvHLWO
CgVKhBX5vJhMYfHz10Sawun1QwMrjwgPAHcOBjUJpa/CWQyyLSXJN8Bk0aSOvKgdI336HxbJQhsU
pwGVfEcfWyJ5GH/kCiaVSnpeXDdzk/dVop19KteSaN2Yxt9lv/jpS9Y+mOKGTvPGtioL6dip3mLw
y29i5hxCHL4YRSJLKxoiCPHx67fwFcqHpO4l830NhV2Q+EncUm3MBom3l+s6qp5C7kwEl91mKRV+
YU8/y8BSdITyzA+9R1RNSpBKNPoLF8G+x9Dmv17sfnEnf3pdAwYok8ieW6LLHHZm1GphKA5NmnXj
ev6DIYR0wNn7C0b3KhIdiXA20m/19foNe+T3cD7KD6bWeeC06/K1mLpazWbPadGLqs7vod/zj8TB
PdnvArkz/g/EEGzJk9OFKszR+jX87nLYnrnKkfXI3kf6buC04PrPWAEbNeJZNE4X1DN6OFWFllWA
sNXUdop3hpX1nDltFSGS6Vb3QWkMDcgWGUxzEWUpjoDVeZUpooFNlYlFtoBdGWuT3D+mwl3JiEH6
iXYE7fIUOEZBBLIJ/AcpyzeLjd/qWD8rct3Qa464nEMHdSwtLK3nasF+6ShqAtQH1vGFjHjyRXJa
69xhCrMOJ3bwZzLdqqy4lSypB4PUXR99oeTeoI+NAyBUZgf04XCO5vXvzKN4fgPttfbzf7g89ztg
7t4o+Mgeg8FGLEndDC/s/YdEVoaK6qkxOwpDO5g3TZSywRltwd27CksHiy1Rq32bOu6x9UW9Ef1x
MI63C360NhXywoeaGpViN6fzlKn/G1TnyBGECFTcV3x8szz00Roxn4Nw2asu+yS0Ug/FuyE6zM3Q
CLgAIfOoJI+jmnRGu6dmyeXEAbzzYPD9imNR9s+wJVtUhEdLTXgXHKsbCA7LUdTNtj6bVQuXM/9S
GFaDuo73Xr5YfCR2VF+QSSAUhmk4MqtZZ8BDv983IFmubKh3rdsampNymUCyV3q1TUCs+HmB8gbc
Jz1fHOVYC+AVny0drjyzOmAv1oGQd0d/7FTDYgPmtorhUU7+2oYMPOkQsIw4P9bDQ/WD6pJvUQFs
oBadDtzkg0ePtv6eeQCHQtzTETtG/50P9GQTSeeQnqsenaHqFhByW06TreraeIkPgwFPxX0f8Xhi
Cg4H3CcHrRwDHjkPsrzzPYljXLM+VVvH58bLDh8zcNpcNtY4hiL3pvbWzosvidv2hQFk/4Fk4A8A
5PjXLsvD24q7wZxvoGgcbgERp9YkW4yGKkvoE1Hj9w7t9Uz+oPji1trJFlpEtbVNB4Q1eMIeFsff
/X077LOxPkpH79f3GgVT7hfyi15htxu2u3Y1EWzfjvV+LABiGtGpvJdG5btx0QMUu592n1qlDSWT
g06WigfzR/JuGpYvbN9d0bnKoEKGWJpb0fyEJmZvx3z63FtP2DITxDSVSudDlHOSNTassOybbwSy
q50b4KfVgamLWChoIj/XgLX0DA5ze2t+9WCkI/Lt6gRYaBQjZ9HmGnmiJjLMwwKiv2dL9NUkShn+
Sz1fFYZco+4uwaVeNOZUlxEsxBaWnfwrCyfnHBfkRp2yoQfprVImFyjiLUXOUgmLSH+VmSE5xkXc
tODMhGeHRLcYGP6DxC1b+gKb47XuCkwFWz0ZRNnBBz2Qq6aJZH4JZz0xQmc41s709fMWfd4NLOLc
zo2edtfgiF1aehDSm+816OJgOPzqb5eliwgdKAZjCvgCX/0izzrZG8ahI4YWy/3IY3HytcFs8GY1
BUx0u14fFucaP5zuY966xSHoRN0wUKHRi1yznMO/TKIsP0hF3Drsd9uggD9zhJLfITO9qz3SzZHX
hycoDZrpd28T2V1NahfU0x63+aPm3v2AJmMXtNqsk7Ev3xkOEZxdZuiVtfDl3m0zcC1CgPfERAbQ
ri5Zuv733hujr7T4GQTXnAvARqk4ACib8WqtMCLpM/vMG66xPnkmfBw8+1bSG2FeiwJlkaZ7oYrN
DPNdsgIgj6lnsdH3zywk+BRDpBWl8/ICjA9cN5Gxi7ZRzXvofCshE6oIZ0GceMQfESKAogdSc2Cm
NRmsjv9fzE9h9E6IlJBimc0MObNNrak478zZUdCaOw/6U2yNh2a+hzGSAvBJSuAFR9CmjdGPdN0F
ppF4Wty0ZfnHhxQWZXfgm/wa44k21WhHw7j22kpkmJ/9NcsCUvkf3SE7vMmNK6J2ADh/ydtrEf4K
jP1dtM0m+ZJFK+l2Qdre/FuhnlnAQ22QAALrJWEGGEFHdb68g4aT6cRaWuIMpba5R9E36XVrq8PF
Z8Cd2HKfMwHkUxEFzxRWhfkumWiv/JXy5LtN3htogy60SWWV8/bDinMJlmDDkgfbzHfARmRtd8g6
4TrW6xBwkzg9zE7tGyqnC5RhE9qqbbiCVOZirjdURvedMCrUIKUAKFG6PhXy+BsQ7jhVR3iQ8g0A
oORsGebeDxIjvakMdzte0C2ORUu7CRdNMsYRZkpf0gcKLeGYDut6a4XVrIcsnZRsBVcvcEtJqnXd
nKdenocWJkpThoD8vq/McjgsDd/hQOO+MYSaINLCUdK18z7v0z7Tomd0fGuRSTHvMaCrIyT3/Vdy
sPPN1ZezZQ4EWok4KGeheDGdMGsnNaquluuWVxQlkN7RKPflVnOxRZIQnBujf85A5otEEO0nb1tb
O9TS2T1OFRdZFjw0U1Bg32pLlc9TalmFUuSmJTeEjI6eI2tGOpgjSYXw+ojMqJzOiRIjjNJpuvQz
muJUmqmfMrUMrfuyoDMzVw8Ng5UwVBKku1KvGvFYFjDPCMF8ZQG/j6qa1MCO/iDltaa/O8U754qi
WFwf4MzepbAPPHlStlojoV5JfIhlBm+P2mmW8ymY6GiQNwO5KKStktjhLJdDR57Zdr5xUVyq89rY
gP1U2TqOp8BycNtY1kzXYIMZIrzpYDG7RTCE/BWw/0hEvHCAbZ84cVtdYsheSRU6xB2SeBD+Hq4t
k+aNRoeD5RJYnO855XKxqxr8hHb/1DeJedBh9JUaUae9Psj/YpdDXOJAUjmGPuYB4o/jLCNlPcZ/
6t4OO6o4p7IItM3k8jVagrFQ0gN23swngcSrmE+azBACRsaUG9/sS6QKBEQxICTzlmi0xxD553eI
mQtNMu7MzSbu/4uCP//NVqSf6bKsdnneomU+5OOEBDt+pfoBJMcKuOxZZGTnb/zsabH2CMU3A670
zAUxSlAnvx9U5VPum5LMKaICj977S5BGL+x4jUw5ob5ZqvDsG5lvDcM4ceP7mVTGX+vBRT+ONIBW
QPL37IdABZ0RS2Cuei9evzQnaU0xXryxNj2jZL9dS2gb7mtivinmYIklg727b1hccuuZzcoDFjv6
uBUgPYZJXZS40g9EN1Al/KAZaA81ra9j1sRBMs7LBtLtasHRrkjckE7a0lE5vPdyy8yNetOpq0cL
HouhtAS4VJfw0kDSPxfOZTPWlb7tfa6wxLnegERPnrWzsBCijRQFIfd3dXAZedIhOVpfIjAKcZev
UG4GhrvtbeLNP5kiHI2VwQHSYmOvKtH5UaGCm0Iw8BSSTjrc31WRx3YtBn1sZt0Vd7kGxQ0oRiqO
Z6VOHKHUbEyKcKah8iKS9cTOhMlJliPvjG5Iht2zVVbGGQAYnwvxlZ/9kKMKofCGhNIdYUze1+/r
503SS1US0/xaQ+oHlH7vOzjZJAbuH4M519QEWTUCAA9XKJLn9uYt/uW9CRpTcA1IHwcWixxS6hVw
Fqpge4RNk1C8kvBZaz2diuiYMnmHPrX59Fz1N/9sdAnxwcGIFbKYqmqtkGCdqaLXDHpbuek8mech
NhG9E3L9tEI0v7r42dC/D4tp4P3sDxcSvOh+gU7UBf7VxHWGTowyuW57Uc9f01SFnHU1SRv9zg9j
ZNaxfxQJzAtDsoyA8XM7tmrrfqjQVZ3K4ma4NMs4WDI1U7vESZzdF8Fc9e1SvJ/EdMARMj3VORSX
PzDB/FukjYga32ThTgWdAtbiYuSq3StE83cjcuh1gXmR07FBnI1ixLP2+DEn/YfnpiG/T4rQzAMO
TQ0p+fDW8a0K3FCHIzfH3qzXgANrHelZQyO0irP9N2DXXb2Qma4xveRZeldGVFdw6SyTLvL4zuAd
22ftuaomYzjV9iwZ9VdmnklLN6XubMYZr/Yh2wQdweelko/s5OS6ssbKC7+o/b/0FMwhTnCrLP/F
CNuvqo89t6yRQ4Fs4brXwiWNnV6Y8WxWkUYoslzaJxgIi4J0RopSSiTi2FwIp5TgqexWAR+U4HyQ
fHm/Vzm90OBRTT3Sy8hS+QKhUuPfcT64R+cna5hjuS0Nme66gpo9ltHBwpfM8ooGZ30vf2YSFVPD
PMpk6F94i/JBwAY5yX90gFLy6Y+yVYFNLmDv/PgQhbtWAWCa0i3+dQqyZYQrQnQWJ4aH5YgDCM/h
bLQpHWR1cc/sbZZlHa8k7rFcHc3ACAg5sNvVkkiwD+spRSJN3r/7PxFS9uiKRKwTzSx5l9LeTMep
u5zhYC+YuJaqbunmB6XTMHtiBqr9AB32oCRYHm0I71dMTxMM5YiRY51ifoR0KR7/Hl7hVjqBGKWH
VbzBBXKHyM+Zpikfw3MXDNTktYTw78ZRF0L6o5moqU3Z4RSBMXn/90qTbH2lfSg9B0Wm3XY9me6U
Ssj4S+dwydCJDcWj+BIB69Zvq7rz0FGkp0dQISXIigff1fku4b2JW4VT3pJmLKDpib/ozbMyZVhL
YWIACbnKhitvloXzcp5TH9JZi6GQPbUWaT0VwgIC9VxBOLe4Jj4WDd+C2QS+JTDWXJAeblGBmdrF
Em+ghAGVT1iDJoWz6sueDP/A087xaBCHCSMH1Uqu3osDjhPZoW2irsLp6Zdp+lbbw8VBXzoPdNhk
udRWg1jrHq3Q7HrQMpiEMtMUs0Fbij6IFVF+L2AWXTf3Em5MBJu9v+EEngBCYOkVQWRQMe85e37m
BIKcjFBXo2g4x9EtZo8cCz6f6bXzqVDZRsQQn9Bbz5TMzJkIMwJa9W1ea+XxDCCoOE5mcd9H0oqk
tPgUbOW8ijYU2+1Ou2mXxCg3oBM7Z4wRAeWdIS6llaUjMczEnrU8WInJUC8J7ZuSbpzdXaOYns7u
oMKtP10q+Ca06QFEXRchkaB3/C3DQ+JzV3nohgG8RnhrsMOxOZ+cNkL/B9zyy4j7EB3/sXNnZgLX
OHkmdCtpTFOUh8EZ0xgeUiodNY5QaNhsNHc2lCKSuPfgeGWOrDE8uCuIyzX+/xoisk2k4T5w+s+p
TK/nRxiGuSX0tGT+1jMucq29KS+SFo9m4R66/jp7U3Df2gaRSO+vkpZdFHpw2ifIOzDLN2VOZLMz
iyzN83J466660u5U6EFB1scqj1vXpqfj72GpLl7Dp4tTr7IjhQi5TB4cw90Cc9Y/G0iLf7mFLHZT
A4OJlv+5RHFcDTxCkB0q82ZlfLByzDdMvAcRQGupGRys+kVYrfgrmBRMqnlF7K612PpFXs38g3/S
W/uUhIpOEG9JHNntuDsRyWTsl2+hmptaK4t5EvOB5ZC6hgnIv3cQ6LGMjRgM6ofDHPD7eLtMeM52
i3fxIniNGeQkZm05QEGh7atOL0mCrCZpylEV8D1yQeYnnKCFmS5McW+AGa4gmygw7voaGMq8R5HU
IgW5VO8V+QgdJUGdbpqNq2hGGNFxW898xOaVSqLeo+ZdScQV5SKMSNW3ouUVBZ13tS2mZTVRgsjU
lWr7KbH5sbOOipXGqSNE3e6bO/DA1PSwEhZkOtISqr2SknAdef3BgK74UFUHTpGygHKZWoAebuTy
m0PqVoZrHrYcagOPNPSTqErJJpcb+4XQuqm6SVPWERXM35ddUxz4gvsibNu64xEofQBER3y8wHOC
wTFi6mwLAPQLnOuyzhfQWTHBuFD3DloEMLfn8ZTeqISJCH/65CSY1zL+mRROpAoCxrXEaq+J5w0U
owsIInP0K8A1TtnXezOwp2tgK1IblIRg8UjTRmxJMsktA8JrFIxU5GMUPdZM7Qu/67qpykEru9KP
b2Pzi7y+nMcFocglbCYS+Ux8SBU7UryKrhyZH9+T8T1rUD3K6P971rg+BT5w0nD8+7QzoKqpxXMy
DMWeH79t2AVxJY41qL+ybb76izz/nP8oOt/bVZ3CqLLk0hC5EwVbytnTGvUZ9L58YhOxS0j72sIy
9gHVqTR2ymqilOSEDo34QbzcfvNGWAu+nCuoU8yfVO6v9PJWYPLNvs8pejFKYOxeHzp1j87/Lzm/
Wx3GadGw8offcA3ozkfpK0sPYlOZNhNiH3877bQt4bnE8dw1ODuect9+GS23M8EIDRYuoGwWDj+G
XdsJ35bYU/QogqWfXqf6dkCavYrizNJt2Ax06rQEOKWW1rwKs17wS/t8Wph4zyOK9c8TQQUAtMcK
R671CWIqk/eIhN74C1mlBq2ahDHtFw8JRVtxq8uJymQRPbk0Kyev6V/LsRvkttw2rV8b3Gv5cxcN
O0wzH4IuNJYmuRoLKD2UbG/9H73palbCVuL0dIEsRRZPSbG0j8TDKemXmQmbfJ6/TNhkM7DFraI+
AGzzHIOHWQxKbtcgaNr4lGLHPQhMFm4mhKzSDNdCizCPp8HbSEP+PaNY0lvrbI96bo96CRIQhVbc
Mp5kDIBnHIEN7eHUy0+0Yd/Ngks/ZOL1MTEFyMo9d+wSddxOdKQjiJ9lapfRS1ROlzDA4SC5Eyqd
cQjeJj1NMv5bkAoDNqWXr7vYz/laJgzFFRdqiLsUI6x6UqcuhIo1onmtB7WuP6PcMW4Rgj2PQXYG
Xia586lYV3hSE92JN/omoqgTKAsgnHiP4gSw7xv4zqG3mVscHdIhemvc0hsb9m9x2GIyPeNM2Utd
ZnuxG+V7tVdKBDyvfVHogOVUqMmhpfeg3FWt0mOWWgELe0UWXESUEIOjLUG1ITuQX8F4AT1bLwNF
308gzApdo3YoqMRedphhFrO/YdT/tvgBf46/KSIhBKgzEJ/u0EBFu9Z3LA3S2chiDOUrmi6O8w/a
Z3b3zB8N65tUgS3dS3vmiXowm5O73/V9Lo7sY9adWL9xp2Vge/H3Ha7LsSJ8GvSpKv6AO/6DBaNl
4haWiNHwqAzMuViMQjpI36mL8oa1urhcuLT/Zd1jqHDUBgtKNwLEUmgEiyPNtOckfBYvoZ/6O3i6
0oL7qwb3g61CDI/0B4a+LVKe75Q6hOoio93Bx4IlI7+g+TioMT3fgPFymWkdLsaLNfjja2B2idz1
z6Rbn9C39TKudkFHaQ6dJnZR/8yGs6q4SxgSVzZXXCFHGzxWi0x352JjqcUS2N7jZ+ptAI8BeSjj
sejzhwAwrDIGcCqJsRSSuDF8qk7+i0nfA4YPqU6wjrXcl8+M2IlxgHG5tRySEYsrfAnhbWGdXmGa
UwSbggLBowElYwaSdyV1GYk0UqDxJOHbVTmWx39dwto0/NcxXvnFW50obtScsbZVoZaM4nOvTwDE
UG4NkJ9UPPls9NoyHkHMh6w6N7z9a3TUb6gkRDG7NdobZXL737Ty6cnYX7PmzmrccBYUoiVZAnK8
7lp7qhsj2sqorZiKD0yyanHwet9hlgvPqTqbEnihXfkMndIijv6+GW7Jh2EUF19bOaNsWUCfcEOP
sFuUsLedPIIXbkMQFMhJlV9kEiz/E6LPCv3hT1uHae2z/YLy5dekpRoXtkYq81D/WsFJBINcjKZf
cN3SKG/LBEehTf/KJXEORmG+ndHJVftWLayUlYxNLTzBBMOCH9SA++VOEAHGj3h4oNzgDhCA9UDR
c2zkSXYgG6pLgY8LfVjOOxrMf1DqH4zQtNg5oxo8X3GnfxaJ7omuVXieLmOvXyRC9xeZpJQ72Hdz
+vj8zNiJNjkJbPiF6QLxfplVqnlQcgwA/3k5yWvvO2ZzlYlaeLpoGS4Y9tuT/HUrnPwFnuCrXhZ6
2QjU4LiEpIqfnqj8eolD6ABEk7x8cwFlTFSGXAZA2SFG26YCUHal+203InOUqofqKdNiZRbvUo6p
Ym0/jvu9as9b4pZm3ejnl8l+z20SA0SJiCo6LzhgxeN8CYBE1ARydZRuzH9OteJVlAEFpDe8n6kt
GWtwFz0ckor00/jgjGKoiXBgAvxSwcOzbCH6HeW3JbOz7mXX+9rUlxtgxM4fUxUeYKTIM5Q0SYxH
ke1qtVKMYgiKd8/7OO5YCAjbYbQH17dJt4O6jPJGOZn7iY+zhsvFDqAtK3Djd3pzKS8HePMaUoWo
1YmYLwcjiNLIMYJrBt6brrMEKQX87HBorwpQCy1V+zfvp03AIjeqDRFOgv/H/IFqLSykyHZfsGah
Ag9aA1P0gT5Zcg+BGKfKTIMUsahr2RjWJWYS7viU8yawmrRHkAzaoILMlETh3hTCamqNtHdsgKXb
sBtSR5OYWzllUG4L5SBeDAePuzWGbXuG+UsUoLCtXq0yE4UOZSYxmE947Qzehf2pq45t6/FSa2Td
IA15ESRZ3/HLRL6wt3PiBeyn507cfNTlN5FOt9DlFh9wmr1lS73hrHyqLaS2X7/SWSBGbGyWnF7B
fTZSJARgXaRm+s0u1IO9Mz8UfByR9NL9RORJtbvTtPpSrfjGADy630kFwKbcosmzHssqe/4/KEbn
aADbQ6HQeI1DirVokHXTIjMv7PuuKxLyNDYUmFKeMEdP2TX3YF+11TIOY98wAZwGhVy4clW+MObp
ye5JjDrURqpae3JpKtwirAqsodZSN7li/omUV4UWFYl/uhFvDL/RhDIYq4iEzcy8S1CkUyrAFBYI
re/rkKzLE7qTnOXFo8V5x/MNCw6YgJZgoWc5Mh5Y0c88gwDKFDEj75gErNZugP0Nd2LLDYXivDmJ
+1E6DqlxzpQmG/GLKu98gQVJq1k1dlrlcwlfZkBJP5g118+SQod5j5WX7lMRMk+oYGFHcWP4IV85
6o8wTaY4E0ploYlrzA28Ku9n4MhwpF5yGjiw1LHz6yR8NDdq4/j2VOKWf39MZ+i8kzysLLeTfk1z
GWnbRdk+Poyw5z5BBZo6vzudTwAhyVYEf5tMcc6UYrwEd6rA1SbNXM0d3kFe7aB1boJzyzJUJBd+
IfaAS0wxh4a/4v+Xp9FA9mwKsvs1wXSwW5bLWePCPTuoCP+0p4dkPteoDilnID0Xv90A0/W6BGAP
KxNr2qCqez37fp7TOh9vRJ01yPog/aXK1qn99paT8v0tDSLwWf/DdVQABSw/R6ffbgxJ2sqt3lcl
ofNn/qZmSMLMi4INbzle1h1YFWO4zajwG6k6UCYC1MpG2GmW2A2M24FdlO7A1b6hWQhTLWrMBru5
T+UnYBXAReeeaoN4dX6pfXadeT4xLUyxKH+2l9dln2lB+M9mP3YNnw6rcRgtuTXHOmBvkGEuBVyf
5lBh+MoAvF1agqhS3vIRNSj03FzZqLgoxqamalg2MWR8aPGGsOos04kbkaQ8byriMq11rUMD/qfj
sTSXffxgyjzJFTlZQXUay7Ylm+iuf4rshcMyD7CesOH9tShAc9MRM/YsoTRI3Y5N0OkyAmEnlWP0
X+UG/FLVV5V5I+fcLlq7vImCdgUkGcmhUR7CVxtEmjW1fSSjOyYa/rlMPkxW94UDLfQ1Ng9hPfat
bwrJW8pLGz3BLsgGw6e7eapTXKVHPRTLaTEwZBLRxLMjYnRoBCAseXXdxhHfOhZ9sFIbaZjFBVCd
l0SePMVzQwliVsxPMTNBoJ2/WxjmRAmFfdbvhi58y8CPEV4g6UUrp/zArvmfw1gjlwuNcWnYQf0k
nKzhJqE+6Ty1H0aTTqjNOZci3c7A8+4GUC7wnhbEGB9ibt6PTcrXZa10MsEAvQH2eYULpyxRG96X
d1W0YgwxJ2c7Dk6jbCQWVfgyiC6UXQk9hIVyRecZ6greNlVINBrU53nk1Qo8rsDkC29prsUrxvCe
aObusiQLs9bEdQ8aJJ7rihddon2MPyr5fcOG2A4yWEWai+/ABKBy3c2pXyVQU2vebJjVgN64VNPJ
ff30XfcBoWbN96RHHIBYO35TaStzHf2SVzt0/35xzX4T+DR7vyePEKinkohhzdXFXeA1feL2L28m
gWSvtnzGDDscyqlu/vYEtEvntaUS0RpHuAvn0MS/p33knSd3LacCHMf6psIkbJmfMJbLs0BEdtqP
uJBf43d5nUzSJKTVmrV+QW8tvfRMWVdJ3EHvcvtYgbQ24D/QuYjW8JMn6yuVtvbtmdnTfAFM7J30
+9JAlss1RMcUAwRyjL3KhLXBr7DkW4yoOnJUsLkd0l1flaz+UTk1dWwm9aBHB007qNF6GwDfuPXW
qKnumbsw6le0WVUqXiW3Yj4Q6UBWOLwqjkVwDw0DNo0UjW35K1LSm07E96i9qo7mOn8R+a1nbh2c
/jIcZzGo0ieAtjPMF/Y6lwnNOrASmzo3gOnfufvreqQi2GF4MCyqy+lkVL6dGVyP3ZXjNHebBJEk
Px4PpXdCrfCNtG2mtNAH2YIRQdr1CG/4UcetPNqZdG/UAbgUvwHLl+TU7d9zH03YgiW2B/tMUGK8
oKvoO03PTE6meSBdpeb2TWRNRT9VjzRJZMB0GpJam389S2txLzfRHgzWUPDQAHn1Q/g2hGfDxzaC
cAa8n5vGbQHTJw/Ro2ekZ1aavDIHP5ZolMECzPgrHNOa8N01roX5KFiMmDt7BNWnD7FNgJ1x6GKo
hM5oKbzHFdmqeSNeS5jZizmNoy+HvhU7HQBuUxhapoyO4Qm3b3kvLZzz/A/GlmOXpxcAQ2FCBnaG
iEJQ7jS1CzTinxGXp2GDj+2XOzp+RxKOx/mhk9A3uZ9mCIJtko3uERDyi00Bs37j/+vStvH104B8
+KNer0SJWhSLz37an9HmGNVzBcrTtrbomepbEC5AyPbjNPnK2Jd5hfp35oYAphqk/L9Bsy6O3bUT
C1eJh2siBM+MRySqcwCBXF0+biRu9++DDFNN4qWYkuyPK9AB6VThMTndiJzbReb8EzY7ukSwe8/7
ND5Xoh7WiNNu28MM5gl64Np6H6dhIbp5xxvvx6Gfk9WwyU5BcvYnnJj+UF4hUYtGNOp4gTj9514s
oRw1kb6R1ht+Lu7nvPrrjdb/UPKUEiFpRlj0vxSSIA52T/Fx+43Ql7gd+O4YM/8AvVu6SkOIY6Pb
zr9a+rqH6pZYSg0VSP86BSeEzYwH+SRPzpLubTAYccfL3p97c/gc12ZllcTrw/P0qlhfek0DJf1W
LqAQUancpxFd66NY4yuzziaquIzssWBCYvN99HM212GlqmUm2bORY50FKqWR69aEW3+2hftnO9IE
Ogez2Jn21oqn9xQneGJBU3MZlEkhMmLUiaG7pxfPmgYW7a9wU7wOmGEPvG4zZ5zcOXRFjSHyU5C8
Ug8ZGEVdwzSp5Eg6ONRPBPOTjbAcbYFh9AGgwfeZgNLlnOn4OSqS1TBmFe6jmjrKxcX7r0z0g4bL
MVYBsULYrX+VJ7gT73QA3lPv4yJ3+7G5Y76gSu8WFf3/J+Q+1WdzynSfDFanGhF+QT+juPPow8dD
F6jxucB2fW8Zyims1cD32hAZsOl8zJR7iwjx9qJL+elIk6bGqVhCSN45+Xhu+R0dLJDdLWhMB2YU
sB80k2yHlwceyZTraLVkeYl5hPyKP/CmurMYfcrTCIqasxqzCXWApo1iZMwk9RnXUkmNkHgNbRKk
kPFFMj7kuAmz5expBnZBI+zm3A==
`protect end_protected
