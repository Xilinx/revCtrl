`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8512)
`protect data_block
td5QFuuLITbKOtkE3oI0mLzB/U3OEn5lA8+gSvm4NzDgr1xoKZ6KXCYimdZuYcgLb1Oo/1ycim8W
PFfdiPDalf8RhWG8Bm3Uye1fGmokMIeViJJFpudOlf2QwkH2Q9nSjhByWCvm5V/7FzruOcyzJZl8
uis+1q6Ca3nhUQR21H8IcHbv6Xy9XdyKOtDQhDkDGI8SOYvdtcIlVOvSvgg1PlHx6usdcjRT0U4H
P6/B+j6sbCmxYTaRSW+MrSFDCMABIOsqlOFl9PQ33XhNbwlnmCINWWiFLXCHyUhb9ZzdGhUCuXZr
Gub6QZtjqCwRLiREU8I1XXrWByoaoiNEZsWHJRZFfYr4hPqI2RD2dxHcIRNwWooGYwIq/aVkF3O9
U4AwMHK79CDET57iRknTfziwrKv3bDx0qOPu/GU0V+jBY5sWup9WO9+2XyGMp6O9lRQx9Tt0xA5i
lWvsSXdN8ETZT0r5moiD3zvj5GceENmY72FNBCJtWWuPqeB/ApxRkin6WsGYcD4f83JEHB5GwfYm
rMh19PJN3oajVV+wVX8QAa1P2Bm149K+sTjXd1E5G9Gi/4JgeoXFz/1KzMqxZpMXnWo4bzottw7X
mEjBfNlTuL6X8aXjBdY7TSHLEtgQ/b0Q7XuVxgqDEwHcpmRGqyyR/broDJSihY3Cd/W35X5AIgir
63MEhGL3+15n8PCFtAolikeYJN0wFFeut3PKijZHtNrIEpyxCLnOdG0AGxAurY3c4xV0Ww1qORaj
0Nz1AbNaCa9fTlK/LO5mpuM+ZCQQJsYrDPB+LK/C428cfPDihJLVb0DO9/5sGSJmYgfQLQ9sfvu2
bWxpDY4DwvXSguGhs2qIiEvqrCtBZVxVf6AeyiqHmWqC22iK78UJPAEJYUY/bQFrYFPiwzKUyD7L
i6a43bOUAMWcttAJqvyvqBSIetdBlOEWuLSneU7t1Td3UdIomIk7q1+rz5yc5fW9KWrmPRBAYiYO
7+eFGuebN0Ei06A0TXhYhfcWvnDjJwLChVeBrrr7QflhKg46J5TR/u1MIWugWYb1pdhxqs4BXAgm
37fFeUeA39xrEl0fmndzWTwNtKYOxEKg9gyuKnsAir8MX6aCvZvZANfEQJpEGmBf8epTsKJYo/cy
k/mnxo6ExV0eqSinLpn1Gc6ACcOTMokhDa45QHGbdd2Ym+qTFfFGRse90ICLsLauGoIxPObZyD1i
K9ors67U0ocrw2rkM6IY8c2bXnY4eMYd4y1NXwXbhrgwxI0pVuFOWoL4uBJwMbwwFXdQlY7+6csd
ezbTP5xguYYm+5f8sh3h5LByn8dxlS2i0v71zA+J+o+dHhqujhtoAxBm8NINMG0p1MmT49X2deSx
eX2Uaov3+kalkY18646K6BraB4DsuVLtSFlpEepOHIPhPcMJE9bRDwJoIEH7ZmulJTa3ngWfAuVi
WTuSSCleyurILSUekODp78X0XDFdTg+xU8i4vF6Xf0O1kN5VkHozbPuqLVo+5+WCL1kGtthk3EOA
GmeEd8Cx2am1nFBD77eb6gQKNSC5x3ZiSD528MmHvshCZoYK9fdGXbrPoYTp847GNQQBdV0guBkI
yB03mBD3WfxSx/apPbWloAMnvfmWtEcz+H4vXoXmCTZzcH5X8BtLO43NrWVgkMBiENvIbOAsN/4B
6kABSw5CO0UjEo1S7wMNDE0etMDu0WbycicQrorSM8ik7FuPwRI4SjqqIptUfbnlAvIzer02/yEQ
Ksji2a+mszSXCkKWUp7dKDEcgMda1jEi0GV7gvSJptUKyL/rjkZri/gsBUgTpzT4eAdS/UqvnIxV
EnKZEtyBHy9tSIQ0nefoOjVwc+lvb47LtNR5NQ7+3xvDWfKGfXSWmCkD7REuEXadUGlByEbnBhCU
O97KHctBBo3pqf8n5xIjNQ8ydaSO3tY49iuqEWXFIUrg4urm7yV+MJ02sSNtiHpVXFgBSJckA750
5ZqFq9M0vsAq5ETKdFvd8tyUNRtsWPb6iuYM33REAHsaUSKGYQqnRQh7LWMVrsniRJQkXuVndvRO
6TWejX9sUF4QyzEl5hhBhiNvyOlvsJ+WLh3IvHY4sGpDRbQEm9pZWeh2AnOeFnPcMKT7gF66tyJj
KgEk+47oAx6p4GVl+jODOBoc2P4QOThENSxyP2VGFmxGgVUPD9XvlRtoKs6qDE4PFiV1GcdIeb7K
4KA0H+89ByY7ngq0a9z9uGxW4Qed0aiXPcGYrpqq2oZevC0F/g+D2RqxYmaGwjGrOCB8p1wwYvKm
34Y06Ync0Dn46DMpy3/AtBZsFuTcEjIHFxhjYw1CzRZvTncjpA+W84jLAltosulMYr0Vyzq3Mt97
urfHNIwC/HdE4w/deMNbbevt20UYw+560mTM7Z7U8LLQA2syn/Ra+boxJcufLlE8aumsGYuSUFvD
+3dWZRVbOb435fIfT4SsSRpAFWGcBD+mw1xip1yplXJaayS+yXz6Z4TwYMnsGA0f02t4YWd903Gv
I5irJIlGIMmWwDmJIBNTFwmrRWBqnGi5ILnCulYD49faXjyuYw4Lb8JvwWWWDozgKzlbrEqM1+ra
gG55fOqURQgQrFhk0eqzOypbBQogQ09a5Cc4dBI48u4Ql9dDLxAuMkwPX/LvLENc1YsBkyXS21aK
76H9Pm1i6zv4ee39/M0rYiGQ3a11AsPV0V5Gk5sihge/sFZ28BMc1ZSqF+JoNyRE+bXj9IVj7lBm
jetyIspWYQLEeEyxhH9SICIf7mfIip67VC36ySM+b82wyjTINuhQ27Dojr9NPJlitlTbdJX/rFnw
H8MmhQzEvdpxvPwMiOLBUI+BL7pPJXju/sGCZ1QLd6DivXO7SGt6VbilyprPppboph2GhQIHl3i2
vUx9lZLlncwMh/YTQjsKLZ62EyeJtvvm/UwEGivEq7i8N82Kr5u43zdI659Xkp5JcqWhm9g6OiPy
vCP75VmAqRpURCCeXPHlDd3tvZ5FhOjZzKF4tEG5eVW7d/sXDpM+tf7i0orKFf9xWvfCjIfeJzGM
woJNMLTnwsB4gHW4WmYf3RREtSDGcQezncKm1ZRXg8idPQ20nfSsvRe6YJutA8kERrC/UqnNkI13
tGcMs+DBLX3AD41tSSk+vdtPJJumnNbLwvdvNxqnSgcmDDsKFjz/UsMAcOnbUz8a9RxP+d0PBtaO
koYcc9H/hc+Bs97OgJlZ9f6qstYJmIcs8qjxY8eygzyns3bg6CLjkeA2QIKOibxB8T1X+jeV4nKu
VoTldRpkN9/+0Pg6jSHbKd3HXQd0McqRoDvQyayl5TI5ges/PSbIdlwDaQt9nW4TO6mJRnltcOwv
O8hdA+XfR0nWNDl/vNvqJVsoKk8Lr3Z4L7RYvhyrwcUxGcEcKNhkz384lHfo1YV4If0r9yx1koLb
zJzJ4/QEK6lEIjs3GrWqY8efqdh3mq7zlwrnM26A+Owmsf2G27skkR75bUQarrQSAkv2M7C5E6NF
Pz+RMWnarsHGEbx7TNO3rd/hFWDPISd3S2viMTMb++hl/UsQcmx0UrZKXlBSKqLtTDuvElXTAW5y
heDbB4kP3zHusEYuhckc6s0qWhJoFYQaJY2EUjgWJbql0VQsWxQT9ythvw+KzCbfW5IXWHyY4MFP
Hk+WZiC70+EO0EsNbVmqNqDaJrJbjV68XPOcdNTqgGAvmKlEWBrBNE8jOgIp2Rb/7g4MUNHPmjJO
sirZfOCloTRZ0xJ8G732K5lkdHDrr57km53TZmilso0oril7QIX6Rh7B9qR+MlKYhQAU19afwNTj
t2jmY9Mskgv+tkZH0sNO5ZIG7vCUAiAYQ/R3lPNc9eWy9FGx6rohhvFmMmTPQxCx/m+D3ECrdrSH
oqxVVPfcIy6xxoD3yl0iD65AW1bLxN8OscBkVAXVWdc07gUKFOkopKGAq+tWNUfErxnL1VbauvWD
B8ZGsRbErKBeIxPPMTVIjvfO+fcgajWeRa9lzQdAf9nIovOTRwqN+SgroAA1ym/1GcmkguLhWKWk
9QMk/QV2QF3NKM3awHd08XLVmTuGn0OAceYDYOLm5ppy5ySfptpuFzpXE8dOm091kakg2/ss3gA1
XKZZsUwO31KAA0iieBOT51fXZ4ay+OiArNlK8QlGGqV8dvueDmIsoBlg+ITcuPrPDZjxi0XgEpVF
sGFsxs/RVbINgSXakWgQQNEqPU7ITOYJ1c9f9gbIZV4zgfbrTWskVyvURp9cvYLpKoa92P8taIx5
4RCmoWoGN7CYAgC3snxE+IpS9HgRW/I72EnzQFQEARTeX+hC/ez3rqHw2zEsWs/xBg4oeaVEapDp
pgFeqwn8Vr0sq0+CCE7YropM55OaoJ6YpX+LNtYEhgSLcQyoFLoINwKvMEyIEI1UtrY16HDYjekj
w3UgloZPsuUCT/iqiFZ9AFbKSEJoC3x04gWj5tZ/a8nFnMEhGff3HeUSHUnTIsMaR2Mtf64eTo+T
fxNJomz+91IWjQwBOalhAgWg5vjVFmI9nHSTY7Adm5GKjQ6NsHfyX2Yk++T4KrLYYReMQimQFo/4
O+KCinUgYIP1FymKHP6NVmSRPuAJ43pLjv7J/tF6XCpTlYSg6AxU1MQbLrfXcesMhzN4luFmgE1s
gCU3qbrFwQmTE8agx2QWnZg04bDgz0FRSetHGZBy9nt8h3/AfDq8vzV+KWSy5uWChq0M++sdP7xb
XMwQB9C9mWsJcncjjIl38hj6EFI+9RWXN7RUKl7j3ou0G7Q70KVtK9dYCdSEVxoF2KRLu5vYQAQl
bw7NNadMCt6Po4eVospFT1yNdV6bJFkKXiDA/Q2LuIun4bBFrKV6fxpaPud5PQ7dxZFWo++mtf5j
FuWeI7yc9tnEukaRJCeuUS9xdKHK+IJMFkX/3X9Xb7yd1Ma5iR+vNye/drJnW3Eprddh/k4VI64/
V9B3emaABIZol2ROsRzRVoeKcKZjtwRkxaAHAXQPszVz0yRhz/uNFKcN2bsW5bez6lvxCz9zx0Sq
1QjMHPiS5F86NXPeXfdztWRUgFBibILvCYzxZfBQYQtLA3GQ8Be0fs93JsTjh70y8bnaRS+2uqCL
YENOD5yG5Lhu9bl3gujs/zG75Y6VGkWmyk+ZeXeXZpZXB0pImarSoPaJmE7rNauD2xIu1vTZ8KSq
PXJ8WGFKmpkKFZPylo4mFvgP7ulZNPbfVYeheSpZq/JLUvdp2vfKbwu2Ewds33NEj7CwgyGt3O63
wldGcrBP3NrEXq2t4WKW0LlLknYM4YUjWFvPSCB4q5QuKI0Lv/dx4xfwfbdQQCumPnWKXQnrYapx
ye63xDPG8qZHqjKa0kIxxvEp3bbMppr4LsByLCYVqi8V2OE6fyb9V2uZXehqP2ANjsOxgn9ss5fx
Eyx3dS1OumwN8sguUYu76h3pQwAH02jjrAMP1cChg8ZjgMIaP+Sq+c5bsNKLWSpKNxM+bPnFx7kO
AHSakYSFOtXuysD3/cMHG1UrbJhKPPDN2YVIlbpzcsfDCld24qxcnyEZX91+SEt0T+kMoO+sRftQ
dxWohk+Tqs7FKG6Nx4wa/E/kPUSaUNYvwhHs2bkbhB2nVVpWeEwUFjVP+H5odl8+ETe0eNGm7Aiw
9uP439XnQe7vUkp3k0Eseu2gFjFnjjXKFw2zYzybi489pI7rkXSGnGVZ9riV1pGo46SusvZCUzWg
jAao7mJ/cwX8OW4NW8zWzp2j9PjbGKEzjVHKqRHe4eO2+sTS05fAzjijPz8hoR/K2FB/Q06MzPaP
mfBHq5AuwZRDNFYp3gMhiTOwNXNA8tROa/WJDDcq/gMfDIF+NnKhBDLvhH2vuMxMCV4iV5TsiHWI
5yFDHfjHm54v3ffUgAjLqXskG5hdK8rZnpmw+TkcFoZtED/IyD2/6zvRn39dQ/x4Ku0v9eXgG7fy
KUxg7HbboaZlAmZz1EJ44sR3fv95F/r1LFwDRPkWw0aRqxlV7XLJaQMO2Ob1iLK8YX3fGvb8J9C4
tt1+wdqwxwcsb/lCwPZ4iVavW+TOlQr8s4lCkrfrDpCryNtA2JWv9zPmtle9cMl35vXpAaGHndAa
xVHJrG4UiXg1bUyb14kIoHfbEGGNp5IoTSjPr77jETWxt3DkoTSyKxnMrO1aW/koPh6JPiH2bYdF
kivUu/TzhL9QqyiSWFTHTpmi/qadkkOWGDR4n8XsmArkKNPHYdi4rjn4I25EZ8EiNh4mXRa3sEHo
VXgnWXZZGnq54Ap2LrS7PyG2lmPj3wI3aR6vqLlQ7fSqW4glLWgnfRN/eaw0jRVTtXQTIpVWQ+1I
AinxDL9lbzJpeX9MzQPKnOOOilFSEj+sX3BMldPSumDZI67zBcOTrn2PtjyvYP6Yd3KzSbRPCZ9k
4USFtTe4IJoM38omdzaniD4xr6Tc0ecwHOu29yxUdiLaC9ZNiPkUCxJ3ClkneJvtO4vacbMtVJ2z
1ySppzp7zQiwnZYxhMBciWyH6sdHpT505+mFuu2StkgnOUYSSOJXOwt39/Uufh+xcBoiufQYAtgP
Molo1uVo7ty1AhKTSRSSPjeNzu6uO72jPH3VyZZKteRwZbnZm/7Kajk57eAyWCChGqW6ZQDDvC0Q
MDY5V/qssYENhk0XujqRd1XEoDzQAwO2YGLo6XPHZ8JGRExOqk6dubuDC2I9jCLDQffPsnw1mvzx
Ime6e+8H5P24AGeNMkHmEPuvqxmXC2kzKP+d8u6wmmWed3oOksbd5QBoL2U/ocuNQRyRverolyM6
WNLPc6WqzOzVaxfN1LZ7GGasVyJLvSlG3A+2BctcTtuBZQ7oLnbv7U8KL2wJNssyd2kpB0Q3FF63
e2ZBOPPMn/o+kJ51Vg35+ucRQ+f2q9A3x+NDXbVA58uSuA6u+/f08B2SKI0sDZ3L7wZay0d3bXyU
g1BE7bsdTfv3QXWraI/a2v9zc9XaFwcrDFy6R83D7sDbgSkOHMyDiWXPdDgxG/GUcAUK0vsQVq3x
GScNhmZ0CY/kk4uc4ihXq3/jMSinih9X9oBoAM0SCEmxi4/WWxW/KyecrOitMk38N0okZ8i6bYE1
+b45FDyaol8VrKKD9Fggw0gNtO2s5eU7CRpQ92HMQsNTTsMAKuYfimyRuWdeRJ8NcZhOdEpbpDcE
+Ru+ZY6DtHzK/1SoFxU0odPPrA8t9++Y8T9dOwY/8WKn5C5EclP5utgkLLm4wTkpZO7naWP8+k7E
LcuJze1PYoNRxUG41LOntZeqzbYui29OQrrrTqmcWGNQCSZkpxB889kf1D4b8s8WKZM98DkIIlgU
bf6Fyk60Hf1dByXUDlLF90OTasilyDMeYGjROrafNQvC2U3v4cPiFHKQhjgAWv8UhJHMSIdrO/aQ
uRot0ofgv4qfK29ds5Wa5NzDvrfJPWb0JPhxsXeKHLUeSFrl513N9D3Af3Z1kuxORW2jleJPtqjy
jdOmVBPZLYZLfn3ZQ7diG3KBRn49s6vawPAcL0UXndnanBq9pQicF23FpDEYhufVzUX3r0O/HNeC
M0YQ8WsJAKz/zIHshNlYJZQngTpXEUTmrAwn7yyBN7CB2i8YPpHOi4MgGyKt1h3HxictL2BGXPgb
2h7TVtMjN+Zze9y8F/ItS6mEjUMQvS2mqjKTlzR2RE9Lxdnv4nMzvFnIi8ClEO5OSKLkoPF45oIr
3G5ovdJHautoH8ZPlhee0mDluz5jZvb5Q4BZ1Ml8QyUSPmKTAdoDH3uYhwAjjOeiydOVV6LW4GSl
37F2zlQs9kS/PDQgf8oYGCMy3TwlkduVTo5VyPxn3p9AOosMmmGX22FOGTkE2iZcqnoidoc2Zkb6
D08vE69g+HijHXJVjx9Kg3BMQipr9GTIOvm2pFgxKYCU7pq4JPIu2TiBccdI/rEwDtY0/ev9Y9lM
aP0tWa/DFeT4Uzp6NYcj/NyzggYc4Ll9V7+bkqiKl31J6DtoNDr4CvULuOUyCmI0Hpwrz11hlCCq
bX6MnSjRxDeUxBdUxLJ8Ux5OARCvLJqEpLdkIkIakhtgkPtFBNFfb2tVWoq6o9UkJlIsm58TgBis
7AN311imSH5DyKTam/4SlBHYpq++HRhw5wqNepCOYVGYolqp5YmmKF+T5f/gcNwOHWZhwHtDnCH2
paaRwH/klPsm7GT4FxcHGt992kKVjfzm6j9oDiNmYCx1+j5Ofckzh+vvGr6mor4LfT81L2hRLuIM
KPpK/DV+CYjL9uskahXflY7XBHNizTyxpe6xJ+JY2JojVRy1JfzU/ZtYNA/SdekqBloSA0Mj08/R
Sxp2pB+2VHp6GySJxPcJPv5FInSt1nUPGR1BQfjOgSikLB2rOc15OYQpa4HAk/Wmvvswpu1Wj9Rb
OAEiA0x600N330qiboYtwH4U5jz8KqO1XyPSJ6VQaT/pQvu3rS4KqM4KQOS77586P3rk60Pd2vOk
++LpxgseOWg8vTmWDeOFGhaHqrUwk9+nWtH9/O189TULOIXx9WmqDyz5+RNIv/yolqYiYO8RrAWm
01yH9hsVOKNFQ+hjWhUEzK8jQvFufDQLOZzfcF/gQQ2ktEQSnJh+1MC1r6504NGRale8jIfrPyg0
wEGrXg6dFsfYJNe5/P6bObB4l/3jksslaM+PgjO59t29M6Y4AEEmxiLX/GYxhZXLFNVdWdWWy/9e
i47TC+uHiDrr6ni33uDYETdrA2TcpWgU79/FiF1MQWs9hEXS/TdS+Z3F0ixZDnS7gXpiph8kEHPJ
qoO2O+0a9fgpuEUQcXANJyLA6zM5KxMz7pEgAaFXsj3toEfDor9/SI/J8/SeNT9U5UTM9ftVzXSW
jjC7t6EYFnUbIKoojN3xwsflJU0qbKWxGaAMGKe+jezrVWSYLMtOs7VX+OaG0P9ufnKD8hO/ZR2S
f3eJOonSB+4P9Zc47dfK+Lez/0FmbC3xT1osfwVvRHJjXtQvHR8PKYvW2KQSuOvA31k1lRK1nWDS
2RNMjnz18TqDk0tSbFe1LyYpOq2z6q9H5Ws1yV4TrllVqNDGPNej8MhwQCIVb0IVkYq1wAkOu197
veTAOiamsVvigEkDVlhISdA32Lcx4HK3Wln8yGKrQ5uoBm+KLvaL2LtHfAO/vQMneHI+oIfmRr0c
4Veez6p1Nq2ak5d2Uy45ZHK+UG7o5LHbJeW2oy1BmXTSZ0VwCBlzAQNbeHL2BV0ZC9XmqNCs3C1H
ZwSku8Ez0nrHeVGTvtG7H/Pjw4R++qkJ5QQ3UE4FgdbsmIyRxiTDQgWSIGQQSEYCK5FClvugxMlO
tHID0Cyk4Kj+P3n0x4R+luOj1AQmmhesL5TSmm/NgWXVw5kpLZfxIhfu1Gbbmf3SWS1caeSoCG6j
4ZlOQvVNn1JNkdqd6S9nMCpoJiq4xBjFUimxFbetABkO4g3xQ4VF1CP+FvbCtUiezhSE2lVLEDXT
iJ15sN4p8Ob3jX1oIY0QJDP3xouaXk21OFcd3q5f8Nmw5kysa39PS0Fm/B4aoSv+y0tBroRDR3Jv
BmmlUDtcx2po3z2vaxuVvLHj+rlk8LYRgZc0cjyIJ2AA3Di28u12not52nT3/34bZw0qH7kmFNsz
eRYImbfpdhPZ9vciIGAHEtiI5H2u5p78EvJpLmz2s5+s/z88riHA/roDd0YYfufp4v5qwmCI0c3U
EvQZB3eUlNBmXNB5sEp76RNA66X51W2whGUKdSEGTtETDaQwBizaxGrIv/W5gkoMcyFj0sIBfqBP
99CHmEddhApapGchY6LcBPxwnGS5WWwZDZefcDLfuPxoY9vjIqHrmpNaUjs5Pl46/aQNA8VMZ+un
hQuiNv4OOJRkGdzzpiUkhdoieeOck5FQ3TMshjpQjRIC55r05PhUfQ77I3lWOjwe9KcuNs2zEBcB
X1sNHp3d9TVeUnK9nq5N6qPlnQuAp818mraPYLTpPS7OsPbOoEePQ9dEBpjkvkVsgKZ7sSQwRd/z
hqhitn9jvk0ZM79Sqo/xgbUxxTBpJFycs5eid1etEWDzggfnbhC8xh71f7DVH2+ImG5RUkWHFrjP
vXEAYsltGNChWhhlbfIsC+QZeM9U1KbgyJtcC/xNPIsz4HXSSDsbHfG5BcERiRUQXvCsgmiMSyE/
f+8Cqj22VNrhkqqG3ehJaXMbEqkgOPii17TEaSEUu4T8vfQ4Y9CtSzDgE6whANa8q/D5J+MUuYsr
/mTwy/yoQhoySZzQaGxkQgafvMGs6LfKKaOQzfRcGo8ZFZocPSbueopbUrkt2bQzIgjry9aAr2kD
lwhjh4z29YMu0poroUK9OVyPAso+bGe3NgNAjcwl2G0kZbYg6lK9xWw8MR3LYbPZmfxVdLRlRMi7
6nKelEUsGgg1OhxVWR8PIwkUKJjqD1nBiP3ZtDh8bS9bOWVLxXiqyLnlMdBx/94DbVA9kYxWMcQC
V/zju10vKrE9A+1t8t/NFF+vySktD4N66S0vriWQPNALtKjRY2Va+FIcW98vPAFV/K6OLkPdSc38
NY9kEFjbm4y1PC6PnOaWuaNYDQpZ84dQqyJ5o4mVcYhEfL1qEU6JS31UTb1vl8N1Msl/pf0il/Ue
JT876QX+60v0e+sfQeSxCfgHq3LTLKuhJQj8nKGkLkHFazWqgiEfRLilV1PETR6BhCT270n5QtSN
14XFLr2CI34M7NnpaPdClWpKHI5ajwx0AeTJLgdkFBJ6RUcPM1Gd6k7wSI+lcjp1XwfLdgo7MlMI
KWv9inkupvxQWjFMh4XnlgywrNiioqJcg9SAbnoqCN0nvxgkrloZJGazx+rjXVpF4OgOs0Q8ALQL
PBMEleD5Nx9R8bpRzQlYtI0E9O2UyjUgSCmbw6Oop5YaWM60IKb/wPSZVKtUgYuhKeAIZLVn0J/w
wQdKX4efpF+OLv7OKR9T4ld1bo90gbbWypH7zZgZ2Ut8SwryKNlaSjbbVl4rIecJPwZSQTAFTOuc
8dz/B7HGOKXhbtjAwCmyW64/xi5qM6yYRjoAcCMPFLIi4VJGF4PUwOy5n15dhsGXx0UNjHgXLxBO
ynXU9rqDYyrO5kyVIdHXd8Iup+mr72zHWS2C18OYQtkc+HqoDc6e+AIO491e1NceVBSKfb8cHeA4
3UdDvERKGZwuElEp2M9ytCG8DfltkCUXZhJrrSQ5N4nrALGVUd4V8SoG09tDES7z6ZAbDXUTGYcc
gZ8bLw+G9rsLSYqhbW0kfxo+Yyzk7EB8Ii31uTVvsVVDMNWwapnNBrJMYWzZxfOROzPK9q7Q71kw
1ZLTs/oOAt3A4Pdk/VcJVF3v+4ZrnGp+nDcZyJJl7nRoQ9fdusEvLiowH8T/ZTPVkUZjT5Rp/Q+4
QcStm54JHN8px1WRsTRVPfAXIQ==
`protect end_protected
