`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jNvGKMNtWEUNKagzcg2Z6WIUWv9gWJV7my4RvssH/ux/cX8RktigUyw+RYrzrXJGrNW7g1x/nBwF
74yzP41Y4A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cve4pj2EfLuhqfhnGnOz5iUJuIGWUldTY5TKWZtU1S3TPZ4r9ymlKXit4YnjR9S0JtAX1GoFuudL
h/jZOj05rTC9CmxzpO6a4qp621eKZhXdyOHyWMf8jPXE24P9V+aRttTL8nXifMfo/UFfsvRfUHHL
a0V7II16UbNY0z/aQ74=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FK+UvGaeunWTo0SP2EhgyPGTZaNb+A6fyrB0Pb4mabhgLBujusE/NHHToooQsIrVtG+iA4L6uoFa
xZk2qbFfIXLgeHkE73Jf9tkvOVSfNHKkwE4Tk/zJ3hux51whzpeHeM/jgYHXV/AGxAjK7wYmqNEp
cavJsaWgLnwe3yjG331MbcwzkmgERAfcBrC1i6iTT7oe42Z8bgt2QuADWtJa6+y6yzc95b43/J72
7JqV+DovmhlKbNR1biVaDlEMoR8wVeDr0xj6PecXn0O/DCkFw3POXJoaMT+xrRj1LksGsCY+qMlG
IfvdA3kKCxIRZxGcAPvET4wf6cGXK4CAVBa7IA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
z2wDansBNwtedB12HDIWNrI0jJ9Of4AnAAv+qKssr7e7NujivlJDkMFVu15DOLNgNtFvyO0niOHn
/kdDAjIwQtt+ugBkFsRzbHtzg25iwcWgxIDasTP9xLaasNHS5B2OfeSNk+sAZRujgTnv16OLLpuj
xCVg+ocyScQyJTN2fY0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dHaEE44368Lqz+gkjyTg7OMF1sLix1urvVlzCGNFKkIp5zxC5Hb5ei+82XYKqaRz661xkzrxnXIz
CLpQVXEZh1wM12r8fA1f5G/ZuHgSsoz7RWoNbHd4G2GQJUG7WVKCnogPJmbAQZpXthW3KW14NIsi
E34leEwjyTjx/frRrPczvVKGoZSH0tKOZiCD2ER5SRLpYvlTJUkcUEXx3CipAjm/wVGV6SSyQJeO
CTF45Rt8GOFQIMhL/GO7xMB3lpMvQg6M9+8i4GbdQOAk3MmCg7nCiIL/ptz2eDE+txQ7xQlXt4Cv
Iz7BX+6KUqHhfTCrqRi9bRB7HwJgifi1MzfmqA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4608)
`protect data_block
dBSVDAWiIsOQDtztSiCUKfDVOQ8T9Vnt/iNMjyM8Slwc8JGThs/+cCHZ9UOmXj6lSwmVFZWPodhx
he5fUQgMauaanjIbqV6JEvrwMWetbjFM+bqZtune/XuTzXE49vduWV1hi98d4wFv5Hqh7P9DStdL
EiXL3+QcHdJ9a62tbCdlazftGpifm0pRgvMAaVanRKiXYgNcqqfXVQYITA0gtkphXXYW6jQxIZf7
tinqy4M6R+7R6beFlAOFP4Co+5LFz62iLoJbROyo2GSv060tNTQtiRsX9wjFwx/vtwjtS6ddRXP7
uLPu6M1FIE3WSSjkk+jmPgIerEsTW31N58Ki25JJBFyc7ll4dhC7Eim+nNdV2So9IYYjmq6YUb9T
uOER1pSEyO7FAqGq7P3N4lo/aoKzdEX6HTLKkdmD+bCTH9GQ9BK3WJ/FiMDK2kdZXA9HM9a9js5l
u5ghx0w+Ud2sNAI7OCsoKGmV0aGxb38VXbeJAldFbaQfuJVA6aCFjrCZYX6nzaZSKUEsXKVsmaPZ
vAQj0cRV1OyFBbBHF5HoeDsFCHNuWwfE997QIfY/s0B62RuLOlLVQEFihP1wPcFKTxI+cUBDQpYo
mbyikEOjafqj3axHt3ficbCdAh3HKOfVafc/kRETu+4OKlCSMUzrmyEjeGiFCrv6Ma2JQg5k2yMo
ccp2RjQ4tcL+Y2pxfLoHBA/MHlGkmC5lGbGQ37bVxAlP/AWxLvP1Z2wA19E59lXGsyo8fwbS3H46
lV1d/xC/LgJ6QRNclRdhLm8irXln0MqtxZFb/fIB9DZSuf2qHffNhNlbJrGmo93lpi0u09dKWcv+
MLBkxTGEpRXRNAP/2fkN0bVcFgxWSBmL4cvWfvJPXc0BBwH5QRk43D5xnJNJku2yCl3AuhMYCQAS
EEbwAmbsDMR6eJS4ZWLS8UB2CuEl3q7fVh4/S8IXUUyAMEPR11BegBKKD3/PT1XPMfGb5aP4m0/C
QMx7uzAPgUCf8hxBwli9X+2kIDoQABS09EgfLlcWznn318IohkLmGOxKGn3X0GCH3Nu+6pVg5Sof
KeVVtnhh5F/AgRCj8Gv68B2HyOOyevkRGeau4/Tem+SPQ5u0zku/Frz5ivEm7fS4lqPutciDfKuN
HMRbtUp1jQB4DNb9MmK35mH40nz0EBb1JiuwZJMI1dLLOfm2eECujBVEyOidBGtD8S6BhSMV2E+T
vvbMdUHOZgCv56qGZU+4e1PB71t92rm/NnzquiRpxv1jLOom0YO09y5in6LSFcORf8bCoMEnitbW
Mzph73s7CziqAHpVrBKMFDdNg+rEAGL83qbXUuh0FjcN4zFcu5y5oJc9iapN3Yp5/mPFLoZFNF+h
E/yJVlawFqI/oK8WHKXFpp5Ry3D4Gq/dXCtjXmxeqXdedemhIm+7oGcQ7WTnVXXFb8O9ySSnSCdg
IRqI0z79c9mQ8w5P9GwuZudeHGQOmxP0nFL5WLj4xmgOEO/JByzI53VpGMfRmPLP384V0svDPWEq
QEqHp18ghxLEgmvF9m+mLFExvVq4OL0+CEpZh54IXfEw0yjgFw+ttTDKrJdQS2PIFhfbgKw+axHk
ZtBtkq7e/4g5YXtY0YkFHsRAONrtnXSlJ+ZVcroTbhfbNrEmXD9vaWIXtb51ghgW+A5ZoP//UAYN
hUN+rn0HJ4g2m/bvWBLFVThxoKhBCiICU7SkULsraS8V+guitnHeqXzpKut9zhHbzh/oMNyT0Cry
+i/0UQ1r2HqNGFbMbYa0svjFnMQx2KRvF/KC9/h3hKbWXP08Klkv+ODQ3hlXt4vRByiKHMb3fz0P
sv2zeDoU5HNQFP6qJrhpE1APLEVL5pXBH7s5EyZDLQyJN24KBSKmFA5HddUvHB2Pxe2keGLRRiPi
KBUbipL2JXXrciAyq3XacrPy1/1d/ahF/Gdg8GZx+hMmGg034QBI/O6wk43kW45VOnJ4s+BQCQxe
KBQPNO1GrsIlyxeGY/DleIP2dqjZO4CYKElzLt6dB8VaSfZGimd/Sr93DtYo0j84/VRoIAe80zxg
eQyOtjIcZzbMk3taFh6vO4cUr00FUT9dV/YcAy0FNVZQ6nlwYnHS6N+W6lb8RavRdBMVQX+nzDcX
1kOo9siHKEuLuvB5R3u+TRetFdxr9gVI1VAtcuKIt7Ks1r1ESmBedN5XtNo1bkuvqyyvGrJ8QJQv
mgdUhSiMQHOjB3vGj25MUqA1pZt8tRVnvMJNB24R3dxrYWqZfpJIG9Hj3bD0fHJhMLVhEa75DexJ
fW908RBKw/mcP1jQ/EIAaNO4klXzBvRTjdvP4tOgi83ymlTmwvaVcKYx9WcyPLghFpmvBUn4Gj8w
3rDN/kijMDkzlDC6rlJq+fOiv759kAY4VUF1SYb87n9n8HowBu8vILtpQ7SjzRh7ZkoUMfWil2sa
+0nSCpMFUxpFctQV4U9UvgSOaeWHWEiEW8Q9ZFgZ7dFtJbw2F+EDHy9DxWdNt/Hq9JrTl+PkNEFd
CJHCE5FLLc0MczLR6OT+94s0GQTtWiL6ZeevQinIwNdyu8ETFbnmMQFFsIDm//7ZpLBRXrwUeiIF
AWfwbzwFr7TYlZvctR6yBjCI33OJKWl5eGbym1auEWhualWKcO5mELQRlj45d133Bdxc3lW4dUBU
Q6PltxAjVt2a+MAIlklmzUtdJPA77YP+ypj1Ykkex8Y6IKHjiGmFFpC+GYpmI2EDZX2qGw0eabOQ
gUnprg3qmlClVtLmTRfNuiL1f2Ru/4MUrF12bYBO5U0Rp5UASVmw3hylTfH59paO9Y9xBvfaG1H8
y/htmbp+196c9nes0zBfkXlbCXzNQ6sc/yIt1MUxCFQSMUa2lIDT5ouZ9VFMMvG1Egk6vdG5Mcpx
1xDmDi10jf/IazDirLGIvykUo1iZK9U4Qs6pELICR4guZhxcWvY12r3RsMyykfHG97Da4Irod04H
IRm4FH57FSZW9TXfgMVsUzuPLe611xZccg4OWzhqE6Lx1INAsIt/1R0ObMSp3OVC2ASrRGGGqeH6
3CDTIee/4CCdMNWYuuGZTZj+n7r0gObuEeJ+XLUelF3OWvwUVY9/gQFZ1hWZuF/jEZemZIe4lN7F
ocnS76dJyB93uGlXoGJ453SH8VdsKSDlEr9AfEVlv0QgQYOW36+zzaTT9UyLV1YleC/Mg2NLUEqf
r6Zm6cIRtReNtXtkpucQD/ezShw5zHbn5cl2YDKWiB4V14FR/u6rUS9s3TbGKdffHOaiMV2MirsC
jbpC3rEIzA/XcuDc6z9iw99w6rBh0iTpaPxruV9kiTkqmcQQQIZ+2BPOYh5I4c0yTXc3QPAOR+HP
3ipxG6OvN7a5XW63L0Q+ACoP5M4NYmfKNyyCOTBcszAjvYdTVwg981jyW/i9kikn8qrkOvvzb1ro
K6Pv9OYRDkhSEwJjjrJ51S6bT13DVr749faRb4aQSlUcFKhbMP3vUP/9wK2dkp1E97T/Qcq69bFC
XNBmkRXjfCsVAuEXbI45dG7jFJNS0JvhN1NUrhasds2ih2XRQFnSKlEvSiZTcFq7D4N7T8r/yFps
urrGgclyuzbtFjDPInYGiId9EuXsU4WwTf9HThL//iuAVR4mQwcxtZygnPJj48yL48GTX7VOt9uu
Zw+WhpPMEl08/BKanvUbs1kR5VsJMm0MarWyZskOtcGu3uGnThL1+PiF4WOYbE0xnkhxLnBJaXDr
5x8L2Up4Zdmd2WFhYMjuszFUcwawr8TjX8UdJn7ebCqLzhHiH63gHknVuEgkPCqgaIdlDRDYwdHJ
v5jkslJp4hTMn1ZBgQXONh451SfLClI1I1jXgf0YRbQ4mpAcQ64agRlBOWCv3QdAtk01HyeVPWws
C6uOf12w5+y9u1P026RZ6AedE8yPsqZGL8r7jCWHRjRAOTc42CHg5/VT5c1wxOrNFm8QgFaXIAxn
GjsL+e+rrOpIpjzPRMUHYbYyBJld2qmqEUo9l+a4mLAjMtYs/JCORBfhRVjTSFJGFvADfO+ZCd0V
mF3fM5X77T8fkjgkhmO/LU7S82cR/U1p3+7WBQMOBZizgnJZp/aPwNSbGql8+eDbjMNUzMdct9FF
iHsLEiNOOFeoKVLczsQWLxW2QLr/I3FUFeK9CyTK2ZeZXOoUMUST2z5fUSzMHkM8JQR8M/jjR7lU
G8BzMi+XKKYEn1dY8nf7bjvMotff94KKZ0aqbz9qBRECyxYFvLXEAXaHZjJz+QOoLBaah24y1vV6
ESJVqqViyM/OixTG7MAMg4s0exC5SkhZJkxK24RmSele7W3oX5gRgKVoodgI6Qq048Q6rdvOEwx8
rRcYKmpLKiYzAvbuTsdwN/U6x8OUCX7irYuFcLSPNMrns8dcbwpbXjTh5XhTmq/X0yyb1FiI7sC6
OWmXdnoT37ICm+QkCQ0u2quFCDP/HBusGMT9k3lKaqubh9WMC+yeVVwzYQY8VXzB9PPNshOy1jpH
rVUDaDLyy2QNL6cXrUxfgAR9W2V33z+m8cf2J/b/2CXIVxLweIALyT2OeG/uMz3amTAeJxLgyp/t
/GZcIKm0F9RPZgtRONhuxX+aASNAIJhf++ZU+bcbHBDRkjNs1NIiArYl0BzD0Ky3ty4iMWuv198T
qTjb06G7Y7+Cve1PXwoTPZpy9Ol5BaSVDMKCJnAfs2duL7A7uzL7NxEFT3XF42N/c/GF09+mKhbQ
YR8AbpJjzjvrGOqgvbG4eqahZfVh9wtoxE6+qOIl52Xt1QsJl4gSwmt0/R9f+gyODWvP7gbae0Yz
HAJcDA+r85pnhxOq0Cds15qVPcDN9ewNxNxpBjRJ+LsTX8aXFPKGYHuYif8bItQqM9063SoyKweH
MfxklW5Pga6I9T0TGkwBsKQS5qV7OHnge3D6dcrpTfoiddpVvTZIf6tTsueXIdJ63GT8yfJ1RyLf
KgWOZjYcLVCGXmWYzQQNDDI0JmNcismJ0mnjlmO3nnRylFwWr9ZqkRODqFFR8dGhxi02Tjhm6iyZ
O30hpbfvj9NQ+M4w9qlltrypts57ZOhyKynpNN9Lt/nMMk/UIUqiOM72pwBlLare9vXedqsdBy9r
HTzB0RsyCKHYPAVurR6cUEyxOKAf/7aiEUzonosAl3lIeK5DbJsnxUFrcWkRv3jj482VWeg73I7B
x3EK7IFBxPVzFLo46eZmoA8CRnRrVbR7WoZhmaTmutXjZpgp1NCsNPzGJMUErJQ9IcDzjZgAmywe
PQC4t73Cp6+JaHQ1ck5eUhYD+2C859UquVN0LbmWn9DLcbgOS8phL2JRVgzOXHlhMmUhnWqqmES0
K+GiQMy0q1DGKKUNLirpCLNUgl6jNjLqVbZGgr2VM6GatOMInzcxspBcdFtJfLUBCgwZBln5Md/V
1VLb01W4tbwsKEGsTzfCRbS1l8gvsBhaPb8x/tCrxRLxZwAqicCrmMCYLkCNcfVBFdP1/1tWZLCZ
UIOYD5XWnEhkPCJixEPkBgZM05g1n/N290wc+HOMmhivEtKdTVtBBqt6bu7gLCyF/p/kfcPZwSjO
HEoLjqGq7OR2tgG85G0eZIeRhRYG3uxvZb1O0WngUQh1484mRmVz645yBNupMUxrljEXav4byJTh
rSYJPTCPu+DYft9MA2YBXQjycKp0Wk5Kh4r37sYZtOQoZdvWBxxtPXrXzw4bfRd8DjldAUPoYgzD
csFB8L7204EWzT0C4xw4Kz2xyi8+wnVNqSEo/Yp4JzOrH3cKqtkqtH9BqsrwqN/S1kXxQxJ5/Xi6
yFh9RGk5A+MMaT5ealaD+dfgN2URwJoTCdi9u+LgFxOo6TBVOGPpO7XKMFPFTIS0TbLLgpQF2rQo
Q1tYi0gJ++Lh/EACzLSDCk7PKz03joC4K28MSM6WaO3w6Pv00DMlhzn0s8rdjehlsOmuMucPOyBT
tsGGYqANpM9Ybaj6ebihwgCrIuYZsEn5PC5XTT57PrGA5GsNDlwU9fQlvzeJZHfrvF8pbDyyuJUG
nqXqcPIbISBIvnKM7Oj7UBkXA04WaI7a6KIWVhAQahbE5v3Ra20pl26pBLoH7UfDth+alM2OvayX
ALIc5TYCRiFOuDieovcIeh+BCAHYtRVbU5dg2CWi0gmf+fa8DUF2lMwTxBqdOJ7s
`protect end_protected
