`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l9rLb8eyF3AgALThasPiNG8/4BBm1wwJaB24bneaCtyp/I0xi7SHB/t0Ctv1xqonweX1MzV/pVKs
tQdRNspPIw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X5KWlL148JabgR5weT9wBUkHFWddJA7h4OZFLd8bdBf8Kop7kg1WdkOhUDgmpNTHeXS4I+xH4Y4Q
HjFAExnYrGUC1wm7p5WVL3DFzD5WTILYoEImzLFNcK9/mSAIwCGj+Wtr+9xrMpQDaly5jC8Sj+rc
Nr34z/YYnZpZdFjSjFA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XOX+x3GXJVQTrGGT75+NpApkQTW6W42cmWaYkzqsNsDYv4er+FitAoIemlb3od3AsSf9WRWhCQnT
6iXQilkemT2DzV4Xsw5A/7I/FZ1E441abMpjv/w5Z3kwpJvNtJvcGvjcX812mAAPcXsPvrB5LXuC
3JiNsCaNzfl0IQulHvHCqzDHmgFxZRkHPXNoL3EbdAxxa3qQNIHMXziT6TfG6V4ioLwZkfmj+nFw
X+PAA+oZbdjyO4IF/qvCl2mnZ/REv5vdMZsnEZ7xmZVfOO9rMWwJcGnuuXesJxcZqnyEOewdy0X4
g5x7ACzMTBvW4JyAsNl6ipSaUUNJcxvmP1Z95w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
umhSCUCmm4WZMMJVCjLiDlzFgH/9KhaxQqdvYM2gFaFK/BSZmXwKtVD0oGzsfgEnaEnfAZpnMH9p
W4FaTz2HfMA8FyEQD6bKpLwcrFDP6FLYTus4W9auRkdWk6MByslYcfESnbPd9BplDCjnq5X9FeJm
J+EfUISXG1WULY3BqQc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NcJ7q/waCn8/m5wYTzYlcTzCH0J7XhsrCXDcbP801wBgwPzwk6W1YaeEGpz6w5sg9/BVkYMZPdHy
s116tGvxEU4yIAoLSq1V4khC1G0CICk3cYOL6Am8EnS97sHVRnu2owQQ8/o01YRhaorvw4ApXGQo
FWXh1RTAkyoxms7xpWs910xGCq+5ztWRsH4I8eissSMkhuy7owGmA0f/OPnBvz/16ynnHSqeTcgH
5zrPaJOgTZH9aMea2bstTOpguVDKDnDoAXUHV93yikhxVZbDx6GaPXUh5fshHVEaMG3kP839Gx+j
prw3SfsWydM2YztaOjt4rwHOeUOZ19sYd2Gsaw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
GMQYRLdIBu3cBPESIImpy7PD1X3NOwgl3uhy287mrcStdm+f2gkMp4Q6NPO/6rHSdrpD/TeCxwVz
GQFPC23L51KK7Ng9wRlWjznNMKef1kDzri8KAukSc/hxprw49EtNN5iBR7zwbEoRPS7X+24vgQgL
opJXSYkXXWQlWekNbLmj1032D/3Y//Bjp5ZCyx/PxgF7tzh8Wl1drdga2j3Q3G8cPHpd3vs5RhYx
bbN5pRcG4QYhd9Nyz74MWT2dRB9Fa+BSv5d+d4CjKnl+HX7hyDMG3wIIjmO1ACmxN/JNrNi/Ai8H
l70nw2Jf2n61z/VM8euiKJhukm+nDKTPCZCYvMRfYTgeGFnB8MsDsRcwAfFiIyPKSifwqc56F1Vp
iomGFZPDcZB9xKA8xxYXJcVyIOcLjp+mIkSL6N9pTbeYsTz5KQu8eXMtyibAhIqnUndMpxQYV2xR
L4ssQJjMQcyFEQjIsTY3xQRQG4RduQdhVk0co8dgi7Xp53ucgje4sA9Dq1gKFBRy7QlWxR9l+AiQ
pzlCuNGn617DDKOKLcuZxGa2VxEhCH2/ru2WqFWmlP4mja83De3mduMn0lNR3qpyYQzupKh1be8N
7tN4pqUgtp5T1qKzL+RZzMsMzzAWI6KIGTwVG6AOJGWOdh7uXZ6y1QlXP0eCDkMkgOOhtOQRgKco
lrag22plSVZGFlxzI9btveJC2Beat4eVq1lhxia+vvvngjHB2ntzCjWzP9/WM1RNDzN1GVlMJDID
dHmQQoysXFPJ77tU8Jay3vdOLHrfttNqM2aj9Vdwt61KC7bL1gXD7zoKcsD5TiKWAg4m146imcht
/oaNovdv9PWR4NTOByHZnhCdvff5ppIgb1EngiitPCRgrcCfRw15+QkfJT+Y3jxtqqLvPWmdTdJ6
zGQ50imZ/3AZiEB3T3KjMRRsBe4EYvloiSfj8q/73OwNO6zrrEi0N8I//aG4DE4e3G1bQwYJx1+R
lzeMahp3aeJOLgdY1UZLmlaC5Ep4YlH1lOa7ixazj+nAl/nbcx+ly5q2cMGXiJLJtOvdcF6qeliw
kwk2TO6xBm40WvFHI6aYLzTClx+ry5AZm0jRbABd0ggUzK4T2Zij/fR/hVarydXV4imJx4jzNso7
CBpA/D43oxX8WaYMPB3m6H+S5OE8PrW3iZWKTLBql/t7+TVY/EbBkGaHLFlG018mSSU0z9HdKRND
nku+oMBqSwpgQpWSdwj+5Pa1jENHGFl3WTHJZKVKr4NIUrA2TOi/RAhCXqeeAj9CsUGjq6LfuxWy
XmDcyUgzsJlxtrQBtwxHB6TorXaWHaZdw0KUr94Zsj6g1qVJ3RSPywnF20DyKKQFHPnPsjOZBTVg
rUpFwcJwHCpHg+fedRZOwCvyBLjESMMeHCeSvJJW9uE92ojgVs9FMsdgAasIdrbI+BlBf4N8bh+3
RaVg4a4vaY86rANQhHMGtWM8JTeve5z0FqhBEHa6nE3IKWOrN8sOvnD5KcvhdCMif2gJ5kCxc/wE
y1I6YwHLAfOsusPbgiwg4sjczhtLmT2xwmbpuhqQo7BjRcgKYV3JceYXcUUaf++McuiMMaTDF1fF
1TVQ8/tiLQfQRbhBHa5uus2/ywdHdU3NGHpRLF8BCjYBNRcqcUdN513KlmPE1I88UwvaXKIyzSQf
ZzhZfZUxidCo+fTCLgHAM8AGVOX1hTTy+OFGLTFJCeh/R3oimUitFquuLLKh0o9zBqzktEE9lqnp
0mszHaOPvW7OaKbay5R/iF/CrmXhcDnR6WDuHEFAn1Alpvu3CiDz/Ldywq5nG+v2YagL9dMKSFse
i0oe+NiMteIbUC3zoEyS8KINST9UmAatxJ24kxvrksaXEEMzT12tWaho3b8uMlAJdVIw5Ps8X4dv
4pITzZMWaT/aJgCMePYbcvi2jCM6g2J6XXMlLVBTnaCRXt/WewYlAXr+nOPQqYHD+t1IvBIQacy7
MFgWQ4qYUXTrolk8DCOhLe6uxEgfNwyXWbjSAu2mEIvfjWT9Yd6bQptzQWvLHnXVfEVA6vRketCJ
IFg+69bIgWWJAS5hJEcdPc+SaGgY0KXZgwYyduyR0g73ezRXR6sm3A3OUkhNd4hfOsDyoW3qpr2V
ZLhwdp6lOidSiWkCvKywEJbphs3YXswUOs3wqFWfTjcalJgBO/e1UY5Sn4E0nTMJ3G+Zaj+GkKAu
zo9UZajNrWK00Umln+6mC30OkOm4lNqzS7qE/fwa1qqqSkwTcNVksQD4rmkD5jEe/Z95VjCFzaZ0
oVWtCSsQ5DGSd41Dm0qwLGYSmTwV81TaLIIkP43+O7pt5S8iaKxGAo++YOo8ANVuYM3cJdyolent
81ddjMK1GLMhAQYoUWflcu5iRLsb3QWL/WaldTfqEMsmxfkIunUx/OlcGc2xnoOPRlgraZ5lv1sp
JTVZrR8CdqA18duZU1D/DydgYDtR1vpfux5D+8004uTsDDLCAZPHm59lfL+/nYPvCgFoRuSayoOf
2UR2CamwN1NJXDv7a5TmJW/X5KLVzSsPNXLEQ0CT2F66/p322T3iAkQ/9SQOm8zTm07njmVKxq/O
DXvPChvcsckaBsVAbzK6liB+zfpEPoR3cImARQm1/Am0Gptmt1YSzQcUT22fZhs4QUq+HhhtCN/u
oTvrR9q311BgvHJ614/OYl3fNzNAg/lWubYmFoaCBAdFvRtXGSVTimlrQtRbDnEVjuvSAbroU4Vh
7yO3lCBsP8+G+gfJz4renEyYjzB3w+vKyPNG7nZdWw19GQBfmJoI7WLwFISi0udMf85XyFbHbejk
CSwWqu2gVmL4E8N24/ZhIIeN0BBb1cogLn67EWifSBdNM6/xkJjr/gG1N3Z6mSXZSwazOyBAO0yR
m63SXbJUeEyjVu2ema60V7wK79cr1ywcy5Px1XAC9Sy6oWtTelHJTYDNX6aULBs+q+RiCUDUyKDG
je+VqFFib3yPpINT4jG4VwGiiB6fKXxvs8tW2io9wYV+oBw+vOrQZDYUNTY2sOhjyDAGWfYR7i4y
m3vm2iat3rLUYbE/4pNC0iATltokoz4tanYXwbztJWYv6YpGeca7Vm4v+ZUV1lPCGg3+ivVQ6+PQ
S3rTENmMJGb2GS15qYvUgLZ/c1NlnY0/JXjZu1XpH0WfJ4wX0ShMdHymgjAfV5rqYZSaX4V3paYN
trmHA+WiXv7qms2kBSLEQt0gt4A+B8+/TrEwMB8JWMj7UnDSyJnWNzwVLpbCzfHinMkSWmtJST67
4tP23btygVba+r4Q3m40/qKAPaVQ9w7QfAggLEn7JPgzIbfqZhHjjg4cYhOtrJEBsMjTL86Fzrp9
T80ybToaeStH1ncidCXHSbLPUgD4C+uwQRHWLnsm9qk5UdcakOKdjjSccM2uh/b5SpQAXzdGyNr3
yveHj78C/jVrFLDczwf7//Q+uTJ7F7AAfV67N6e4WsPcvraxP4r4aXBVDyTne49jYrwEGsXBocpZ
FX/65kYqkAygwu+IAQY7MpIdcdg8ERZy71t0VXtdFu8zjiJzUkdFAudiVO6ZEsplcdfG9PiZGUHB
vBaWt0XDzpHnKPFrQ2gSRVos1ewJ6XMQ50Oh6dd0oQATjFyeAh8nE+s7a5s5Lq4ElAIaIoR++2vk
sPNFN2gPAQfqrL6HtNfLAp2AHJi8Aen5jmZ3leIiLg9OAUlDEuiPG/I3Q34QeW/WuD/Td1++7MEn
Q9XQsp3t6Q9jsSghJ6muB9+lY1yw/Uc9OdQQupGSCKHnMXITNdUjvMMeDWVeskNS3o0Vd6Aamuug
TysRKVzHu29mn6BoJmtX5/Cp1WjJIWXKh+VIITyQtLAJ8RYcvVckCyPnrrPs440IuWitM/hzsPd4
PCJy0wsC9lVZyVgRMALDmftcI0j0fsAwgcqSpIgGy070YabvrZVboTAV28tZ6q4D11pjpjsFCj13
21f/YP4HZ6RWJWcPjpqjLHEtBJLVR4gxde4OxzryechVyj2J+n0h2n2o/hnRERfLXYrxflbNr99e
GFDTT+MakVZ6fFcQtbW0qpbYVY54J4p8jQ1sNjziRDUWQ+DvaldATvLWwyMI/368hz/W5viSO8NY
+XUkPbsF5tDeQGedZzhSEonciGzW7uNxzH/9NJPIsWfmNl4wN46WBzauiT4QIPel/qSIOFU2bnef
vtahQhP2CJKfFDkVMzaTKKPtvstIr4W+iXgkfCprTZ4RBhcgO6dHYsQjJsTDDa8q+wFbTd9X9rf7
IWYAgmpFrMwkqvULh645vCFym2eoPohAZ2QpI8LQeIZwF9YQ/YQqFoT5qJXkIWYEQJylY8iHXCA7
I6VlkEXzHgRUCwxus/2O/7s2hueX9Q4rnL0qvnTaPBMRzdUlOk43hJ0HNSyCkOxz0eUCMmVGnIxk
Qriy8GD/OLlHfa34CwPv9+mYIePpxJ3BeOwFteLU+Uh6QTreSc+IJ6S1+9C8D2bwiu0kvHvc3fLG
jucxzyrHur5Ua59PNtuEFyEPduyZPfpPDCofaenraIrEH2qehmz5wG085Q6Or0IFDe+HDBZTMelo
qxekbGDnvdwJlq2om8qq6F5kzCnXz37j8weqP0VRMTyjQ6OSjAukjCMUtgxiQj7O0n7Ytgs6kC6j
eiaW1dyGB6Hx+8m7b5qNebrVJRV+V34tkvfne4DkrVZdPwVSbQ1L06iVH1iXkr0vTokzesQQtzmt
6ek709XFtk+CECe7RsgRHB4UqWCKld4VxxrWP77uOs+DMQCWGoSclJI7HMH3heJMUufc8nz0ABak
w4cPBU2llS8IU42+/JEwt+oxde8mtxfON2Lh3/k4u6ajfyI6G97jBA4fLT2gD+5IW11QJCHfs0uN
EK7wrcBu7JWyXyVChCYJSryUyZn4IWuy5Ve6wMyu7uM0M44SqiBPujDuC3jSdoQcqmbnDdWLbeAL
nFhK4lAo+TU0+5+mszBg7tXaNKTkKP8+y7OOrus3voto6rytMyZOT+su36nvrl2En5Z+v0sj49UL
4HT733djRTnoNPJsXJd67fh6ksbgFfxG5WBJm6F6XAmqGLWrVI/XEdGrKdsvfSV9uOu7Feh9N5Up
uIp5t9bDvv6JikBp8mcXxpZIroo74uOyfHBTEmgECarUkQGHvs6ry5IFx/6zkjN25TnmuFTu5EU2
YvaeWQscNY4kYmn/+Q2cprPFDW1XxetpwHGrr9wJSS+NujIjjjMJbgVv8r4Oc5MSKGDybz5o9iV4
wrBKTCJX5ZFoIQluovXQk9+UcHaW3UlaPOh2yS0GvJF59mqP46YRVeJWa1wuAnXF6X72/xIG81iE
xcyVX+s3aL4Y/q/2Q6U3VYegpCMePezW5xpvoCXPhdXAlp1gCYMRFoeBjObca0Aitm7pcHj0qYfD
BmBTcej4EcGgm9rflUTVmCxTFNOxjSGBMN4JYfsiWpTADzEW/VY4/Of3WEOm3NWvnOqju02/dOYp
/idgTPqkzxOv4k0fQvGntq9L2j4DQ+c0UH8FFesTbFbUbXnmBbNf4ZShIYyxqyoYhUha6gmOPcQ0
LvPVodsyu6VAgNgwIMvH
`protect end_protected
