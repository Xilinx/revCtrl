`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 253312)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbB/zJnlY9bLi0AUFrGn2gHL2x2kzl
0IsX27FVgcMWfMlKehto8ZKyKhqi5agZner6cGv7npEsgqK0Jdd9TrzqwTaLmjme4zMM4p1Q8+PP
gi5sOqBSvQOdQBEYJVW8Zv1u9QCYR3qXhstGxCZIPkYRP2DItguhFlFP9r6l4Vztp3EBO976fI6h
NyGIWQeshooPt5R0QjtEJlb2GFxS4FaBJQPhbEhAuu3FZNuSJr7n5dDcKlJciCUIDT2PVRsbNKGn
NyWzNyP6aIIFhQO9IhdznAezR6aqh/j3Jw0Y/DFoPJmOw9RWC3cIVoYEgXuwNtg66reUHkw+GekL
nuzaGxpZs6gb44D5+k2eXmE9+VSREFj4U7We/UKaD0UyIz99yVbwCo3+KPOkVcbYWcFgbXbe0epj
um/X3P14N1VdkggLifmp3+MQ+JdK3q9wyoMJzl6kXuNGQdvPJFak9tMb3zrQLD/97uG6UwGPssHj
wF8fIQfaL72AECozRBx1KZzrfSyIDkSecfH0OST4kLix0yEG1HupXm2xVSqOj2YscyJbDZTeADaK
xA+/yPjUuRaXXDKdvzLDVBAsJqFux3+Mpw3wqQQ3yT9h8LaGb/ZZGvf2eSMy6nnWWC5PoqwWE5pE
vSmScg05svgxHfur4+zct6MeC5BcOJLFYc8EKOU1tCEiC3e1LtHFOGDXupj6Yeq6WTP8U37lrzVa
wGAPLw/8uhunP82m4qL6p1l1hj3lY9yklMMN9PC5O1moOgvS5YKpQoaq4Kd20v1ZGAU16H+BRchJ
4MMtRBRIV6MTW/F0EFfeVxhZvnEadFCMIf0cw+2by/NkC9xvjk3hW/DGZCuh6nEDxumksS5v6Iyp
s0DfWtK6iDKQe9CS01wXnpO04s8R/wW+Srxo2cYRh3j/5snQ76RJQHEckKJMz9xZz3R3tCBLNGZ3
/mkWQOVFC383OqLBdjOepG7diywFCAdHj9Ch0Chvwgl09kiBxRDG2KHL6AnDK4NRCIX6BTWn5PLQ
16PShb5JA9DsBv5y1EqBiTwXgqv23fx6iRUG6PoNI9ZjP9IuacRLgJTatXL7u499DndgAkUzglmI
UxQIksqBxm3vm0eGSn1fyTZzZ25pY91osQfGKClgCDH0S7YExSm5WAS7XCFSLHrAV8Zyz+dmh2Nz
I0tptgb0RATjUqZbKADQcwppL0ew9AyxBZcBt6uJeddtFcSfu20nXw+OXUKCJQY3ZmBzn6x/kAGj
3lluWw9daxyeB16oBRz9k54p9BkYLbnY8+I8Z+4dV5sU7GFkTDNWi3C9+5ycELBKbY3VQXivsIPo
Rvu18Vkebb6A9O4XAlpgpQQ5j6q+E9YXLjteFXdI5/j8mJm3l6Y0VwXdpJVD5jVcjsvGQLvLfkvZ
dduWKTX5CtynAlHVIA9QfUDhzxuZa2uAxFk2bDFAmGpghOip9fyR9kmw1yaPZ2meH/95sGvwP1WR
A2O/ElhBvn9rwb87laoMBCMEq0aIktP69BGhcQsrBEtJlc5DBXPQmKAz26i0NiCcj8wJQZc8wyU4
VoIMmfjGI7jx2/Gu3zZGB+JyKMyWz73UP2TnAB4qt9rqorT+APK2BQw+MVz3MuhhiPHRQuTbAxNF
C5QldaWfRYrb+rc3FwdNBIFB/mFQeNei7aX6JWnL4sDgomH6hXETP4hflYauVsvSYvdzCXIRPcdR
IqO1zE/YTbkoZM9Pg5cwkebgP21QBGV74XYiDIhAvphciDIGTF6JnkGQMpjdqZB0ukxi5Fo9GbKF
7Vcl3sHaAd0Hl1avl+vfRSo2ECGD32zONvbwEalJVLHF+cHvIcsVdVW8dqF0RBqxcOmE1PPKXAkb
gd9jjfengu2eT+qwUj72inR/UfBY5z5x/rBF3A46PvgVW2L4C/AT4Ism2GsuKIoL4SmKpeKwxI7g
wVGS10ejIAtd8FZzs8kyu/gpl9YWteofBweva8su9IlAQq46DTdlzjgudRwyMF5asRdi8O/YGWZb
MyAbeVbe44jnRvZZY42pn8eETuVh7905XcBWBXTBM0Df3MltfYraR0kqsn9yb4e0jc5xq28xzOnK
XPnBg516mahj8LRpjP4mjJ3u+5aFhTXje835UDVJutOjqF9IYUGaH0j/fEYjW5lZLo0s5VLS/8mz
y2KIK3LdGvbOAwV0TAYw+1xxpcEMtq4HXorZBfzYnyAYfuIxo3R8LI6cqy+0t5ug+T1+iNczygbY
AjAilH28Zuxrzk4LHgJwccThlU9ZluiLJ1RCEbBkPLxulTzO7sPL7YEYo6bOicoO1fZbegEcTsEY
0kwoehlhRdosI8i1+d1Dywc+4VDfEgVoETzpCUwbFU4x+BSY84LyDdwNVmPzgW9IRDQcRrtFgbQF
d5x2FBdc1uW8g4iEvHcS7VMeJj64Nqedn0QCJJY+O2RJ4VCXLQuXVjEEFlxglyn/JbMKUCTXXGun
miqRZPrydWR33SOp4SC3/J8UfPjHU/zv8jIHMCTWwjlfKY19gYgFbqr3maJCLoUOM9QIkVtRY6NA
VwOaGLp1BzDh1SnC0tivHq2KwnIcpO01WtthM53Vz0RS0tTm2DINrkXZkvII9ugAnW0+nnInAdnM
xxqzcR8BTJiSuoUInCpI7txOLxnW5Vxl9nP7Eq4oBz5BZ8qFEWiRQpsOPpR1r+OfAv/acuwNYJ8D
AvG6aepQakDXl5n0tYemscmuXvi2fgmS5oeHmoepOqD7lGkkvbyfT+i2CnLp17s8n1yY/m1Wr4GL
gFei9ZmuAjBjNmqCA8aQEZ+e4+1ccINKVnOrQdYMHPz9BjhpIyxpzPsvxbX4CaxD6B1nnlBdqxKc
X/QX2jw628OIRUaFZeCUjrUTJMUqSvs29HGbGRh7tRRXI5T/rXYmDRtmzFn5BUIcwl2jU0HVGX73
BBzJpFI1DqYBOlZGV5A928f6/pkn6PlPLXm/SECsV26I+vekd5qTOcAM2yJn//etH1Egp2yVZcWg
uGaQWHkZWIB4JToie8jaUnQwNn28fQfzjfY5S1AErgYBoJnUEFQFRz0ay7CK3WddXJfxsQdGqCQl
ymNUu93sl7UoeHRWMihIWSKuFetSRexUKGCI2HE+TA1fJmnG6FSYY1K07jIlFWcLVVg44uVCQnO1
P2WWZEINqfGV7T7DcrMteBZ4lWKPzwDfHIXhFuLlLdTJ93jGYGd7SDQT75icRSh8jwsME/RBB+va
5QM77XpNeuDISaROcxGycnPtxmXZEr9j9l9KQg1cE69WMoECJuCPvClN3YWm3Nq6OWV2WoCNsLmG
Kq8I/JeN714TZKyKoYynrVx0RZdYbzJamiMQ2s8esf3tswkMO7Y6GXCCooza03O/TuRGK2ekZZhM
wORqyUekI3CAECBb27Fp5rIoINCtzhHSYwztYJqvKuGCt8h2vXDTeUiEOgYQXtQKoyXq0UmzOPt1
BFJZKxCB+Xslt758mQderJg1YbKepvB97eaEOnN9K8hpr1FEiqtbW8jwoV4bnAR4np+Xgh2miur1
p8oZjpPazeRAIEArEO7L8KtaVugCF6/HUE9cOizAVoWMIkrc5uuit3JR0Pcf0gbfxeefxqaPubJr
a7kLihfXhnkWZkq5YeoeFNXTfPF6UUzc47f614E6Jy4hRJnKciUxJlMdmfnK9VMrmdUkpCtTYQEq
6saPFQ3pfS7yTJzo3I/dC926nGkRpJP8s+oAolJIUMRGbEVvthZa96IDZAVg2May6YeresppLAdV
AWiI/6GW4/36GP79tZlBbG0FpNeCxyhFonK4ZV/cn2gf4T9lHEybnSMvNw3qUPOw22d5Gnja/3cP
F11fnUVIrY6r/eR6JC9/72ZRlgIANIXkpudaiSAsmzcBgzloXiJmSe/Mn8e2CeG4yWaLY5NhhkLQ
IRZAv2FVKLq3Wx8068tvccobPzuOQMvEaq5DrlIQ8uIE6YX7mz/F2AEqz9WvuVAoybGvmpiJFJXo
ruUIFG+Psf0lZKKysB4Gre5K08Td//YbNV1+f8Z+tMRODMpBA4C2XJPzBGjVQWqqkaanDGDv29L7
PUy92hrN0bd18MBBtTLG2J/O9otoTUtyTqOFY4DYAo0LB0hKkEClSaGX301Vk0Yqxslc4Egrm8PD
oL9z7ZE/tNCW2FGTyYzhMRMwJg5VqkZ5Czd8vwYHAKO0BhdMoHVS6TyDOVWxX2jyiVyKvYhqfeYs
sSuJMnYRC9QsXekRFCjlceTYSZyRcdqGcTOvEFUgL645wwXrjLP7tFZwSnz65ziGJm/5L5fA7vAJ
UOnTp2a3TGD2vEnbRScToVLm04D13d7I6LRerBiVF+L5Qf1rxYU5SUohKtDGAYniPI6YjYiFwA4a
WFuGm2ek/QaZ9nlXRLDHOlmt/ymdkc/admEbJFl5p9nSN8vXFuhPpY51VP3EJr0IP71bF6eSAmzV
xOj/0bS9cu0G3xitCVYi1wBECZVBW/RuB/0h5fpN0gyvjlxBslVSz5gi0aj6iArE7OdwUfdUpCZq
KJhDI5Lugo+LUzlMLNuBlOcLPlXF4U8mHSKOGwSKDBqfmzkWoxjBN3XMVDgkDz9OVzvavmqmaeDo
LBClVDRsjdjblCVjXI+owkUR8HE76RKZJBaz2+grvUKwBclc0Vn7eglRxPpZjOq68h6HviZFAbKr
ycxotyOZGbQ/PYsU8gYiH7FFx86Hw3G3R/r0wLifhcamKfwvnfa7KsQMvDmuRnL4noqons7VSKYE
hqu9dqowVFCK0c+acjHm6SMXv34e9k2w709hHuVpia6++KTvCdg1rpUVp4CfmFZZQ5Ea3IPJhn9l
+UjkYlNOrkjyfnr1WqxqPtyXXW9ArmWxiaTMPn/mHRdHw0GR7KDH8v2a/y7uGwUvu/nsGM+fCBXg
u+GoiQHd6+gwQIx1qEbT6T3pMn8xB4xwXQ++My+7i8VA29aTaCdVB1H5k/jjqyD5MQfx5apCTl64
TmWp0DVtR6UgaRc0LOiHdwuOm1iZzxwZLqdeupHKcLL0CEi0jzC1j/M2CG5fVe+XAjvjqhYu3wVu
OX+vplTF7Q8nZJFtajynY3lHBw0f+TEld68E8jLSH0SuJk1hQc9nUtdrmNCFCJJKIOt76zM2M1Q1
SiHP/DGcw2IFggs3L7tyak4rsFp84zuvZ1GPhVm/p1sM1xAY1tT1r0OzrA1KIjO/mI5b476igbVy
gjyflXkRX2EtNveMzogfwPTGJQtDW1QzeEUb7gRfpnMeJ5B0qyX3+q0actx6fKmWDBWyVw1yCWTA
a28N2X8s54cFyWLKaB4p0/d8UkPI9bco/MIrkP6a+lJWboAYlHHm3VrdDpaeFXGUCefNNenQBn6d
kuvlzTimzaF3wXbutDvSI/IRiGaBXR2/A8Wk3oilLATUSay0CJbL2JnK6OCina0ulaRbQxVom/QT
JysS4sBcKjmT1Bxhm6IdwlhnIg6tbimZBGWPNPZMvwPJiVB1NRD8vw6fNtyqlIoBaFJqZFTDr5wM
rxlrikBPbn+IhdslkKfOqaAOWOmHKjmtxwWk39oZdWSVE2maSkgcJ3XTqtcaP4py2ZpRiOy4A2sF
k4YmhM81grVlfFfzQincV8Nhm57ghktyPZ7HyBapnO2cMV1/C9weU4H1GxcwqYhCMGTSnrdVwLrt
Il2dE3bq8SCbstXgnsebYvyDnM0r/RUGsTt+fExfv4Jb3e6xyPRpHlGf0aslxoaRI11iZYgYCjuN
I65wCqcHYV6+Qwgbgg9iF6aKyq11NWwxUz+GfH1rBLyYs6sj9TiwUTpnYxkUzeNg1nNYTl9XgTfQ
K+l1O9IyVWBp/f+DN8fzgyxhmyPBW2LwYdRZRnAi6l89vf85SR/m0PogC5RGLEruQblZNVww5pCg
qv6J20MzuUROs7PwxCnjq5mVrBIYVQrmLlZZQW6uABKMUuzWwCnRSp6ppbQ9uXvzzFKR9oFuMN2R
5lvE4kvcOeQE9p0BtPqxutsrV2jhzoIM2HizK37qQ2/S+P1hkRyfYZ/LKdX5YlT8amVSw8dsfeFS
RKbo/qZmkOFY0JYLt6LdCSH3Q30DbVuBhhwRAD/8D+K5BBTGNNLDoROQz/yTf7yepcV3EtKws1wW
mcY0KOjyeVUD+ITpwqQUCZghISdwZw3CxciMZu6eAftk2bWNVApSVsiW4Eh0WrluXYxqcjydCqeS
5VUyo2JUj/obhWh0a0CU6KRmBcbbhL2zNcj6AZE8QoXsYMCCtqm5dzc9tAZPt+Xta3ikBipb3kiQ
qjECo/HwqiXh0af3AKL+/FUydnCuD8cvhqebm0YKHjTD2uVlGGIyJxZ/UKPomsioKhlkxcD8N29h
3g97RTcCBnsSmjkPGambbAxMr49xU4teAGfRwJBGUfD7vuJeJa0lVnjHequhzHXZvXAjVAdcVrMT
frdh0n4YhO4yvdBT6eJRaaCaaABq0vajKtxcm/nSGs9bPXgtBgLZmIRAH3BNIdFwJzYapX2+UD1Q
JLlMAmDdAEk5mGWCNKt/sY1dRita3mjKD3VKZbvzy0a5HmT93LZ3yxEWCBtoN8enum5QbbGIjayP
8LCvS1UrS3EjhUpgn5PDDDatcV7yKnndcQ7ERuL+7wp1UtW8X6equmWORcMHokhm3yGt7AdfN6SP
KQzSylDcjo4LUhHrdt1MHHZkuSzPRWBsm16M/wRvuHZ/Vp5FOSZ4Du1zg1w0DDOVXUFEvzZWNY2Q
ZiiniiRlS0qlRzmklaf+yeMbJ1dVK5xS/vNfAcNApVA4gvLvmQIrd1Otk/MldPpkCKHKu6oOTlQJ
URY8cFMQvoxwLk2Uj1k7ZMf3/yi1BC60g8O+XBcZ1QcqrNFN/G8bUqw6K5mFcae/PjYTxLhPLhI3
rFNaKmTJw1Il5tBLtDiCCgxs38kZcsBk6GH7ZksCwdiL6UHtA8pZ0YCEPe6w8u8kj213Tf3ebwTu
LAi4G7Yc5yGrBiItgqYh1tYQaVbt3iKEa+mZxIL/2ydaC6v/5sZQMyMl82bTAfs40b+UqVzCCpHq
K8okDhK+pwo7i0YuBB3uRdcuVXRHM7c7ark7iq7EuEh9DSJpGDsLWabK8ThL+b49LS4fsOKYILeR
Z5vU1yasOk8fr55lCIxGwGmKCNF+haPHzb6/xKXxYgYSsfSvH+wCWHtR5GqKiDi5+kLGX1KbgrvL
Oq5Zt1XLEOwzvGZHepEjSI3RNS2J0P79O0OEXQit59Qu+3nRob8/Q57CKq4JKZfudp3nQ61H2XNd
CNCDylVRkhQVJn+J9YbSRcgRc3pWiXcVoNHOklJrzeanWRylZmY/J/NwffIPhifZY9c5U3WZNjrB
VbxNYqSQH3LQyMSekw6d3zgjSB8xJFoXY1Byv0Lq4xPLTQeL7J3xexfUewcOxIaFsKy9A6ulv3pY
7Py9z6HM/EybFWmZj8mmQbuX7kyt/V8hxnzViPkKTYfkZ/A/o2/FOxSg/R2/pkDHTagSoa1C7kXk
rklnWsXhJ1ggmqATk2MLurQbkYDyC8qwUwxPl38OkIvj2U7waof1vCE5Ic3auRzeJrIk1FOPa2Ez
lsX4YOwCt5k0Kg6fEVCuQpJjNAXUSzmvZwhqTCOdaozv9Ny/pdgKT5h5TdQG86PjOL5UMZ8rvNB3
zPX129Hoqv/VWT5+XnpvAVXRmvyEunR0OuVZTdkiuBleNQIwvRdNtNTlmL5cNN/AyP9Z3Mxcg1N5
CacuHpOKek0uDopGvUGI5PHBhcDuIj25wcU/bU9zg+1Yb5faSOV4AfaABKgLinAdOqVsMw4sH8Qj
+pQswYFeP7kIMN0kk3NS8PUPzP4f2aeE55/CwveVNEbf+WCLSCoxxIevt36L+P9mylDVgG/o1xWI
+71iApckDHpZz57u4DQy5nx0PuMP+v/ritLzN6eEAQVZiUaIr33990x+S4ZRLyXntkBUqugYKVxi
zgp27jU3s8ZsyatsZQVoKGi7ywUbb5PvxWqgNeHpZPt8gV/dKTw9lELQPOOz8EO36LNN8wWuEPMB
7da9KrrO4s3E/MmsrAbbmTaPXzFxbLGKY1xRU0CKNvsL9QpopfWUDrpQKJHWpVTnsciGaHdXIRcH
MUQcYWqAU75S+Cd5Cl8suHk2P96z/UFVxm1HiIT21maLy9bBCuCnnzIZelllXvKXnrgX/s2XM6y1
lweeDfHpSZEJbbbSSab19p1NkFFDKCLH4FKh3SlD42nEHSFD+3klRa50H21BsbA1DGdeeMN+XP/E
5EkXdx6bWqc/AjzDoMkhu2rvWNlB+htWW5jK4qACndcTPxD9+HKr3K3HFuI9d1r5hyBPzw4gyPjB
qNa5FIDO/lgzTmNEFn7FE/GnDkP1YfAIsFiYg3AKnGS+TxDAKp39pw8we5vzYqYOBFWmAHmaGwZz
3bYdegv1U8HdjCcgsMTpVETcpxC1gj6aunfNuSVdn5dRQcHql/13FOCiTGLOt8ZQ6fjxLeb02iQw
MCJmrTzQVz5o/sUIZVOZDf3p3e5p/l7hJ7OYolf0F+bxpYTf1HlgN4YGTyt/8tqYqAtpwmqFB2xA
JYzOFVTivhShiHHK7VEf8eJERQ3MXDQcOvPgNAMYp14+SSzDZ1UTWcDY26M79cF6YH7uhyi4+vnF
2nQMfTeZNYSrrQQ3PR8mhVwtSRgJOk+6TFIJ859o6Iqg6wsqJyoOkJ5IGOVEu9nAnHQBs944V2cC
/E36PwhlrpxHtezg9mDJ/REtBV8fBqpXpGaFjrdSYVdrWxHLBbw516XucqL9FEPh8L7+KCljZ2+H
ObKd0ATTUI7X/IJHZkN5yDPXALybzntTi/FExvN3yCJufDVWwTmQub/CK4QVhPVbTHy6rk5YD3NF
ejsKUp3puDeShgc+4gP4E3mrJ2CzNko4tNQMX2k+H/jy6xXFnkraVib4GdoPo0D7qyQmnJMyjj8t
M0UanTDepXMHrdkFW/AD+Nct+eb9PqDda4Y0okYg7vPuF4SovZSZjDqaypNsdNQSgF9Yw14tjx9D
4tEcNzPKAFEuFnRwDHW+sEC96/fG3zTI0MDEZAp+ODL+iqxFlZno0dby75yvOWXiyuMKNRklfDg9
YEQe4KPpNYLAtq40fVOExTfo4sIP1QshwjEz+NYnt8J4Ug+AB2B2jEmnSPONqXdLCp6rt5TfD48i
fzWrNB3G8Iej94nlnWXjiXOjslRAvXG379yY8LzWijAyspMscgU4ZxgKw7DIruIGwidQAyRtarER
jUXNcDM0HwU5/7vgTylcr8zHmRsPYjq5Z7UA2GSzhPl9HuqJrmIZ4ECEbc17ZrDvFoAPNQmlGysw
lt0Wvh6VgQgfx+qNgzcJgg5V+0LjbeLvnrpG239hhMSl72MoWuxUs6Hx4HiZrwJQO+X6V7yh6lFB
i0/ocp4c21zLVyKmyjW0Su8D6bwRbHrhkcygUEMd/AoNm2FjfvyoPrTYAjfNFAGFdxTSGQ7QkMB9
LwYGsLT7eIZxh1BXcmbggVKAYjABDOyifBni9k9G8Q43bO7pf0JjYTqVLI8Sl1emkOiRx95E1AgK
YdQEcbYSCRzfwyfdAXjNIYPPHIVKOQcTm4K2UhAnMQssxkGqg08R5OKLuoKqMQLO6pGusb3aIfDE
efy5hkrI3qnk1nbjhTS9pxkif3MLYoZEuMgDPmkYI4sj6j+aZirtuAV3Mjn5BmPxZ1EFz9jdyEZH
HN1h/GnMjiOVfynxg0drisqnf/pP24hJnPheVW8B62ykhMYce/Pwr5ZE9TPDc8fcXkre3lRC5nIO
dvchxUGoOSQ1Kl/4GhDXL+oKgdHB68lIgWkmOSlK4KyMhCIrzszB4WT0ZPw2AXCuzT5HR69aDWoK
SH5SllGroxn052L0cIs5eDablJfMsA85mFH4JejXoOFbuEE5Wz9a07sVw94XxmX3LSqCgllo5ZMv
gqU7CPIJHYbgx8XOJb0WfjJYyUiT4tb0reONpi+3T8kJG9CcTA5TZBU3ozLxoS/yOyB1GsagJkPA
AVMgdzTanV/SdTn03mrmYI0MS9ByHVAHjro+yv+RKxvE3T+jbSdNSsCnalfqQIU94hZln2+UcUiL
i2uGUTq6zyHcuasSqvsQUwWYbpV8CMcqDiBKrjPwuj30olhFrohYOWHRHFGVESWyatdRsjF5lIEF
whMobWu77BbFVfVJzaiBD51HfXlSPh/T0I8/C6Jp9pk2TtEKKlMX69eVlicPNws0Ny2xrXAjsR/M
y3PIvNeSTUTaXcHFu+7LGJnHDuS0Eo8HlMpLSE5ps0WZdltFG95pmZasyTp7n6bJS32sSXBReGtP
Pb5746UmVRogpmjqgzd59xSJB6a6KKUEYSQMtE8QWWoP4PpZRlGnGDR9oR5Az5dZ7Ge9U0h1Pol6
PMZMR8rcoBXNI6jIzlgPIyC4EWsmr7rhhcb+I8Oc2y9JReYtgirxa4E32e9HqgolJcmvE1QIHTDf
o25C+xjrFzKVADTje3nAjFIxUTeQ+7HmnBCnTlX3n7QZUqlUwk66r4+Wt8qac3KzedEUus9c5zTO
DhhE9c+YbnSWfi5/4krGiLNRghFLJ/8CCSalK21/f6GgnDnA0mbhWpiNE24gYwmViA7ZVEiWEUug
lD7eZdPLT2vU9m+mME+Rbpdq4bcJrhGQufFgCyBoIwpq39geifqpR0+rxxZLnyJblGi/LKWbNGfi
2FvLB9McL6Q0DTYW2fYMh27AwmxF6Is/Io2MfeLKamo94993I2RV2038DrSMuGP+jcs3Z9zTJHmG
Vly830M6LDn4dg4s+LdKzKiO1xu9UIpLHX5XX78SrPEARe9UNQ827TeLlg13/UYn8RVG1z8B0Tmo
EBb55G+dfoklYTaLB8/HGqnlvtJUVESBVqxeEPHZ+RVqOSru7nRcLHDOpyr22j8ol5NgNfvPYPK4
MkNGYYWEfExOUqBX9vyOPdXvoHiXqJSVLmqIpq7nD2B+l97UbAMJy6jTBf9hsB/zF6gfMBkzki4N
0NKcrKaQnz47jgbhrkbiQ8KUQCgJO3cTRUiYRg+r+7bRgtE+xjUcJuo5dKyyM9tEmz72rFx6tPys
mhqM8Pl+bdY2d4MneMUCJzNNSDz8W1hiOP3Q5ZphNLtiV10cdVbhUWkduDwrW5nAqN61kGgwZX4F
xRCjZKZfjJP0kPkp71/qgzdZSfCYgKZEnLI0uSc5YrS6HBX8eC8zsDqRP+n2Nfy3exWgypAzHwNJ
5y2nW5MPZfW/3l8aBXpQX5xf+/rO1Wf+Qx8MyowNyOKmol3Lk8fQ/qQDfW14fbKUzDN4u0YjJxj+
w+zCfg8tiu0jyJZh3b3Q4NeFhvJ8P1+ZIU8TmcmzuTd5JhJk33FSMmbqoEx8+8I6X0Nnw/dWWCI8
ccizOUrOndkQij8Gh5Tis2mt6v8yOu6YtkzVrv9eZ5P03Qvrm4oDh95y46j4aU/fq0XKokVvKfM6
xO+yMFuZeCjFLa2L9SYX6CdTwJkHPQDJi063+s+nwITfV2jQUk5XA2zuMrB4LTAWX5I1AzIbXCNk
H8IFFm1WvTSYfOiJ1uQ5l4IbyfeQOZKMTgMmFsZ4pk0ji7LWGI3r3fesXgZ3tFKxNJtljuo4LPbi
E7KbkOYuAQaPqwlmUpn07Z9NbJfe1A6SGKr4hQOJwrBHtKBDlCHWlR681vEFrSx7UKOYDXOZpfyu
RWdMYFhiOVhnxtCsWm0MjmrcWkcvKjLxyvEqvfIUt25Wh80EzkSzVrOxk6uQqUrcnzXoDNvD6e3x
bNdfk8Y1W7DaSiPwInCbKvPEwltxhW/4zArQwfRuQYLUgwb4ATdGoaqGIvwfpi+cALPuv1mFfQrp
TY/o6u37gYvH6YwyUdcejwhD72WF466/g5dLEg+54zw2arAB2AtKRZG8Fmavm5FXlRMBIzoMZJdy
aNUbQfYgUwssK+A8rNDABdrONsHSWybiw2wD4/rpJIzcOlGCKViksrTfU7aQ0Y2YG9n2yB4Pwqk9
ogdUZ5kq4bq+i+bfD971YEP1tdszimxOHTdAFZbC0rBFF3f0NDQIoCfCct3CU0OyqsNe50pSMlBs
14hUaIMWxrLW5sy5MJvLHystyGm1XvZ37HA+2gv+kb7LEiCjjLPA/ASi6vxMsiWPCinJeIMxa23O
tCcHZ+A/j7k7k6XIVAtXSoUOOVknklQFE75NATyhhpRKHDCp1CSly8ZzinR8PWoeLUxWwID+ReE/
N8/L9mqIjF4iJd7H8nqOenw0nHsTI6xzjYli6/t6suR/ExkhVNE2uxMOmG+5s8L9MoiJlzELY+Zx
vO9vQfiNq/D8jxot4wQTHaQHQ0FAiit4SJRU+dVmy9dtLZjm8+WTqEoQmzy3/3dxC2Zc7VLO1UAF
oasAXIFaddYvUq/ynHWPZ+OweF52KWx6lJ0R4JeGOSmX+izhJQiVaKk4jgc9evljhpQtFkQWqrMI
yPDTDzar+wa6PIY4EvfgVCKK7k+6ROjhn4QfEvEGRZjMCn8vdmKTk/ftUd2ukaKJ76xdVoSQltb6
ffRuppfmV9+NaWGAzTU/iyp0PASOorcCA4KQ0cjTGYcGv/b+YeA7EfDgi7WSnYX7L2LcPqFDG1z7
vjSGBCWtUduoOexrIrfPos7NSiIZvs4GZdNoijIDOUReIWMMyy15M1PdAH4QHRRFPlxAQqVKQtet
/1POQ3Adgs0jASk0s2AnUKGdlShnN9FoBFd4iWK/2sd4UckC/vdhYg4fwsgub27fMOrfOFkxuPlF
6TWfcTJ8+M79v2tSM5lfyAA35e73nBaMmq+gSXt2hv/kUUzGTL507JE6d7bNJeVowkSoRSJDzTWj
YpZodqfHfStB0klts7UcUDOun0hYvmsGYK4/YR0vCcUg5T6id9breDk67aW2wFYavpnc7VACoTT+
WvTwTNa7kiV2NBa4cJXbShspGdjwOBQm2xIrLaP44G9AWnSA5JR0eamh1kh+1Dp9EGXGXaNssU0T
mg3lrPtzP/VTULc/a62DVuLw3kDVC5sVYLmxULPJq1y3rs+LRScHvK4ApaSrwcst3Z9080llk7Fd
9ziPap4LZilGCbWCJLC/dkeSJxYfMBzFm+ZgL3nPZxsybmrKrYvpOIWCR08VAECuqJJHkDkmlGpH
O/MR/KmXB+o//tbMAxKoRJJPQbH6z2QJ6EJIIFrj/hMPa+jeXXyTXdp23nvEPlFsFCLcT2cvUNA8
10/bnnansSkTWl8dC63uiXV/B1rNRc+VolUr6IBaDs9c+71ci1/ZSyX5PbtwLT1C1wLaD+D+tLLS
uQKQ3pqcPQW73YQN1nxrZMKcMY09t4AbEMVcFl7JCEDuqonm9qiqZtsocNHzdnck+2vyFCQ9fkNI
8OV20waYtofCMKq7RsssLwuZohdluTxL5Z0r/EoDofK3P8kQLMy3VKSld9LDjXLr202t8pJHsFMq
D5bP2Zvl0KuW66ouxKeClDLhAX5HaJ2Oi62c0TbV9UUfBMV/iysV5GCjjSGCmKX9sDYv+WOcEiNU
dOQbrvEHxotu/xkCXp5mSPH/Rm/3UT4rkTO3BSRIr3XVqgGeUEe4TMH9dKCWgzQOLS9XGlXVOrcE
1t7w1zdALSwGKLUu0vCL9IGYC3sr7jH6Q2LgBw+rptXQXA8Or2OQ9eU2Xl3eQv5HqQda5spBk7z8
FiIVH04/VUWZhs5x3eaDLLe30ILKysSOqu/lT/HynHTXoJUSbuE8q8r3ZraCvU+v2MADsZidu9yh
sdWCc1RXaCc9sf6skV+7Sbr+2XNTm22VHg4wvkKa3KxaaeMX9w3+8n8b80PRHDC/Op8p1vT/O0Hi
n8z2h5a2w5GCQxuVQVyPpgBaFBkUNGEV1AfJScqexI3l6VeqMLXWm/lO+39eH193K0WSgMvTuzjc
Sit2QsGmb0o9HaA4i3PKkkzI5yFKaOR38oQCwIrOGXA0+LU8ipxPLcGWi0/nBAD1MwRe6F1kFf46
OrpraxqWj9TnkdeY6fAZDdpsPMCKRnvaXwo5lNi6Y6cctwyO6qz3560y2Egpu1AFnpUh1DvBYtNa
VsP2hwbMWD1hLgnP0ceUHF7+x4MAQKYuB5fA7kybDXV8GoXq1rhgXGq78olYeVdXQgGGfgpt4cWH
QGBFVRuBxx5TRhtGQ6xn/u0s07PmWKhz4WNr//cvWiZToh5A5wRKY/DWtLvDka8k4jE3d31F92GC
Q6DrSSp/F0hXORLJw2QuY+Nhl+G1BCMj/5C4ivNhh2uqqQlN9ryWYY7Yyg0R7ku1qwFxOqAvgeXQ
tD5ty/HOQp5tVdTjQYx565PtBANTUriQ3HQkbl2jHM+W2QfBGQyNwST4qNDfe6RzS2gkrAQkE71/
+cRcdKdz6IO9MPPlVSpKOAZGz67sQWjIjrWE0Ym1lXi4oyGgBmHSYf6kjhC3xbsZk9rR+B/3NL7f
4ZQfxYUYw0WGteELKFlLdLbZyMRicu9xzn9NgMwixlpcWiZAZFVPVLyK27YuVMLCNDNmIBiG4aP6
XuTm9jz2qA+FjeeS6FyfXXgYUF/llRBFCazeHEDqN14T82ojYMoUrUmJJG6pyX2VyoDqlLYgOex8
+Pp2sJLgEMs0rHGt+yNpbLW+pacYojiwtRQzLN1lm4h3zQGNLBUC9b9ePTowsh+T86RjOV+3E81V
O4jjztqPZ1/UVeiHkare+oBwoNBgdpA3nmqFUgD++7iVmvlH1FBCByhpxZy5U28ICYzCzH0PJpUb
U5T3+3E8R86rINBvRxXufMCivRPmAkU4mW8/DuF2aDNpzJ35F4+G0U+aJX6jnBU48AsXx4E3R7po
tiuRtTdKaoDmmep2aKluYm/wF3FYcxwDej+Mv2nhUdfdUtBBP4lfKYnY1qBxlWWd2LPiXGUnasbI
1RhKT9QGu93g/eDDT3t++yfMzMXMSosFzAFci+ALKjlqdmBxC7rF7aD4IHKtD4yi4dsvv3RHosyJ
ElzLDjkZc43wbCrgCXI+sDpH8Yp8kMWZECaurhW+PsNwbIKvzScTDXzj9ymGp0pp57EscRE6/3H5
8RegZzpwOuAMJGWNbnDBt3OPJTjesHox8w/psyRt9NpuT1xa4dJnQtPktii97mCoOlXpEpYgTsq+
qZ8mHuOdPV+js0n5c/+4HI7o4L+awgqtS820sz+5uktpz1RihK3hJbLE9Lhq//4LRQX95wzajW36
rXWfeVB2LtkblSXF+SICddoUF6zFY7ZWsXnPbxP4y/IJYgXhJC26veGbgOPMAIldpLPooH9ldZTc
8LPtk0Mahxue/891OYt5bYXquG/wjRbJaO1ND7453VjwLtxokLhuUqb/qfrx/19a2SyRtX3TCwhY
1Oyi789p5IldPHU9ZGtaKEvlAgCfkBXDtprsnbaC0BU4F6Npw4qA41EKS6jVPVABIQe7gsWF1C3/
UDrfj1PiPpSy3mzdJCqRmQ2VGP3JznXy6+hTPXo5GnM03jku2iiTdHjMywXx2Y8BTCsrdBqvevZS
5zzuIATYcrg5Z/wszs2H/9ZesN+EedAe7OkthIfG18YSYAeA1q84NOliaYVXAPIKe5otTpvGCsUf
6gqq2VDRicawujXoKTVtXwuP5G6gJaKOXmW5pIbe+a2x/jRmZSYT8v66M4KaZz3hHo4BeJHsSGP1
deNc5JocT0HQwBdORF/ZPOdUlTaWx9zeiyejXjvTfZELQBwaoXoXFj/cT267ADhMasCy/ywuOgwO
/rbOq9kulifK56cpoD1E2+5fryhp18JoSDX0knmzSK/QW0AQqvoi9e54B13UOLdBUUaeL8fWrz4S
x9yF+8EMDo2f+BuicFUddxIiHsCdUqtNtqBPgMIj/OSR8Pp0S3AMJ1zQle0k6Tin0Ss/GK5+2zXf
JdJADLMf9ZLw9nVGPzfK9o4iOJtiepn6Bgv4v6gshk/PeamV7nXdnx1PUZvj9EBpKARSezNlPr1i
aTBCvT1HcAotE3rqOlDc2hWjgIA+ZI2G51soQMFu0qCMXA4uCgssvnLs+K494+O9sQLrlvpNHKFF
ISWSOFkUxQtYUGuB4yxvR1LgKFacJkpuZOIDHTtMB4/qnkKv1wFHIe636w/Y/7KqDMewjR+LN4zg
XQep/zpsE5P+Xpsgg8FhXl4ViRw/dCNpfYyZvfCoAnR6Tbn5w6CvoRTc+KU9cwZA5u5nXpyRm2ZT
t13GecpXGdJ6PgVKJcD2oVEoyWHWCyBx1EkENUpy+TahVyyKDjsoTazUoRMlMsmI1luTfxI3k82i
AfvbihVKY5EyWtES+fBQggbHD6o4yJgMKJQGxiDQ4AIrh8lNAEPkTe3/XcCS+JAjHV4mLbodMD3t
XnHH3V59DIwGZt5OzaKDfwxWBTW8en7IulRhJagVxxFJZ8E9bultPT8+ZIGpBXyUZjvRjLtkFWVR
T/oiA15IBm036SN4T6hx4Li560MsSeXn2GPLHHcBEv6NPZJenHYoZ2D3mf1pwIyFHVk30XmvGppz
iXd+eLqtyVSk4PeaoqoQ0Bb4tFC+iuYyKvp4MW1Prd6cXzzWGqjmsmeVXVMCNlq2EXh53eWUuHBE
gKc4w3RRAwuHtASOlkCUrOtSzwiwwcozVLykk0xdjvPkyaF+wiNyeH8kJ+55SVc4wJ//GyydExFB
DdpNijnZDaoV24u7OgYuD/f6YCYF5EluW7D+2+KYM0yGJ9UswlDrCo+3qyJygmnXR2z+AT7KzEs9
O8NC3rn+a2OhtmZE2Bx9IPv/Gx5dGq/TMaNsrTM/h8rsbcfpXpIqAawQaPVVxdzI9DFqceNrtciQ
0gJuu7579uM+tBKnn1IA5VNsanBflruc4goQf+Rk/2H55vbSvDLqby6ehGWp8ifJuipyFdH3KrX6
6dF88NaLyrDff4fl8OOdBmrwh/U4Ryh8yKm4jo6DloG9QMhnfUcYTYOzNa3q4szysiGD4gPmwrsF
bxdcnLRMEfIynIOvoZ4SIWl3NZHJMjcXLOeXs/KRHwNAAnlBBN/A0lu1zaWUFzCYU5Gr+ue3J3Di
OPnBZlmbArymENLjUrtNKAHGFkBdH6mo/8xpKbvn8ixXe+RlVhdE9HVn2RJqJJzzcxMFxe9BBO4i
l5YLp0LnWN3iAb8uzvBjcsgtLyip2WCjoeR/FhY6yX/IpJFzzd0sHl9glaHp3xl7Y83ZsERdMtfi
o9haE0JFL+tDrg5vT+JZGIRygEM/dkbAKSYaHNGk7w3R+NXRS+gX1VTEqj0Jry67bq3nxgGkfPBK
GROKwoghL841iTsOA2ksv6j0psREZAq/IDwuxeCVpeyjF6mWw2KOlEz7eUzM52GfE2Oxd4LCYjxw
8kVkPRLDlH8VavFUCW0GorpLI6LUs7rLfvMLTSFSHtWPBdSoBdlszhHNagq1BtTxMbwJfoCr2idO
EnU/fhd+OHzL9mROs3+fMTNWdTqst1GMDMWTox0wrv862CW+eYbvTEwNl3l/j8kHWfHqtpC0GPi5
cXEpF0G0kbOpcMEAVErkWa0Qxd3y79E+eqcAViwhQXIAcscXulcO+zHxivF1Ve6QF86BzuP3PIhN
YsBbYkpmPLAK7mhHC3G3i1zst8XpPMAKAKYe2679mmvnEztKi2GETGpmQUpoG/huMu4qWrwKQ/DV
4rBhB4VSQz9T7yZkGxLqCemEv2J2L7CPHjVZCgmkZ8lpFA2OI6nXra9tZF3iXAHVrd+CelvteI+B
i7syLDEIk80fFluuGnsLGrL9Z1DedgjqXAIymti2oKopKLeXpCjz5gcy7zAV4abobjw2bKCPygoP
MYBmD7rQbiH6mXocEyKsRAJd67GwD4wbKsjGAjaN3CTeHof3SaAbWOe60WlssLn/PPZZzqyA3XsT
HCKUfbPtJU7fwiLNQBB+CGoopprgrfoJeir4G4dJNWqQqnkMG0U1dGXh7jBdXob5/+2FtB3uaiw/
c+dTCCJUW9+xp1wTnRXeg343JZHRJG+P6oiR9mHVDr/zwHyKNXrC2uRNSDROxyTZq/tkKEXKkzMK
6KzHl+7mhlJNeFREM0HCt14DZAmvSFlUlx4nSiqkb9hHYrm4zertWn53DV35J5Kfv/an2XnfWRWi
mEddazm2mPldQwIfj+K0+N3daAHuxwLsnEJzTdsJzzG3GAs7fjr3CaLFZ1P+vglE6BR4RVvMWqWx
4T21H76QggqY+pVVbQ/qT205kN3clwVC5xrbbFuO2mqtvk3EF/9dvvRdjtZ59YROirsMzIcOjgfI
s8yWpHR4/jrRXmojKnkvXMo6L4DtsEODKGDd3RR7fiwJYbFu5o9U9lyPB7Zrl+P4TgAJ4VauxWMD
Mx7QxGAJFtJxQqxc7nr3L7ghHFxU6cxBeK71jbwOsbp643f+VnEKao0+2VzyoaFr+RGg6xKQGAgb
qu/kp/SpN1KwGqaEJJazB1N/2vK/+EMUrqVMbkcf+IDxcglHZidKV2axInFqnGmspGaBRdXGxHjC
R6H9Qa/Xxvhf+Sh63wAVXhWcJNc259UNIfB5teZZfai/PrkqWcC+joxmjtdaJj1GbyS5Yw0RP3XQ
d2J8MYhrYZ0L8Gd+zo1ZoeQjbkOuez/sSIkIBksAiMZ65RVI4UcIZn0xawlGsXQk+xiAbBeNP/ig
7F3zD4zkD9rWg5GXLePtopZXwXGGvzrnDPn1bZ8aTO70aIiDQCWPILBr3Y21Oo3bgqzcu9ioh2p7
01A48bnOxvY2n03mhUxGE1/rDPtsps38RHInfurIYXnEWzJmdyeFmwdFiDcOsrF8VTZOqruYFbc8
Rz1kzjkOt6MWFNI3aROpFwTHcC3kdeQi0rp2mSr2wFIclc6iiSn9oGqujLGGsZnbVKgRK596nA7N
arfOGbaSM851ZkTSncJNmN3W7ol50eFmZAp782tiVymASlngzYf/6gRcqyKVmMClmcLb3QuA48g0
tzAxYuVIsQiNBtUHbySE2513GmDJuEBSbioetnhgjNc2xroS+suPTkqNx5/jawy3eofXuLP/pDVB
2u+FCmc2r4TT3ytp+EPvEJe/UNA5746UEWJVQ94hwFfqttPFYRkVtciQpLaSsWni9JNZF/rxEVXX
cvucKOwfblHVYaZZ4i+0z14W5iSUxKEB27YsJCDskWLFu3y5Ze3S3WS+n5KC8K9v+B7DIILMHwkU
ThuhE1hitF5TVdemajkQ6yFOJHvQBVDIy3OPrhmRgQ7h21bm9NIbRqgCb0Yf57pEzoS1cPGUKAbh
7qFLZijrpHlBQ+Z1ca1fqTeFw742rkSH9SggcAXdjsUaMFtNrWHr+UlxYz3oVkKaWRSXq4RBaHtx
fs0nCrxeVxBK32oXFeAoh9nAai9DrQ+ngW8ZbNnUPb/BLFosORZL1rHk2WZF1nfCFF2K/3nFeYk6
y7zRDLFHL8c8xus7ZNMyG3gQlRAlX4pbnLwvca1nAfMQpm2xvMVoQLuuXcvog5PebVNYbCB1I8uW
2lxvudZasvRQ+0Dwg7rYXkBgX55WwIxMMz5/B98pOPcJE1ONImRo7vCJva8JQ7bdqB+A47BfKGPJ
vI+gKre4d9dwiKnhjRfst6/NCfHR2x1icO3M7oE1+1oCaCc0O9uuOYN1H6s5NjKcI9VFIsYho1mr
4YAFcU2yrkuU49WFCZPZQ3qW6jsATPgfjTuL9R8mqLLXW3pc3dZJLCma+eo5HEr/hpJs6afcOnF9
GaA9ECNqj7XlRGUFZCa/3IVnFYMNIQyBuTZroLjqUgreQky0PMYEBownUnQ1ti+WP/b7EqP3ryx6
s7m5kgTwjsmhA6FgfKrSUTXprxdc21MrHvC3xbwfTQQ/3vTA15r88faT0yLkG6dRs9of3WkWI6sq
6bG0I6GVYnPvdDMOYPXDHznksJrC3PCp4f1gv6q70mPNff5dsSQXXLq/9PLhiREcBexJVVszpKlI
oM0R+fsyalzB+JaJdMcr7M97PM9GAD/Ru93NdkYAJawaNGJWYWJxikaC8mXtRyecdYd2gRRjaRpt
do7f4wio1Fqw/B+rbmwJASGc3b/EuEvoBWM1wji+TanvxmM1mqTkEDXkcG3Va+X5mfnm0Qvmraes
Ss0KfquSxiPr1AwyJaWrSykQPYu188rM//eQkEJRsLJIWl5//6KqgNf+gLxsaexUhHW8kAkNZJOl
S0wVushBH+5mFvA1pFtiMDdLHtwztJ4J1L8U/eMzJGkP+UFbGE+eNDhmzzkCyzvs4EyCtuExiJBq
Yy+3CbkdvOoEfCJtXoh1be9ExqGfzIdy9Bx5YPLJ3SEPBA1/1vRTx7ewnlKqidxR8jLOV4sCXmD/
vp395d+A43cSEaGpbBsgsKRPbWMbjhLjyqT/3kzyN/KvnETKyeinCanqNO9blpMO/Hc/UAms5x5f
IbqlqXrlxXyej7YrPwTSwNnmBwdd0/ifd6uknH/ToVDBLS8FR7Dd5Ob5FDa9VOzipH+Zu+4HvgA8
CoxfXn0aq8dIcO1eJ32vbUbzDlsIuBW5fwqYEn1bMfvbipQK9Lhq6LWmmOI3NwdYHM5+HBTA8/Ui
hAk3Bo0/hIvQn94fPZNpB1cvMkjPyLdwiLj8qEdFZ8yJkau9ATfXqOANg5AerbKu8nUDYQ9Dowdv
E5qiKkM8bb1di36F1UHgEm7rEAy+4hNIyWYnvGdWkq0egugON7RUdV4cklvxdeuv7Z1yVAsoguIz
dlS6yA084WEMGJTdlHnNtbF8vnpx1MvfHECpMH2eyWiBC9d5wdtr4AHj23exZm+4XJQwfiDIeKtO
yfVDIAytuYuKS4Flsnewx4hWBb9IKEFAdNNzwmax4Gzh9N31mrtHGtYONqfWch3+BWRfJ7CIWbxa
QLSrMIHSfRiOpBnl9pFOq/RELZll7ha9C47wbbFSd2IyoJG9jY1JSZhyve7vqlYhN/TS/4yrXf4Z
MzQKjpW7/j0nB5aJ24TBik+GzaawP/XXGxp6F27GucSIcnw87IBIjn6s+SFJ3pIkix2sEi6tFEvd
G1iCXLRw/j8W3h0EyWWJYlRowS5z3JC1PN5zW0EKb5D169pX8DuDAkFlPUbBVnMlv+SriXRMrfqW
SLZ9f4Cbk4gG9kUbNL/5ZJUJNU7eIPfreJdkiok4Nbzf4ejDcQ9n3YlDxg50EEWeMZERocq4yoe0
0+h7SwvoZu1YcQEOjOcpF1kyG0MIhb5mHCFgoKT/1ecllQV1hjxCscHp83ArcaDrRK0oFmKPPMfn
+ppMYxHDooBWgO6+Mr3ssWku9z7z1qpeoUwyt1pcSf0pDnM7DrCc7Q9Thtws0hbgtZZdTXvzreZw
H4/VKM+FkhM8h7s3OPdmQpKpgmpD6jEYLnyo7QOv9FLWhiTH1aSAv9Y6lbVU2YaH/qRQeDbEcu3U
orYBT1U5UBIvLc6zpBTmoxG53ohLQh0E2ZJ+IK1cFeYnn2rWsWgaapF+0l0WnoktSlMm1UjmQoXK
3Jz20KB4i+2MZYzPHVgnTkE7wiw1c/Az7MwgA2Hmp6BFu5OX5NqIVdcG6fmvOBJ01PpA0k+PSm+R
klj9B8nBW5MsDb5ndIUDpNbnM4bZxjo75HJhHTvty1Iltn5eNILmR5/Y30ejJ2zs4yDbKRYshwVJ
dytU+LJ8Rr9ZK7NG8B6J+Y9VecJ44roqFyVbibqMTkSfbMjVG050+XNS1ZTZP3/A0MVAvvMXtYHN
ui2ErgWq6JW6le2veXD5tkz9TVt6JIN4RFJg/6tE3OPrXQhEWGmQZEKFhPojKoNL1u6V/PwfQBAj
0vibWTPddZ0X/nRKsT3Tk1zXzLLlnkLnsY0X9I5Xst0YaQ3mkTmX5GLKRYoDlG68xmLPTPVVIgQg
6wVeaytpyxG8vXA6X/FAs8rLMg7noaCp1lnZWnvZ6StgWBkRbruKVhLfcOEvKt0zwqPAhmQR0geN
a366PtzIlkzEHrBZWdQPIDSrp/AVAoh8L0F+MEnJZ5QoDyrf3QdmjIj8hdMK5BRz0yiEUSbY0oRD
Jx86Zxda5SbcHlBzXIptFzDK3f+3p89bnWtliK0qeCte6x5Td3f6sQr5JODHE7xJs9l2XkboGo6u
gXMHWg5HxnwkJHPIvTrMIRQYW9bKcWXOowhHbVqgmn0oZKj1HO1qs67z5cP2QNkEGriVmiPPLJWw
unTlJ43hffiyZvNBBbSTDCUrpJ2ELDN1Hp03ydR/x/Yn1f2Jc+bhNByaOq1zXsgvSfFKnQGZ1c0n
ZtKKsKZlE6GM3AlMJLY9wGL61F3REwRkmYlBrOyZ0RII64WYQDVmwjKygS1KUrU83W+zCsBLrF0G
vEubFl89hVk46uBp9p/nTLPS2c9/S4L5QNTRwgV33gO/7YCZxJUNQgKCMjz3S6cgCOAa1BuDDCYX
8BYMuYfFsH/48yZl7VMk3nySFWdh8dZ3StQHJOtGGsD3UzAI7FuXqh2zqEdnqpqL+8CKe9evZKjT
QxapiUv1vSf8nUmGPvqX86KQdlkLj9gJydrQfaXYwc76G95jQno5Utls47ZYdHnlpW+ML5OoET1j
UrR1+77R99g2H80OzQsu/ZGKHgg3w8uwea8j3DIsPaHUCdZ2ULrSfSrbT6MaK8eqToHXV+zGpqlF
AjO4K6fenO2qv5VF+1eLy1g0OYQIIyVP4xLL4gO5YNBIHfuSfccSB1wWtIUx0Hos+T5Kdk6hpJoE
QRyRPLJaYu7h3G/nubqA12lT7Rj+9pLkgtYmHJvwPFHUEEGC+GLuT2/bnm+SF01fRRAqGmJfGZNh
UDMlqkIdoMxbvCzNhjGuvaiB/Ri8Z3ppap0HXZH1HXXpYSrXTvukWVPXREBSs/xzgbWKhQYs4Fkx
Ac0SRTBf59I7mm4HU9NJQMT6CgYdAX39SyXte8Mr/w9mXnYMWZFXMlbRGjXNfiC+3+Z92BGXcqEv
kI2WwC8Wh2LAIyLWhUQVBxgiGNDQHrtnf4ny+IB2DSxkl31uHDGWOniS8D7zedMGN1WDE5zyBlI2
2+HpPs5Y+GIhIvUmVz9/8DX6LMFAC7eYIR5QHOVYKy8O2ou7a4iPQ8CIteRBWy5HQHGWTYeJeR5a
Ck4X69lFjn7ISKDzEDeo3Rl10OJASZC6Vft/OCwxJrLiPl5mBWzTtZlVWhELyIR9ZiMTlpS/CAcv
p3mCjErj05pJ4dbwMsfZiDdh1t2RI/aN8cImmjWEKRxKBdlSqNIk4wW9MPphgc9U9+QWK8jS04Lb
1qTruyOUaqQrXAx1PYobCaZxjLVn0U2+gPZThtij1A8pUALZfCxOASRNY9lawvteilzbRm4YbVco
VY9UT4WRbEHc1/fxO1xKniivC+BiawIqcTeUVuFWnBQjoU1Q+mhhoB8HG/QPP4BkvgotWBPdrxaX
CY7i5JOEqIWIdZpAYv1tDpjYhYaN7TjlLLx3Pdzbj6nNxC1qv/6FEFK/913UY37pyVCNMMwmb0A+
SzLlVQkT0uGxFrof7st+2kHteP7BY46fyQsfaXSYZn8g1RSjDM8tQ5D5CxbQzdvk0YqlwSMV3D/F
rLvQw6OAw/7nIRodxHV72P2gsJuAzvEwwEz66W9rmOJLaBdOG7q150LEuZIhJt8C03+vG/mn1EFh
3Q6mzdD8jF4FDxFOqxSt1DyykP9dmFmB9mpk+uuhTDIE2TKwEBEuAgcVXb0ciYjTDfsPPsTLj7om
vkZUXCw5dodG67Ft1IaHsNHfVKkXx2LQLQU+lTy/o3yAlNwWgX6sqjaxUS8lLXgYoXn0FKBAMIw3
StrBrSFjKKRNXbOrMlddWYuj4QBHg5UWo+zUcxCG3/1AcafHAX0Y9+lis7mM7io3US0Doe3D8h8d
GTD/cUkXJHi0N7ZXhISnDhX2CthyUlkMzfcrAIlbRtLQgEw0/nU/tVIaVieXxJHJcpFQwFvFdfTw
tYenHmPpEgRu0voAbbw+OVpaoQWFnw9XVPpPhf1xyCsiOEUFuaOVlaqjg4bozDwvHyctn+zU3BBL
aUd0RNvEOOAMlI8Mg/IATCm4jiqoG4KZZoA8BEKoGYKDNd13Qndx9s0OcAQsggJ8VABmGQukMeG+
WKadjRig3qM/0Ttjyn8RnupyLpd8JltEsWtg3T1MjwheCg1FjClJxKfgg6jCSbnEncuEluVk9gxM
BsnR00nQUL4JEKxdO0tPWV8csrOCBL9KNvIBBkFjSFr287IqOLKQzp2J8GIOLsyUXk0z49UmNs86
Wvr8ZTLh5UbvrzF3FaCQMFrMp0aP80QqXXz+k6u2Eysl9QGc3OOCHva5yp7qsV+iN91axWm/jTdz
L3TTH5HoeBP9ke/AgXDvzw03/HxqbpDhq6hIYYyVMdKhoPXftI1JZtOgcjkdDIPiPYBOs8i6zfDQ
xRzQ1YCuCHaMv1Js3++QcDZ5lWAD9Y+RLEAmTLfusV5Z69s8SjkqPSaCDM2dQf28e8vpaTVg6VzW
nkkExhhNqweH9IivimDBdoGy47WeXP8c+qQUxKI1MX7OaWMiyY0S8ZmM8E3VTla/pirPGGkYQ2zq
BvfRGRRVFhq+O56fIg08S/qTLroPdYCq6Jfgj2ZOCyBnAQ3xfNyR7U3QgiKVSr/eERocJ7TgL00o
+LfVXRagPFx0qd//l8+sGhQ7d0sWma+3VQ/VueGd7NSuJE9DhQV7HIiBY45DyQHR1nCizwZz9h4t
V2BcF4Q2f2ZDQH94PVg5dVE9PoCCxZVG3JUNDUtaDK4jZsNyC8HimzhkHtb/9X3ZCv2kfu66QCIR
m0AuzCWAqWKwcF98wuHHXXKLGv7QqC4lPZw9VnE1dBEyuulQ1+z/maHsPociOixza5a/jb9nKULo
EBjfISfENOBBVHUWnWhXXk1isSzzQRJDaWBLAnyYka6c7c+4Lvgor8LXdHSofPRezGrUaHUitTek
ZII4WDnt80joZC2TQ93n8r5XA1tl+a3JlO9RxudHLcBgFtaMyTRtD/muMaDacTfJGTbfSZpInWgk
nW8iomXhOG3S5HRZgIDsIgxOIydcz/XuOQaJSHQv6dvMkKG5Tgm6RvMYyxvPiiYBlNg7uFCE38cR
US8zdZ2QJ9NXnNPAJQiksnCETVZTmutiPFq8LoZbWlHwnd47Outr08pjor6tyCMffLMxuNv51ivM
+XWUXYYaCJfdbTCHsTsRUzSeYypEhWESF0sPCRYEVu45cgOfeIdiUIzt68E4Bxpv5k1nQ8XaltaG
eEJwn6c88jdJLcUqAPUBVrNHny/3tDxRW4VP04zZX+RpRj8fQggRRgNAgWxckK4Dzo3R300yOIg8
eA9KuuOB34c2DvKCcRthlZVXaOTKuFiWegqheO+wKqcWLHWocbT5MupFT7lhWQldHRWTSUu/1wZA
Jb2pVjtS7CiSTa7gNz0K03FfEMVMHYZqQ3N77mye0dP/s1BNWQvOwnPv37qJvQRiegE4PRqhjObp
yMYGmjBlUTanBnD6qgyr/KllhPSozVsA7qL0L/dR7bYf3P2MC12jsLS5JnqjDQZrabC1SQCUnBGC
Wdgm7UM8AAAM6X9A3KsvuQiRaAoV8jSXP2zI+jiCJTi8mRZj3ZtPM5nRpyUnPlllXU7PwmkNpash
JfthW+hBCaKdYA6q/1drvYZlqZ4Zbb41vsuOWnNeNaomoJJcAuQ0ehZnf9Q9/Fh0VMJb/StkHnoh
fhlpa6h57fPsIuUhvR9u/if45ZvTd6wO1XP0rNZV2plzUvOLhXdh8lMUYnPkiEpi/RUy0WYcLtI8
u46AHidAZ0PvF/tNwbX5AIzBU8A5kuNUjfZs5294v6v0ILiqa42/4bFU1klzw+/J79/3MRagHh5z
RlV0kOOD8y0dZYASiCeBFdejbcNZQQZRs7biPs8fKkVrHO6Q1TSoHtbZBZVAQAWgUe64l0IhsTMD
40uXg2mqOvmAagaTa8Hu2NMkZAwICIZSd7MPxltYUqEfe4HVYmOz/8uEctWPIvq2OGUt42bdb16U
SbCRyXE2NK2zac4sP4UaogBEll9dWc7BaM4izMSYU+9NTk6ZpNt482KU/G7juA9fTVXC3cWEa3yo
l4bejJOJkYLwr2O5YDtIj9PVkxLwU/Y73f3HVKrPXOAy4Rd8kj3c9F+wnUUrsRf6L5QITQsRAtey
dfwVXxpbvVz61QfeCDE51x+Hs7Va5GGk8tW5eKean2NG/PJd1dF1epoWOxv2+jsuOEAd36QiujO3
mU2hZBT7DZnyExxOEE61OtUvhTb0X0uvNZFGQKUe71o1jJXbxrzYSXp4mUKRDNAmeXGM1GFyDa7k
1L/vjNVeC5ECb0e8dXsQ+woZPyVbvWXD9Z1PqheyIUZA+IN/r6xpraNjTXyUWiI4Pll6d5gBZX7w
JuOqZ6j5A50vvC8fofgR8rsd5NQgcULfv0x1DBEegqO2Wn5N8SDJGHmXYAiFsGoPVuMyxJzxmRgb
JsIaE7dm1UtiBeMdBpHxlqJHbdg/t4MLTVGNJid4lGon67K6qSPk3Xgj8elYmxbg7+MDzT1Nc7sq
/hCL7DiaHmbQ4UmtxBKIJTmIov+1pNKmLmNF7sPP+tRDBX6XYXsgw2+VW8fIrgXRA628FnelA9Cr
3dP8kOTQ3IokCYsFA5zBRkQsUa+4F2TKHJpJ5ylz1ZqztQpQI7uZFvQHwYPpLJ4H2d0Ou8P35U0S
LD7AznbmvMKs93DEmPsBQtDYoW+sHEhFz8tgp0JVUFhu11QeNrMr2XYbVG2SgbT1yo/+PrlmNlH0
kxAwcyOHFC3rMdIoCvbCvUjAThkD6p3GJIsGq7BTqkORf6EVvZS/sYFUXltf1+ey8OQoV9HPUmD4
9g6/Zfh98ZFQzGtTes4HUZSitDZLWgnocfKCWqgKYnUgYChWY4eMWBi6MsrC5a1boMcvxUo3gZ2J
kcj8WDPmACeTQ146g4XlWsIWwyav5S9G2MgP3H45dneJlBJd9jE8yhMG1bFVCiuJ/iZZUy3+fx/6
GQ4KXFE/B2BxpVOT2xqsY80lahWQJUulxXpnRjP2Ekr8i2KVvHA3PMTj7ZCPndMOQZCAvcHgdwfI
2K2Li6/BZQRZf5TufiFLchposlcQShCi61yFNwA+v7CIbJ76AtQtIsT99xYDpC2iaS8P6Bc1mXxG
aB3OoyljWxKUmMIQTpS2SUYz2W/0js/hsiCuEQipx8Zl1UBJ7+NLtdqhuzh8+6Zq17ErrDuIXkJN
MGR00ZQxyJliQ+y2V/224AoHt01sxQRCgTayXPDTGtecHIdZtiCbdw5P4JkbCUYoEgpFgpTBOaQd
rhkfTZ6A6La5+sHgOwXhT7x/sjatDSb2Umx6GLV+oVMm30gesC/X04g4uNUfPCp3msRhahEyMc5G
O6cFxswDxH/l0GwLsxAkUTwT4URFT1YSYHT2rd79ePMXkrxJfa7tZSLdfCRNz/XjcqtNSrQhy24H
5fyYuK/m6+thAjHQGo+WRq+GFHM2Tf0Fq+WM8l4jDHmG1KidwPYJByP0a/A/df21peOndFgI7Mjo
0tpOM0LSU/5ZCb0Fy0HnzGmYCweCBkKBrcgsrvbmrBy/bMMgeDWI5ohCEW67xW4OynbQwPY//89C
ZLo0EsnMBXlxARRlUpQk97+fECze1uqGOUH9/T1LFS6SxRg09KecepbCbkn6xEufJXA1dkoNn2u2
rRCLVBi7O2EgUSY70BxKrTvVKhX6zr6vBHahcDa82AUAAeED8I5Y4Ff2Yg6vdgYC8Uo33Df6FuRE
PudlkD7K1QmR4y6VCrbmu5ZceOEBBcJ2WmnUwviGE/3Q07FbAuM/P7VIe0BDP8y8ix4el9ujchz7
BYylBGC321SyZ6SW/EqurZYX1/inqJ/5dzCm1V1439pkCU50SdbiankmMtJWnb0U5W6Hei4Yez8z
5XqpQCLenCAQldGSEBKABlmlZEwSjgeKDxGu7GUOCMKfa+E3hsJshTQs3M4G0oMPJeAVmPxzTZgD
hHGbp+/znPRaWnxqJzJtVYx/OS/9imfW6RiQPhKJtJbr9lhrEHV+WWbZM/xPnfUamI+LuyOyKBfc
8NW6tzTzrvtGsHGJDforSp0BInrS+BDo5CpHSivbfWb3FEgFpadphkNkUgqt9ARb1p5C+dP/XIu5
oZgcnZMxCYnx6l50VF1kScelMzxrbdd+MlcwTP3J855Ny9LADUGHIdHoHUZLFJHJ1z19B6TWRljT
RbK6uzlHbAf4rBm4a4B3M/HWPncLfIefJuKG7wcj3QfPtzbafDt/RI7k7YdNqVtibxfT1rE0A0kC
wvFb6ZNSBvEkuLUxGdyVzYZ2i5BGB2MrtR0SQujebrNCD9j+NrkysPHSUnQGOepguQp1XdvDJNH4
ZhuBFcO2l+VZHrM00rc9Q0dLXkuCUsDeNyoUiWXqoNkYMO6eXsudw8grAydcIQ37XFgxWfz119PI
/l/fzdpVUkCH/6NbHtWju0SO25EDC8rCKYiiM33+PaLqq8GGX3+S6UZ1Ss2tcmEXJA4qY/oqpNQC
sGHZwJ9JoHmz7ZsidNTKWiirdT2Zk4kMXEhuUroP2qX21jvKaaltRQBTxT72p8EqcjR5z8VzDdP9
XXKWHi14jC6z/RoqJDJ+sl3mSDn5lSuBpXgRgrmXklzOmhfn2W4gHNIkyduqFZqpTs8Tz7xPxRzf
9L57KJfFMD0o+BGK/hDO7n4R2sCqTExPmYzRaf2KjKchpY+UZ+yU26owUKoh0s2u9e5E4B8DejYY
HD41zQ2nxlWdQ9UJVnaUH0k5+Ay/iIloLduIMxuL+snG1OMeLRzsLDIKytnesAbf4gYyLPvVvLVl
WMVUz1A25nEDg84pyDypDKaPk/xb/CkQKT2y+REUhz1NZZVDmS5BTDbAD753R0giU5QhuwMfTHCs
PN3/n7FBEyI5nNy+2EFecOTABDRg/VwwnCm3SljRinIluYgot6URZMGiyHLMehmWHblkhovToHJE
QUOFlzVufUviXgWJckRzVsuwTYMPVL7Zww0swZ++CtusGuUnH7+Ixj0r7UP6lnjCzTkf+/z2McJ9
qFJeB0tZpBlFfS7Lh15WE34G/DMNT2moZRGsEWRNDEGxWkuHroKRmHgjii4kTAQ44uSo/xKiW8ic
kHMatk4n8K/jVt+1pLXaN7EJTTwFPhXQ+gzZGa/dZ+xY6SvND1JAoILpd68ag16ExAs437JPnuyh
eGXWmuyCuPNZ3LPqdrWr57aDwC5nrSz1YXb1Pj2vNGsrIf/kTsAW6ZbieWkr0dnyHUNschf5Z5BJ
vI9bgjo9VKBLlGVT1c49dk1dZ3+j8DY8dTnBuXRlt23boMV6M6i2J/n8S3rkyo4pF0r+NuDB8V8j
h7sNS50858o0IX3ei89WDYvfaKgxA+rDYWpn1j2X1g8QVGFKqHspCndcPxshURvk3VNqvE5Q7xEX
oj8H4q3ttzHS+a+NsebLmipTAJ8bCcaHYEPX0S82hh5Tir2Oq+CILeOdkRKhkk4q9fFz2dz2iDc5
K4tlu32FAHGGne4z1/Wdzj/mUfGlUumk03rKZQR8aJSHeDxuQ/9Jbb/3Aswg/gX9/5ZcMxtByA2e
XUqmHDLhApaWxgneQIdbU1V//rtOe/9VgQIZ37gCckkOpXba7c5iCiOPtB/sg8+9eo5huJiOv3rY
0Jmg3ISjGA4/dUVoRdJ6/Sn2KVRAUuCEDGB2SuGLjpv54xLJu5ih3Cg8YrKWaY1Pb3r3MVs1yYBP
Ojq6qkUCBxRYRSG+E8Hz+VxbaOzo2/SpcMAvzoblGRlpElAayGN0aAtGPbmtZUKmCRbYy1CJkfIq
DNxQUEx2RDt413ZnlfYGBWOBehV34wtgSu7Wfh1gSTfmaBqmPiq8q0lwMzkQradkCzmUOqLh8fQl
Nq7oMNebxlsq6O9SQ/qJxblLJtCYUuZqBqr/OZDTmOJflddDQTGynO0+/FVu+e4zDGAZPcVNI1Xa
N9heHzd4JA7m270r+wQPcvucUG7o0jMDeZR+qmau/v2p/pcN5ADV1+xjk7XUJumQbDYqC6m4ICLO
39/bOHldeT3/4/irzMkF6kZZA/8Crj9r8xGqBuihWorMLDGTJSFKxiLbDupxOFGguCTr3gQWs1SY
uCaJj9KzQS90l9nk0gIOCZ2STHhJpHwAhoBQd5EhkLQWtbJo050GMau8pvdnbYNdLwCHEdg++xp1
r9RmFvIU1FNoPlwo034wfV7yg2HIAP6BI6YgQIjLIDpXVo3ixcdAr0WFlJbZfZ0PnIUWNaxUVfLk
DxO3OTKNf049knSucijEh5u59yGwrLLiHGkFvV8fW9ltidg1vg14fYQ9GPTDWZMtSRKrhFlwCiWB
Si+QATn4OcIOgprlKuTE5PRjrMM8KjcCzFTL2nwUj2TCTAT07NHEKIKnl3P3l/A10bTowWZc34Uv
cWVrcqt8ogq5jWGXEjXM86VD1STyGiV7cYI28VmKIukAottWYGboHqh0rUJXH1NAi5PhvzgHlazo
ew1SQC7t3JG8s/CoEs8LmXKHeKjmDb3r3cddCQfrDwXQgrI6v+YAQQrvci9QjuSyOdFh7IeDJCk1
20X2qiRxo6kxe1yQgtcU/FLvc9MK8RtmGvBc6mt0qpYA6p1MZdKCpb2P/YkUPM/DOoL1jKk5UwzR
8Rh4iyOoFNc3kDUTm9DIrYBKsEl3w3oIg1jgz0tB77ODSBB0aAwn8ngwHB+F2A/Su7dVvLp0ulpV
0+VUj1566S6zD4rscRp79FLIdOV6po2hsGV4v83kr71NMOzm+VtyfDgfYkVjlGbFBJ+Ci7M1QomT
XmJk7ugm8oXxJw118STWjngZwyBPL+WTjC7Sl9n92TNeNGxzXqKsXe+2ItfdMpUqkA/2nSnEwujm
C5dlf+e/za7C6ZQo2gOeTbgz8ydg3zcZAhaO/ehZhk1RrccahhUg5CDfk1J8NBWZd4GS+tmOByNv
xU0y4bVW4Ch9e59vKL9lW/+3sgo3RW20g4yTPfSwuMX8THf0ELEExJTUgNMg6aVveRDamiaXJcYt
2gh1hjtTeMmYppytaJFdnO+KS9oEG+/vH9yHlmjWBz+1Gb3K3QUx1EHDeXSvsk2uRDt9o3iq2/sa
gCAfnpV9MRzXRxCuGmX+oVIbVpgf/UnqRBYxcnXC7g0aBdT8sWjp3I2Opz68HdlXzBBQqlS8UFty
4T6vdihD17BsSkzjQAFIuvfaLlHsS9UrbEMpcyUf38F1j/T4Y0XwMSaEpFAnFebgaZDlEe1HEsi2
IR3oi3mLZeiKgVBmFKGbxRkGibBAae4szu6paSDt9Yt1XYHW6f7olUJttEqA3tXoA9Mky0nM3/2W
THVpw9Wr5WpIvRCj4hTpQVVhb1MVf3pXZzR0RaSkLFM85uZYX9m6mSTm6t6YlNV7nHRnizNKV21G
HI67yW/SE1Nykc5QbBUEWGDJvUuo2144YZIvjz3cbHQZSEe2cGneiA+1Vx2V7UrsacPpOaJHTpB+
dyGJrNz2b0PtDLsDVSC+zwJkXhfcOqw4R38L1CImPloubEkhyoN0QNO+te5C25x2d7M4nCGrHG0q
kun7xmeAsJWhFTO89qEoB3VYxKO9yP/KNc+D5Qgd957qSHq6LQFOdC22hL/TcgLH1XTXUSobmzPO
ysubD+Edn/8adD9EZGyEw4qpqup73Hu6viA8bH1sT/RmfCC+8LVv1b273jM+/X/MTGOORy2ALlsn
JrYV61c7FcZ5VclMfTtTkDNdJbmjEAICslPJlXeMW9k8pA1SvY+1DsjENUALZIKWxTmvlXcAXyms
eHq82WNw84AicWxAg2Lc0HUJ75pKxvwEquVVN4YI8WSTq2PSZDVwRsLbfXLPp8tMn3nfOgIVXKIw
z0t+uptRJag6/Dne4EThgBVh0qThBkI2ch+Vb3KRkMMGQ+clnM6paz2qCV3faVudhregkNAeNBx5
Dc/5I0P6qmIZehBbR4fXIY9vbB/IN8vAu0bpr8STYXt6I3kLSLmy9UpBW+ZeaoXAWoJuqtpEK9Ur
8d0l7XSGLJyroyPHKpvw6YVDEe+RkXhpGsUhonY7fIeVuTjd+EDiATW2JilKsr1zJugUGBfdIPwv
wm5yiAp+JIZ+WAr0tPtYukPa/boHoWOyeSXHmRWtHFt7xUHbW5oaiVLkWMKdeYhhUPxheZTEQlEo
P+Adc34zAEb3UTnXie9BV6jQM4VB53jhd3aGK6eiG1L2O8IAcb/Laq6Z4U8JXGEaf1pV3fdFAdbs
6PIwBjCdGt23IEe9L+I/6VOUDo3Y5LVLPUKKzLlRFaUygg8VCL4pdVUG494a355ZOxN2zf5RhjOB
SIbWBd8Jzan59BfN+qtuCiMya0K8upwzlTxEkPKu8OjVKNi9nNOy6W8xdnIaG0BjCD1LG+snhqTQ
InHc/KqX3+ClRSIr5bGAKlCZWJ5k0WjW27ulAiudL1GhmkIiXrjePahDYCrWSKEZ8WUPw8HbsMIz
ZAXC4/laorM/O/j5Sh6+/7UGZcvMh2BHf9NWBcWlqAvf3bnBrjLmwxFk7UiWPtv2W3q1FblR7kQ2
LIZooEFkLkQl0M9xyhYppJ32zwClzTxhcoZZ6JqtcruBLSZP6sBJMvVmEk8JQFeYHQmDa3XVbxQ2
tBzn/GYp24CarhjsovrMObBabgS4LRNcfko/SqoVwagq2MH21s5O4kE86z5LeOyVNd+8KjmrLAOz
fCl33PAHpU/obxyOlixAjRLVAUkp4hZKr5rYb3MkREFSpibyxqRu+jCSS05z0uEnDrfczBrB6JWg
nl8EGiw6rJ9rkzBAlF7s/P4z4VlpZOuvdLFd4pdktoozcZnRmbXpah1hpcHHOG9OuSXE2EwVIMfe
g9r+0UmLGH86loEExv6igGh4ppzSaifmPXrtVL9woPAjrD2Qn82i0N6lo0dKk41WSSFhvwno3gg7
MXiY0aJ6TWGamJdkLQZN6lu5gBtxSHZCD+/WvDe6KYTMj4UFBlHGVPufnZY4Ih7G+oPuCQfcBLvU
i+pqxDJtyMI9k9gJpLQYfr933EEAg8Zq0y7FNetJQzE8TBoTW7pgnDNdRMPdHJUnL0jI0U2H3t/K
wZzV7IBC4vV+WHwfEFnbrOduKB7dtg1CU8x28IjXM056aoWqURoKsJQou+IcYYQI90DbOuTR1NaG
69D9+LQLblMz+kNEex7oHrvKBmYjXDk73ombwaOAzRFig0kGu3EqyF1iNY4ZeJRuYCLXwfGmpVnE
VuiAlx4fGv9tNJfEVCTsju6pctSOFu2pBb1IJPEOZO9TqSAHyY13j4jhA//MUOEcXZvdzzN+2o6I
ViJcs+3/fOHgRJd/Zxc40k14EISMhgEb0WLYzjKi9Y0wpfCXyjYRrfUHjIR80L78YFNlGDzDsv9Y
ICoaaJZKqi/FQ8BG1/n1On+g7JXBMyTuDQmX6kWHInbRe9+/iICZu2/nF4aO8LpqE+Y7TRNSrfOL
3T/b0Jao/6bt0v9dJZtQiFhMB6Zqx8Q/R4EVmasjhpBT2O1nv7MHIao7cKBfBfd2rpsegzogvdEV
fFzyGJ5PNGa8GQMkbVglYXU7aFi3NDJN4tq3mAiy5uoj4BnS7UsefmsSOqL12W6OT14AWzoi2CYB
TCejKy8/gDRARQ1o/PggbA+JHkQmRxEC1tMN+Eo5r2U+I4PkJd8X+0yTrlUyJubuw65HUiyd+XJ+
RY9tBV4XaBxRT/ZwFz4hBwLvOs8yvG/ZNTyNT1HS2A2j5RnQJY8BVcJr1pgf7wtOnNPTNyUmSQ9r
lmUBkwKcQhAdHSAUJ7h3I4fLoofUdUY+WHelovLPxXtmFprCWYCVtj96tynR3EtscOl55s3K2TNJ
nMQEXGaqZpahpDzZPzEsSR4bzwklxwibK25KcFxYQMG83QIgsdSBwp/oM4dXfoQOEUeqgUcGB5Wr
PK3nNzLsexVtDiCPleg+ZGMlcq5KSD7HAXHdDWmsrDo3TroxQZEnSz6WWLmIkz8N1jFojDvRmYA7
lrMYDZ0A0xbLiuEJAOp4LVpcbXqqy+x9grMZDQa7rzMqMeWn3c4Dq+4Lj5dWWr34Apfal/ZHZp6n
rEP8Ce6UVRu1gyiRYfqvKl1DN66++sDJWCC7DU9X9XX3ywvisIhwCV3K9e3lGLkDtsnPG1jxL4ml
oRfu13qV1P8emtEHfFp+y36FXc6eiOgprH4Heh4o0WCmTUBfPQQcSzRAqi388p79b0G0sCV9DKJ5
ql+Lm6zsyIDwtwy2tCvIAWzS9Q2MbM1A8JpT+BJtknq/jag8vb0+1qcnH7Nlu2FvEmw8wrR1Sijm
xWYQRLCNQDBUsDVvlyF/EDu8ZQIX15IdIXlzo1FS/L/Gy4lk+UPX2EnM9DTtDRWrTIYMWxvqaI2B
FKNEsvjCOb8ujrHubUyrc8J9/+1v1r6z4jwdOWsoTOJ0IzKr58gg0JHu3K1KLg8fyYVBL3j9j0IQ
ygCfH2EKAUnkZ87uAKzsQrasOByICEELlYwSstCYTt2j+RnFQy2BiO8TwYN6OZeNDHim0uBKk7uB
2EMIx1FnzzQ24KMP4ehBxi0rwWPvguf9iUm6ZXp2LwkNZW27SvUumcbVt64NQgtw+rY73hWOQKzC
7ftGUYFu7Ai/rOlFcv+ZJ6J2oBugmPoq05felQ52YfF3A4C+aCDlzu8coxrgp6krPfq3n9ytrcxd
5/JmrybqZVzomxotWo6/zE+WjXjUJWko6A+BzsclUuV4BkhvnHyWipnQcDx7yGLL1EJQPaVbknG8
tEueRLGax36ZwDKJaxC7y5OJchUe9u78q6UhWNK5tveTLVDYY/UfKc6xiRZWpSoDDbTWK0EVfa4M
tmx2TTGKqKcYvhfojBpte3rN5iFHaduridTjsgNIvR1PDsUdlc+0nK7qEOrBCvNG1sxaTVlAFfH6
6Vjfv7I73a6jThJZysE7wjzLoc4ZoNgHLb+NYSKaZcmR56mboyiP2+7DnwgrqDMQXtbEtF/lFIDW
yPbGhYbXXDv6XqAa7LXx94Z7PXmASHyacJ2RUwpbQb6qPSLaZFR35oyoyBmJzTDzkGMc8ezU24EM
FE0K0J2qhsRNCG9KC1HDAUuqtH4MXuwSfgpR+/F5m7J0Ell42S3T9nMmnFxlg7oGhqkjeUPhuOMA
XADixTKHNtUhLU0anve/EDFymtEGYz+Ls0PHVjWySMlLZDaQFmhG3bx1a7jd+QCEC+mAkWJwHlaS
RwuDmHTfJXVpgg7iZ4jCNfobd2kz0X8vxZh3BKL1zlKWVUIx0/6xrMZTjD+CjFjonzk//huSMXZI
sTH6whWKszuZhtBecKiPelRcrXHuK1T1Y4vhAjDckZemORiyf7aFj3K1DRWYyHHY8o1jmAEDrhUV
rFLWCyHRlXD5Z5jtxYMC5tIGu4z7hm9D5akd/ZqnikjQgVav2ar4Tyu1vPbMiQ2YyhcZoLDmy/UE
z+0rM4QYPD0vin+ExwfitrC7612taAOOxJrAudxaetgGRjKlT3bjahwpC2jBu9n+wKosjf1CCGUm
WaLAD2vuK5kwa3s5925GAGa4Qz3TfEVCZ3YiEnGR9fdjm7xJviSWdEjKuy+J3cq+Dv7Q3d+DWI0H
OINWt8h+B0d+8sZxp+mPUwSPFHNUGdtL5x6W00MqYDo7BjKDKWySLq4W4fSleVO1eyUQJjsIIwNM
z+BbgqllEtT40loEculj2dOdpK5URh889ekpIVCmeRCOeWCRBFESNhwuaEmC+syEX49MydQ7pYMP
+RKd2EO327U6u9De44w11+2nwz1+MOSUs0FCUyv/7OMeNSLJFsMebIGw96M/wyMAJGMUNxgitHXR
zjR4WXsBTyiGmOFDrOWFGLd9VNe6S27cs1lUFcAy8foFcjtdj7hmu6ZufCzPQV/oxHetcJdiWVOD
RgDyrP4Rf3u3hmgTW2VMfbM85kPQXV4pZ+xueNI+rjzL3C/nSmPD59jIW15lrS9fX1N53kEtJC3V
MOVuzXVrSzdRyTnL4v0CHvEGJzkwQI5y7kpHdtvhZZwSWB0MgpaaiGGjRlrb5fUJ8sULgGUQRgjD
pV4Yauq3KvVrJkTsN9jUsqgoNt638eRpCaJ6AVLDXNMuHc/kGOvfG+b6vihpMrFo3dYiIHWlSk0l
5WdujVvNwm7kkJZENO1g6yYThpxYxtYoim7snnRb6ap4cMWSAmzcgdct2hpsk0sWdB45RDnwsT5Q
yZk4qF5ajUrPX/k9H/tVG9fcez2JP8zHZL7kSiXVlK5P7VyHyYWOQVGM92CJuLIGlhoK6o6jdKey
Fhg1w+Dv64CIX5DkBOBZZTRLosAil0JNE9YJvs1urVxTN0MZ3fUBIRyKbKP6Dl1ipa44A6Bpw1hl
VngWHZq2J3GNAerKM+oTGJZaO+6Devs9Jx9VTYv6/Aely4KjB/17AokmEjUN4aULbOTuJEP+w20y
Q4U9ppPNYY/G1dYDioOJRWY3o4+FbhU78oC5+QUbeqvmtlzfwBvvcltKrwPAPh91RMfk9EWQeyPY
a053WOnmq8Lh7PNaf9VTgyyCR+LJzJyOaa9mu1lf/Xi6rYlp77n7ePpcWweUeRiVAKgVmtNhJJ7h
0NkXnb1t6b/GqFoQuy5zF6ilO8jXwcDsWIkYWAvoFDBPA9gukAhbcz15uOZxCBZqYRPFKvBLEugZ
5vFZFo3xNDw1TdHrZuTt06UTuUuwAA/eZ2NRlIsTThuvwfcEsKSYMD96OAcCRO8+It6mpZIQg2c4
XUpL2KFKWgfaPO0BXvHAwRabNgh0UasUGMJSEhu1ukGwtDGu6/jCZaxvnFbwySMZZvnEv2NZECP+
Ik8pxF6Z1SRcqixpTm4QKhHSNjI71YmdNNKRFIFqCbOpYRirXFIvzCVNGXZivcIG2R1/9zSYet5X
h3wEv6zkH1Sn6nNUVJ13+tIOCrQQwsDjKtWqEHdYuicL1h+act0l57AczoTWUyx8DEZUE/TiiKwI
du7Q/MDnwtZQ2VhzBGWD4XFERBO+bFRFtwtQqOf2z5TGnBkk6EsoTseD4a4/NPWnbJ7DJiUZNVsS
RbVFHHcd65ds3/FNMD8PrpuUzjTvt626xM1iqSfdRqghc0DM4MVppXFJrhqxhqARu/rnypNvFYUt
X/1lrNq2qud4O4eYczaoIaXnmWGayQoVPX4u+pdmM4GlXqy04Mo+Aqq2qiO1LEjH0ZhWzY9gmt33
D5V8PumhQPvVcCF14sFg0AbTM7lF755yRLItMDSOlUbgeMgWRtbvJc6CO9SjPIwZgyTvpBkTdUaa
nIbl6PuwUi8YcH5SFewVdnxWnn0lA1Zj8Z3GZQ9iBdA4dcER5OxgeLuwouSTT9Ct0psfZpCujDkv
XaWeZnH/Q+ftDoSJrMUBPJaDKA24B/yKZPfzgjN5IKWcpwLsmQqpOS/ND3uDQkA41pAwP8jus/e5
PWEeifAQ7+2ZN0W4Vv8BMVhe04iwW4kD1yYycGDbMxC1kxQvxBLPh+2W0QoZK2XBWKqVmNDFsV7m
P10bP8t41YFGUVA4INOtjwQgp+tG3l5ZfEHXw3P8Ai7XN3/grHHupez6xKv39NpC5gVeUKS16MnL
Vi+Xa8HeYbdNlyPsbGxfqj59DUpAkNU/CZwPqtPcrTGSspthI1huAkVPkOMHwc8Ufd6tQ3xxzbEV
/0AlAlpLHaVFpJToHv5GLKRQAXQCmdAAaCEilkKI7BLKxZSTEtsoV074aQ+XRP8a12tEUhfb8BCh
8lNGNKbVr1knQ1DiseDO5lw3yQXJjlUdmqTmCjGVi5HwOqN8QsMGAzR7qgCEMJjl91Bfoo0FVO4j
BrcTw12H60VQFHxUwfsFG0YeGLgR37adO8hRbhZBI1n4VNFq2lxkJijEQU95zpr4JC/WEDPsMnrM
CwMBdb2XdW/otMzn/t15z1GRHxVCpndHFB3AGOW8D7RdEk8xhOZWro/9wKaiTa9KXdtklS7bjoy+
aBMHOVurxNdjNhQzC9/LIqBaAJqbeCmq6my3AtjMk6byGaN+98+Tk86y4a+dnuksMYiFi+ou+cWt
11zJ338Z/5yHfX7MaYG8qSETqROWf8u9XoikdYO01YGipe2T0h3z4oSu65/3XDJ8gSPxI6vjSjMt
KVbX/fbbs7drtrwdL5CLKdo3S0CPvVz280by3WVtrvd/98o7o2APDR4JUDX/ZclqOzyNDgZXwOm9
/HsmO4PDk6D3AEHiC8TgNXyyRXVBZYunE6wKCp4Jr8H3X8uV3NE3VsbfOCT5wHVbuwUkAbnHX8aX
91eVkWAqU32dNLj9VaEiWpNtrh94C4feFhyg5g+NAdPrbXfreIwc+bkmYmWOkN6QGClvKmTQgosw
N6GZwuX/BTFp/eYzCZUh8tO6JuGbPACpyYpljC4ISQg39L4SZGVL/1+kRbW0VT8gn0g9JfjLsa/1
4qG2WAb2t7PG8fC9P8+kRSnFpRuiM0BvbWaAwXyxuH82/aso0/cZ1AgMxK8jeRbhv2zCRf3LZmmK
6aFiXqcenCnYZHw3uivWB3H7VpXk610txptp4NzsxQT6xUS8wnA46syeC+imZDjr0X0+e5JOyYYo
a+pU0aLRZbrbVVT3PHiR01LJTt8UKIEbuyn7TIvqziCQVLZ1YVYBs5JBbBEOYt85bQPc/WEefxGy
+5W5HIDIUku3eHtcRrMyB50IW10eDSTM8Diz3PiywpjP3U8RqW3h5ajAUd8HipmWUfunScOhGpj1
ehlaIOoZBzCKyqMvNrdtDE60iD7u2GRq/7DJDdy9qHLO63crEKdZoIpRwymXHPTtnIlkxmlLOP2r
ik7Sou7cXMtFg94xSnHBNf9YurBBN5tNoknzny2LzbaGw+03M73skexbOm8x/+6BtWlUkVUmzoAs
tEQw2ag900vk0AsNsCLfh4OcxyyPL00CGvpBq8pDAoW3fuMKgCDcLLgUc/2Mb9XDqm8I7WMn0+JN
Fh0BSE/uZ4vNMDzDuW1NRkFZBgssE4A068xZ+UZk4RB/nrp9atc/HbckrpeYTbna7+OZYrQBVImU
Qb04oJCMJsUB/MIsMFhG4XTNwPUky7XdJ8pvp6onZeFFdD5vc0jusQXCqJFBseFvL1rHC7RmwaTi
CcNkXRmzZ0FWbZyVC/1e3eMRIhSMwZQtoK1VVo4JT6hFXnN0cTX2kuyRjr2+YgiQ4NH7yLOfAQBr
wwGgLa98NmLZGUWxyq2NTlzqhQeEHaxP7kZxAoMXcMllG5OhgNZDh77yUbnTHjiD00bm3IH2yTqV
AveAk1Hcn8JtNn+mqPH5e94eVJat7UhP1M9AXHjFVP4dZiH/Qhh13H7vjuZyCwxzkTvxdz1924C3
guqQs3+OUyjBVX/FfIh2FzI93E5FoLOiAPtcfD5JqcSoCzmIafRO2LMINmzCuaVrP3G3a4D7Wjxb
MqIZbEcBTav3RSSAEscaONTxVCGxAV+/py8q1ng5NWsFz9D37BuG53b2ZkpONzuIxsqtif57TSm4
lWXSFfIkiA3ZhWypFW3RcTe4OZ9eRE295k/KGdJJNJV5lsFAanrBFAQcjP/J2pwlpimQYpfXmHnQ
1EKeuz/eNtZCXtlCEYoOZhPTb3+v8rUp7Kz44TSWnjQRYyBjnpbQVaMaswO8KZFnprAdw1TNBm1i
b9tqx+f2X1+R1xdVZCJiBY0kLK5rlcUXiofPzKFt5cqL3xdlP0gt8S7gP16NVLN8d9FuAD78T9Iz
padl+udGFGGjTW1qCyfKMivb1eccnNZgDE1n19ttMke5YU/AaLOKUq2s/saPH3uu3rpbvkItmUoN
4YHPK9Ho9LfyAauyPwPsGkejOvNsXFgXXNhxhla/sVl5MeKnoVUJ6efnvwDoYGywkNaBtSMQ1Yl1
ITy4M9f55xN4aLNjINXqbuNZ5ba/qhs2f1jwSS5w+57YDzOjjfZO8IpHW9B+1HsgVoHVfQGs7JGN
hHgW2joC8NisLyN0qUE6KJhkWnzL0wblPhFK79KksGsvd28ja7rndP7sSXq+PSsTHAZsVDmEsaGn
1r8ZJUJKf3ygAQ5UaWGyUYd6urN15tpHys9gzwxud8vR/TcsyAAswSVrwmPzCuWzs+aatUQzJyDd
TtvR+DhXNiNELaz7Dt4wBeuz6MkVtHeX7rVUmq9jhuUkj5I8qnxbI+Ed0bCNMhU9vp8B/rtl2XeR
yfNWECTCYZCqQ7sdnIO/8sujAp0byU+Bx/Cj3c7tVNmiSBysLnMWM3gkKQ/B+TRQo9w19Y3CAFa6
rPbZQeCWCmT0pkmcHKUVK3LE77d93vqXyAoJkFMDnuRfOBTWeNKgpbeJEMihka6Ivj+BKe4JTxPI
Y0r1z74av8yZhpdBnFz/l2su5NaLM7nSR+i7JFqqTpG3o8UxkPx2GlGFrIgERWZtYs4H8MR4uDXU
mP7YTbAzlYG1vstXnJsttJu68ql6vs3yvc1lEcCX/3NUCZJvNfV/jhQXYYcpy4M44y9FWTjRn7YX
DJJfkQRf7tTC2oUXhKEsmnbVducgFhcuFPjK9h2yfF0DE4xevOaBI6H8EvFmhu6h8V5ueqZIOpic
VCpSxvy5i6yiNi++TVE70z3fTnUPwzFPJR9R8jVMS3W2J8/6BU3D3t4YUdL8RO85NS2qdUJl35oy
AGGHZQ6Aq0o5pKyp1ylI2KQgH5eIXpy8bGohySI409OnQ3Wczgou8d/lyghrLpfRdSO5jmyzjfN0
QnanjUuyXhVwYWhkihjHmErmClSmn4Y948t0vLhwn7lbvne28AYFW0Pvpyk1e2dX/6chgHYsT38m
2RsW9uEl+E6af85tic/97rT1fUA2386JmqumRM/MrnEhbwwrZ00spYeA8wE2r/ayJ+aFkPX7bcZY
aXYStbbIliT5LFItXXhtDDMwbxLb/ge5Y770zaIDS+kbNmKonrMh7s2m20iTejERyl5OFeKMYAHh
srlCyASk/vCt/IhMIQC3HSXpxcfinEDesnW5mXuvfRjivS4cpWUIRFw8z200GLEZcsScLQtsQ3EY
RgsKW7y0D0iu+Drteu70yEYN3ngsq964AR7WFP5EpDeSW4AlTkYFNMwC2KQP3sJI9uSzr/auyRW1
2GACR2I628mFZif8V4SQfxhPz/2JCI8GbXjKP2btHodMNdw9dGMppmhmkp0P6LALHPBQLw7O9ZjR
S2A8NUv+VAgV2G/lxfCcQbWpBPyO9yZ27/4oahrI1XsAJ2KuLStM8Rj7DOI0MpoiMwy1RAysui5p
J4I3S0Ev49E66l65aDOozXdCI9+AeKzW4ddITsG14Y1GgLdH0AEbjh2mJF6G9zlublV0P60FRfTz
s9ktvE4nbYAIlx13+rClT5FvJgnsUXpmg3E1iWcoKGPcgx0cTeqKgQqnqbQJUQO0T94pTawzNY/Q
/LzpzD4/O9NxTDXdgBXlXOwiWL0AEfh69vkHSFo7Zzs+GqfTqLXLdaAqheWM3cQWkZ1quGMZddWo
09QSvWCkaRVZldTfH/LTv9MpoEBBloVa3cjkdsvOn6BuvOpEILX5P0XWDDG04rx6Ps08JVW/pEiz
q3metHVmndFozL5k1ZM741ldBXkUR+EMZ3Aw/JZxES0HwfEyKzDXmi7pjVCJ5ZJO/Sa1hoHG+40m
qITTZtblorMNa/KbIHeJ2CnOMyE2bgwht0pefSAzePZrEwJlHjXWs1AjEbcCVo9coV0s8d3ZRYWv
hB4Y2oGGE/8XlfgYIhILy7kRLpGRn0uVP15HlrCxsPJryYvLpTcIKd0wXx0twEerJCmz7Q3e/twg
Xgr1NgzVHBb7Ppy2oycDDdnMOLc7xyV4b+RxpZXS8ANh2X8GCvF9xBhPf5RNSqHSfCyx2h2Fnh3g
cW4WScyabnPCWAPWBTESQQmCgpwr9x3Meck03c2HD4qXV4H82YhuWcYYqxzz3o4kpp+c1Z9fc/n1
k9v/IUMUkc/OP+ImSRDUieZU0Aev6C983Gp9carU4iinb7eOeaWLzB3ELl7enmVmrVUUgyuprVLc
2C68gt3IodG/B6hhxgOGZFZh6/JRPKJ7KeVLRGzU50cd9wAr7eTZg11qShoM+3xv8pUSOWfqFWWf
LKJkNRl/ltrPXWRwcWBTa2B9xo/d3MFI93STdtyxiHwzUcmriJIfdoCcaypO8fX9Vrs8ECD3hlpL
fcEoxtNFR0klXYqEVlNsgrXoEeIS4cV3I3yxJ7XlMWybVUTb2TDLU1YgopF7EAkCfby2bV/s/WoB
5G5huMIaTP79LXv7wJiMzpdrQEFTRysi8Kz1GhoJF8RLKfY705ZFBH/5xUs1J9Zl3pE8Hyksr9Mr
Py7CCNMt8iyh3Men82G7iqrhWFn612ENDmiSWrejjnBzefk2vdo+s8LmDEXCktueT8I0SORtsi3i
zsH8EPwUCIE6rkj6vtmoiNMbIwj60XjjA3L/onI9LIgYkXXBbA3PWA3UuK/ORYHuh6drY7FiuQkL
2bRTkah0MSQjibA7yMmITNJGSLX4V2rdM4bnQv5DiRQlLFr0mZdPzx4+bJUJzFIbSE/zAp6gqM16
ljco+mTkMb/TMlBsoGN+Y8nHgO+eCUkb/evH51SOZGJVSkklbwSO4TDaMJc4rM1W+vtccpS/oysp
fNcWR7IhqN/Y0wiSsSofva1FMC2mG2jQCHyAcQeba01PH9XhX5CB9rSbHZ08sQQ6atiDnjA7Et6v
D0o01DbZadX9o4+zqJV5hF2Y0qtBmpkslYBY8oL4xV+QPJdww64oMbW+Sd/g+mFsFEfD2CvCzHDz
1lcWuwNmQoYnFfmAqzhZwG53etk75fjrQiTR9ykQ9v9PG72dat8Y4Nj9Se/w0nb84Ks6640pswSp
sh/rtmq9Wct3+fHxAlWgQL5ENZacPWmiBXIVAHoSHXPr3eOwRAJOze2BMM1jQ8FIK3w2OQ14Dl4d
RpVYO4niqK4ncrJTwLPFPG3C8bDHto0UQbR5PVVD23frXb5KS4LT8EMJ2aP+B8XfMXbYEBoaiwop
8+IXKwenAzCM9SwQzRti4bvnt207ofWHHGCUJtEODZ9BLjEDJin4BF0LfSLMnE9M1Jrk8CtTET/M
EjsgWFUy8wVykfjSeUiqU0F2pPWaXfF1fbetSLpVqD55gkiDDGySIpmWxmyY2DxPfLJGWDqouC16
94iiR69nqqjpX3VzdCTHFLHSEX2jga1ardrZnR9zE4YQ9nq9mrtSb2v1TzwQatSfKFO69iPHu/g8
rJPakzv+u/WpvpFO5qSMQbQK7N60kiIbE4j9uU0WfO6jKvundQ2nnB5fd9ZTnBQ5i74vupUU3Z35
+/RohY/565QaEIB60r0p9spqYmDqruH5xGXsr+6xMnsd0ckErKLj4tmVn3wR169yN/74qImIulN6
MjjGK9PN3F3lTMUkrCVjWdF7DnK19nn7ejLpKIOm4c3P9jJ//H4YDxrUFIVN42brdAV9du9lfUBw
cwt3tvKN33ex6b6rqX31Z/EpeTRCYRI9OV0yYiQJnDqefZY0FV8lIDZHvHJykmKn8HtI7T4KdEfD
oCSaaiiH4tYBIfsOwyZYBwoM5op31E8FvrqpcdfJHrNQAsJjDUub8+E+olX8PMrS/tlfjl6aFFSV
zY2LuadhDAjwtMRRfqtHG2Izq2prLin/gVi0I4t/Xvvt6lWGs8YT0TbbJxvF+YAFw5MtkjT7V9ee
FbPmS7EwImOG+BOddBgtXrXew4BBpIIW75XHscZd5R6QWHP2oZJnH3lAQny1vW51orpCBgUFLY6Q
y7lYn2+J2etRAFhohPsRgeKgj+Iv8CayT4eQ9pa9GQJMOfnqKYo5JHqf+CeCVGCjJOzfaMzA/h2I
RhMDVTl/ujKWLKzXONTyYjBRElw7jzzcuMvs09VNVj5RgGTUaiac6i7cDlkw3gQBTGHeqQtfFU8r
6FbkX7o4HeB48pnK8CoGjhTRzjyP9YDxYcmZWy4l/T9PEe6OTOxejXUQ3h+cEHysfZVCzaUlSIuD
6DJ3nEFmmi3VSkiXP+ZJdl4AXgigdJ9bqzZNuwijodMv65kg8loZaRTD2HZQMN52VgHsqSVJHiVv
ay2fPYa00/2/JNWKpooJ2aYtNR2R0JJqVEyTYpRXqJ4fzzdaiPKkRW3qfWwHyMSyeJRWCr6TIGMJ
XdgyYt1TvSvQ2GCVMUq4w5ziJfVSDvl6gGLFGDVtvZzbGMqmS8HCPScz1qFjAFqber0ceLPfY0xV
hmOXunbedB7vpLAvajLOmjwhxeVTD2w37ElTY6i/pxTCFlBc+cf8ZnUQx/p1vJWN63OkSyMbbN8r
U8cbxe9Ma5CcQ60WvG6PwOME6N1d6OPHdrMNiqMU9Jb92X28wVT5EIp+yW+rcAdBmdwDlOF0AWbG
aFTx5qv+bbDedtCgfmrlskF7b0S5n4npzeoaol/NAHF4jLtFlHfFUxoB7no4Dln1QeK19MrKntIz
2YIIVPKORG+suQV9KV+vYbpxwaDRXZ7s2czDsWG2MxdGTdP8L2I/LwreQN411YTAZyHst4edoUa2
ccpZXYr63USBJ9NsPSucsPSlfge63Q6B3qOhL86yaMj4auTE7CDs7yIt2JUifs9aNL5MrC7XrKgq
wWq9mpRjs+btDz/IhE3/f4xjjpJLD8pDfRhNx4X6fHAQp5vjBh2cXFTHYYIKDOS/V2FgG28qZ8vV
3u6c6ygLiwlPygMhGpJNcsGAbKNyCQ6beEF2UURo5qQxWFzbI16Pu9M40NbEPlgE7nTMq+leWBf8
x+SLwFF94eqC6DTMPyed7rrAnKrU9yDoU6yo+DPqyIBoUyPc6lIs8U15VrvVEwMq24ArEAEw/Qe4
tfUCnsHS3nYNXikb6ZKCYk3UzmhS+LlGwW17vMr+hwOSdREuD2m9cWaVY0mClClEOE32cJfuxTqr
wLssqB23GEjS50NUVCemtk8nWCXONAcsi8Fa3Bz3UyeWCDIgGvFHatcZC03X5f+OHwK51zlWsEOP
HLbqE4izLlfNd2Suc9R8+yW/0ngFURHnQlb+NYb4/ENVlzlIZW1yoJy4VrHBVVnAMiUNyqZhn82e
KRmOp629qa6lpF2Jf25i5ca75KYwKXY/GP/KG+nGHmUmV52FVYhU4HwljRrgdHlnELB9FaHJt+cR
kGE9NgX6/0UC8+kdLSU5eD/zXmgZybacgAkkXiYJwSDAvH7SXfxeJV0E/MoRhPzSj6QA3ciAoE/9
ZnMK7lbCsNN+TJociuUl3izV5ubMm9ry+ySpTq3YM7N+yU6J3OOjoDFHdR9B0gsNGaDuAgjBmR7N
RQ1LY6VqS5IxJY/2X9QIaYZQFXPEDGGyWSZIWZfv94ISfTztmTKkL9U90QFFvY6lDvkx5KU87/fK
BDIAMWY2xWulDC9/IVr2cS4RPINKS0taCDK9pFoDAceoFxMJpNBAWAJiecZYmHG+Qy7SAiydaWtG
t/N5JjhowajLYPVlLy/ZMo8MN1TgZAMdUB5Hn0cHfu+3advaX//0NAf02W1tnACQZyFpDJIYXefw
zGR/9mNiyjtJIiTropZZjBOX7VdsPEAcFoi8FyO2M7y8pBiyzYsMUHWuArAKJmWblR2hIyvHZFqV
Qrv3TDhG4Fa1xs+/VUMrdCSeLuz/sw9W0xKQMYZE4hGIMNlrv1XQ7BN15uEVom4mifGb8/pG8o4Q
h81ngvArYRlJKQz7rAqGAsMsr9orcgIPXMQ3JvTCwUuvd17mzf+HqSaGNVcqWWacCN4MalPXcxBb
tkvenvAUpK0/JJB7DOG+KkltplURRwIqPjcu50VTNy8MY6VOVdkNblObZ0nYJlaSozD2VItxLX0A
3aK953h++5zdFGtPmf0SVcTnyHtInt8cRlEUbUF2D+1ENgorxTNTAUClQYGutgm2T186RUCFY0e2
eavoyY5mLP0kUPG4dxZQJWDz0Wr4+G9hKzKPRaD/67xSKoGEA1YEIotRcOkFJBM1q6qKzoErmoSz
0jikSDdwX6aZ62WyvzIZ1xY8gPohAOaH2Rk22zktRM8Ll0tRF1z2y7TG6brVGTD+lMOS038/XUzy
xdFnrFQXsFW+cZGgbf3otWd5N1rftM7YjSnz3VS2YzH3wG410sHBJYMZ51oWxRtBb+4w3y66EvNw
8xcMy/3zZuRdQBP/1xb5LCzMhSgIdG5w/5Nrf3n/rh+BDxuvpelwo8COo+D5ER5E5FeBqo718lfq
Lx5LSn7mInX14HGCZi15bt+i03cMYnepA8Boc+dhp0Ztc+QAxASOtM7X/80VnSwF17UDIwajprOX
bYmr61EqqbIyXi2FszCvLGTNhM+IEOs+W+J/arj+GKnxD3dR/HBDZzrpY+kYgkQiAljNvthrbnCD
l3OnGlPutgTOn66fbYKTunr/8RZjrZ+Hfj0vK+CAcS7MrnNYA1SSTvn3q3ub9Zr9EPlRnycODsLC
xMdOlaUQl8SQXdHJ3s2zUIty4a6fKXn3DlyabmZ04ONUZylf2VyOcV3meE8Fi29GHzzlhQdBCmVC
J9+DQppx1H8npQY4Atr+nBvFxmKz5Osxn5bzT0PmZ/AI5x0DKeHU4hvsSukfIkm7hQyhLd6XKfGM
Km0wBDxBudOc4TmF4SVNLmqJQJv6t3NGHPL04HEgghhmByOjVu+VsfKhsdSAUzpVGQXHlxKIseXj
nNHhgQmVKXOfwNzL46sSszq8gx1yvf4BjmU3qcsYlHnw41dSCQSUM94sZ0GkISbWVAvS8EEPDlJA
yUWZ4OFf6NePU4UxmQfJze2Mij4wEyLDOdUhMlVncL/fKZbh5IRK90ARP2MbdEpDSFzVPgP5NzFg
ZoOAIcPhtHWuQ+NVFabx71Pos8xIm/jW2nZT4WQB7w+hunJNVnh/dXvLSKj+PGVY7H2u4E1Uyipu
Q/i+CvrrjSN8ccyF848ysl0Zc3K9cqT1JaJY1Q0PMvjVnn5m0pzh0NttjQtwcVKS99HEpYLkTsQB
wOAADSlPEnJl5LPZz4KFTHvCeUCFiG1/zymgIznXv3DU0CHL3Y40fQOR+D5LxE8bGkAsfk8eXz7J
2F3bJlqxnBxlAlucuRqyOgyTBKlwj/Cjg3YJmNAllUcJkjKDf+lFt3UhaxZaNIb8t8cHYhwT3CJb
YhTeP9uIL/IM2RZbQUrsOfMIVjjwGFFEZXEvIqd/IVtGXzNxsEYjc+B2hD4OVagFKYtiwQrMcunm
L3TgJyMoQn2bnuAeSFdD1W0aJHseUFujoJ1H8mxyUyiImGiRPqMmWE/c6Yc0De27cLLb0kk1u8bp
qouFkg5pdj9ZWK9QNIFFLzRWVRBOPaqRyQt92ZXBYIWVPYCj/n5EB0ZZ4Zf2vQS13DSf7BZ13Tj9
MlGRCg++jbY/jCEMQAe9ZC2Ehj4HqUJSO0lVRZsQVNtHCLFAGfVNhcNzmA6j4OlwivLVeP+zvZgv
Ew2euN3tyPKcT60cX8ERzU1bZSvTXOLfU0KvLJsZFzAJPen/egUEzPvvOwXYNrXvS0tCI5qRZH/s
w8Z6/7vcB73feMHDTUut/+BjuDaqehnX27G5Mqe2ywIbNCYsvQrTgg0i3/zdXZoeeuqOy0mNOSdo
PLa9KDWcd5lJ5WQVI97z9dkO2Vq3I/XfLcLgVCIupM2jPPoMUHqPrjjXagTfZlmA1YDey71WdXxx
9KZPPZhWJ+MwvoFfJpORXSKpsV/v4YDv1BOtFWRjXtKWlxCP4x2BZqI1h/vaii4t2/pZAataqfvc
ZcFJ2TB9MK4mFSbt6pXRf73NyETSoYRCdAe3yK5W3jZRq4TTQ+Y06CvXmifM48EReK/aNXpJLKT8
ChauaPQOho4DJBhBnvbRlx1AA7MyZ8i1FiF5Ag7wjRHN188eEsSSc6y2B2aml/s80aJ0kvnFRPML
HbnHCdjP1DmulJXBYPB9qpW3l820Li3g5HLT6J9MlmlLNrHxqsErbWSvz0jWYQrj3uvTPVfsGTTB
IhDywo0pyJTnF0gYnoAK3ZeSYK6VfGxLqx8ilow41sW8jg1bwybuwofQrXYVyRWV50Z8sTyku1Pi
90YjM2MortguiHgkQKjT8vegYhL18p7oa1wy5KS5In36L9jkvdK4DXkV6btIgDOirGT6PGsuRRSS
CmYtz89hGyWjMbOPZT3P+8diYo0u/zaUEcaq27CqRjiiZvL3/IZ5LeW4OI+ua0r9iy9Lp4Qp5Ed4
/u7JvBQYzaB2KZ93WmAcy3P22Zls1ent4Z/GOpWEoY97vOJBpnuP6uqMbAES5qY46nXWHbwTXOJ/
kmAyojAHeZTbOvUVVcCHPy9FCz/0HLaanamEUygtWlUx1ADsyUoLNRZuugLItzBSbb9iMorIZlsg
PE+acG7iQzkPi3NIN+hAtQ3k6gziLxw8xN3c7697qp7MRYsevFVg+FTRiEtrTExQC/gfrWsakoov
ME9dGSLF7bvPfRapxiMti/lftVr2nCeaUIi4nYY4AjKVHJel/hnHG3ZsqLhP/FWgZQVbvkUAB3vy
BJNYb3iAE+7jG70vXMV+iCqXGWftBSMpGErGWQrUsHBRGtogiMuqcjcj4nutjb0iAxnFpofvYj/L
TC48pO5yGzKzounx08P+PxOihChNMAB/e1wHfbi3OZDUO1nh1WeGxVOq0N/Bj2R5CTfQeZKDqjgy
VI0nFCGA34J1QX8D/wtWEtGaWxP4IZroq/b9+eD1aqZ1h3tfnHHAQm5CvcVbECSisys5sS7y9WfJ
QNjiUnTK/QRAIl5PdazpkiofGwDRBofoW3sZpJxxyXdtboNAT8Lp4qVDmiXPHdr2nQK+IqImw34L
lHSys5uM8eMp7H8TTOchgZWPSmvsq0jQYw7LbkwpI9w8yHNARZfzGRI0N28YhABjHpEVQglNAGwx
RbDQEdZsTg1CjaTSKE5Rd5lzech655FQAXv69QX+OtqIeT5N+9N+WY2bPWTLtpVHiGVROuAVmZ20
WLMgyEHhSSU0CDXXab05p5ldFNsJHr2vC2H4+QHMIQd7VYAAOqBczb3/1qlYkjcCIq4+TZE77UZK
nMh5SE9KePgxiwoP8otggacTOL5PAvCgGDT9+oX3g8gYmhXv5ocihk74v0AqzwCmdvv75WaVWbQ7
EFv2o1VsbyawN25/UoKyKR21uZZRVz+v+zdGGP7tXDZaMQ71zEsBLBKQK+oqCXPKuQO/seMkVYLx
bohznvwwaW31EMY42vjR/objm8o8QbTymEmkcqfGY3FAYStC+gHi6iLPRnm0WcVncnjIH/vDxSow
zVklgI9f/SJgFOrhD+zkuEc86iWru6bRqW39DjO/w9QetDJSt+EdPhTaF1vjDuoKkh2J0HdPbIg+
j3ych2DS7WHTmIWHa/9j976wGQqbL9uwR2RJrPC7FxqdT0Vi8a5FCqFpIsopoEHXRE4K12IzYqlQ
WwV2pUa5nz4oYuXddXon9MKBd+yOElHb7Y1XZd/KbwE1tAgllcPN0mTnvrkVwdDlSg9UNvAdkGtr
Rh3YePc5gXH4JrA3I/BhpwgwwnnDR2+pMXDcoZ0kgUUZmcDYuVVgVnsFKprOajMQGTk88Xnmrm56
GaqxRIVpfmedjGgFbJ49bH9tYdghX0e9dQV08Q6NdJ/6lmFc/qrUswP9tCcQH9ThkF+efBDpEz12
1M/e9ACoPjKd0JLE6UV44avrocdcb06N083KoCY6kllUDYFQYilXTTs4kSJ37NWB4bhK7ZuDiiEN
4+x4gdCKSf/TYmNPn1F3nfsNThMA+zDEvncf6oB3q+Zo6AjJKn9qeSho+mvU4CpioVmJY3JY9sW6
V5qm+b+2BZl3IBIbnmplfGg42KnrGRidvxoxSINJPdLPQIzuMmCCdwufk5EwtrfutMdbpIB9xXeB
jZorIPB3wc+pDTpOXKJJOSQdiBw05oehEPY9EfpfyyOq3uK3RXCj9UXtCaN0UgLACj1bEe6JCr+S
M8Bkln7tfkXmmJ2JUgpCPCiYM0J+DCR/9wLAa7Oixgtg6qqtOVPJzVapt/opDFRk0fnZsrCBYlIw
DW9CpB3yxNr0Ixf6aVkYqTg1lZIsopiwlVdR8NkINqB115b/ja7RrBjxfbDJeGuQkHq5U/IAHjDG
AgXxroOvRg31L9cTzjtrqk7896w/hoaw6tortnKLJHfFKRn1SM0K5xaW2DakY3upCYaLHFrr58Zg
IaJvW3kkHbiIsGQcaH1mKadXXghZ0eQQ727j2hoRJYqx3bnUw3kvSQZbkaUAtlWF1ZA1jkZxAIe0
HUSZ7BNu3kkUt3HNItYSH1dLEnce/uY8wFPm4JFmSwMLwuvVPUCA+Qx+miYI/pH8uA6tNcxFSInh
GaicPY3cEStaH9QBw4AQDJTJkm9+EO3aiLmwbvfORPJ6BOTiC4g9aqkPFpYUiQUYt5bCzGbulLLD
TAqTZv59uhGGJRc8pxeOQR8D9huvOGabj/1Y2krvSJbSXcTL/77bgMat4CBenb9eqnoU62M78xSA
znH7gehTcaNUdTipBiz26PFZF4h3Sit0cFs4HXPa9TcMVD0qy9Oq65wR7AYmwnSV62MZlUHOGlhc
yNvUoDLH4U53luuZtnXESuAVeIoJoA75rz4seLl6kLV89Zj11GL1f2HZeNQ3RaRo7GV4nkFOuH8k
6BG3bNQXqMDc/NYQ8Z2QZL077R2EALFzLSW6OqcmXTYPqjpt1eJA2fR8zgWJ9NyMeJRe+XUZ56d6
ZpdNCjmARs8NvHzJ5N1MlJczUKuuc+ZIerTGhe+A6Suv92vjOGXZpvAGvqFZlojYy5f/4UCe0uiR
XwKVeLLudE0IcglfNkfOomD56IrTlJjtGr32+FqVyIEnyWMWFmciNwNZTqRTYfxvxfzFix5IYfHO
JrB5Tcmukc/D8w5hEpW+9LXmG8/0kjenJR66AR8RwvGIe+Lk8kCba0D6/fu6i/3C2VzgvzwIfGBa
Wze5DVkZMl0RGtZWqommlnW9dAhHW2NYN72Cq07fd+lJ1FAC7Ih/Lf4HZc2qfZzpa33msgccV/CT
ZZ/lDJqJo1a8szDhLKom1aONY+LKPuZYz2DWj779J5LSsGkRjC12phuZVtcMvH4bIjO5FsZIIzP6
BhS1mD0dttX2KxFx/1V9tjPKhVMhDcam7P0QXKaa+IRL09NkM3b4B8VnGmEDSA+QVpl5TNKhU0KS
i7MaYfhprTaWFfGu+pDBQFa+S4JJzcn7CJB/QK0PIhGFZWJKZiTftL0R8oRjBKfouI75Qfe0+yqK
rPVzkN4K/QGC1VvQesHLMHpA3wnZRijq2u/gSJ26wu6UVaJmBO8Nu97rIwaVSIOFn1Zry3WMSVIa
2dNJY+dxh7fE+RnWPVNiB2FkpNy7rTp7LY4oJhPkVDcfzQzO62Vb8MR12pPogJ6mnY7DOsvdsLEM
f1eN9+qj4oOv7QzaK24gwtmaEwN7qgRPitcJN5+osHekfVwfJSvbm1srzkAkGlPnyIToEx1laqLU
gKgzsukQLWCCMgp4jYxi0I1fevMTK2dPi0ZwwnwfybgwhPokrf0IaUaxOmFKizSCfY4S7qxPc+fM
crT5FdzLrjRAmjuSVjYoX5c8okP6e3QPD6HG6a8LdGFiz4Tw58yfQK2vEx1eT71w8vdgMF6oAdvk
WmkV+9tGKe7PxdpE6mG/76wyJBQdklvrLAsG5XV4x6HuZprS9tDrdKaavtNhd4DaIvW1wtlhMOuo
jkW615l3ivUoGJw9km67Dl+1tdqm9WzqNDLFZcNqbddmqllujQUNNRExoy29uE+7yc8JwBuCYtR7
b+TotRjfz5s95rfD9ewfhyDpwID07PvY1/MtID7oa7hsNBxp95Axmsacqpq8v4S5cgGzcZtmC7JD
38AbnfDrhj7iYaK7yJoINkhUhTsc61pGt8GxXQmqGpnDtgMsMCfbZi6oRcuqKoqCMfiVeN2bBv6u
bPkg9udYSLqUfp3KMpn5uYi+UvxbEJRlU7KFmdrqoA3sQPMoBiGJ3r3pbmK6K/2iZHmhYpl5VBYj
lRC36384of6YqNA8N3CaaM9XUbUeyMS6LKQyIZVWG2gLdTfCyRV3xgs1xj1OOH7MRWyymhDN13bb
pGh8uVVFBDAhUzRLFQaXk+zu8fLAOAqQKIZTRPjNVswN/9glk3ogsRWvB4nseu63Zrg2E83N4JcC
3hVECA4K2CxlredBNOclC9cp0saEwpcUX58b7/6uHBEVO2Jfmb9vDClg5gEwT5VhZ65qSSzDlk4B
W+LJQwhhY9no20/QxFrXLeRgjmOVhZaaDNKJ+GZliL6kgbw3O+c199KIXs/OtkIQ4ZqyL6FVRwmD
7Z99L/AA93C/j5OSGEinsilheab2CyH+gpJaDQ7gK8icWRqYXKlO9nIi3H4yCUDjXkFeQliHtzgm
RnbjY4DItMTRCOd+j2qbrUOFpyqYF+PrgEnEYsT4eFl5BlQ6Ph/xUZblBHotBfghUbPuI9U4er5/
mfhlVrUeCR/9SCr6GXT9PD88ZQ8s5BsIOZcVmInzTQNNp9CVDiH9odnEVujggfVGNLVjzVNrBf4Q
vMiRDt7pl766Klr3bBUIbDlOYaQ7X6vNhdWx7mQTEXUiCqfyKGzo3BowawZxBiaOZeinJ25YLj4F
t1ijmCGFc7o2mdpys49af1CVXXQgofIPhBmyLsFXIwQca/uGXPSbkqLGFuVWu2VXUF4NcTKQlIIz
2M8RJa45V+mrzK72qKx4bu5mIwFvAp3xeaN7cyNT2+UelWeV4ZqMcmPQzw8aSnlb0T3stDcvTfrm
hp3r955SffYwChFE3jzH/FmWr0pBre2EpJ4YgyR4VdVCwF33Mc7IW8xmRO5649wDotYSvkRG/maQ
KqOh2IDmBTFd4LerZKYB70xsYqPK4C4nhSQl5+jtGHGMfXtS0RaE8nwKH/71dWY6drAAWGZoQmo6
AvAcVRE9/YyYrHKUdb1ZtLFfJVAkJQyI9me/YwB8kfCHesvFUCkH/Wn1ndq1kyaxe+C6wXGKGk0u
zum3G0+g6GMjzPL/j5lAbcxTBHwPWXQewXB4KHw35+6jpIitkCfMTnQkxoKaD9vBGd25qLzv5egz
hoa1pddMgh68GN2huM5M/aZwhHtURi5Oi0yGLVcftyQk/PE62xmmLqea1Cf8qpyPBeIcXvKdfHv4
pXtFAxATEG1vWNWvkRun76OBrE6gClG1uxeydRG74kY7F0cSkS7LgP1Uv0v8V/kAseVERxyI2YEk
bfxGVAlvRwlC0znNe1XfLYLyc/AlpJdxmF3EPSHFqTFs3MMmlYtVClHHd2WYqMhGDmoh0e9QJmcd
hHqyZbqPEIiWOk7FuXSPzZ206EUkOEclS9qIvzIPcCooELou5kDfr4XCpiTCoNyK4FBwMIa0I2mu
QkDc2XZOBGXpgkbHIUFdZAqa8axFTg0nVWxKhWoGoIyuCbxOW55pcZk2jUPhyhEV2ht//npwglcf
fkiBODO72v7KwY/s1Ui0H3N22EJZ270+IE044B2osGZHYzXvQW2mgXzklbr1IaZhvQeWoJvgX1f7
+w8ihFBar+xfBwSN46vPIa0W+cxTJSpdxkarn7pk1xt789Lt9WkL0nHekGxBFA7rQJ7jqMb39RDu
RWzL4ji6W1v8jVEN7wuDxVPeQdZ2VHMH5r3GY2QcDiNTQYHhUU+nPxbIshNkRmCMxUOi08KC5DsE
zDYlN6qHcFJfc/NX5ryh0zzbLboXp1oUFUjMP4tPvukne7/++AVe3aUK5gqAmhbmlo+3VxxqGR0J
FGNZieEorE/6ZYfw15UUW0NLyfylWgIlrJvDoxWCDzfU2f8FAsMAVo/8Df0+PIc8OlJxd0vK78fm
82KFsmd9KM2xK5HqeVLbi4wPGkLv/ZggiQkAu6FL+JuLA4gZCQDf2RMQyC+G9YM+Asr9/5CssDtt
Dqd841yre3+pQtZFlp4ktVlVefyDsN54VnaCg0TmUjGUrmOyaL27dg1vzaC/UqoWJmJYrvbghQ3i
Y83fmNQXgIXhIj5HOTxFU61Mu1vlO0PEnDVr2+ddDRMIZ/RFN4xMuJ1irw5QJCafGvtVPOggCPGy
zHPPKnd2m7coFgHN4B/fstiGhgQ59+OUW2fZyWlkHD9K1h6QSCAWX0pDDW6+/LuUSWuFrXG1szAp
UDxf5OIq/WZz2chdg+GTM0fjBO6A4GZX8/mssB/Mjs/mf0bEUeqZ8Uoap9yxXGYwks1nS/PVB+z1
iioxUsbu5+N08gnrL4R3GRALiVIcBh5EvfY9sDrZyT+QunKe4DPdNkt4IPmABecBYjdOMGi5LEZP
84GOXtq3bnqabJEVR3xpI5R1S+If5pqSEqxyPVzIEJen7ce5yHDxR/UugyKMcpLb/8Kf2Hct0F2Y
wopezOrY4+hYb1Q6wuyFvqkyThGqTjhu7P/Q4a8y8Jk1+yGGeYIfzpAMLbK7UZu3Yh7yDuFnkCck
sAkqFJin/tV3OPCZjZsCIP4c8Aieok93O8x2CSH4omJv3J3La0/NKHwCsUPmmOQUF5NGVgDYxvhr
lYoMGpD9r8Yr9v6FNkdq3XZH/tHnc8rI3KU6vBv5VgoGOQ7dIxsJHgsl8yewYBnvTh/+ClFymd6R
wFSpYo4GrU2E2SyzV7U4huuJEDAEaw+yCS4lydcD199q100R8hxyVP2bcFwIcmmS9oss6zihx5E6
8UGGz4lexNG4YlkYR/Njuav2H79Cm3T+fzSNsUm48U9fpiZll7HWr2XkZCZYG/Up8T7dxxYqH9kl
/0o8uU3xMWtB81oTyn+lswEV65PJmRLGsrHzwZxwrbMJJQ9iviZG+mhVg4Uj034l8vsq24I5SxgI
jbHZrs9f1WdsCOH5pLu9Svntoz6a0fUhMhe6NIYJHuEmB8TX4jn2B27f6Dmb/1ppAUMbULdGYm2e
Auxq3PX0j8PMSBgGd/gQyefDAU/DaDwKfhcfmM9ZZLMD4h8tiITBq1GMxmSKH86B1z1Xm8Fddbbp
8y5/HZCQgwoUXEDLKkB6+cJHg3l9rmPLQmoAdJr7Fz5fDfapELRnTMtKnoDTOr26pyJtvEePpNRb
yeYXytKYwQr2yCE3h1hcjM8FVVC+SphsIyr+NR1SmueUr2qboumc0nmt16Y8dW/fBnzdyInxaHvI
O3j9pOdcYVWeUYnZTS3R8DWc10K8ceScQ5EcHTvxlGB3PCRDKLrYrKQNl3eMQDzhAMwTwLkRJGEU
PnQis6L/8G6sQITlDaYYltp63CafNRvDU+SN0UtVAV8a+tmfLDnSx2LF1wiHyYBX+RieruNdkCRO
berr7qEKzS3M6hC2erEslhQJr16rA5mu4hCBL5KAZLqDMqafvA3JTgUN6U39IfTAmnCZja3QWOQd
IozgC8XAU/CbwtWaHiGCMQTtnHpxDCqPOX31J6FZdJqK+GoIg7kG+jeVICNoFP7UlIYKdU7FoQuN
xpHHNvAp63GHYnnM+uhXa4TqL8Vkgyu5txAgv6SOTHIXvGtqjQvW6oXejlddknmJHaI/r7ab718D
wAiLLy1bBoGUfzA29re2FOLue3B/F1b1nwBKCG7I3gsjl3KGgmMDjsGCoKqIxPtnFZknBNbMHFaq
2q5R+wAsgDyBw8stn0vwDvUVJp39OQyV0z3VWihDw7/kor6tE4GoNzGS8SlY08uRSwUfBLmdRrGY
+u2U2OqPUjPRAEXGWkQY+NHErrtGPLdXkFAZWcbYgxi1x0pk+/ZabWZNMnVaHFHOnExJKsgCi2PJ
acs84VM7FoeLVpw59BBpTgV5QLClCrAwkvUG0z9OkoySOagvdHzOc7zb6PUjGb/vWzJxmNJyTCTd
oJYgyrp3PoK3M7gjnSM1eyCZhCZLvlmm6qEtCaWNLzOjbiauKS0Ykn9oxSWDl2koPoKfKFwakwaT
0t5QfDtwZpc6rj9LYLE5eDbf+bXBtP48fEKdgr01wZSyFXq05sbVp/ZmnFzOZtlwrJrtzS0YLEye
vjnRiXfGdER+qK4qB1PNwLfKRqwKvGpYLl7PVi5whBvnS8GFj6RCAJhcab4KwbKZfSoZO9NWRbhu
q7NGKdRczsCBdAGo/9ryUwDqWF6TtNjX/QJ8fdPU0IIjNi5+WFCe619FmjabABVSiZ9oLOMYGBta
AMHpNlZfZfoAuozBYSGGDj34kARmR39ieg/rh9uD7oumSvLylzHm0mefQpyxVwt6WyUz77Vo0CeG
45ZMub3z83tEjTydnvld/zmynlcxg/UJSMjAcjWYQjd+AW5+4ZG4TSy8eJ6QrP8eYM7PXqelHdU9
rwPaXavx4hJ34MUxbtWA3digDtveu7RXT2PIk4glc1EVW66Cbi3QSmIckM7WxTQO/lgbfbTJAw55
GB0iin0RbWt23u2325IN28MdhZXGhI4OCBJ37QFZQLo9AOipQREbhAtr9Bw6xMJIZPhX5y56I4W0
0DpzxV5pcH3HviUAx62M5Ytn/Z+e83RdAk9yiJIsbw5EJYlRxudNODh98VAKi2VHuiV22CAhUG1C
znk1lwruEoYp4wks2TvDnJd3E31s0pN6jKAmVBFE3eS5bMoiTrR9egP+Q1a1o2NqfMK+qS0G/qJH
i00PiIY+T8w4ANNXPoPmhlO5gaxSDLC1R/jbr1RFrPb+5Ei0laC2XpM8S1NXWSdGcaePdYKPD2ea
UvfngD9K1mh+C9NN8Ik55Bhel9mBo+DUUuB2/qt0XFGQZ2ujlvhTPVTo7FFASohHYG9XHYIajVBT
mW/sK+c2cPcJLqXaBz3VCfBfS5P8I/K22ExK1orWgDvhtpG9KkHk7YMjAsjbvwhuWBNxCcmcot6y
lewTeM8q+PcovJo6zeKJwv+OnWAlA5cadQxJhXYDrsOyXkjugFSZrPniV6S2K38hwR5vQwDbn/rW
eU8vaMF0VeJz54mbAgz3pMyL4hsDRbfAt/3T/hB/MFLdNua7NRL8x+ArDNq0Tse4GqnD5L14madm
/lw+XCx/AB8x5eXxwTD5Q8KNz6ad1HGPydMBmTFrWgv0ycy3CymLAPur1sP5hHsxFmvUnUhNa9g4
hQ2ooNpB6KFIR0RrhZAgP9VDgmakJ/IzBjlV8B4d0yCGPSn+pDjcj5m83JOJ9SDTduDhfxSzguu0
hcyuW4weU+rSw8bL/mQ+tkw81Av9G0uNOcb6NQdN+KDaL8au9aNNd3KADFZuoA4Ku+NMd1K9FKm/
hPisybKS4vyM8DOrJN6fWhb2iZXbIrFgcrC5z8q79/fScu8uxx0PqkU1PoG9cqhpk9FVRK69PFVt
Q2x5K15wkNqApGIImMn/S5xDswezeXAQl3UIBjGAdr+ZYLxfTsPM3/HeKVJJV3CfVLCTKOErHU+N
dNAljYhUOgHbDTebL0gTwjA4+BsIC4ffiws/2RrtLZJkWarByZrUfvkh6YvjPNC+Qr2T1e5d6G+A
rt7jxOTl7fQMnqCtm0f8+TlAItKw4Idz+zJMqM3tbHZaTHIYK9ENcrN3vjtZ0C2o7e8QWO+faX8D
vERuelr+GBcDqpgYpMm+xDVdjpLGzSdD2kYqlnY7mSCsQZAOp2Vzx5/+bEtcAs3qk5QOxZidrKRI
5ijDRun86S/7D0C5Wgdf08i+L3gR6gDn343rKtG3J4/itDtQtKy+QupVjedwDyFVWbOZc921ag1w
Wr2FBK4PUngmfWC9WGzO8xUTrQmvirqgBoORgzor9gkHY5EyfU9PFna3iIn5trJcByoAOC2uyRHK
90++qQQBWWp2cj6wVjfSmtbLZFLfGzz1iPForMDmTgh+hpn/zhvUJ8TYfIsHD7QUi47FA07c1oUW
wow5eh9V8M1v+gZ9xuywMmnS7Lw90kPtntb5oPtrlieqM9/ZyoKmCZfOd9qEgm+cXIHl0Naz0l3S
Pbn2NxfvdOx+GsblAVdwFtGw6EYGLDiPfDo8UJsffM/99AV+3rRv6OfISGerTmkTx3Wb4Gwc46N7
bKCc0Rx9k6j1XiOUs5kTgjN/8SqBG4Dl1jSOQbVTi+18nk6PDgStGL8FPrSJ/vPUb4OQl9w+TZAH
w+uFOS7K8g+njhJT9tuH7TcrNC23aUnHkcBoVDd3Josv2SUt2hO25jYfKVZB/8KfbNyk2nZtOtEr
q6YuDWJPhz3OX0InIDEpHaFqaFHUAhcPn1JIcoNGc+V7lTm8xk0t1j+0PTao7a4BkKR41lgmkEOD
hFoFsf5uvkdP7I7ZN5PqlXhb8D4U42yOgLDtcePa1Lby3bW1durliG3kc7U5qtCUH8tugGnWsgIL
sx/d5xaX8lSIu+S8eq45hD1pa4Ql1s++a5dXsgf/YOhTqw4wCF+Hbmi5AI3XnoDBbZGf8OG/fTXr
Tl9c7H59l2UI+mo5rGlWrx0N0x//i5KhnGL8F2/PmBjrhls2jX8bgiuwvzzEnnkMaNJkemump0QD
/YFsi5bo1YxCNElJ8CekQoFYCwkVaN0I1tt607C9Z9OquFWvJoYc1jJYrMF+bD6VwPJCMJo16Z4I
fPcw42kVdmfuk12/MZOCzREIniRgGu1z/Jv7mDOuoN6+/D18ZPyCFnBVjZhYs23ibdO2LIz1XetB
z/An0ZiuSiJE+w7zQoxgwjjYHSPCOq362Lm/fRBQDkIG++RfPu4KVQ7MoDv8JKIsSdPZ3migb7/9
Ch2BzNpC3Njmvhr9HL7aXesGV7vliJgMrb1srReuPusde/5FemE1p3U4Su2EvzhqfHb1/gCDpuFg
m8ntj4MxEk24UZjzJRz8QfSVaay9mv6nJ7WXfaexGFPqTwS7wasmq1daVbJU3qAfF+givjuJ9rk+
JaVFUXbz/3/lVZv9ErptOBPwU99CVpSPKDW5LAZic8mNilNF0qsEGFvvBbOXYDw2HXjyyDzVViTg
Ix7PMbT2JC1MjmaKOEjM3syH+S7lmJAOZOsZJgjKwHHHuPNerCBmFp6sAYTVuVWpZqFXe90goL+g
cbK6MoiLnOt++ebh/7VEgTDscfYArcJjHnX+guhQOE+V7fBQlnlHV+vB6/feNWfbb1SaDPdCKm/c
m3YQE6Zu3UjXzkzeKCSoPcBl8pXScsuXJitPVffjsH/51IYFJk/QIP2i0VH+Ql7vx2eMLJWWoE2t
O37TKV5xaIB33KJ4Na9jgkGnr2WoJn4d4F1Zh/johIwupDTejcaTZWWqrKyF9py/SO2G892Rs2fS
tO7ljM1k6uEITzIwehoVwmD5q52G6FW+nTqV+tUEp7xAUmjFFLfhx4UBShPBmGAj4SwtkynB1aPI
jmw0aEYDa1UJT9W9IliHsTspdQTb5QL77zGI0GNuowYY9nEGTTJao37YqqU41vogpM+X04ZqAMH2
ASepGYgbUvb9KdGwW4zEwPVI7xs2gqt1LOKhsYNsC+WwxgsZoMnFvarzcfQXGQwYzmBv1kcupbcw
+Ok+Z5Y34M7iIqHEXn0XQoTnVhMKCOEd5hLgYMA82rwBY20V1q4WJ0+vI6O7nXcLGc59ET5HqvfX
YfjXOx1L/5SrxA0r5q6pZtuC2/iUV7M4xJED2qM5IkWmoOwOPjkXJMkyZ1J/snXKv14CumzrO2SN
qYeUL6r8nvAOngjEsoAHeXvHWVX9CulV7UtvFp6lUb6vgopliGMxA96kAAvzjMszu/z5V8QH2v9m
ZE3WSXntiH95l3ihC7fDdvRW2nXgUFaqyxoUZtK298KVNWLLVA/NG0xA9tUfauBcg+MRmiPvMCtF
BvCoQ72no+nxF0BkUayVkMGGRxb+/rLZ7b7aLwElg2uWqYoDfMYUB/qbAVDOggeLzI/wT6xoHrIc
7m3shzkGTE2dK/VCNL4WhTDUtPz4f8rVKdGWlVRqn5vLzTF891TttxcJEketK6ns59sozFc5/FDX
xuoLqChP9daS9/Sp/XbWLLOMMY1QZOl6h+lubw8895WiXTEB5o39I3LPEqYb7jYXq+5vcHWqp96g
zVgtlWDQPbfSslkhKi3861CJF99Dtf5tGTLLAOfNyZ/xZqBFDoPafXrz5mbcqvgEOijC4zIElWDY
NHMY9+EUXOkkbp+5JcytOGiofoUC67skpehjzLpsFL/WQ2XvymfQNkbtLHFFF4D/XnAX9o5Ja0Ke
jV+FRtrprv+mONZX7zlwFgNNmciG3f+jcZUtzWW7mMMcM/gX49igWFGs+DS/b3eHfODRePDFvnQN
d5RDJ7E/7j4UgJIVogjAKM3xM32yasXYhhhwqg2dtIsOosbx4y10bDEM6DubPaSFnujq9LTOMACT
e9T1SHjYpeGtJlR694ksqJ7fablpmpq4WKSnJwPUCcu344vvLgZPsMCozxcCuQ0GJtVkAhWnP6W0
oU8V2wKofYqdxW+4/6PeMx3Zroo7gzP2xUvLqB5QTPZdmTHrz6zRgUFGHIfLwSQT4jekZx2JSsZK
1xgDszszLCk/ezNZnDaZsiE0l2NLMW9b2OrtOMh83bACFdXMEy4o1Gw0poSkrn3RbdvDd7ssQOkW
JJnnQGknxQwuw5IggVbYyoIYNScxTATPsdcr5a++W2lMbnZmP4nKZG8sox3YrAcE0ajo2p3jrPE5
OfibXDwS+eMg0sP1LfiMqu+ujvBxm3krdvcTqmyWt0s5wSxkJOW0nV5547qtuGWhnzzU0EurW5gV
MF2WjzTbJ4l4MIzZKp3uerKyCbggVSLvWM+1A0PRWeAN+dLRUcZBxUFn14BaXYnnWAYb1og8+IbV
FTw9V/CDZ1rzzxPfyflAeCuqjggfBxy+IbFue+vJ53gKOau4ymn/0ZNUXAHMTTYMUUCgeu+8MiaY
mkhs/zPHCtN+LsIL0CWPAhUfrB6EOyi4pDBcH/dByEhQUToVWlWOW2fyRJe3JyunRKJAoo1VVXp7
ngETKvXTPHDO8TZwf3IRjhQBji4ieI0Aeh8P+z/WRopO7TaulIvrpeesNHu9yBmSHr4yWHTz8gZT
lyuYp7MLcZccVM26KQbmXyo8JOldCA9RGSghOE3GHTDNo3tybFMZbktCoo7vhC/aEFzByYswx/ks
0QZxa5z92+/pasF71VspbU2mm/8Aqh7TPQgu2RHhvGOISC7T72xQ2oNmd2SonaBpgyxx7qBterjM
hVIipZUKMYsWzoU4Km+XPRWeJyifm68S7qEQOhP4UK/HPsBvT75YOqNCZ9etX8LADIqWTO10bP4r
yP9I8WSBxnjxejiFw8zmRU0sJkGi2E7smeQtIpIrHKXGV652EiD+hge5xLcw5vYQgeC1hZWQOUWr
EY48F9G1NFHh7FQrfvQqXXDauTiwX+UXezlXtf9xy5gdKTB5VyU5acTCY8y6Q69y1n+A5o28QdAo
lxpbnL4x/zX6eEuMhcX8DYAaxWAko3fRxSnL6tMAeMFKoKz3jfBK29C1vWWC6whBYHQIkU+Es8ra
Tw3OeFZ6KJH5hpQydChGrfD9Ph6LfGdrgKTEv4PSKXeqrJ6ohXn74mX9zLci0T8nVKb7oDYYmxs6
2ZqJgg5Wl7oivPtUCj+gUqrNU7UTscWxqagoTV3YdqUBMJxF+UjH8J9GInWP8scAHRBA1DdT6h+E
XTeJqtp2ZgipjoFIEgyEAbEp4j4hTrbVRl3/UeLTY4E+P7xsahHhgkjzKzaDvOjdCkmdFcU9tLNF
rfZ1FBFohMcb9hIch/nJx8TuBckBcmaHiOlQqj7FtWu0Kriaz3saqHt+5yTq7pvzI/eSANA1pZhG
2XpSAOuli3lVUrVF3n11GJ5IkmhfSuizuqtMHi19368Ej7ke/sC94QNRcHzpC0JqtOcJ9wMhFAcc
CnWQIFbfnCPqxT7wGWJHQLXl3BvvuUrmJqtCPVOxwhpHJMEe7KBdhNjLB/MKw1YZ3kQQ3fij19vm
I+NJxqZEQPvUdA92fm38B/zFRvwCcGDOrd1YHjoxZljGLYfrosRHPPKMfFqJ9Aqwe76UIbO5xqAO
EKf5+6K5PsudshPfWhcoveYDZwy6WNKma1/U3CNvy4ITiWakf6G+JIz0x/JsACKFnHx2AzVifFzZ
OpomaQJ4dNmgwT0cXwJlD9KuNCIGRZDqtZ5K5xzFoAnkkdLYq++4sPGZw2IGMfh/UoT+u758mBF7
W0j/kiomWquvDKrA8UV66zk4V0xnLR+t1NkyrvvMP6DPkOZuaRkIhHzAu2viNblMd94vD7DtD5hP
e3v+htI0aKxbpLOmEtd7dv+kRlZftCnEhVeZ4dLBAo6XFyGzjY+vh75W/Zg5VjSB0UNZTpaIQHJc
GzRRtZW49i4ZExiWJWDxIDB1/u6Roc8VC+XckEpXMJJakupRsc6bAEJafDR6v5AZ9ZMx8gPwComA
ulh7GSc//63Z57MFEFS9wY5P6NvKsME8SXPvR9xA07gvLKw++t9O74hYZZujckbkgudINC7xrP6v
7JdaFchyuBh3Kg43e7sifSHXmN6hqMVCZBaqUgmwIOfx/GsnOGgg9PhSPmpwAAKy+yFBRP7jEX7v
zg/0PGRVaiQL7RX88LxMQvBZH1E2896fDeu2Ya48U7X33YcFg7rZHwWOV/PeuFT3pR5V4RZOdN2n
4lnHPir3JSEJkAAYomIyHOvQuXNyrhSaoFyvNDUVR0WLNgIF2ve9dadq3uEmlWZBTCK7dxRvuknT
yWma5sJH3TAv/F2qo3hVYL1Eoa+CvqBQGMXQrd9hBLU3XbQfFf2Ozda1BzamAsAn1iKoON3bPAsk
+w4/VieCNWypqvySc4ueeZifnxoHFOjNml+qxtzAckj7Z3T1Xe9d9Gq62ut2CKnM7LJW3U831Q/T
eFr62tj0mJRs8OP+Lom7Whu06YOKjVogw/RZbFy3UUrZoeunimpsZ76cjk110qSg38YI9y2k9vsi
2V1OgxbMZoJVi4gv5xPVeZKXAusHi4c/zDRs8aqNun4KhUA7bpJ5YP2q98agpZ1yJGgdcAkzsTod
GGvh0zTjfX9IfQah7qxyFaIvnoUgKEhOIdqmbX0KcO8XM1HYhkS63JY301/llAlU/Us+IlthgZlF
4QDk1KgaX9WYP+MAdhagUZE06zAFhuHOeztLKeF2MB29mqjnlh0eSTR2kuPCijPzDSGgPEYda53u
8ntT32RrPLr033Cw4zmVI9rZU09sO/cEvW/i573KIfAtveU5RR8mb7DzDlKDA0jvv8DETTq8yQ/m
DOI8Wj9mEl2du6AFhyG3KWZyaDqxqU7d/ZOWF6f6iqaxGyD19h6U+okd41yu3TZbAZU9RNyxzRit
rwYDmF6Zfi4nfxGsxmPEYYnaf4o8q3xLmcLY/0U9V4DmqCB8xi19lgHgLE0vPTTbf13LnQZQY7bU
PUsTyQ5XzhFP/GoUj9v+ebMyE2opH0YrUFtRB6ISUTKotpWGhJCyE0HTn+BjwY+96GbxdZZoPiqz
75ccMZR25c+9wEkSxQ1gqEOQGAXdWSvoatA7j93Bn+i9cf5fMXLCPWGBjhtrkopGK4rf2ReIXBlx
/+3Gs8afUry7gAjYqrk/ezHst8Brm6ElbasKn5aHuXs1/t1I7rn3XXtxEjDqW7qsY62KTTyZLYqM
aej2gU5PCftH80bnYk7QGTcgZdf8xPwNk7g+cbI201o5NvxCzUmcdn0N/a0tIF65sD47c12rXq6B
Csuzd4uSuHHbGcn5J65Mxpf8eimBmcwqw6gPnMNIGv7PGWw7hpd2Lqvq0jwIPr/4TH0ZpsHChx/J
XYXmbpg6K1NDvWvMdnFfS8ySfLBrW51fufaF66O0AOmHkxaWHZqjrZHadQA4q1ZtRqof3MuIHnVh
YwtXvWGLnmBOGi04s/c3aeYOlHw4mQi38sTiAcecYj7Dussi3CAcnGDajq+cTkoF0HvKk/D59+zc
Z5o1uCUvgvSoBEpMYXbimXqu9VznEeEMZZLY7Nrdl049AYyQr2AB23gzaMgoiNYZNYPdO1zEyxaU
gwT/s/g7IILvu7iDE0agmY5qo4yWOYtHCZWte53N1MBczUZqdDbQyXgRz8TrXzL9u13pkicTmqjk
Dm3jQ84YJS7afM9mYgi5T07EHZHIrrB50C3o4oSGWCeKDDBWO8YNFX0acJ+gqJ2V7OfSgHw7h5g2
uFoWMOd7HV4IBnrZFU3/jvgJ1b0rRjLCQHxg7CeIclNRroFeMhbov/93UA1GQzts3RoqGrXT45FN
MRdsDvrZn39WEGfbS7rAm4lT463IbcagzBrC9Fqb3Cza6mw49MjqAHUeiQXaUj9qi5CTk/BAzDLN
IHBotPnt7haIzcQH+PMhLPZZxBPAMAPeapKwvmvZ9p9lku8HycJfoq65F0HXL9IWMcAGfT45VCLl
3lipkFYeE7vBn0n2CX9lJ/9uWI77gTHXvDygI2M7NbZkOZI/HFVO6PxfmTmKp/gafvezsEoVzBTY
UhmBxyU8OH9sT8F6DJK40SBhek8s4iMcrpigufynUdKqIxQqBhRlnE/5QfAQpIvN91eAUymXmCo7
YYH7ozrA8NO1qWXByk9sTq27WBmyihQ79y2WbKTEofAMk9iLCrANzad0BUbpwJ1LBr1v1VoJ3/e7
9g6O55PXAbT544JrOR2HYplXUvIiADezLTunidbwv3rAbwjlv6g/D6Ikx6jiRuMMimWq4UmpCX3g
R0IG8YOMDu4Mxy8E2EgSOtjbk6uZqD9vIsKpp3OIK0LCGqA1YD7TDT6BJucpZzfFvqrr5jWWTOz6
UKRM5NrNmyHDD6rXlqvwqCzAHlLYUc4ad/g6mUWynQfDCmSQupKrjm8VrDy4QGMBb6SOn0yYsIml
tMROq5e9lS+O/icljcpsr0Z7ZYJq3BIsJWrRjQddljWixj7bajI8nqe8vm3VsNcsESzLKOZz1Oz/
AVDNVoB9WwxPcrTK9ToQihZ4uy5sKEqrP3VVUWRGrJiL/Xt9f98Dsshbkw2fFDZ1z3MylHRSPxqP
WkuwL7BDhKnt220eo4gQb2WOdfJbQiMVb88vk+7lCfY6bsNgIF5UYVhzyQBMjGyQvA0XDnhfWg+w
L41nSUjHc3rch65/hVLgKi6Q7KXUCSAlTq4GwBpJRlp2ah+oW5veRuvAAkOZid792jFjFJRZy5KV
aVMdURT7YgMBK3yPRPhPZProi/Sv209GLK/rvwJwZnD0hM89yAFTv5bnnSeeq1pKphTEDyEv0AG4
n9bWX0mtFFF75GMS/rMWTtTwDZgt3KTFPJmNnkegC3Lj+3ydmSkaY1GBQhuc7uuRwPMfkcpVOwRo
Jj3gz4etazPS8aRgiFyHZ5lwwlNXaO3v4UsFoI4MrQ/T8huYDi1u4iLEHDyxr3FKvch6XuctpA2T
Sn+siDrNkbKHj5HoIEo32/7nKrr/vteiFefvLzoouhWzU8VX/FvVPDYo6G05dnxhxW35snF4rBNK
FuIbquEmZxAs8IosRymb6EVsmVybctZxayyGwl4e6inXXzAlPY9tHIsmt59fmgAHY1nmx9L9K3UO
zK/fOn0uQlUJ88EFcDIphYWPZmvLWmT3lLtunmThFlm8NyPMcfnaeqTrYwZ766T2/zuwe2z4kCS1
mLtaL63iNngrb7g5nMFLz5H1xSoVrahS/8n3V8q+H7klb9nC3WOuFbnYOPbDl0oVM52IXFqKq6XT
1vc2r6u6eM83tAzzb/+WLFPZ5/hdKmMrLca22Ot3lkDjFakKSDpMhvhrNNJVnA1sq92bi3rmOZuD
97vKnO12v7FfMlJ5o/rgdC/NjPBJp36IYq/CYEZu3OeYnM2PISnId5xOlYG4VigBbew1ZvTAdYgT
g9jvc1tRKlB3m1Le1SBN/x+t3Q7pgj1+0EqEBKjx9Cubw1O1Zjbx/X5Po6ypYNJK0XL1clikGYJd
WlqHN8c+ugNjF/zWDeIv4BmAH0QZplTLN8ZaZ5dSoaUkKoLmEw7gr912IlxXqpNX2adcFGUQrbFk
5JonOxATd0VXPRdxFDzoQtLMt+Up1h0/QRJ0vIlbhNhV+2kQFAb90ydCPJZ31iRbBjKfxsubuOu0
Ye6E2jBy20oPvMiEVCETGDfUY+Q4pAPAnxAuRHGP3+6Q9PcsOiOX0bTIAMfaca3XpaiDXPUSAFMg
3qvuiCDHN1pFKPBET5nqaX5CRpQGvjrvefAlGXbeY1u6X8xLQvRe64Dm6vFzj5/Nt8do10sq1+RU
7uqy72fX4pEFmnv+2g938pUYV8yOz1jaEhFN/iTW/N38NEQ6DAhTFDM5sVFIC2DVHvzylGVYcmny
KRMnoGqyR0DCkjC/LK+HSpA7M9ppKQDqbg/zD8EoQih0uknMAIwQnu/hLw0zXZemL8MfykzdMZgE
4wTrNZxsBDXlQ7SoJ43cFqSwGMkIBwbeibC5BrGfc6Y3nIG23AOqpDXwlZsR3UzZLo0Hh6BCjALU
ejT9P/Mb5fAJ4e2xSpvQWVMN/lUIqdV9kj0rAYu+zIY5ZYhehjU35WQNEXJlk3XrxA96AvTRU9Ts
ZH3qEg0f5Fq474u4EsaMqRQQJGe8DDBbUpoOWQtuwzblrhS9QrHF9fN+uQIUfa2ln7u8kvKKRoyD
5z78Cw0lmMNVKcVzxjPYn/x+Ac/aQt5SGc/FPF52mEgglNsuQXrHc/MRYXKg7B0DsEzTzKLcLfyl
rVad5MgrLZRlkO0eoWIBvlC8tttV6rS3XXBvkAbbj0K/SVv+grRKYZk+CiLhxrSjBhvBW6V7ou6X
00BJfDkyEaQNXVnrnY5BFteY4wwyJs5QjJtktcYS3Ra64qVao0juQKFzoUEdFQaR4jbpHDztISFn
COZqqmGJxfZ3zl4J2OLKAQ/PvCOBX2Y0bj+pNxoyT39sTyw8wVfbZrPxH6NfifTeibpeYOUqHdN5
3PvD+JJg9wParXcRzd4MuqfP7S1YopQXG3ReZ3FAoZ3v2U5qivF/IcLPivDj2SiJRBYYrB3mo1u6
T5XuRly16+G7w9odvbFIJ1sIy4XwRIrex/7e0ZVa1fUDyJHx+sikvGvQtCxAfSBdkEKAvdgwXUpJ
uGmBSCP/oDuFdz6xBoVxFCLAQ889TEc8+XePgZ/H+CwegE/R0SfI+IQc9QUMl04prFjAZceji07V
UNNMOLY9Dq5ZKLnFEstn1qKrgOCKAFM8NUsa5GrJ5+TAcI5P4ZP1/UGzIIYEcgapEFKgUgmC7eiD
g3Es4l0PcCP61SXZyuLnx7prWqnJo3eD9VKedPLP1TT2DkqsFn9yocgiLX+bDH0G1Zo9MCSOqxla
e0GVtiwZuMRI/EEQ/uxvxsdqGgAbpPC8v0t9QJvRniAN4A32gI/y4phcEZcqqWdKQefoCsVzwSl2
mIi9/ZaTMLBpo5ZhMx4YWF4B0J1/BzJ7j0J7I5ZH5HuI6Tc6y6T9LHAt0xIYCph+B1VouC/02x7v
jKzhMmHmMjM01NRSChCLGoAS4HjNCRvNsjmRJv645DPNzIeA8moifBBBBPRSiwpaFR5YOtbIRlya
+DOqqqp8AUQWKxvu8terxa3+nW0VUED1L0q8Wv1N/6UgRFmdyJV2N2yibFnZqvdSgPIPg6EyLb/e
lZ/vytkXKJ1uWl6o/f6xeGBk4FLVHsBIRYzSkn+ph9Lj4+1OwrQ1r/xEHD6jzMVg3btvrCrw3Sfa
xLxTVV905XyjHojhBnMl9ryb6CfCJiAZZYzy8XrBDVCujm3Da5tyQ6bDvREux8jV7cHqJlc47+ns
2v37iF1ExR45QGzWVdUAYSMGFvqO+QgS+uIDpJsZCkMhU/5eWj8RJCGQKQWIKUZWCIvwjP4OP98i
w5ye5p3TvIPNTOqyJXtShSEVQdAMurJ0ZGn6VdPzJQzgQMe4a2TRXXt6P9lGVoGv3oVLH06aKkao
H8i3Qqm2iQZawuLyVluz0JP2O0PZd+GXx4x6ncAl+uZIn2SRvf9dqRJAlIJCQSmwNq58lkrNhKeA
gCYSGje1nq0Hpcw3eCV/0auvpS9SEnmLr6q7ryJrezDaL0FFZuH/j7jjfW4APSL6Gu0a332MFKqn
ZUVJSfDpj5hBdJjpJzg0GIQHkQGbbpqnwN+ST27FSFFXcrLj4109Z2MTTLT2Dqy2lbtApfetADav
KzVemaKL9ZdfpuQISVIbsoq1jLF9vhN5upwqBy3uWDWC5XAHf1dUAFchKwrnM5JEu0Cs0Nkadnav
zxfQg4Id2SzVwTncJ6Hto7PsEazjpLhPGVlnCcUdVy1Zfu6wOzgK1H1aD3zSakAT182MkmS19gEA
+sa9jkJ3d+v+W4yHna6OGJEtwSUhgB1gyfq6RCO2hLtUU/iRRfme8MxeSc4FVMicJfLerHiQw20v
2psgEyRIXPA2KzKTeEsCDDldmdmhHisp/YcAUFlDSNi8sF0xBBnC97E9FBLFrLJrHpOp24GmJDPb
Iw+kN2PVNlNT55V3krNvhrliH4AwgtMhhs47/Y2D9ByFC8voiHZ8kY6M3tO1wkL28AhAFcS4Em28
O7FpTWypUNyi2Ee4JsCgqchchqZSFml/rAO7KSd4NuIX5b4QeZoLR0sN5E/6tyuYtZ2WSGgofaNm
K3++rWY5wuDy3FB2r5UGrPqEdo5UipYWjNYIaIvJuThvLQCluGvIeGBK9kNPh/ZY1R1Pw1xprfFm
Ut+2hFrTabjMhjHk/ACL2VxRFyF61aDJvNmxbvRcOVyoLghfrlInVB46Qx/OGhWv9or+uNe8PcAq
wf1FGOT+Kz9FcgeIiPAjXkLU/8dzfdurPs2xx0ojVQjJJtU+CD3YcccZMvt1ARIyyflitaogIDoL
Xaj42+u8jKtVH3jn/TjqNYJAHXJPXSzBRV0egn2bqdDwIqh2b25CuIVF9d+2kjVtdrad8Ch3aJw0
v1iqc/CI9aLzaQa3WkdtNaYXOvoePKxCOmEWvHmJc14AlnqopKaoKzfIDVfwPsrqE7YALY5piwd4
Guu9mLCn6XBfvMn1ChonJqEmcZiOu+TKKZ/hF+KFrzZS5eOhxvLQ7Na1l6uYwViMN2aUeSPH6rGl
aYhTip/bXTzW2+yAtWZCZQj9+w3LX4iFcQJor8EOuf96ZoDbt7vjLesV1zzZfX5SkgvpfiakQxK/
EA5JuuFm2OBQ58kJtc9NTE6M3HC8H8Pjs9zKTZ1fx7B9dlwjeymi9Pn4vRSVinnlZIG236Tw6LnZ
yYrQy3orILgsX31woU2SQxnGy+W6y5SaoQtwSgkpxYS6XBewRovByyafD+1ifsOzGEZVsIDrg0pR
eIcRQErRSIWDfEZiaHo7/b7BZivtAnsKf4bQnlHRSeWcr4r72bsSLT9cPFBOt1zBvZ/qgaolRpme
+0fgZbzUQjjN9ADebq/J/5CfBlVPZGhHHaC0YSafNOGpX+NSGDUv+Qn2ExB5f3eaGwOpKzN+oHAS
VuaooLkS2XWVyTA9ndELSkT3UygXZ74lGeRpkmiB2BHz5/uR9Wa+yp++MoiZom9quWZ7y+hqkBhC
FCooYNKcJ+c5Tw4nwx9Jp9rglpC1ifHmHTdFuZBqstMlm562t560ZBeLMo830bEvTGDS+WLPwk0h
iIY7z5ZtDlkQoR3cCiqCOVEzD16lZ8NHpB0H8pgWVQo1p8XVrk/JSM1ezWmt7rw310URtIDQXZn+
gw7HUUPClA/GoCmAzFdPTbnt+812tBNpxwhCplakwqevbgxFVqwqzURgwqom6U1uh4tmQZIjNwPd
5IRDp/V3VGA90UXDEv27MP7AVUqMDzX/of+G7yYexf/pss3HP+YWfc5WVzJcAmdO7WNOEXIkR4gp
qQBM1YJ5PylE/QnHMYNFC64RUfPZhUUHN1501BHz5peh4aH8WQHP3BnF2Bl2Cuk5nhwkbUICqpWk
wQxLKPKG0xiaDR3VetYsmfFPS99cGGeeI9EfkxkwwtOkRINMoC4jBKfGd6e/47s5VnrT/T9or+vL
EJ/koMz2kylP++XS/7OZanfGvoPncNg1nw7rbIJ0VfDgKdlGwYlc46zoqGpv7GO5LP+NCRoWwqYz
eGZ4BHJDWT8UM5wHBzyEo3uVso5GLy2JHd8coJkqWV5WlI9cNH9j3XOZqJuBnA2/GWWVT57j2Aiz
MpwQAJfIYeraXR3PARZl24CcaPRNECtvyNMimAFzIxAcfS1kubKZuX8JaMVUeo946XDfhfN1N/1G
d9ERcbMKvFbLRjk5REV9WhhVG9L9vwPYOEpsq60yU1JcGnIlpB5/d6Klz9wvyry8mZOqttZy8sqr
0gOJ0/ciRYOlU9SQU6Cu+BTjSjgAUY5a/tqeepCg9J78iYp26gD/xQJKBoooYu9asN3QA7uR5i5C
GbWFqKEKZ3slCT82M+24uYbxljfWULdnaSj16RDjcYSRSf6aIImhZHi2bAHc5RNJz54sGTt0KDi1
NVB1ubVPo76+pZPWYg89KUiac/w31jBbZihbyUXzTTPU/u2bg5aC6VAyZqa3qpeBziYlAP2NYfq4
XBeqsv6UHXdR6y1M7Ad2gWutUJWBM/DB0e0Rx/cDZa4Oid22SQZHNey9dq0N19RvYdSoDqoGuEY+
kJb+TdqS3KBRfGoojI1WWjz3jGyNlm0lkIrtm98P0NatKnJfrJ2LDaJUo+LEaFm4uYfEDNS10lnv
gKT8SnDBCE4oT9DyqzNtBhE/h/Gi1ESWBa+am5NvIHQ6R9Bjp9N56+UDNsRLVYsSD/fVeeiA44zX
cjRXtZMgCrDHmWpdrKrYCG5h+iYD872nxa5qY7e5PmdZi/9Se1vzewnjPeDxJ8NRwD6Aqq1/6CkT
415zJprz4su5i5SRl/UG69GetIuFYKsLAa/28GAka1NHoBP+fDFKN3XEyD57EJrTx6nNbPd3f7lG
TRPeXHn+UEzu7Qbw8b9/dgiZL/DhINtRS5iNtBZo+eG8ylIygPRAQCexbZ7dmq5QN5u6dagsQ9ur
p3WS1S4uIi5u+uHYlqiaeSqeUps4nS2H5bt8hYqJ6nlmEOp9k0k/ffoU+PHGKrhKkovxyxFMQfhL
fAppgquYSBd4uIthussSTdhlt2vzvT2b4KXNql9CaAD1QSEsw+/cb3P4zZU5tTMVsrnDAf16yzY9
8RopyKFl2NJvG26TRbVTElzNj8CXJyiUp+2ecz5V8DgDy6JIfqiyZPyPXJHAhGzakliMgAR/n2N2
/AKmKNLVbsGl5ecT2nHifpZLrfN6Ho+VGX3wnr6dYk/tsfdotPAfUpjvsC6CgzIx9UO0/o5oRPC9
EXhXJ0iAqYQkH3ZRp7DtfqsoYtVup/ovZ9I6cPkMJhAZewP0mqm7UNG7rkfiJwWDI4sfFDhuFH2G
3h1Jhtm57P9nJzK+HgMgKHEDchEkFTVNKK6n/5MteHfQF6MPPCjbFuE7PlTnpfirin6JRyM6nHCU
/4ZPB2WT7yUgVd46srq3j3NsXgYCHF0hmMxmotA1oCZyDRTf2e4l+TUT6HvgNiQUABVRyjh/rQW9
bpP/5M/6hYe/bNlJob26xzPR5J1Nk83/0Fl8S8VPSTbrWDDTQMw+ng8ze3rM4NuKXMhIP0RCgac8
F9SVXFybwh060Jy9jg9p/7/s7fDYfguw99XUo9nvrlLfYpvzsaUF5KTVcza9bjcjy+GlXQQgb49w
UBBULKtq8DiadeusZ8oaS89Kvo4ZvQUZshWL1E4eC00GkzI3F3WuupECCeet28KGMYXU8svXrU/M
eEIrUktuTjiLQW+HXMnrxks1FJzgJIfqByHi8D1gjKlvwt38OK3FLA7eVyNQFFlGKjxV2+EBBTut
cmhpG2zPOjoZSBsl+nDgsGzM8lXJnFOiEB0TnY3LlwOAm5dAgYxddb2gll71wbIvaoDLpn0ZJBB8
iQyJCPZKzgwGkktOOM4VavieV6GY42gZBYFeB2Ivs4f0U9Ekaw5h+160Ppu6YIb2De56QY+g1/Jh
7D98fLDTI5PJMVOOhz8rKBj9wb/SjWxGO8K0Wr8ZOk63bjZc1+aDBaPhYl6ZbKoQXlsbhvqdviaX
FZh6SLpG6yrTGBCWsbO+RbehJUiKHPb51NCmV3uqbFAFNXfd9rLSfAML5zOtIDXKfvRd3icA+ss6
0L7ji7AZYrOLho3PCjE2kobvaYAvVX4xfstJTFIv6E/mBb1d+iJPAMK5CJi3sydyU7dH2DkKKhVo
lImQYqLBxL58WrXXDce3t9JAWX6nf5pGN7c9Qbumlh+c9Fv8/eOuJFWRbwAZCpbojILJcs/fyADz
MfcFmPyKkgertWSwEjT9+Q1TPkpEpWvEJD5oz0ZDhtk3PNYa8Y2R0TWJpRtgSqsvAvRbPHv4F6di
IB6wd4YdPG4nMhUXW5DdibZ/2wRp2sa0ijjGGSfTluijyYk9GohCAfdUcWgXAy0mXzzVhC7MYFs1
u26s7NRw2XnUVeweARtVHuyJmH5ZkiIJkRLrHx/IgE98QmfgHbHRYsSB6UK3YyLUb0fpGmDZYdd2
sm7qDGqlvMG5eN1j7JJI+qPYXnmwheEq9gSN/01BNdiVKJAmtBtGzCX74QS6TdymQGUC3xYHxE9b
IeV5S2t4PZ5Wke1QkrOqnctvUsAlWsP+Vzx8AMizNZN9/3FwiY05WWdId6E/3Rk5IVy5rrmv5Wgc
hWQDGn2r8FoXLuWJZ9TakAV0hOhK0vN59TVtDCpKOHyX275QzMeXobPwydN/nF3fRBY2AzTQWp3N
STfZx60r6rs0OfBNECr0TiXd9fV3LAdSp9ITnRFOzyFWHd49xVrxUvLiWWYt/8BdcX6hWuX9xq1P
X6Bgkwjb3e0zArj+pzZE3iPdmA0Gt2DT8/ga+OOW7xnB6tCSAPet8Ldpw/UL4xpQgiSlZWY743nD
R1Yg8SF1TvNARDRvm6qkCEMMtCp2n7xzyBXc6doeHQuz/QU9S+Fjtv6EyPe4CDTGddnTcSCCcAD1
l30NWwiRtcyMzYtLaqsSGOqrPlSZz2o0Mgp/prmEnn1loZMgtCHl6wT00kNHt4hPCTISJRSIPlmW
38pMlxxWh5swZ7Ur1+gWxn64wdcVeGCud3X6QVfk8cMRorPLI04i3om+zTAD2rzl+BXz9V+qvPpC
HdLuDmCiH0//MYFdM1xVgHY6/DOrBMOGf7qvNk3GVFHTjz44Gl5HInL/TOGbGnc8Nhgem8yCKbHY
m2WrtJkonLNFv5HUELkHXkVoTL3PqKVyCbwwKj3J3zsN1Js3hJAVx0IJMI4oHECkIos9jvmZgiAD
mNFzgetlFCxzEyTQRy4U4ISifZ45LfVLl9IbN5EB3crGGtDjpQTRUtDHJuZVJCduIOyyFkdxJbQ9
YHvJvtuw1P115EQmis3VesPtFxgz44rVfOS4TKPqjYoCti7mjOBHPcbt1HzF4Mn08stwcVGItCBs
3vP1VW3aLZzh4Usj7/s5cTqnvL/tBiFMYoDvgDCHdUFSvlAS1E8qaHpfN69QvoaSWdwQituEN8qy
sDghjvaxaeeivEdAYZBxol0Q0K2YTK+PwOS202bdPVXLsVjqtBf7+rs+sS4vG+wEuIfeJ+JsemzJ
HUS9pFGY+FgNDnGr0Jvty4Ac0YWpF3bDUKoHJhCnRX5RutuKthrn/B4W55X0gDcKUb4Bzq76m39c
07EBPetA31s4423keniqaATzhbM9pTZwesuONoPZfmonrcDpllYXycewvUQlR/Vd4XrJlMHtIO+F
MCt4/CMq/b8yp+U5pPAOCFukDPrKhlM4v6brKqQ9psjKuylj5qXC9evWuU/8kiMjb0QYkzoNqZhP
1CV+DGBSbgIPpbrqOpybhEj23WlxQBD43LZlsNFplKuhYYEBrv25SkQwh7vnLNsnyHx+eQ3VckRN
vEuh0q1XOiiyiCOZ97UgbMuKTJ72dOO5x2RXXmb6gJJiOoReQQ6rRH8rTPe5/VF59T78SSlDuaFW
ahWN09B2pyJyV8V59e5HZ6PIT9S+zskoOI9kt248UTfApUTgJNqSSVyJIIM4cW2deJ0zqxL4YVsl
gw0fBFXoJH1DsRNNnSmScMcyttaIbkS95O2CEWCxHORwRLZHkzG7afuFDC6LUt1sFwwtP8XktQSP
OaE0KYSgk9VxG3xyY2DIBCtwA8pv9rp86sYVRA66/BDi8hNBQMCgG6WKg4PWpVPAdlf4csBIs77h
8ANi0YvbvUbFC9KZyJqUX8a6Bh45d1yVewpZ2+eHgLHnT7VzjqNUCVuRPolsngBEUMPYJEkWEJqU
0ORR5zl2IfHCwkicF9gKIWGMbusxCNftkH4ionNJL94Rnl1/7MlSKPsHAHIZuADEfQLT/riz1+9j
M8lWPrDYL5hKUtDck542MrwJtbKbj17Djdven54TJMaBXX3rgAdtuDedpHnb3FWb2sR8SLPPYsoL
49U2JOusmEp8gYij7MmYIFnSaEOMuF08R9btZxyBuNxZ/Hp+QpzBsDmvHr8vKW6BRs7+4uRY5aFa
YYKPoFFJPqVPbuv3QSyUoL78Im28fDZRf2DHT0QZuouDoQso5wq+x1F3HvqlhszP27V+ttBJQh2y
BTUtssydZWqLc5PMM/Sdl9XuQSbv4WbykL2Q1KWE3IsG4XfeVOuSq1Iye8xcMcMY47rDDqfh1EBa
4+/O6bObHG/E4b4+Th4nFcjWLZAKY8xBVqSJ3n+Xtx6rz8nNjsV36plK6gB0vuhcY2TSsvbkZT0G
LX6+F26Objek9n+CA9yDORXZQQTtr9l3TBgQslHYCKCZ2DppoKlfyXImol2yGYYg5UsMnJxqCL0W
zAn7IXKFnQCKgaCnaf5Iy95lyRRgdLkbQWURWG3qFqa2dBN9MduFTyqx6o3QESgZaa8bddEqmsXX
9J1WowAE9fkKnJbeOm67huXo7hpmcC8884JsgWZkJ0q0w8fE1WcEsq8EGvdf+AvukeFPxbyUscEw
eNkpFaOza4vIHuWE0lhU5vYYCdiuNBqMedvN8LsqueAzOLbGtid8cpRcZ8XFFG5plCgOTtaid+fO
syS5t/3vqsXW8ZTtK2B7WojUeekg/3GY3+sFfThxuT+Bm61kbqEmAbBFhIw+c1VI5zWmH+PUOo4d
Z0/QswOdsmgsEoDNzVHxFQc+hIUy4QcXI75STHkH6ZuhGSu3q9TdOBMA2j3e/wOaF1Er4OWErWTR
dmsHPfT40y92peIoBZCJU/aGmxBfECFxoqpVj13eZACRg/9CEcVi7irPbMmimSbsocomh3IdJ3Bn
yx8ql9BGPBn+BFn7CkVNHjrlR9H8gxdSSSiz8DRf0e+m4eZ0nXxxQu0yWXGwepkInSuJ1bDridep
W/gI2R6f1n5SLpBKAFhOthTa1LFltZhythaCIYbFuBg6vrDuOO4f745Shb16CHI9SO3VvwfpeXGy
dm+CK3QYJh9Nknt1eiS9OSNQXkmEwsfvAYbu4BOwuKD1yvFHj5GZS2FR3F4nc4DKh3O6xF+yaogv
Pa4/UNaBfq/Nikd02151bxF+5m9tJMAZRC+6tI4YLbOIAdxVt6AQuQT7xcLt70+EC8QUF9iCLyVM
cVPRRwV5K241S0zzIkGZ1g+h8kW4PIPWjUTtdWG3Q4lpe19KZ8oQ0QFaVls2I2axwRS4zxeneAYN
BB5DyODKkKfj+FRk7IuDyZr+b9MVMfsI36lUuT0ZUFvz2uZV3VsYuOjE+8iXmEx5izcetbuIsqPv
Gi/AlMFNpEdQKw2lIcpLqqhQIu7zmHFN1ofb9zKS1EYBU4rxtSlQy39PBmtsEkclhDHNgV9vsn0L
zGsblIGFeoUV38YqnYykxXq7pjDVlJBvAiIT8JH2JJCGOHMGhY0rO/RRSE4k2ZuHJmOXpYpHYibP
UU2/2fMmfocVz+oJzislbeqsf7y6Ox4TjypvJlMn3mgSYBdIDPXVGuoKREkzq65YE2TYg/6hz9qw
uJ9bY1/T7ya8/J+XznZ1J8e6xvyi5gtEnI1zVhLegqgS9HQjFhZmeen5BuosICOOPz4nPoqa3+f7
jEXAyfdOdK691kHnVsQjXvXgjcNQgLC7R/9gBe+1xboXhdYyoGE2Igt4VaVKS4EavmAzHLVNqlEX
EUd83fv836snJs0+F0dJ3p09aUk/aVVqEQo3P91yBRcADz6k6zpPBrFeJNT6hV4AhuFWQ1h5egnl
EIuAYCtgM0yjbssoAPnhKa9FY21YPWjBeqMum0+eL0PxLORrKwW3/GbPwaLMvLtUJtKEi+4JMplm
mZyVOElpc3BbzX74wpvUxLVb+3kjwdsUiBtknW1lEiUdzPSWznpas80yhYqFx/RWkr/pVYD7lssV
AcHseZ6NHnVgkgMZ6N+YWZXiZe6GhGjxWEeg1WZurapj83wytd4iTdN3hSkqUgffMUsIkFaZv0Eu
x1dHtFv+6GgoUYAPuoTRykZfS+iHxQtv/nfdsPFedNawoREI3RNM78y5wMvjXJxorHjKhCnklXlD
PUnqyzcd5Z6V4l34HHlZ8ILEGJJNUmgsJJbS00FJPOTBPTJQCInbRHm69NQTrpts2MMjrryOkoEx
7qOUz68Ah2UW0JCkAZRzIvxpQ4PHSiHRJo3eZ3ZlzUL2Gluf+STmgxcA8W57WrYdsSCukGN/uWWJ
4C6ISx71fICmzsARkSJQYufXRDVGOVp8D3l6uU3Wv91uJ2ku4TDqgvAWVdXfW90dRTa9FQGVucXb
CBYG19UoQ3973KqVmGUu8vvpda94G36Oy4wrOwa/YQaKugRS44h0VRhf+nwxXbTPC2KJbkal6cUf
g+to6fSM2YxlkOoKap+cgqu28hK2h3JBQ2MoJDzSxRkOhP7ZrPfDdyDqFKcYIs8TMyaaJgB1D41G
5IFpaEjLHws6J7KX9wUb6SjmJdRx/FdQKknmfPKoIgk96m7ljzsOWzDBCyBUBwpldIJcrNoRD7CQ
kcT6+rI381032amx5sC5JHq+pPLPKpONMAfEH96fNAlLU4u8NL7x7uZvfBSQNSQ6Ot5QcpWjIemA
bW3LiZd5Isi5KfHb77442BpUlf7WB7lqOsH0y2SxxBg7Mzeq7KDpcAEkeyEjSpocBjjFhO3taSXH
c79a9r64QMux4/HNVzJfqD/qM0OWH/Vk/c0vmGx7xMnYQLROoISNiVuAukWorG1i8XQLf4G8f7WG
ske1mG+7z+eDbW2Lt0KMQxjCvnNIX+WnfzNAmvwOEfFBnfwekxDD4qGEjgGO7Pwd0TcEFvl1f1K6
rTPXCc6HOdfhPGJH5nT9PWihKIj3/9zIyWwSkRwxB/igVJlK/r3yW8DU9Lea1ZIHLwKYyZA49sgy
jipUYACvTcUU/EiXZJbD/eGdv2XniKSb60tZqruMESNHb+DDc1zaeI2nJcwFA1NIyWEpaL2nSWKv
QVIMqJcJu2yhvH66ahO+gtI4nUOeVyixcLC0X5+x9ju+kyBmPsok6GTkuKzHQIPP6ntHFBpZNY+t
TqyoFxAxFbmbRA1XXPCH+C1ftTpCxNrnEv7gPuvV/T9RMhFnvPiDX3x8HAjMPKi2deotHHIKMPmu
WN9YOl7dNz1ZVPdnYXg3hW3mpGX9JJ5Hfoa5KZsq/0iuqDcP9wEOcvrr1hOBlroQbjHnT6j0q7NB
bJzA2JqGjqA6ny3wMVpa7sUPehtgMR2uHGPZeMhxXjmVPPZHfSC/H1i7p9jOhyckdzpHqVt1PQ/7
mUL9z/KsUFcIYwX0c5UagmQB6DA6knYWd2koIYPOUXe+7gxNieq4lqffsqpwBLJP5htbRdDzq5Pu
BOemBdUfMEuMI+hp8NYuONb7guzS6RxigkaFcUVq6BMrpUPZapTKOsEEb78ILHdBuwGVKf956Wa7
Zm7ZQoIVU5LZLbKwIpJDVC3RSYmnjQKx5E4gnc71P91fn1M4R9hF34MazUP/RZrMmsxR3GYfaJG6
dvsIt265ZL/vZQQsX+BP3acesHSwR1XVuYvZkfo6/MOWPYDviF1XSBIh3jqtyNOPMdYyt+6pCKM9
NianZ163eWuoI8xD+PcQLYHaPjWbVx9RhYIOY/d6UnHhffTayD4avF4MKkPSOr5KATtsZCnadQ6r
REjRG8j/sR8CVQNnKKs76wiVYgkNqSXPH5UIRnUgsAoX+T2qTLoKz/vQeM8OZw0okv79A2MWySR+
r/NeAWc/pRFD0owZ9hCgrfOUk4lfysE3A9+rIIP+7DHx6GVSf59CX092wRiBOUAu4i64+Za+1X+x
GzvdQdRpX94Cyp/TCdCzOHg1yuEZz+xyA2FYjFjvNEa6wMWaJ+ndYqLOxfHHBx7T3SI6pGr6ni5y
dbxBbhiD85pHEs03aLqagaDl8UG8kTNc+7ue73rhvnwjhytKKPItD0ZVrLtifNvqzbACj5QScvai
k8NidG4IaVqoBbx4YbWS5kNYipQdwof9yi2AUCOnU/SsOHeI9xtVld3A9w/ZO0t1i09nCqWbU+H3
ltW4duXOJJtLI4jhZKwvolVr3+xDS6nY8zeBI80Lc3yHitB79npK1H+QLYAz8J/Uwy+30/jSsfZG
5fIflp+oJ4EEVAlaJYlviy5jUqbGpCn8wUjdWCRxLR/Pv0stY2m4DE5uwUqjwCaRafWYqbsblksy
66JL54E9ZGPmkBP8vbP5d95BdfYChsUxh3ppr/qLCAjVWJN45eilMr4Y6Sc5HOzE0EWUCSvNT29l
XWmnYXCqh7ZiMpccYWaEPyQJnO7hBaMKAYXIaHNrPrd9qIWCr/KWn8E43OcwFL7qvSd9WVAYbhL8
ZLi1wwsPxYHpffsmR9k8+jYQoygcI1uxwvshD3kOzGG/xBxO4hZcIjja0hoOE7zFMBG0qYOFvH1i
ePsWuqrJ80cXcfsohKjhO4VZQGKMw1R55DA5y5hN3kjrzgNh+3HsuhDT9Qj3pEkgxEO/wmJGc+Hl
DI2cDmPVRvbmFCRKTnfvfJy1KispDq+pgwo5rCw4i5X/4GjIh3ZBpbd/S5lBs95vttVieMvH+V0m
PB3q1jhR53vyXQHnvpGuMfU30hAGWt3r3LYfUcFyPhPI5kzCbrb0j1XYt4Vuk7JzoTXoCy50qs5R
R+lBkjtdNmP96g788wb4KF48LJRyB+8JbvNxrUmciPm2+70gEH99NjbKFsCsmmfXDKfLy3VU/ijF
FSadkpkQBthFdkbtk8yHJV8IIS1ild2kzfRwseJ4ZVP7+Us3Ob6vOIaH3C7ZL1bhqickoapWnXMJ
EN2OpeMLR6lgvtQBV1LMeT+05WnTVAuaI2f+I2snEjP9dny4inZeXH6SogHst/tFOlPFD/x2ceNF
DNQmcFdA/XAlH89h/nj6281A5avl+gUcJiEz7NH1UuskTh9PxvMMD5v1SZMDDL2h1tA91ndmcrmC
yJ3nmkh9JwgHNpuRXSCIJf3Y7NL+Qvf6fW54dDAJ0uQ4GsV4c8nXXoSVS2t+D2DtgDMyyuDNJvp5
wFVY3Hxl9TF/yv/8jj58t7pl8lJO7vu41Ea8AUftisW1D/+PmiG7UTmM1Jp5d7Kd2PGneLPOsIWs
uchx0RGi7C+xuUU7z8406Y6oV/DJicG4i+ocYObg2iNYcm+TybnqZqdZxR+rZEN4Rd85r2gquJ61
1aYWW1rZk3IR6l9EZq7waZXTN7hFhdgGePFaO3EBf/69RTnVhHpQQvl274n9rz6dcJ8tiDIKrr1v
XkAzCjOlML0yofYoN/ByZkuJk3rNK3OJ9JtkOIDPSioZlf+jksFey/NaK8YwdwIqsYGJxlo1FJCw
gQS2rQmh3M9nJFndQs1YPVQbcVtULemHuKxehz6onhPKWJ7Hccs7RYU9ZSZuXj9wfWkLdNsVHn07
H9D4TT9s5LMuSYSFq/RuZbzF8txS6G8e5QpIfjE+hajgDVBoqeJ3L7o1y9DoBlXSA2T6uryE0oSB
9Qgk7vDdlR03hltpIyMrE1liivWEJCNDJ65SsBv5okgWi1zFNPrnf2Lo5uaEP1/u68sC0W8sKZfe
TsShINaqBXQU2pf1cm3xSqvMDDW3gcTplFAJtBhu0keL1Cj7OwAOTJ4sKd0Ps39njBheiMttO87A
QOh4fexLZLsZfqijaYdvpegYR0Z4EV4d9cI4iImdDOf//cYH4gKB3ZrF1rz+sWOMO4JtScd3HOhr
6U3DlRICi/1bCuE9IT4ypSCK3rBLxeQaIDiYFFja6+H7PMo1ZtNFuX4i5WO/Pr4y4c5v4EhWnwoD
l3ZyyuUfOKAOn5NSJlPBSYMaAuSo6A8Bxink6hNpLQ2JQepBwhZQ2DBk2YMq6ElRZJ0UVNq/s6Nf
2VZbSOwlv5AVJQ3McTKajSwOrbL7QSaoMff7PMnHPZjtnNZURudgVd7S6OkdOSs+HShzkRaBbPkK
i3qlYeQNICrHmFhFSRw5Z2f7NaLGmvJAfHxzEoAjJOXEoZTreNO4iigfoNw7wwrFt5+zudlm6Fz3
vKAc5b9g9/qy0IiaW6Efyf7tFbG1Qdz5atA+vf0QnzYyd63YcCa4RsAwXnr2QgUIn+eJNjigfD6F
vRUisGCZaCIDvv7P91JjlowOzcQYOd1egID49kvhi+mHy71s7Zzf/0otWqCgJJB5OQ7SC0RDEKbC
t5obr8zQ2YXEve5GcpGavPnSoZNQMWnp08J1DudAcDoKPc0qm9iEzSdzveQ6XFP7XhDJM4g135tv
fz2JFwREXyDB3c4TlsEymc0q3NeykLEwGBLvQw4xvy2O79WwdQbsUBQw5nYv0+0jsW0LDpyCbP5x
CGOwx2MUO0s0uPInO05umD/khIyfWhjQ0KGHJ46I7jShUpwzo2o2RGdNnX1UhtnlrNqckym7RcLH
3zx1goYFZ3Whs0p5kAmffWDi5Rd0W35MpQsUpZnttRsHDHbcyEWotHwsg1c7Tot5l3YESkDb5joj
/AXJR+IbqLALaCDR+IQ2lVMhAgrNce4gBBMqOkAQ9ym0jeWaMGDoaYH7PebKa5GNslFgHZRSqDbA
wG4ss7P0kntI89qM+utMmEsUhmN0rRJRYyQlwP4D12ux7DcPMpu76n2bdvzQdhRnzbvfXmgSHOGG
zMZ6BTy8e44Og7jGnFfsVRT5Pc9Z/x5ddAzu3VvL38RcvK9E8wKsbg7/ZmHhcAN6LCE5sg7WOevC
w/N7sClzZFd67nVz75xPhI0XquBfNcGALUWT55HtikFyFYkBYwgGCwNLXvoH8GIqVjASPRd9Onld
1pQHYnlLYvc7Zdm8aPCjNiIGgn8okF5wbxoXKcalgasNvqA+6N2EHq+dwqKSHu7fHz8tF8W+zSkN
/SccOiQUqJtXpt21DIMRwvTMAhyGfWjruaX+sEhuUjzPAU2QmDCObNm5jagbmFNlHzdht0hcfI3/
s9RPTOOJ0j8EemsydEMdh2Hi67PABji/9+s4ZByMp5EHHriUmVZdJD1GGM8FT37AXA1qbeRPHrII
6AyO/YcvG+RVaXBNs5qP7547q4U60lj7APh8F2JOUx9sGNJ5pM3cpBqMZpmOlewbUYRl9wsZA6bi
C5dghT7NUHXko0S3hRLFcTggojbD/xO5N/TvKY8EvWK+4u2s2qVXJJieCFSjvZ86UDrcVuMachfY
ofjzAdtDzGQrmkJs/Aehe5+GONtFnkISIGmx+3M66wnPQ8vxBNA5/lmraDESj7tKmIu3c008cDz7
S62Ej7B8AyU6SgV/3FdAPNw7qmDOi067i/L1i+YAkSO8T4c+mx4/GN5bSpxWwyPDFc0nerEbO39e
F1Khd+x8U+0GnnIDdShecCvnTA3GPbaleisaXj4y3Bc8WvrevAJtXc9OqVEKlCD5kDr9+1qRLMiL
dsg/83oYYuBxTPzBR79HzRKUKoHm/i0vFncPyHJ17ZymmyKiuAwnEQwuLUEhDH9XnjIuyMt7+ndS
jme4hsLbd+u4E/O03WEC9/ruUAtz/arkYh36M5Og/277y7UWr0tRZuZU7tB6Mjp2ia/t0UeUFbg4
2XPe5qAqqIuSXUbbyH4SjKpzC6bi+zTmq2KM+3wQqtGALo5ip4KkBZ77KRVCobRmpd/0Cs66EzM2
x/Zh9xSV6RbXFdzMTPvw7g4E0o2lK1iloISvyEAcir4N5LjldTTKYR9tiiW9mxmqcZEA+QVZcMsT
tbOuS2Vwn4tponp/zwQKl7+NbhEevyk/aXEXEbeTt0Pf2q5jUkxpUFPd0hKGtBdU7xghA6jN8hak
3smHWX/GQpvipKja71F0r5VMgjL7HDwwYKOVMnjPX9NmcbdLXCA+uKwe26xkLmn2MxzuEPREE8X2
c4V6lgOYdJdLEk/JdW36qUW78PPAGjeVzyFDIe373ecNeLsBAwm/Ltb3wvdc1KJzLivcAFNjPI/j
OkTqLbTCds/qFQaXoPMqDMMBai0ttA6fyy6EgOGezC1BAUqiEX7kGjtRCzzrttXHnlD2UFdXDzV1
IiQ6hSfYRrQvqrjwidvCnoWkiCSjmoR/i+5nhuA+qJfeiWQ9rRbK1cQ3aT2g4Sag5zncnWjSeANP
ubpN1MWIuCjhoTsMxj8aR+H+tH3LJgM/MsV4n4TZ9VvgoUzVwvBh9oLArij4+lvcLF/+ZbhS4uQV
unjB8fvyC9DWgotzSIuINHzWQuR5FVCYuw2LEMXn4gTdesVmIx0B6te2GGOqC1ayoN5fV6Z0U4vG
wIGhgVzv2Md0VarFx9i4wzCx2yrXa3wLWv1xz5HbaBWGmvDkhATcvguPXUdumksWbw+PqZL5PncJ
/Blyt1T33GIbldPAaRHW+LEAxxTMP/8v+D3GOohUMPD4NdoPjR3l+NdYtjOXWQYFwjWhClrY8TML
ttY5rA1p3JfmmLs/TxTEkij5adPBLY8NpJkGvUY0cHPwDGpGSWxM9nn9a8TM+ye0RC1k5QN8tPLi
nVedJrivd+eQFkZZNa1FVVLyfMw5+OeDqHmmNelXQa3VwDP7d8j2nnkZPxaLo2FRehxGBwnu/HHx
XlHacfksJm2vPKSIP2pGyJU1LkAZjxa9J/2XMnhabdJ3cE1k3w5EPu1iEmbEUpCMzToiA5f7UtzN
YZ9BV+0lvxJfNwtVfhS+En0/sJzk4Tcb2TziFvOSIVf1S+z1+dxNFrDAJfwAneCQGiSfQbChvfEH
gHjFFAmFFNOsj9bheNWEcXnwXGuyJaMSWcGhMRNbCBQdng8kVO4ajMYchxd4T1PVSg7bjG3wr5GD
G67YhTFFMu22mAlzFnLchUalmtV92+rl5SGxHB1fm+9sNGg1kFQFcpdd86qRkd+hesKKsEAyg3UD
sKrBx/tlawwP70KhyuHecIEGHCQI7madwzvQyWzm/eJScK7pz8cCHu5R0NHkRXcI8xdNuhT06zc1
tJodLRrP4JDESWUG+TMcjhuUnwiU7xfGMDG+hYTWO7aVOhFgKkhx/i+VgH/GGzgkQcDC4j0CFzFZ
yHdERrxFTrGmAMvx/Km6sVQUkGrAZF8mASce9yFoMC1RyegL4OmlP0Hx9uSrh0RSnPr+GtyFFBhz
ytPeu7psahUqnpEj+U9scEg3FSlPbc6mcMy/Qay5D3SPRRV97HwHdQky42HDDEAKD5NCmVMhDKUZ
JtdODaWYbqhv9eaQ9GrIBvcWvexacOrhMciBZp82btHaJGHtPrpTBqk4goWfqvJKo680xQbZ8Pf8
Pw/IcMDv8TyQqJpQ98o+d5u6daIzycvzlxgEGejhLZPs0MfL7WK5DyMpO9W7CkjIz/Zk8BR1iCdw
YBearkc5BlBRbdiJg1cwmBENrdxM6cm/MZTuEVfqIdHouOmgOsaA3026m/fFjj4tuOS5BTgPtqOU
GWvWfIkGJ2Mmh5CW+NkYgadiOgeYcYKlxv4ll/znNDDufnrrYEzqLxs0EqdnfitX9BfIaCM3sOGi
xPX2XRQ3s/Oby/rUwLdxYWFyIJkBuWsXp0pS8ki8SAYPeOjt0MSE1cLTGiF0OdxUHUYhQCCKSkTG
d4MzfvRYUmAktmsSEJ2r1RRPB9lNXgZZQyxtUjbOl7xr9rwNrRoTYTVsmyqday955oZ2vNzbeBqY
xpy/rplPahwDDUOAEAMfYwXxwCO1wWlSySy5vSp22kY//+yMcARG09U7v7O38ALR5xEXMnYEPWs6
P6fjgNlSq0UXbfoDC1rtoHtltRcjaJj1QWyROLRm8s0x2v76yh6oRNMx0XOKd2nRVHm8jVgMIh1c
QnjzOjMWHaXE+2hj+Gx8vmdNVRhLAtbr2uMETjGm9wboHoGNIhqzsqHsQQtnDUxcBDMDTg2ZXLqG
i62UxG9FHEzkFg5II8H8UsFzaXxt7aBsbhuwV3V8J1/XpLF4i4slrYkbz/8AZsSKOCj3OvRVX5sB
WX0il7zns8YNlj0ORuCK9FZzrcLhddu82riK+K4nqmINdqMkNlHAv2k71ZC/vIJ2i5XtvWwykS21
lraymBoeblWLBJ4wV3gBQZjkgcWTorX+vcLxBqgbFLmypxUrBD1FoUXhpPARPi4OQI/dhyNAEDIA
lQ6tFdFHmHffemc+eipU5E9k0LN/zRXevSxtpqyOJd/6kKJ/H6V6okA3rRruXSxFR5lLeJ0+GyTT
D8AXYxJ76mdpOKikMHD5kKo00DYaKuhMBIoOpZtWi39HY436CMwpO5byZGTA4BEYw99ZctzaiMzl
X9JlwBlval8SWkbVhAVTfNGPTh9LRg8fFbKSnmIa/MjdcilOhtckvrmYghAPm3PgLm1glLQBHoQD
2X5eAhzx1BM/3ndoiXEvNRlEoIbNipNIMupaSL+k7Y/yCLEZKEVYzknftPj5GRWAoEkRWj2ijaNp
u9qJ6VcJyamFSZuDgToAnwneKzJyCW3znhDllgaj+wuATrxfKnGFhB2KQN7AsnZLTb4cHAjrotXA
ToB2acV+uihGOQWWmRjqF8rxbGzsvFo7uu0jB0LTwCG0unq0YABXEE4PdHFNm0FHUuy5901HAmF2
JCmZYVmDmadXindt18KTWM8E4mlll6oBr1cgxsEPAggqzvMZfM6TfpY2Jm5C2bE/WWnuFOOlzZOs
VIUFNl9b2lyKyOAJWaQRJ2QkIkdiOZKWVuLnCgr8vuWBZE8PXiCSoBjM+T0desMBfhSNM4ZW46rH
XEUcKmA/NcpysSLlG2KSogEgNcn0gAS6L7BuVd3+VoWeDvbFal0BQ3HKwTkG+vbnQUMVIVUZgrg1
GuCFd5/7Y0eX9tXbvFgG5MlxfZGFeCvkRJ6Kev6yNZcBXja8+jOZLOWZDYBCv4eBmxi7SeFV/Bzm
0hurmSKlzQr0cIjQhx3M4LMoIDJy26YSHLib4CCzxUa7TJJYY1+de5FLxKCakHDnXRUJS/pgwHpj
hlOtHQmZCQvSUaku7ShnZogjTiZuJuFhyDsUcSrsIWp8BndbAryY5doVfA7HKVc8FdEPHlRowfRr
JLnpanxpqKznjDiB2ETM7GdjG6Psy6z1vFLPVINAwBT7SO0gKrx9JXD3NjH88ykNg/zfRXZ52CtN
/jVc9gxUdxcjNWfztr00mbTEB/sdqMm5JANmqLwYmPmizlFlS34oU8EZuMu+MoUvXiAH7u1rA9PE
mJluGVgMaWqwmbJKr6sknd7bNhXbVD/bfXOt9hbcW93uNTkvhV0DfyEsGQchsfTu9/AJHmlAZbCH
IDCHVhwvZY/1FhQ6hRZHZ6v1rlGMR1HTLASTCiyUB4gU5Ge774Od179XqSEGg03ivjwMhhcV/YrO
Z3LuWhaSr6tZ+k0CWeGF0vCRv/OL1jiu+i73Rc9RFpDjD4NbG9e8Wuehj3/WpY13UdrzvIUMX7Q0
WIkKPtx+KA/yTgMVcN87awHht9SJcOkRYrE96MSP9dF9ZoXTiVAI8PwqZOsD9kOeokITwl+/b5oi
w49ITBfQ3T+YTKc+zrRSHQgfTqHmb++MlMhUy7PTDuZ3i+6nRn8mFRxVCclm6SDmucFQ8sM1LpxK
IhzQ2GRV//8unnr0RhWTRvSXfMiYAKo5pfvRQsl3v4FPQvfQVB+If6ubXA0x6HMGcq8bI2L+hy6e
AYbX6IxXbnIi6nrN5tE4FQtnnatn+HxlbS1zN7lq2yOZ0rrSF5SlcgWE/jtoEgKl2zqzKVK40DZM
onUQeZ+x/TypJupe7cObkgSbhHUkOhwMF1mwsxhd+YBKd81Q9tR8Pf1Gkwd88jKLiLiqHkyCZ7iK
kb/q1G3YhgOpu/eyz004Ldjuw1vMIKMkGpIu5IpuhWw946BUZxHBVw0wwLRGM6lyr5JDDND3CkNB
389UUbjBwlkd4jecKCKTUV05UJx+9/5wh4WLhqp2nK8+4Tbu5Jd497Sti6W/dZ+tV5OmgukxeJyE
OIMre9WP5VRQLhV4DcOt5wRDsfp643ZP5BLXFVq9HtQUegv+fJpkpcP7t3BAahDnnikr3xMKRacQ
e3DvEa1X2srFwzKCX0V6UMhRkXDtJ2ssfwReJGvKGbJRVUpJoP98Mp15qnqfH5/6GYB4S/lGIR9z
G8U/rwT86OOOO5DVUhvFUVACvKDIfbPlfPPkVFBcSevftMaGUIdjTdABNdv78r6oPaHBsH1GfIyf
TK/9cb4Cv5jmMj55TYyDWBHnZpndgpu3Sj2kcrcJcoI0YyNIOktBm6sOcjxSM7hU8d35owqAQTRA
cxZgGx7BT8QexygTmaKkQdHgub6AF2H5XYzjS/8Lm+YtNYeh4bHtBfGqIQXqF5z8KM6GYSnqZ0JX
1jo4ej84cR1di4kINJsH7YInM7qhsY/vDF5ev8QEj1gLoQTW+S7OfvkF68zaNu/LM8o2K8JZ7vdz
aQF8Xn0l+6bqgX7i5UGPMxSumw5fP30udM2ufLQ6v253ZcCzyb7pUqTe00A/GZgHHFXCfw3OYJa7
c+Xaz3fTlW0LtAXJGJYrYw+g76dLl3TL5e6ZbOJd27jCmsFJH0hzozOftA6FYLwDpKkH7va1Wkiw
m0wM7K2ZkMG5aHxCbXpPpaoTBTDAdcdMh67e4ua1xMOoYepndsQbrsT00HCtg+ckrULiq9EOf2AD
OJR12r4IRdw+15FO7GEE/AiH3mLKB+rm96Wv/M+u5q4GxSIoawHijY+eIKMkIVfZzmNr4q9d5ssQ
bW4iw3GcAdWuZf3LLLtkwB7cUH+xRpDYrUS5TO44ZK9jf3bEhx6/sJhMV4VPG2b5fyKO8wPgyScX
YVfrZEZUFg88K4YPNRraX+Zh+B4KHNFkiW4zp7ey2UZ4N3Ze7ImP18kmlkVL9/0tBzODoiQ9OguJ
NilKIT0egqfxpoNH3a71Si+VIcOXKCuwEdX1GngUJL0b8p2htDprgC62qQ3BBqmK/NohayV0LxiY
2APsI9dAjXjhrm7hcNFRnguMZUur5NKLWUWJSl9To6Ju76tPyDZx/WR33btej4Y2HikShTXbrx49
d8dA6gQbIa4b07OW5XQoneAKPMiKeyT9mLHG0DtrC1OBuwvlCf/yyU3z8kWhcWzU/e0wMoKBOvM9
m2UQcSbxUoTggjYGMeXQclIl0ZOZiephpXi4SEWBsM7pMW/zu9yloIZ09Hr91ujJCWTP3CChgaFS
Vqf1IB5sJKX2BJ5CAKXq/3ELDp5p5Jfe9NNlnt0qR44nMBBl0Ooc1hjhrNkmUw4pHzuxmO7HtyT4
Eh+AYPelrkGWcJDiWI5FT9yCkC/zMXgyZBITiXUUcqfmj7fZcJ1lxnVZjGgFfg/JfU5FHFttLL3a
uMFR4m+MIG3M5PmX0IIW153RM3Wh4tGbEuFJTTFWOLbPWwxu/O5l7uc2kExYRS1eHo/TLHECiG73
lHs8lQtchtCwU65PNung52SgUAZgYgRHDNl/5p9CoDYiJR+1W9GNQ06vZvM/lQRvfgyCl5As4Bu0
VnhS5QqimYOSbAV688flDliM6sv7yx625cmVt8i0jQF4bbsqicxgx463Nv+NoblG/aCrNycEUYlt
nHQbqRTS26bW4p9Nz3abNQmR1k2p7wo9Kmx5aNylFFBqFz2hd50uKeogxjSohy2vZgYCcUmMvXVq
Vj6bTuEe59jlXz1bADeV7tOocxnICZ8zfm3nuR5zU2q3D+5jhwIQUapZ4Pvi3Tjl23NSm2OPi8ze
NtucWWrqPf58T0ART5/TUPmgoPNFer9At2znW2dP3C2MulauqFz8qXnx2nFPXjrERHozx1ViA57S
wl03MSiBmccgXoob44WBlhoVs2DxD8P2sxUgqcFtsOxGg1z/Wc+vdy9T6Ywnq0GhXM77GN7+YCXv
C3bqN1TizFGjN3QMZEg6A1ufZeTgtyJPbABaJHWH90ecADEkX+2KkDrBYrOSL9svtghYD9jeSqVz
4gfcG2iwaRXCUi31hlWI3MsPcnbk+OUexIqwWC0zmGvVp31fOVKgiErLkw9btqPp6G8ujrzE0pZO
gdmBTEcGnxKVq0cI/TGlZbrWyyj/EU3K5EHmIa4AlEMmwJrhH2xHSiKBzAGEjWJ2Osn092xM/+R4
HcOzEL9b1O7wEGGz4c4Ny/lHP0W58XWebDkoK5g9yEhgPMg6ESUJ9kUXNG1RIhe45A1Mf/n8xls2
lZc33Ootv8VU7IgQ89lgHBJxpD8TFsLc/hTYOVtw+yZdWgW2ltHD9Eqi/6jH3NsTZWDCVHO1ogfJ
RHXI5XfarmyWtDW8R08t8OFAq5Qy5kJDPwv4INWJEodtbQRAlFXkaCMRp/am1TeOdv1zT06sKmCL
apYAEPKNEZ1F7MWcXnkSj9j05wUfzROxJAzyiuTtp8sj1vnpbNUeFdl0LqXf+8n+W4ieglfzTUUT
Jv1IeBZJgIZrJbiufEm+OvliFQRvlOaEQumdEhbB94zUD4Vq2F3Ugu2BvgXtSByi9mgYMNfiV7Il
CB1U5SHRG1NmY37m8jT5GF+2TzEgF+BOvqpPcxpzm6tQEQLwYf5vu9n7RwoOFZdJ9ykraOY0Aa/9
ScnpZ+ekAWhpVMypMvZ9w2OgbkI7Yac/wLU+ulyODlvdIlRTLYGuHoF0u44SwZ2yfWUECad45SnL
8eTdMhqB6iJ5EY0Btb5UaMLk2IDFVEVpmCYuNdkHG0Y5b5rfuLkyybsZcvQvUVbSpY1Z4mzDquCt
bfQleEAlP4g7UyU7qfh83wCS/EawU5J0LD5GMMsbe7LGkecD/kAaxaKr5MDub21ztBhKX3oYbSQy
eLx8R000guZ63OtCIrCKk+hhbm+B+eVQBI5nDs9Y3FCQ37fHFU/GX72uLqFfABMxitQgzRheef8Y
BdxPwIofGPZp9/U5hDVrhzmWJ4hHEOyOR5uaHZfn87dWkEmFV348GIJXaS09sAsy0MjtL/vnWgYg
kJvIlApREJjJrFxrBorUcEnSYxYaDjgYHlSJYqRCC7T8g2EVYa4Oc/rTkD8WHi2UHlM0SsF27Smw
uj1ZXmRhzGCVTJFY0DQ3kuwKsALnHQkM6CxKtMmNV/T5J6gIcHXWKbSAqnL92ErYdUcOefLQDQb1
eZ1Q4xbeZfBkk+DwRRW4zTQ3d6xgoVKX4mvY4vZNbJZ0xAvvXtG5KYqZFWNhy6oGo/WUYj5/ygSA
lgp1voxUvdsJ23XPhEUlz4rtmkjxIp1rJ//MDMC44/x+23Wk9aIP1xytFsZBX03pxOX81ekufjad
qwORG52gB48QcISQ3/vB0HR+Tuu7lSraXVz+9kYKTkP0t00z2kzNSKrTNh/TEAZxmkq9npekzwD5
oAqpGSRpXpqlL3MIPVqe8AtzWsMMJt2D6JRCqYh2HgOtpVhc5aEGLfITigP8dysGS4ktdiGmqg4G
7kDm5S5pKIN/UkyZhPZyqKmZm3Z2jc49EK7STdDlTxDzY0+X612HiZE97/Fmdh6zTyT8me+3DEpT
iGVyjYhVfoqxqpDJ6sBIV0+BdMOjdUGnz5ill5VX1FWS/O1C0O0nHwZyK2UZBrHfUMlzDprbAXlU
P1qPJpXNep5dO/aGVOpQJ7JBbmo+df6MobeVxBvAoQxLISHGB3ZyUN+hjmCsAsq7SPcaz5zzo0d+
yNf3DZTe7PVzU99/nvgtrqu8OoTU2wOloE+ftBupjDsx08mrNOzOeQxwdthfUTYV4bW1BVaoN5kM
/VYUt0Xaqk9Pz8/ci7NkmTwUrIv73TsAQZnibp6g3gNIxT2vyjyV5eE/citnxIJN7CNp3BR8LI1j
mbNIhUeYqRyTGL+/PfwZTZv4jo+y8oV7Q+vJc7vajlZPLYUk3AGAJsfm69/+KensyxXqQhbgnpGM
nXSy4U1rhB6teTKytoeZJ8mELPz5He6pZIwS/1D5HAo394N/KboREDek1R0YqeBihg5nk/8dkEoq
K4ezbybY6RXI1xmXyIRQcS2u78kADEzjt5MG5RHT0HrKOHwvanFKDqCy+FrmHfyzfFypI91kiBqC
xq4BfgGXDj51I7AS3lxMUBbXQ+J6vtCaVwbAKuSMZYRbAxDDuupvpk3r7UzOnQddPBaGMYwIwaxi
GnHBngSkJaapKYFYxtJDgcljS9ue7sBDYnuJ+4HZkYdf4ra+f40M9s10iPYbFKVL1xvbQoBCftJA
TSOjKhr0dULLcJgY1ULL4v3Emvyn+sb+qvcRNzd2u2flo65D/KuRxqdQhI2Ay/Nd5crnJvCJeweF
Hjl3FusAJkwfvYjj7PbhZFIo50y/w7xZ67KAgzDmcww1YaHfC2hQi2A8wnJxxXiTWyWbUBV+tZLb
5Rk9pAPG0o3cW0n2rcPyBorT9Ymtxcu46myk8HweX8xt4j30XGnNGDLOASmunOc8rbgQBtrCeIhT
pfHd+qGb+8sxUrkaJJf+rI55CFdI5Y8fKyggK8e/hKunA2XCTzycVkdJfViuRqWWC0ie2aaEbyZw
qu4oaE0HXpACO8kY/prvhmPAUezhwVxuNdKxWXok7pbi5s7fKEJxlouGXAfeUTGxvO6BlS4wFOyc
XOZb+QHp7oJenquPL9uxjqyx4ByKUPjW2gRBaD/xGamGUnFxw2/kex/f8sDnaTH/P/kN7yS3w+y2
AmKaN4odLkWKfenbvJWFjOs8XWy/MF4vwk22doGjtV6lXoa4+B/j7+/e3rfNSzRUeqHuxp4Yu8VR
rbwVpLZrxZMh22mqEzJwWQWfMRFsLJzef5/J0jMrZagD2S8T/RrVrTpYpthlJc6kEmU2O+O05rdM
LESOPDfDEuWfDfkzsvFGyKK2Ci2x+Yf8ZQLAxIGNKsLueq/scJZCRxSJgH/sRV2+XA6pDPYKObw/
/CzERc7/+Rm95cwwVHLCu58Qy20hDatRa6ydK8baH//W2BOyrH0GodSWvSVokzxuK35n/3RpS2a9
T/FasjfHqt8IgVfrJSCQSdj+DTv1F8Goxvq8ihG6b1UfRMJhxpKHOqNhRHSxibsb6H6Ovb8H4h7e
rJVdZKI83HiZY4CpEkbIL65//TMMjE4YHU+yn79zA8ARJf7OsA/fS2DVdURGBWvbYPR5K9TJJIDQ
URLPtMKt8ohygcRT6S4vKfrnBjBJfC3Hu9XZJxtDQYrh23fXox9GvL9O2dn20QHNu6KkmQiHDY1q
CrqYn0ZMaLcUIQZoAXKbW/YQDyQDGK2NnNZMvaVUN2NJSnRUTBjt/uoamElgJf7CVaYE6meXsNVD
cK0jzoO4iDQuNK5NGXap2nkRJv5XBZVmzKVN4yjVKkR9b7s+b9kQlQ7odlnZuHqBrDZ3WAj2J/Ni
I9HiyUeCzg4VZFeioc7nhFnyEOj53EuVaKKlGxmZKBXyNyVygSxB/FPqWutx/NPuRcdNo0ZHZa97
ZaMZtuVhrtPYFK1ZyqQ4rdVlG0Yy80513AvCLn2f1YkUTk++fZx2LI3cGJxSix94nEbVHmKF6MCk
zlcwElYl30gqC5ZTuVwDLOq2/hqlHl4NUEg3NpMMMgx38Segp6wV+TXztC9qlJovzmx3HeqBC0DQ
W/8tf9oB7TF4h8azS17QOwN2B/zH/SXmrLb4+BtWX+XEGPIhKkUpwZu1Mw9G5q6RRNDV9d+tpy82
ChiyUP7PdLRKsAch+9jLJNlPBRRe+5rtshn1VhWcoiIT/joz2agF8z1Xe+wMEfFHC/IHAeU6+i4c
m0mYD/aIOqS+8mZCGN4yFw8Dr68RYBf50MnZZFNlySg/9PR9L1UWz9901rjMRtGzaluzkbNOJ956
4jW+N19S2Xb4IIyVWaIhjBjkNDPjSaiwJ1BVzoq1Img+iRuT9RUOK+XD4fDADA+FqS4v939wQIs9
pv1pBmHuGWneYUbw9bzzgsmNils+EjygFMPWlpdDuzxHGta6M6XNr0RHZKizoMuy+qBts7tTRiEj
PH1uUuf0gksfM3iUqHS+eH0vLRPx5650ZKKwPIqwExbMKduYLXxHQhIAvEF5uuljctCtNbyVmalT
KS+KfDejjfog4JE8u4/k+3g3Xdw/bPB4vbVuoT52+BrZXHg1F9wt+I/9fU+mTeGO7vJF+PkQ70+4
xZx6jezEir62CJj0AyoFJXlefEMdlEXddmPqqwbptAx1OFiStMElYdPC7+ukpKKqrh+l4dvFW8FZ
EntS0Z2XtvkhuHBJNhxeWAGS2zffjHnlJ1kWSe6RKjG9CxXPtxge+BiuvBq39T9xdxUDItlNsYsm
w52Wyyx6N7GfNK8tgLqQ3bYpOTvFobVQeq4YmoobyRaYcLeEb/V5bhVaIy+8hYLHu95LuXi6cIoM
ngklm6RRrR9O8FqgEUGQhSJW78KR22e+0fCVcGCaMDzJDsZaAQ6ZIyRiotbui5Yp9CCWnA4KMpqf
7Wvs7bIWeaoRq1Qj3+sRRI1a4CuGJUzb+G1Op9F271wWvBty80verHQ3+JMgUtd35pJ+PlwX9k8y
VXV9cFwyuyNqUHpmwg/B7/EYsFU/afejHwr2gzUQ3svQDIyNiTOTfFILnpyy1CxXCoEaGJsXwsm4
/X/3WuklmIYmToswpq4fvZuKD0LtJURtJjUzoJgNmpZxkqaHl2Od0a2Mm2200NgRd6LCfK/3S7rD
vQH9RTBM2HG7Xcis9KWQ79u/tZ9C22xIgMPSsxsCaAps/+bdj9ov18LNJii+84IDOIvjvdKZaH52
Rzxj+Ao8zCGJjXzMLuuguZ+opxMzgQRqSLkBvvONZm1YOogddY2++IVjiIp7+nmb373BmwGtvH1C
tyl7vHRt261CxRdGvF65pAUX5C5RbNrjIQIePi8g1ur9V+ul7RyPOU6VO2rDYGGPaesJIQfTWKj2
L5IRUNaZGQ6q9oAaCf+uMCw2zjuV1Xlf7HIwTvWKk5lGPGRmfnuUADMWxeFSkoSrU5I6TAYmF21w
jk4xbYSvOS/aQS6K7049OEhGbdNausJCZGlmruUOvR2hnbMMeZ6rNnmba2JNzOp3jtfe1QSD6cq/
Vs0X9pn7Ld+u8lH6mM9Jtd8pL9daETaBedM0F9Ue89Oz6ae64F0ZC3MJCI5cNV5wAYWe6CWc7TxR
VjY6/1hJJ0ZSe+ATFiaVgeMLrAb57FQQ4/cogbTguJkOx2Dy3B6BKNGaoTw4xo7E1yYfIP27b6r1
Cb1ZRd+GuY/iW2SCCkvJ2E8sOvZNrDTLONLKVp0LF+remlJuoUwE9zRzBGYUW2/iZzyPsxn17zoj
ocOA5RFGk/4ivE25BcRlCaMTqyxjeIkAfuAXA3tQxdoJ68oXnVgVxInzc2nY9nAReFqcncKwcUDW
bRYbmKQkI5u4+8Wyy5GJbksgPAVcdxaq+KGsX9q8OMGXXi1WCvr1cNIsbn1Hbl66Oc0KgV/GEonf
Cdyw3/I/e7X4z00z1v2IuSwvBf4FIAiEEbERj4dSyAOHX/Iiy02LZlgRaz6CED4lW5kIHyuxXqXB
X55TxUmEs0lc1EIrraTd7IgBfTwrEwFEwylLugedY/nsxfe22k4GZh5TSqUStG4HFHrethr+isSa
aUrT7eECpqZ1wgJxbMP5XASgzmVM704jkoY1WS+Z6L0vb4Vlr0yvH1DLbz9VLFAs8TFMOtNGpoht
1hlGaQKekVOG94fxNsmDHagXpZ1VdgsTM2B05Kl4A+B5TLmQHdHA/JmIsz+rNIK6K5AleGxRPc5p
EPCjETuhABhqw9UxyNXWmsv1Jc0NO9OWfIyExtsXI04EjFje21r42xlOc010UoDeF0chArY74Oz9
/ThLTu4Ww4cDpz6GjYHks0cTxmQpAjVRqd44uDH1F3HQh3enAFcXHZ84N7cM8BsmJxGBcnFDuzd6
dRJCkiwQTSQ4vVIZFSIR3tLehS+MJ++2Wl2wLTCsyMJQqFJfLLpI/R9ZIEYMs/KgZIhsRTWq6Y0D
y+VBAwzUS3vBuB+/b3qY02gDuEBD/aAWR+Pai2nMutKdZITj0tuX0tp8BHcAGbCyEEkHHM33Yhd1
cg9mgAVMtHEXPf/zGAKFzexKCL5xMhRu3B3KCaovtzEMA/9ZPxiV0VXbeh59gd3Sl/HtczvCfYSu
1oS5K1jq+id9m7/fdWgkil0cQiOjq5vnM7nAPVF7bwgc5ERyk6J6rYJyFiC0Kot8KXETmHiiA8Vw
0Y1cH8XIGCT1FhUBVPEm+2PdKD66ten2fWnYou1y+wDC+x67a7Fkz5g/9Tdflc2FqIma1NFgJBuO
oLAPEr1EkYxzUuZO2Lv/VPYsCG5e4cxVnuh2MH04LAxxZR/jnFwOZqAWIRSDjqZQaRooaa6od8x/
iOO52Gk+UY10j9YsDWhZYYkzO1w3Grjf13cY51oh5Qy8QxpFK0yzvKdnkW1EukY7NQ0jdd9Rp4/p
nnZhXmMDRhLtjRzRsaV9OzJ/rT6/bSgQ108LA/LS8DLDt695F6K2sgNPrX8oyoVVWfdjWH1wJp/Z
E8fZ951116i0hxEpSBubrM8jrSWCLOuAjoO2RNO4KPSienba6gXjooItEbcJcfu0j9p+sYhCfw7V
DoMeV9cuIzJgJ7L1y+IxCg99OJh3BTCf08uCcOBQnzZoCyDJ5iZmaBuDXDTtFhOXQcjiLzsYGuPF
tBYFHvdByqyXgKW6zCaKHI4wgifqEJ7SZ/du753jhZVBshs+ZuZpfI0u4ikSkW8iuc8iLFr+fzzI
UMJvn/esI/F0bDQG6TGvkVdIZH3wPYI+bPZ804SKN5xhB+WiEdLnDSNK/ep0w2yqP/xiNhdTQ1q+
EBlBI46jKsN/i9LHIGTC+Z1YV+bguNJ/vrllHHjQMluIW5jPtX/OXu+sl75yHb7t1qEV/pjfHTWm
MF++9SYDC6ETygN0ZyfDj4NgijYFhw1ufGQBnwccQXguOk/VyHlSeGMkTD9l/qLwOd+fZ8cEmTQZ
1InqJGFT+1SWzV+KUdcdfU4DeCqZH4vWSn9SzrxzorwLudgNalKRBwO+kavTr8L0nh5t4JbfVdCC
DEx8kckW1Bmj5fRTTpePfjI6k+rJ6qcMFFatWYviFiZduSUSOXxhHlrHs9Jv8Tbh3XuRE3PPHDs/
aLJWyZTvFDmrRoUshyn5dWNVpX4/5E3Ph8p8XECNRQQxHm8JJIJhNelJ+lM8E5GIyeXft+IPr1HN
lzGj+qHLw8rESi2oaqliMdFg912ES6OpXx0hqKZhABhsO70/Jv42icGX+gXZxXVwGApMDnzWvSw8
7TfO44zmRqfUk+OAp4fUVtYUNSWh1+hu8WhHi9EwfHztmTFqMGnUzeiQ+CBL+M/DvPA2fX6JkxsL
474uKFP+geY8nsu88J17ebpXHesXcWpLThLMmJd+t0l1clqbn1sxEKsD6P6EWT6xd9bs3T5KxwwN
qD8yPELabAflQYTFFo3i8jKZdNpMW9Zo+vKgR5KEJ5tnkqSaUXCVm0al52uqCmcPxjLBwWt9B2Xp
oI7FFg/Fdy/lNeszKj0HSdxwdPLNsw2IfSHIhWzed5+jd5BxWBMw9DScKP03Qkd2qxOV+WANV1g+
/a4oGfZv4TZp4ypntfkSMoFn4MTeTdjbzwMS4Kl7sMR2Zrz0yod8WAEqWjG/d5fTJZegqjHPQrdA
3lEo9ZmluACJiEJn9GlScQ9CK6a7FHWkYuraWE7ZI8au790IauBs48gDPUNXcIMK4w4ggbV3QvsK
in+9hKahKZ/eGpEH2FmMv0OcGrJwpYFBWQmTF4mcROSmRhK8MtJxI1A53UwgjEGpYHQ5sto1hF3p
s0aRyWLwK0uXwsDnUctgXRtxAUx6Xq95ol4ka2fiOmaePbZsjaRRe2x8DH2EvVb2jyMbyV+foPNL
+uReFMgGy0FYTwiNARAEkn3HICdMGHlNEKVs4FYfLNLs+qBeXB3ZhWnrHJgfwxUkT09MVs0MxF0I
Kb92Yk3t9I0gncrNO5fVmyZVweGDf2YdtF3GaMqqamyfXVYTixfMC5+pZ7H/5vlQGS/ktqUyRP9d
1y8RiVDgN4uN+TD4u4fM9xYn5zU1jbz8OCB2oAtPIBRB6zE+RFK5ChEUJ8xiCexihSQjS5URM0t9
npRLT5shrlFfS/RBa4WZ5L1Mhz9rgPos1+OYBM1e+JjCkpWJ+WK7oSggeDokeSGNFMPtDLLakkzO
aSTdab8F7mIDLQM2rvHxZp7LaWV3CPE+gEbm0oNpDZrXDURkfKG2hULMiExE96ttz5uclfn4kcTD
x5WomM8qKD7FRJTggY5rMOjADotUCe4p1YsgS5PyEDKyB4JcUJiAVCSdPhoERzw+hqVDp+Nj0OQt
CfKwLIpq4LzDM88Gu5nUORvsiO7tqRXKy6WvGUv6OrG5coKwkr/sRSnRGMJTL9oBhHOHPBFW/3QX
7UJkgX9+jfgWSQ5g6Qo/Eb5hko4Z5aIgz20vyZQXrGKis+NqQ7riMVxp4FkdE9HwmT8rSXa83a3Z
QYRULe+W8y2yAXOryw7FbMwQ4t0LgYay6D2jkivvA5FwhFO+QnFgxqlXcynB6wdRyOzfdYpWhDq8
svTcuRWYQC8CAGVL1/OZqnygKeQ7mnSY9kKTkPAmcPuGaQdO1EIvyy21vFRyJh/ERLDZpD6J8X+p
21dhwGI4fuiwjpiwizuyWlOTbgKY7ZSZpYGyyZxme1ZmQxi04NoxccvdXPfJtqBc6W9nEaZlsjp5
WuGP3br7vDFc6/SmTLFNqSoQs2pVFRcyPJ2mw9C1jVrIfMG4dWS4x/U9mcphiL4oydkQ2k5eXyBj
Cqe9meGL1UqSsUW1a0t1vbB8LzykGAEX/zkpwFROOj9A+uo0xkuYYCGISV7Io1TnwxqnQhbXGT1e
3fNHYYMrjmuPa1dhE3H2xNbK7x8B2FtlWyyljPcZhT5KRHahn2TZ0wGIHBV66RrsvHHJA66EeqSO
krSADCN1DnLSZvPvDRwx3rxuz8DwQ90UhXoWn4R81l3++BADHya+k5tb1ZGgdb8WG/BWY0LrVuuu
UpJgVOax8dY8EcICHPmnBQfitUnqimHOU+bNwbktTNRJBnZ9B+P6VEajhtPdaZ6GmlGzB/bxyEQW
KbKAMEDhTJjJk4WpkgJxYnvRlOZKW8qdB/B7srs/wa55kS+Q5UjUXNuNSJzTw/By2ElRrTZfjaiS
896R32yA1NVa+kU+KZUY0OXvF4slU6MORPC7VROzVl+ViFqgQJnGntdA8nrThYNF82+vucwkFrEY
NOLnmQlMwuC3aD5sUpcNq1twInIAdKcMYNnsVQx24M3fMwqSxUPFCr7Yg5n7ikHz8fwpMwluYDhY
OT5JBM/1JJp+sDm9wfJIA/5kOWdWtiM8e78SRZQtK+/v7oQn3vmEww2UuB2TPKvd4aHHxEsNvpo0
wCmXkd8Vc/RZ5+yCwKg1UDnr64eHXqqrttbbzgk/lVkjOFKBSaIPPUBaOP3AXn7Nvodik0WXDUTP
9NkNz5xKwhHhpnALI7oJSDayksyLjHCvx30Ch2MrG9P6tGpVKRBkZSQblZs9syheWfxzPCoztQTW
ebhVKPV01/akgBaa3rYDpwrBae/o8ajNf32v+TxFotu188jKYZmsTHJN3v+PMYc3StooRSKtjfQQ
Vbn+sN6F096ygm7+2TBN4SoQKOXVXoGlxz8H/dhrDWU9GhEQmorKmC5pJDSzMpKB41Lljuni03/D
RdW8ObOnG/CgiOo9Sdo/bJGLiy+SWJnA9ZEQDxDFPne6+shGLUDy2c3utTfm2pXT59b9Gx+Hx64z
xR3ruokzzt4wgd+S0zTm3miAxCQo6RqAJ8oOK2uVGoEtCkwn3/NaOgqLPihUSCg+KnaE08g50pJ4
mDWEji/UvrN99NJHCUEsJqBFg63lcyb6ef8pm/vtDCwSfiIXNNVMofZpjd9FsAVnM35awaD0INM7
WSjPlR7wZQachio+SVXMmgNPT6AcbjS1lx85BL2KTvwfAy9Mm0OBFFN7Hoen/DbJaglqGYBtx6TM
bqINKntVLayq3Gwdw0aqW+Xrzc72gjnw5RDHDLR6a/rNq9lTFuq89yu8b8wbm4adLj+XWhVQL7+z
hcXulhPCBsZUYuBAk9ZPr6QA//I4Z8TvKe+2Y+23kLDbxbk0IJObbVXK+OHP4nxG3FRh52taNWBC
AG76ffnHsptV+I8QenUI/7s+Keo0ebEBhBtif0MBgVDY/s/KkW/xIgfPpa0aTLc27yjhkb3NnM7S
9r+BHJ8y4/2tkvZ0KVa7Ju0r57EMTgzt8+L9SIHtdwu4D24+eNRWNwHXgzK+RDlCaH7yVyU50lKy
LXzF5TeplXXo1+OcfwsJBSWGrAwWEoUVdbi62p7qprUmiwd1vreYa7EtXEanaAsPZkb7t6HxsxYG
aa/JopF1T3c5Q0CqW71RMpFu/T1vE+wsLWVlG8ovrES50yfNOu7DnK9IqJv3Du5gUn+qsbqkyGWx
97+zm/ZRYR3v7M/gxtRvW4DghA3mZznTj7BosYL8C9zUGmTaP3ABWFxW3J7ERen/us3ZQQT4v08D
nd90lFJZvtX+Wd1YGr6Bqs2RcCVVJT+4uzDLnb5udYxWtqISh8Zp3CXfSPapDX6TlH4hn99FpcaJ
BdDPwkS5pg78KUcLJnAIHC98kGNTARkmdOSciwG8dT5OZ02h4a/qcAvO+Do3MfeISTtuabuK1M33
4VMqQ1prJ9I5r4BGCRnp0ypLdQBf0GeSWt6KQZv2HhN4JJBurg/YFzfmGpdWe7WBhxLwS+aGW3x7
QDA0kNL/b1Gn/f10QpO2vYW4hxQ/jo5Djpz+clLdXAXPWoULBnxXDGJhl+FBHc+Igtlt3CNDucwL
s1fJtsoBJZwPZ1imr0waaU79QQtyx6GMa8wSiSP+IrENe9BZH2aWbpi3ZwA3fQieYGWNjYyljYph
SbniU+eVqWtXinW/DzU7q7nl7S2Tnr1bI/ydMqbP3oFpYzGXbiblAt0NIN/4TRoMfZF9shlcKbkO
WapyO77GyeOZ8+sSFg1Of5EKTYmCGM9tsSiveN5PD9PICN35z8YZADQ/kEBdTI3GS5QdVb1xoVuP
D8dAtwSobZsmkYtQnQb29aZJ8IpAmO7y+fytGmNj6dFj74OdugtR66EAlvnllkEP2fc1Mjjtshvc
YWcui0wf72l4sYJRI95xd3UW/XchF4cyXL88Ta7XhKZSiHcwSklhsrMgTr0qEnvtiO99gUM101At
uoDii1Is3zzguz69fFRYNQeiStHi7xuis83pjpXymaehYc62KOAH8aKdvSdDZyAc9ilJ+iKhwR/o
VB67C1bYty92vtsyMjW3ujEq5MDBPmqt0kz6B/YxRunNd79s8VUwowh3ziXT3Bf3bHij1tt/ySdS
B3Eqq6QCEJ7VTNQNX7k6S86EP5GtQ/645MNIcmSGhqMRqJ3foBGYNzU3d468mL/ROyKjaUGQFzjy
g1GZJ2k+f/EbjBdR6xRQ4nEqIOa6aLt0tjU2ivT6wZP84EMKWbE5VphX/zayE1NRmaZO+JExFKIa
UirqVDZHF8P1f0spv3eN1iVBojKQCK/2VnTHzlAE5l67PLQuirTkz/6lk1ND7d8xZebN/Y6Y9E/y
nTdggt7G8XRdxqi71gRVhTHnxq/+8RCYaC0VmPqKWGIGyDPHd4D6Jec7kQgkz6ToVR487Of4gDYk
G5QkQP4Nd0NpZKos3Vy/7Vmf08QkHiuFUPdYfFfKSeAYjmFlVNHxM5D5rG5k5AFVcpkv1KoUI9oj
znIr8CKcBsDYJKA2RVCIXhpGe5Yj4ruih+FMfH5HC7D0AYPNCBJYcPDdpdOKYS62bbFv8sAz+ynh
2N3fgRguWTy7TkKiR10OBG26DUB9SdmSOnqrhWRL/s37rfWrNLdxESsgMWATcVb+5zLOsKY3DIBh
qn5LlnG9mOgbaQaS+zBPaUQdPnNYFh/J5BsRQZv8DWuucLhNFY/KAmje+7Z/LldhtQ/VgvojarDE
zkUWJ1c2LXLWCSUvHVNh+Oqyxel1NNP1bhJEV1j3OWDprZmhyuY7BMnXhmmzJan4W8cgZChvfPHv
nyFxAKU66NchI5NEtsqi/5Az5D3tAzsWVz4U1Luoiqbe1wdZj1pQVw/+CecFhESTei4pPiQuG1aZ
90chdPvsxYwl+7MswCorJkxX2gPp0njqrWBI1bkZPswHmF3KFTUp4E4dxcYjZIgB99VrHV8BVSlF
dQgtDCgsQoU1ADR4kfdWyWFwcVQPQ2G3k/D8bs8+KNA720bQq5H436jZC9iDP9vZZpogsrAzc9Pv
e5eBuABU6+/jX7mt+obxOof65T0c+uz2+36TAsAx+cYv3JiWCAQA2Mr/FqRNupy1GzGB8Zd0ZSmZ
YYrjwu0/nB3d2DPpajjRsuftQhetpIzby3vvlXpXpnJNIbgeiB+6aysaL6VVMnPlE2ZbG4qFB/rN
CMff13w4UPK72cPqZ3pQze3wwTENQHAlhX5mbIcNdzwvJWMeMiv5VlWpaJoUV7bxrPqutlBwUxkc
BoXyUEzyi6S5855HFY4Ae1I/xjLL3J4iksJOwCRkIoeKAMIA5xV5o3teYC4m/xBlpxkJQQu8MjIY
JaC07buzag0csM/UURAdMXNbcHruj97BH/fUb7dBQX+/umzf/d7GRkOgYlrilTgaBzmvb+hqHc6K
Ir6FDDwRmcjSkW6yTkBJGZRTqGQT80OdEBx3FT4R7ICvT8KhfnudXnHoiGpsxcLM9KaIv7JFZVHH
h0FIn4ONt3TjL0BJp8+IZktqUJvHU/LxjKy+qDQYc2+k4+i8mx13r+l41FuTP81pYeu0C2DV7vV/
hImve+fbvxnxTWi8QucP32wKWRFMoNyzHo8ZyL4d57ahZy+7AgCtUvsgcsRjmTV2TppYRvAHSqmp
Q3+vOci7VTmJezL4bLOA9+6TdWTrCkGxtxGY9XzvFcAYpZJRiE3lG8oobZVklcJomSGDtvl4LDaG
Lw7KkFXssrF3n19xDP82adP/uHD2lMwFQTqj+Fsr772wiJdBCJr+LYoo2T3V7NOLlATUF3iCi5Mt
GKtuBohKDCFS9PDXXHxJvqO1YG2a7ICF43/dUj5wnlWqCElldi6N2qNE90kae54ag36t/RxdzHMY
PFKEwIAZxUei0hgX2lYH5LnJN295M6rd1V/5K6s6KTVDEUz2C7yPW18WYLZvy8xNG+UziXuXlyHq
B/jPiRbqTDINg7h+fqUfY6Th+c73XDPGB4KlS8UToiRGx0+9quY1DMF48s+2Ux1Ci1+qVuMPCViU
WqKbE38MVPH8vbk2vmnO0dPXHeza9/EhLhAKJn36f0D/RM4xQra+R8BL9Naq19WDZQxofRZeSgTe
a8AtE+4Gi4u6G7zrWic3KFT7gS4Kc6amu2/gXOEnEhe/+dltjjtSjfeIvykWz/WXiuij1MIRz7bJ
N7feBaA6neQuaCfKdbZ22hcfp6m9gNqhZ+a5aZPR/dDnxyKqkTIG7tX0pryLbxeU2vj5VwZfoy3Z
pX7xBnaV9mT92gATKcFMs+3vKnVcrVfcud3uWgutRP6OPjZXUbVFq6hqx2/TGSe5jRb42SKKXURb
ogBOZmO4RPQhq/i767gFl8A1JbjIv158kzCNeVPKhCOUvyvANBPmsylC1psJ+R2dTk2kTyKFG629
vROqp9FvIvB40HD0EjUNzhoJHM/6DaS6cerF/SdDa+qP6LYOxw0Mb3TLwxNTqPrcwco7AVgSIrsB
TU8CsKnz6IIb7Bmbw40aPdYJTj/kqmWWn7ImPdXAzNYvwD9wxg1vHAqGlamjTEQswjuCVaicVR/j
ubmyi520XT8MTKBoTVtpWIsifxeXv3dOHRBlfwavrxQJ6N0qfXNiUMmlVICmcAU+lHxs2gpPMU1f
Id1DqE6TmempbvHgmQdy+y2JdvhAk2GVVRmYjUN+iP1bT3nbq/MlRuYD39DQWMAp1VmHmvAJlkbY
Hju7cAErBP1wQGkOkfXyYNq2p8uP8ThafNVbtxHH/0WUu2Y+lBWT8BQR+AqG9JADpK7DLaJpNimj
d3zF9Uxr8hNDwNV9G7LoDgFLERF7QFjEtuKW9fCTLbrfJ78Zsfw1Z3VfnVwbCsv+NqwR4HTCRgz3
XmOzt0+ePwtCX9QWF+dNSrSMcCr4eTXnRL2HcxgRajJHFVeZ6G8zuhMMjdeC7+huoSFDan5pxXEz
HtrPxpONccbkhlvlDZ8C6uPZe3FUQZ3hJCX10OIsqiRq355wMluk6JtWnD3isCzTWjep5ZjR29Ic
PrJLMaKRvjaZ88Wml2BNipDIUg7GETcuyD+TF8sgfAy9A4nTtKGEm6wTK0Tu3Fyivmaw4ceIcH5G
3fh0N0gUCXVCR03g2GGO2xTfIyRA2t0E7U5D2ERSqDZTCp8+vSQj+Rk9HbO/rlH3xUcDtfA7bZgr
pAwi6URlVUkQT/vz/xMcl4sFPmIUygfszBrBXLcpBLId9yG1dMPukv6lZVkebmfVPmWcijXSQ/Ox
np5o2Hnt6n9Inebfp4HWt8tsGXdQfrMmCX3kBpASeMqTjdBXtR5L1AHId7OQ5lA4+kAPhqiu8jkB
+8pklOb/libI2QVTdD23EUAcdUQ8TgN1BROjnDBKTqXuQtmndmtmMlafiOga/osOSP5X5Ooj8Zdz
1uhfF+GbdXyJGFgbNifeavEvLSfFZIdsnkB2gU95R5PXP50R6HFQxm1b6axr20UyC887rJ9rDr+H
U9fe3ud1aD6XdehmTdPzzHsa5NvBfRQZGXfdC0Cuf023kCgk6fI77QTwFEcm9SOFZ+AZ1QFqV0zB
6OWH6/1lq2GmswLfGYz00SMHh1vSphceEWVpAmpCeO6qdrjR+jpm+HQ9QKoAU0OXrpO1B16sIwt8
DwRco7UqiFOOl+au2pdXvWdXObT58X/yriOfRz9HEw0sg7mGJEK6N3hZ8FjXznchFIUm5DYgx1Kg
mN/zapqbBIindX3+Z5LPLGBP7mfLA/QIlaB82sJ2IRvMojWaeEoujha4YLcDSeSltG04OEL/H6dA
cho3bRqISUqSD+VKXBPjWA7Nrw/IFKkpfeCcwYOYz33JXeK0uHvWTQNAu8D7lcpNK4lML6o6lQOw
VFmk8CssWKVgP+nveg0PU2oA1wF8PUt7Xax1v+dmzQjH9UwLV0cCRs68plsFihGDBYXj0dpEduP4
0Yg4RsDiJSFBQ+3gqSrXI9R4qc/yfMaW8YvXGDNG3G9Hn4NRwtIuCHaJ3W8CtGmtNzRvJf2V02cR
9FGViYCY6kitnTch/pawlgPbQETw1UgL4uKVtebGYQGkTHX3P8+KtmZqHGzfgDyFoNJh0z+qxikM
eU0JZdcrWpsAuKASM3q+DOsu7NrGmeLUdZuzulTXIWH+vSgNpl7bBupdZvW8KfaewDuJDrK5e6Wn
j8H8UJxNrBTuED/817N9WkMb9M+JZ0yCisGQyYtGMbgFcejFEd1IwtvNiCk+vIKtw3gqEzs4kmZc
UBz0jgagw8JjkYFlx4+pbW5YVH00ZTqPrBkHMHxe+fD6S5pxcWASd4Pq4aPt4IAy69qfhNYo+UeP
W00J8YbSV3/eev5uY9HaOQZwAGVlt2l9PHoq3og7XhKuFL7/6qUNSGpI3oG5Sya4ZTUxFRIfN+Ef
Il6AOAh2PT3RWcRxNMyf6ep8f8fZ/0oQyfdtBjqKrHG96BrGI8cKOoICpbaBUpsXbJL8w7y7U4iT
QtQ28VzSxXUMZpoB3432THMu3shSCTcXLYClHhEI6evVudMzDtAay9fdlaODxd8lMY8RZL/pxDpS
NDLJqwU2gq8TZQS9/VCrbzkUTHYdpiYfAKkFGUFLDGMq1P0eDCpy8+yVl48QYHsZZUX9/8LJyyqm
WEoUZnn23mK/BrwHJbWna1Dw/afkhc4UPq+7UfOhuYrEo0z2vGDdrI7vQWZu1yvdnydK7A0YsQjm
WrgYq7hMQaND7fdWJvHOllp9Q37N/0zIi88/6W1ttVJKKQ3CPL8beQ0RmjIsfAk9HTd3FXDdfdEa
IIZxeLW21JPi8S0T4XmERKdJdEOfd1q2UowWWfoxHAc38TDXJ7lu52KN/qYpft0XnmJo91lbDjDA
9OBPliwj6Ww8cQt/HvEv29RsHE/FhYESl+fFlPcuaf1wCIti36D+dp+wbpSAML8w8D+TKuKE33Xg
nJ29zg56yNKXbrwiNCCDAz8lQsbFTpFsfyPFBgMSJahJrvEoZYtByGdyu49Mt+ETLSYz5GT1j3ma
DBiu6Bh+cruhurJW1AC5iU12afI+D3lny6aUmEVGpj0puRBGJIjxoEldv1jZDj3YFVbWW6l2Zgdf
Hs2viOUSIYpp53Z7OF+YgXcXZG49wBq5woXEMWm3Whu3qVwNp0Y1SD66jgXnMiioghG3eNkzseZw
cEwwLGgmI6DN5aNAIAzSWx8AwXumijnWc5IrqlMUQXIityHQbVMoUbX7FKGgvT7wfjSQhRAHM6Z3
qWMjXR7RMs5cEnUkY2nVve49PQ9LHaddBJnPAnDycpInRPQU5w4vOVIWqeKD4z93w9TGCKHB1Ygh
NtiWJ47KaWUxzrAsSh2vFq/AK8IjqkDIxZ+o4H6NuV7ZQP/MC14e/Qodkr6UrtT73on7oP10x88c
mkLcnNwpQ5zKTNfUOzD/A4DYt9FvC2VzUBOjn04NVy/G6YPKGzqfg8D65tchrWq7hqJz8xiTCq+e
Ncx6KhI2AhZpOJnf/gDfqhSOORUYnNzJ6hYAkRobUsRUOXDU0OF1HOtWC4+uL3P3FQK1u7Nr/n9X
V9YVfAjQMM9UnwgB9F3IiCHgzcPutuBr6v7w3vdGjxUrZazts7D1jfme0zz6R0x9VF2gx8Y9G+i1
XQy/nvnwXIh5WS8TyvOGjZxIFQT/ZmZiLvMR3vwxXtz0beOUqgLSB2BtZh5BaL23JFxatZxKegCW
WXtnnnOf6qh0b3K2G4zyZBSMrciYSi9an/z95d0Dj+3c7P9PHYjlmiu/YkJg6dPkQkEaQtbRJVq7
vecsEp9AnLXizR5+bBNluw+4Vn6aETqad9ifFadK6HAr08TjeZUki/UXAIRg8cFAlD5QSVxVwxgv
VjtG5eJInsCsY43wokDJY3kVmJckLl6+fMQjy3LZueL2dG+XkmCQbLBTMOXAmIsUO/KCBy/gQFbC
aeD9yHCWLnYXXanZavxYu18/1uBGyMZYefYDHaWEnZ8ZlbFmyfW8rrRcPH10pGbWCpAsCRioe2AO
r17avJs4w/TVYEVDIbAyK0Z40HbqtkbpdccV73jjQS2NMo90kVAShsoXgU27lhwe/VOf3PkRdWVP
+YAT3XWP4Hex058S1O6uynYk12Kt6r9AccvoE9M0zjdQZ461xQjijRMRKLDqYbnII1YRdaDmSsJq
4v/7PvZGMXCFBlUiwjab720S+WcH7vTwRcQ92RYYC1JLzWo/E0ypiBs3i/NdNiVI0Hh8yq29tZ+i
cB4IOZlYtk+i2WEHm4wTrgfcUeZzVbxH5jD3fncXSVfygXlFo0OuJbtr/OrH0h2HtdTaPad/UgNq
HJO0WMhFMQ3qzMPFxzFQAs9NNLoG5tkatxIy0oIAuN01/SVywRxZSe963fGaP5AUiT8xHFZuyLSg
7P4dkYCrd6va2QamOo2Ylq3RvXINuwx+FLcBKXPeauGo9smyxXAanra/CBxeehpyjw+QqE1mqxZQ
a+2wjOO6/jjnFX+26lcEbwP1PTA0eYq2ZvQIEqCjphg+4K2LTU3nBcQad/D87i4q9YzYfZfwZ0Dd
MHqz9yojJd4hpybhKwki6YvvDTRFLJUsU0KjzmCP8LjYTHJDoxIygXhu9/HtsCCy6o4QkGeXNJC8
LKbnw0VQgDunTuntI0i9X/9daz1sdy8k3b8rQ/WoBDrt23KsBZjsjPhM9vqjGChUGG/MbtrHwRuM
a6HF5D5Xa929yncuOyPeyQ2W9dxtxovNaahwu3pPJAS75/OgFUWwHO80pKbe/B6ec0bRW9oWCmd9
P3GkQ6DG9zlwA8NkB5lHt4Vwo7dw/P24qjMSv0x/+x+EEbSL4UHMitrXlFu4lskkXfGadJ194+yZ
YbtNaAB3RWTI6ofzmf7fZYEqlYnBxiIEZ1xn+bPvqVPwoaFmnRJiBSAervudpmm7sCug8fDjhGWH
NXPy0YBzwkpNkcn737GTEkv4prFflSwXiW7NY3J+HiG06CLcQdgoS55aNojTksk0Y069++fQK88o
YkTHqZdZ1VvQjMJ8iZzcW7MF80/ilg8HrXoIXnW5VmqdvKduPCQpCq4gF6bRwCZEI7bH2Q7yauZi
NSURaUEsuRmUV5ow/rEyXTo9bzRtr9nvRAvoLwJtpixnyEoExQtcwKeErDUpn6eL0/KLqxiPk07p
TtQrRPzdi9k+B/C+UNa1+QaJKzMVOzJkCgACeATEzbWBMlRuk+NI6xPOPmPzvCSAau5LKdIXoznE
0iGPzTmKall6PGKAjVsbyc027p5ZQ/WpsU4/SVxbkVXtnCFoFKahidz6dXwcFQQlEWxNdog+AJkQ
7d0wbebLjhphEH5nmufrdmUhTLvkKZ9KPe8S1Bx4Io6f7gdH0BjsM7rTzqHnJQ4GsaqlM6Y/PtuO
Z/YujmIY3N8vqfmp7dEsLcXxT0FiGQaMTjN0GLbbtjHkRnE2+9y914I2lFeYwsll9FLMHONYrDA7
XSOV+Hfs46fjC2ggUQTHlyocC24jEqZ8UEc72oybUf0UVVW3e94j9FmSc7fgn5SwpG0JfRiKqU0P
/n6+k9uDLFJDJfWsi2jebzkbXFkcAillcl1ih3znGY1pV8LMYpeJTD044VkozdpehRFV4iC7gz7t
0FHfWRsTUv8wezkRm+jEEvagVt1xU41OX6vYjNPiUi8AY5b598XC8/uT3iYhk7lJG/OGRkGPXjZi
x9yFkywb6iqSWyl97/dNGD9vqrUPOnUspMk0CoLw+VK/VUoJCjzXb6bIYmgAKfcMb/DtwQidUE2h
xaUri879H7S2FVl5LwbvaAfPlDD8VgbwKMKGdZ1tB9fEfHo9ab9FJ/aQUuu/QRPtlqqg7lCZUJ2V
96UjVWAlW7mWtM8DGoTOzRgKgxNiUvYgZNr1j/wweSGTuAK+nd7Db/hFk3wDtDPlpErHFz5bC3ln
ZtIUwU1c3DPQDEkYmlFGd3mTZaz9yWF44dSbvgjB39X1YUdQbmyrU77gcOeV+7FHOt7kO01mQxRX
VXXBzdvvdIL1CwsBPKzJm6c9r9MNPDTZIZjTF1OaJBcxbPxKbay4tu8pzvYW5443NADC4rpNqgUF
JmbPDHyRz3gcMftCFI3sxL0FjZQUAWTwMSVek6U7M5IaO8V394Xz7XgplWqXr+fcLYaqQFR3tHX+
JCAgRptXzXqGadst4t+c0NBf8VDiQUaiZa+WaGJt4bbnV3Y8LcV73JxrFGzY/8TQ72gInwO4tKui
6tnUVGd1OlZZ0ExduH5jQOwTfdxI2IfErE7fp8/OYFOWMlRA/MKGqxXhq8v9LL2QPpZ+px96vgJB
qoezM9uNwzySd+GJd48MTpmxicUCyjqVA3bqwzbo1F7ku4t/lhLvGfohMH0PTTkZkhmeUL9JUNy8
serepGL3OJDQD55QwrKhB1aslWAasYlwix8Kmt0BY0lJ2WroK2bbLd3j6atufqTU3cGxkOGYv+Mq
lknVVdYRI2KXsdKq3ufcjLNsAvzQWWvAx0KiYVafwkPkq2QViDem0lhysDpA7omKH16seHWspR8W
6cyIc5KNYM/1UzlfmegFYRFPY9u6oWj7ZB2kWLVUInhoTVhdXsK+nZaVbA/XKit0KEwvpI3AzWy5
voWYBISyORR/Zy9zG7M4zwzzwHn8SXUrIi1uuEvR9wSJOMw+H2FBm5ZSHMOnlpsXWNZH23ypZxT1
N1659eGLzXG0WwlIcVTPw70zPSVTQ3gAuCdOqH89P6+k9LXv5ywR4UzsEdB4j4KK0XKjayIVhqqI
WZ1U4A6KLogpuPoIZwfrr6FmXpyaTuvkI/WhPmeffOyLwIpSiISyiJfDLOksxAYBlL0FP8f1hv0Z
n/DfqvsAw9yKXfrXfn+lYLfRP/iam99fdhXdm4LeAOq2LcLjlmIOobDJcHVJeQCAjsw3fe8U1VFC
MXkfzrVhoxf95T/oCBPnxTj69Z/KHsHDt5A0Pcs2asqRE6u7ETrEAXNgRwzCkWQg1ma5BXb3OtSa
PBwUvCOAs3ssbxH0DAjIo2PnmVMeeEzGvunctM6GkSsseZcAQcmYkLEZGac39EbLuj4aWEaWGZaH
uP7ttWbYxdtqp/pdUGzIJwp05z4pQlffcxkh96/eAqLSM83v5nRtBsw5WL+k7WVv4Zqrl4Hb3iqU
oIPppi0oLAvO/vTvIWFZ2Q7q2tqEBoZX3I9geOANrjDPy5/4I3YgiNQa4aYiEyii86xbnCbYSlCc
PiTYZe6EFe+vfJq3LowwtkXqlU0HFtek28GG0EbwB9vPVi6YAfRBsHWcTUckyR9tWzeyTNjW5NaP
jvXRlJzFzrd0NMVIgFRl0PCezMekGdD9tsWuhyzAunJjD2PhgoZX07C+ReNaLsP6EkpgUBjlFRyO
VZAXykEgO8D51IkHg/WiQ0tcWOGXf/pnFftMQ6FuFlxhjB1wTv9tAhb5rkjHsQK8CL+1l6krtZQA
3OAUF/MZof4HOCYnLG/zBA/Pv+gpPX5TmHoWtuk3GLL3VpInzedX5/7w9JNQ2z/Y3pzcefsuIjry
BVPZ4Du2b4r0I0JeBTPo7Qj1sroNZjNujkvBDuo4Ft86FvD5u4MWeTWO3MSfmi9WNfJ0zc1r3LUJ
r7XzfI6MemJ1LT19XEEvNBKwKgYtVMMCvKsgCL7hdshOag+KI7HONVGMyUmo6ZupfRCZvZdmS1cn
BDwy1UBPt7JKTIeakG/QJzCILK22898T0GHqvDA0lI8zuoGp2PNCJbahmKi0HFdsiRtYiTYS4u/V
vFJPEec3oJJddqhXS6jG6+6X+NndoCGsbVIsAw5Xvsb3iK+T2zdjfFh1Z66Yr541LQ7ztv1HCXP2
Z4D/YUGhYwEA20hoRgtxY3+jmjbZST04W/iHYaDtbPXS2NbPrLTLySpFXCg8f3GoHIdMI2CwFjoK
WBPOWNC2hjDPceki9xufVZAUzKlSi9faiQa3DmlgHXZVVWcemNIDFDh81blAc72I5eU3OpNfoMO4
2nOpouIz7s0NXLwlBvE0+UpzAkB9rR8q/NKKtyFqxe6J89euXWgo6a3ZBmIXM7g7h1XyIXFG4nqq
zO4M1xScynsqvL0E4G1MYBcXThfnHaq7jN2zm8ZlgpwewH6IAUopICF5jfO2rV/mwoMHZ90QtxnG
iP312UzI1OupLbMf7xLdjBw94k3p0UQoE3QGzOL9myhMpdejdFvkJqXeA//f/4gp9Ns3DMpu2s1r
aAuq3ExtdaD7z8raQLO2lxJqSuglx/ColPK07HDhDRKaU7CkVOCkwauuEeE0cf2BR+EDqd4I+x/B
HE7xnlBULtaZaw+5qZkmek5MgxBKvV7WVEfwRaA+e+tirpPPPJgbOx36FYcUwTw6SivhY3kozu8y
rnYjWvUlwfWNeVlsHll9fPIhS9n8n5mWY93E6RW09mZ900ibpIxqHMtnT2ZCA7tjKLZW80V1AZNA
3GmQ+BnnWl4paOQ/46ar0a1QFzfaq7HTY1WJeM9KPCww29x8qv39sSt3d/ptbH+hdIwj43lYALn3
bCHlGQX04eF+JUqaIDDgBsE8OnHaE+Hk/5zE/Cdg6OUkj3CEogvzYs8hyFtAuFl3c2X/noPtmJQ2
0ovjiTSxWnUkoCW2b0dFraZrNDJPv0qutf55oXHmBnNO6N8krcJrYVIrvcr1dXq9cyX63ph6smfq
rX7P3zoYacytR45rFxvs+Wo6nNM18GNSPoNyVaBV2Z0GybCrnf8wlwM/7PXflegbWWuqxpytS1o/
oljR0DgSL5nA5R1nPQ/Cc1MaTXqkEqKhJol6oK+MyOcIi2UTxkkcNeHiebC+IYHEzBMuVfVgomzW
aAkBiiprFsZq0ERFSwp62HV8D5f0bCSTQ8Aib04hCO5GV5ImJxKl30hSvfPmCKF8e6NGjqjQ85yz
9RzzZMg/GNj90kpBBdz3jdoHa1IjKfpHDgU80t6XK+p73XkFJQ5PR/URHtQE1kEeqyrfxqmdJwgX
V3djNWGDrLbjUGil3dQ+5Csss0uoy0WctLwj9SfG/ZuCP8fgDx5PL1tJJcPkMNfJlB4SyxFuw2X7
UszkYNuq8mBZcodDxi8VkRvRynhCGzNwm8L+Ne9t7flrAjrMHAgJRytBJjzcyKRgUi669+m6QEed
5E1h89TEmuxnkqpYzK6WTM7KJfGBqb1EDR20yY+rcaUt2quqnzD4omg1SkxtMEYE/w9c3xoGLUX7
D9/EOjAmoTJYMjMBMWdBG0DORiDKGGG8f2pCpzA9TMuACemHNr9t30s6ktLuI+V/HdE8RauDEUZn
VgDsZV7wwtgCm89lmRrEY1RPYWvkzpcPVQmwhBflscFRjAu7C//8SM4qjxRruS3iXgCnohRFfPml
6vT2SPGoZ9fjWszon2QAriDh/cobzl1e6NNGRSnXazRwyAEss/zDd3dS8bFPRFbSbNLl62gE7aZF
Oq9J8erF86HHxNjQQIONDXVYvSMqgcqM/evO3mPfa051354BxV8FpFqt4iCOFkk2TTiJxSIakSRs
RlLWw/bgAB58yLOd4V4WPGpzXsyks8/TLaoW5/PRdDWoo0c40+ssFphIL0MaxbKOYJgFAzb1KChn
kpZhVv0LuPc/anv8I7hrCA+W01jviw0kmNEC+tLKmAzw36KK4dtmpexReddr1tFke6FBGvAEgsou
mYm0E7xDOol3h/V9xGztHfFnZsiUK9d0bL9Epjdc+vGOO0rdzUlp7DRgODbB16E2FZHNgPEobNFY
jKX4zFctjFxlhiqowHjjFYh9hpn31E/weqiYvOiMP6kub+UXKevTIYVfhlVZzESuTzMG8JOjoEQj
5T1zUv3RWuEIWQ/mMewxlBKX1jLCtdA29Fld9laUJk588MaWq8QSayAVHol+yU0ObklANHn6irVr
eoYLRRgcLWPLOIRD+u9B7KQP/aqqkqKMS1+/XluHVQABg+DHhxM1Y72ewQZ6JkcTlKilMC4fxOVG
ir1oe2qxxmRYaRJa/mxs2WWjuC417DRynHpD6Z7R04tSCwH7Q+TRH78jN3qwfKlpkhpJUhAzSuLM
9VDBL80fJmYRmitcpQemwcN9PDAHae3JIhM2q8/HV7vmynVwKFXwp4J0lM+snPLPyJmG81JI4rwX
LCeE7yDuv8qeHmRk4dJkogLTJXJ6yhUIX+69sekLXuQ2ju64kuUWop3lqKx1XqPgldbHl6l7Jce3
M8N0n4t7Nsok3R1Rvt2Y0TuSqkdTKSfFnSPNbHkd4MV6vMU5qKrUVwtsn80RU/8uoAOD40KNO8t2
yo8ALjkzyjOKJp2trEl8q6IV4gz3wrwfVyTR04eiy33yKo/oTeewupblURN1gYWpCg6bnLctBWn1
4TYkwY3x/pc8X3aLATRmeNzuio2dNL3u6pIkb8dBgwUSxcIFbXfXnXG5VcBaFkoOZFMwpUpWWtye
ndkAL3HQ2IlyXo81VMMDT7Wm1lEStcy5hBhy2wVhxJH0yvGSHenDuJnoEocU16xD9l4fv8n/oklg
L2Jg7JIQb4WQNRACLeEmkHCWpEEzrSYMvXCICAwdeL1FGUspBPPHC7nORlBoR3X1XO1KEB/g3BSd
/PLHgzNctQoFYuzE0djgdlvD2pFQoRLSJF/s4ug1nHwezEs8qxB1kWQNYw3JcVhPP/yV7zpJuLzR
r4OMT/dORnoOvvlRZJwUxUDHKpWFHTKkKH9TogoQZlDXRXg69eKoRdc6QfdyuRATpGlzkAoiRNgQ
0teIqwZsPLL/6sYvMzK4OpBp3p9EGREvLiJsgyBFwRT5NMY6dXIXoMdREcGwsrvk5ZNZY0zoVTk4
0bK2fEk0E6TQDIsfaPOmcDr7psuazB5R/yo40nMRqHDAKSb2Oojm0waA/1xmA/jckcCeaM2aJlpK
IDTXgdIj0gIyIK8Jdh+F4V1Oi0lGdwpJAjkrWy3zSBRuOy45eRM+4vREtSftvBVSEJVFrJU/fUJf
2pFGmmYJdpCPYkBGyDE7rnGsHf+X6YQUULs9XPLG6X6bR0buB5OW+K+pXtU6XBYrM5ZobG05YyXm
t2wMwiXwBlhnXFTd8kjm9lV6QuJV/RMjy/IcKFgNRKdepzDrD09K6jdM+eWNkFbVnxAQ+nn0pSmK
v9XeB4xREYJK2uDW4tpkoMRhQ8Qb8TdlLjX3DcNUNtKyCfc9RdQZK/EBHSHCsvQkOIYYiKl2tBw2
y8uFoUAZwjyivCz1+a9jn3S/ejCyGRDtM8EgffOUhwm0vgSGcRUCfjqufpHZF7ozNGRrugX2gPb1
zhHElhGCy6WWd06QoFEqmtf7UhJBcewlSrUwO+r/pRRrBxnx3BZiuHAG7X4P0IhtCLF10Vy7siBS
YFjRX66Ke1Cg/CTjDFwXDnljv8gDSXPQvJSaFQqeizibqGn1CX4og9uXxozOHT1zNS0NqMXrki2+
rAXDFis6K1zNN3xzxZN0chX4eRChiXzRNdTGDGHDGs+vpbrASSArcG4mWLvJx6UJtKan+Ruf/sZo
mbAa3L+ySF4GV0rEvBiRN4e+VJmrPn1lLgI+H1JxKTlej0/QK4CqpFCwvYg3FuCV6co5Q/VnPFCM
lnfAoZT4loj1aaak8XykJIDhNqHYfNhFh2vh77I3lf75z0TWDxTXFfY9S6O6vYmKeaRumXrNcWUW
6Raq0pGNiaz10lnv04uFLwiN4kgbVnQ9yXx+O4kwOF1zwjoJ5PN2Wn+rko2EqfZTd28Y3AvFVg5x
eWJma+VRFiwKGB5vS4Tg/J4kyL1azv8nP1P2Kjb3RqjftoTpaZ8mmS6tH3suFNNn7qdgEJA/dCtf
O+Q3BQcr39GYYnLtzMM2fKIvFM0iJ4Ko2i75VqYemetnK4uR4YLzV/IV27DgrPpEgAaApB2FaCyv
PUrsVrIjh0P77JTO45qdiSYhVb5605kse+ZZTzSpKbvlP/IffUKcSub8sWeS3v2PTuR/yUocgp/A
zFMzMtfhPUjHQaVtMUV8Bh/Mes2UoqqwO4iR3OAM6rwjJi4gooqFm9T55r6MV2Dtqymm0pYZZlZs
7OYPKEgdkBdwmSbmBTE6TcaC57iJIA+YR5mjt1EWU7VVeip1wSiyuyG7gM4bOX5f/UrwcncY8mTY
MununCdXXpU8JBQ0wjaG0lvCznqdK8pexoz/Fl1UUnm716mQROXiT6R+bKI9hgHHsnDMHRQH5/Xb
bz/aUqtXirSx+Vd1jLk7TwxJPZojQRw0kgPk9/WA3ej3LZx9a1FjUI0gCw9REI0KkEqRZIuFnoKy
DFS9ym26dNTe53g1E7xmTbm8uOXbDdR+cRotcmVW4dWN5cYXTRlYFWfnzyzVsVnYbF/hHPtB9KB7
x6NHoOmgcYIiBmtJ4T7A/ou5jB3lH1Z1GdFNagvcpBZ27t9JHvPgza8BnLEuPIAIt1z8cIDqupcC
NuE42xI99PD12oRVgzjv8/hz6HoEfdSrUXvrhAjknZclq52yUoVNU/cR4A4t8C7rIQyt0Sj9t9NO
UVN4hoBxHEjoR3Ggt+85uEv1O777gCUflx158DX2Oll6jGeNkHsqzzJI7kPz7uomFakwnhuEgEy7
vPwRh2BRFd/ENTMexUE0oyad2X3cwQubxQ8Jt5ble6/a6y+nZoWiQpbada45UkfctpeNM6I3gr0g
kiYs3CBKq2z4YUJ6HBaKDzzQb7bWHv4f1SSRp8U8rqG1rnWMBzhHYU5kFLTBJK9mzCnslKp/lMq8
r0iG+HQXiqK6kjsgoLIFs1uuEUB1sIKV8VHPSEEDrMczV6+TJ2Qh0GQ0aRL1ztVC9H3rf/QDhS7u
EB/KJg8AuFR1uivB/8PkzMMbRJ1UlaPlzLyhV1lwJQ8lSVzXZQHYo5eMWQNTbn/EIF49fEMGJrxs
WmtKntl6U8S1Ri/3ToUGkPlOfXEF4sZNwHpDuLn7i8VA3yzdt810LH84J44Nllzu0CMa3TdWeNp4
Z7LRVA4JeLFRJWXIfBOxVAYRMfPwIBxtWDpptRCRLOWVXbU9G+YFV5vMjANZo44xLLx4vG7VCnCp
1uJuV7TEcUuMw2NIDj6T6js8bnsQDxzywTmL+SEedp5VlOORhRkJgZMUblbajwuYdyiYelPJgLT6
rBlOzmWCOyokEruRiG+ftLflMOphdpWhnI1GTfC3x5i0rIMf+gcG1Y/OxeNZf9Tq8KrypC1Cch2f
T43W2+7gkMUf0x1qnk1G3T65ky+bFA49BrOWTOnH1O5UT9d68JhdKbN7rx+v2+d3L2rVF9a1Bp5S
zjvULgBUyPZ4PkN63eVHZR4tjNKPWPFORpT4vjNO+egaJw1W+nXDw26Zi0a0V295yWs1WV2QCMH6
uQdcx/btfLbvGjhY6kAVJeP5bzvSoJrd0fAYcw9jtCtMb2M4W+J9SXxH2ERBPzNT5DDenTKbksqP
FZvGzHDZ3vjftEYX/dqTAzRy3pM+piJHw8zxzV83z2wL2vpZjXDY/qRdggeVKNbhWu2hjYfLl7W2
fD7TNhT9b9c9em+7RlaNxD4AttgeC4aT1+oFEpgFYdb5lDlwMoETTZrn845Qn+w9c8wlXt5Pgq0q
rsuvGPhLvpihGYO98uxD+tjPgRvV5Ftg8A0aSUBzDwlYQmq+8/4eW2wxigcXpxJm7M7dguXUNpH2
JgAoUM1xrjdRPVonnwkRGOR6KvIC+yXcOpsLe3UcrfnrIF/dKKuW2BLEHu4scgaC2AKUgecUglJK
cQXG531FTLQPDg9D80/FMRQvEunZm9rkCAn3oSS8LCuUzgJe3SS78WiyAEYXzyRDbgNxgnluIPVU
zAQ4V7GlO4IhhUjhefgJJb6eSGc7BAWnT5wVFz20zXXsSRGitoci7XF7yVoTrYkQMtR01tiJgwCt
udTy3wsY2fReZ/BfCMcStwy8/HiM4T9/itOzHpdnGu2CEbWiuJyqpHYlzvtEvs9nSbZ2fScTR58T
4viImH1VaGwOo7228FkmkAkQE3LM/9ESfDvPfk9l4y10DgigbpGyUYKcdTJGzTGxv6UR5V3908Qn
qemO/LFg9pJpvkgD3NMnC6iGok1cBj2jxfigwZif/lVtaNpEkQiBC/UtyqmPRBLmR460CUEQMBUV
QdA5f+YCfD+wgD7X1m37IpXOmYN5BYEQJWZQIPbs44oNfb6XKnk3GC4+9IWols4lNGa4vYZNieqp
gHpbsvzMTkUADbqdWemLj/nxHM0+mOuDEKm15OiHJuVY2VHgZR/6VhT+iLu7/UD/r5BiDnv/ugqA
IXJrXswlvIgfUUODIHuy4uc0uD0j+1OH8jwNZkXq0tT86hl5hq2U4Gc3emcZaYvnEfldkOxN5GYy
jhhWMiqs30XPU8jpFufugtX982OWQIXT4YbqRn67VtvYK1bA3zwDjcTBepX5PJG4SaOEjDtlKgoY
ESwEKN0K5fhm8y5KIDEGIUt0RwnkJGlzdQANvqa0awaDFVLMa0pMVqfOLvGK0GCc/g22EjDC5f7N
6DUfcpO33t463grtUI/FouuWWqRwXqxGkdf2EaWy+7vEYsSZkiGUB7iWABbmpDsaxvEyQ2B5omV6
uL1DR9nP8qc7ypZH+bN8gtYm5KRfgMJ6odeOBfxBRCSCDuiRy1YrDYM3SIc8irHq5nu655Vnv6l5
GXu7/8pI0w3JqB2lXLcegWrc7H1MLlV5xCGhQDhrIwNI0fDbnZr53iCLXbkiZg5cSslKH/hclqhl
8bjqU/+ti0SQs1o8E6Vf+5I5+eJm7/3dcRYRdWoJk2EG478CNOCuqS3Q2NSGN1n1ETUosECBEtQm
KcAXKV77UebiAY55MAtqsW9ezK1XY9+edtHCYETaXIeGmFx+c23bazpRiSGJWOCoXsshKUuQn02u
3UHgKQ3WIuNIw0a5T1fyJDwOjyr/SVjDTQDeMhdWM8eNCZdfR4ulLVbcFRCh4O30FJMw53Ujk2RO
Lnzzlra2gYbdPvimvqheYFBH8diXr6chHo82loDzQXquyykAJqvVXOxylx7a4iBZmeVtE1xhj30a
Vdusguhd81InlSIInTAE7cSwPkJYBARRd4iiRTRjC6Vu1MoC2/yk0NVlHAOpxdvDOqzkQu4c+HA5
fnZ0H7P88yoccVzw/mhyePbV0KLH/NcA90UvQp5d+COJ8sLAChYeGpJCDaAO4+To+ioUZqeG7l2N
OpRVtr57IArpjoxkSh0OVLblBQo/HiR/gIsa2hciLZTG38USy/5bKsupJpTAwMzKYxqsZZfMtKvE
cQrJ8dOKQCNYmSvLBD0bAUBUZ0hO/wQkn6CCCJ1eL9pSpD1ZOTDQ0hW1HCHELOMlDvnTD8gblA6o
y7Mg9ROHdkNiibKLJgahFoRLynFp/e6Xi4syydVNSMCtAy0K+KUSpBmvcwRzQr3iavfaXulsjUdl
926epdXhtoaEu8Rz/S3uWsWJPMN3QZTGObIzvBdNu3T1vKVnU3fIUSxKI6ba7TKCGH7cwzUnf+kz
vkLEZcCxjSa9BVY3EsGeSEwi/8Ys3LapaVZgXcVFJ1Cp+GO7bC/y6IDIxw7NPdjHj5Cx/e/uZKrG
PlWBa6FPh0rbtzzDRL111JAlCXRtjbTyU00lOKqF4wNSpLcjx26e8lM6yjNsKJ+rxe+paC40CYkK
Eycw/873Pnn0OA6Uw5fEdWt26Lx5PutrGmcUkOnm6F/uKSqEJWsyUa1wNOwYhMeeJcVqxpnm13Ro
eOYrco0gt+Naba3ELyQtceX99h72k2/iycJfET3mQaBPxu6Oy44+fG0ieN/4rnPr8AUbDvWVGWpV
SnT1kyVjaq65lyQm6PCJPOzw+3AhCTu28cBT7xpSWmp4VoKCgVOcHCR4rS/cSJ8irmyWgePOtHat
MJEQmwOK43NN1XMgvAjtKmWjqAqY3NXowozl9htvXMFr/rgKh0CoJIm07Qr8HyJgOjH5TGOAXRED
vVDFadFB5Ucuyo46ZsPH1hcjnRdjRkgaloToUh/fcp78SpoQmmQmLkZHAa5gpCJtOmO3Dd4QWmC0
vgpj3Uh50/T+ow4+7JalPbrxswHXvsIy/1bJwiCiziYOezNuDavek7myGO3T+CRj4O8jGVS+MByR
iNwOkzGdWWXd7bT63U9EuTSxZAofo8IAo0BAxzUUNNiPjKBigNReAtzKJVzmp7SXUK8tdbuHzLI5
Tf1f7S9doOL+UdxLG4wKrChr2Z+uwY2kShTWj8aiJeYgBLOjxrYK5wJ5cN0zVZn85SsP+rglAyPQ
KJqjd0kgTLcj4TPdFCE068Fd/tdplj6m/cRyTYbUjcSI7kToYzYy0tYoVTEdAkr00ouDloFUrtk0
CzMolchndwCJNGJ28LzptZ17MmX0vjnITuT+x6G4PX/GJ/4LS6bgDPheLi80qzomGOKYiByGgRoZ
LCkbY4TrI0eF001N4iabzSCV/YMIIfsjkQIE0v9DiH8UNzkL+5izHyd9Br9HhUK2V/g68Wsq/3l0
ZlZyPg8/z7vSDo/Q2QqL7fxq2ZlBuIfR46596geeM2Pby5J5DG9BiM4tGwEdMOVQq9AawKLiWjEY
J5nah3Lt5Qdj/3JpHwQrkbsJas4y9CNNPiI1c7KOOo2DNQ1GXWE5uwCP4vIX76xkYyl5QsvcLmFT
ag8NY1pGXpGlUGP0bsGWJoa46oNJuAK7czGnVvd/5VbnQH9xWRHLvIL7zeLjJQoCARJtyPzVZbk1
3EcKsKmZp0F7jJz410lekuXtQ41g2j/yoXcf41G1tbAVeuDovuhTtuFrgA76oWbFA0jqt5vLLIwj
p9dLuAA3IJ3874kr/XwtzKmqLzEjRO5KQVwWeV2I9lyN/BxeawzzGbcpjVTwAUcJqrJE625QKBrE
1U4TJRTpzXdjnrsmC5NI0Z90umjqVlnYde+fZlEGMuTtRU3+2uacredeONtJ8musEp/whwQeeP7V
DsDbA4gjGyHyQVJhjrbRxgbvlrywIyMFMR+DLXNdD5/B070sWymrnhZEH1k2ovJJaAc/Oyw1KBX3
vek6flFnPkkkuy7TINhLX0m6/5bodGda0EtZbgZOQ4k4TOVbdqNrZ991Te6HhkjK7kY3Yi+81yud
1KfN2dfZzMiAf3wWcgzA0ltI9a5F8V+0zYziA0EFxQX7bmC6b3qVi565TjEAtXb/OSrgTZJp+b8h
MnR6jjtBQr+KKAsbOgYPN4B/eFohsml7VwiRPC+SdjmzOPDnEIzAIYFOYtammblrG+YntEKsMB/0
s0VJC+lVr4WjJgOC6ayLa8XCTLtfWxFpJm6abSBqQ5Eo0dxefVP5sqQAXRTOtrBBUli/iCOBgOQc
eQ3G6G7+3YEQAoS6fmvp3MeI0ubZ8UVOPsvAJAXuCUqzCFDIjpRy1Ho96T0ErkGxv8aT4Ng3mrNS
bAujlV/639/7l83whABdYBoUtXIH5mdulWGc0NeSdz/FwKCRCVp2NAhhovxtFSJZRYjm11Z2Tc/I
cEhz3Ji0/qVPVJU8BLPPq2pjyEuz/aAUdSwSH6ZBzqIvk1A4vygb3sqDofqd5xKj1D6O0ByyrG1a
LrtYm+0WnAjOFJBw6bfqj9RLV+RW77XQqutcFRmqptLnM8AkKMtjQhG+6VwT/vCdl03YZyuC1onM
AaUrWnisNtgLX0zJ/xF5amOSVYop6FY03Gmt4Y9JZOnhzpe1W3RzFOrCcgTt9lco9779ps7d9rRs
2l6X63vhi93Fl5iJ6sb3Cx4v0A7C5ZFskW6cBl0IsdDbeKHntWopeihyyjzfnnxE1cjC4mMDctC0
N8UFFsARHMGKEJiweb0eH0l59B963kfW4L9Nx/uM7WF1yx0eAkWuenIKemv0H4x4/UwegXz30QLW
D4/xRqSYxEfuz2qt4Sv8sNKLHAdU8WrSEiwSuuqg9Nu3l0GjeBC7oYVZR4wp8ndsb0wTcuEwoM2i
H/b9q2qi8DV3L2c6wCSjhA8hAvWu0/L8IAwWbRAf+au8TgvQjJ410RCx5zkTHhFJVrs70T3TKWWL
vF5XHwde9nYUWU1gOo/JMPgN4/NOBD22IH41AjeZkDbN7di2IhsTzp6y3YbVb5dfpnjsPS486J4O
4lXIFSnYUomTFWPm1rscQZHMmdPB9487cH8JGiqxwpbsVgGl8g39ZQkpIQoJCATx8nicnVqekLDL
PgkvQFdh8aMXpYDX2FkoqLv8IAyqEpzJLwgrBT4uYvEcHlDthhSMITYyC2LrKNjDGPdT4M+S5dO9
p1DTq2cWZ9uCcwusP1xWQq1AIETEFd825ySld/fbbb+PrbFXn1KJmFhm11/CAc7vL6T+wkd+ypiM
Ar1Yrqt+NdRViQVk+vgeEXpNScdBMtoyPAN3ALdRluYcWx4PJZufNhGnZOdmRmX4I267aSOrdke3
HBWe6ps/UyWXBJics22eAJFh5MPG2hwcOsL0AjR+jYWV74E5xIV0Z/xXn9EZ9zmE2Sgs5IfHwUTZ
HFMU0VUN79pfVI+m2kdkbtAsKArE9T13Q+9N/nHP+IP79YtRVSyvZG6HdFz3N1yDY7Nwt8lEv6o8
CmQkf1qIzUfvek6zvLz9RSBYHmgNUSU0j43eR2HpSa1ioUTb+HXIxbN29Pfb782QPLDyDGJ3oZH0
XNX72YQ7/miTMxCVbc9WFoGaIobnvOpNnOI0gfx6wwpxQB3ti/QmKi9plo9hlS6uyQ3bjb0pzTeA
qazYByG84HT+JSznRAdOjTKy7fH/T0wfIkHg/HDYzrn5gEKLtj5BYvbHE+lONMV4XCpw9a9Xk5zi
9Mccif2avSiDFfNERExLpRiXFMA1B/CPxwQet72KSw5cvvTrE+mKUnL+zgPfaDFsb1eIYuJxhOo5
AqlhK+0jjIh3itAF4QMut+vo6kVlekcjlu4bvOBRgc0AbvvTEdvFUf25iXRMKruLXP0eXpxr+CfR
Vg32cJNxIaH0jMbloBb4W+g+oSqyiSH+FWeWLqsg7elxcimGuRWXnt8tbmWUHbbQ7lUxs+MT1Wkh
GENilhCwTCGaxk/P94a80N3evEVIDGVMRPeMyloy9Z4+Zc3ke51rDBCWoLRy0l5ZWrLDKs3N8cx2
AR4wH62sKtNyvIceKIBe7+/YZQnCi0+pZjjvUKROpDZvhY11ySm60XW5v3hCKVX6zwtdkZYtG72I
7pXjEk09khDIq1MBwXzcUnXLI7X34DkIFICPONpmhEtp8+fIJEVUiCEvb0FcHnfCj5hEplchb1UQ
y/WAGVDFFZ6Do6+3RlHKXkyB1BP8TIoC3d4KnKYVUANcwUhSvtzdUJgTPU4Z55xln4QN+g2pzYZz
7owuLhDHcuuqkprWi9kIchCDgMuSxNhCIm6MSkCJMDpJhuZJBA9Jzg+nnL6S/8x97ozGaiKPEdbP
pAqnKuE6GKZfRx6U0zzXGkjuZLm87x2xjKDt0CF4Hi2JQByac4QlE27mfLak1+9dnCK+sXjX/Btg
KSDU6omzaO+i/nT6wb0f/ULu3WyOaaR1dJupX0D/ZJVukA+zuvt02tyRgkp8pR14sI37m/VCKo0x
5EhTKjiUVa8jDP8qK0G07Ml4FAeLc0bPgrwPf/UreQd+MiPp9mOCaV3di9UeJRHBJbw0575jwIl9
8oDrmwNWJcUufnAGKunVrpILKAIWVC8fZ4mOL+W5AYoVkJfgvL9tU+hqlhOPPDCR70DBkBbuq1BR
ARjMqnz88WWROsQU8JH/vWr+bco+F6ZDts8po4Dty47sqJavTvlemhqpI/F5eA++HUF4P3WHwsrV
ot5VQizoJ0Ws/WuPk2l2ZQpl/OiPYoz57wf9kueRJ2r3YcxRyooUupoADbvipJ+4DU2KTSq0wXtR
f3oBWXC4ftPTFf7RI1ZvhXqaNtQTO2iHLSNGreMPHzEosGxZIBTam49gVt1B8GBTnY7eBprXaitv
/HfefcAVXGG0inebGrsa5y6fLzBkksUN2y7HSi4gaWlvdI7aFLsrslMKMBCh6X4AxAhjrxlERgVO
3E8rHDwrwWQE6kDZr6rrkVKhs4ieGouSyDaa4z1d+88Fi+R78KJhvis4p0s7ebSs6/ZM5LDWSogZ
J4TBnpdNdZHiKVcK4UcCS3O8wrFACHUUzKQMzQQ3lnIB9r2scgEX2QLlXVP9zXDHWwzvEVlVbsjU
4GlTCD7ZyQT1Dr9kb3JuQ+yI2QVrCyUuwIVykYqfifkbjWYBZ+PgUzSjsgHjBhszpDut3yA6jkEr
TaaQULN1BYmdOFDVfvSMkBvQHgjek9KY+6DPHbtVceGtWgcrXY8pfn+B6z/Yg95ea/NFyegitc9w
ZSxRC2i1eJXGEEwW6/XJtLETsFao2HtQyl6b/4iSDX7wYj/NXhe/5mj5yWUgpjcusydb0+ntxY6u
58ewp2hcQX0uqU5fWmJA6H+YnS1hMncwSrWQuBtCizA8loog+4SC+DRtRX2UE5UR+HB6LgMWAbXw
o2NHHOlJw27xIPtc9oOK7cSt02KNQwWiroZ4XRHA3NZzFK2V27R7LRBTOmRm8FPEX/mlyKpJq2kk
N2hKdE95dUpKOHQ2ojNBZbfa6pkm+IBdr13N+oqG01gU5Yaq6wOYeDIHqe03auiXUDk+vHgu63Hr
HlE+pnr0M7JtMMGr/oI5fCc5Y9nvfulNdp4nCQovwlTnLsG3WbQfbRoEuyxnnziZUM0CWGUy8HUG
6QR09fE6jv7yEAL0KcG4jqMoX0rKOk91se7i/sZ9ZzQ5VVX2EvwXtsYIIZGyuTrcW33mANRnqoOM
FdyYQC3wKg4TxLQR28f/5cSxquyq5HuI5tGeoDxXsJeAuCyKIM+tvysdQtXrw1Ti9VgLAAmuB6tM
9fDtDMpQOiHedR8dWdt6Eaqpg+Z+WB4HswifTbsn6brKRgYTCa718YC20a7hcz5W0EMiS85t5CTu
3cFvMOOBYQqKiFDlLQIqhPEVJiIEvRkxp10Y+WCetkxSowqd9E3TK62U+/gTaOQBMyAMbfOganJY
JqwWq0oaFKVRCje3swgneRrucwK4OTgkDKbsR/4MzlehRiiEHewiKaBTsz7YZLkhdjjlLJ0Kzohe
Z0jWGip7md3GVgZdwqYuuA0LO2/FCyXPpQaPpX/N6cm0C46/KZtA8eeDEHlYshyp1uozvRE4D0CP
EsftZEIzT5ZRzkvjh3BDueCfL43yC+3BxXkp0nAuMWrgTTwLqRQ2MPnC/sLxVN6k547Rv1eguqAk
q4qhOSnYKkShqMcsWM9KV3ghQIAnj0Ipuuoo0903PeeWgq2nZRSvnsBlmqCm+fnArXi34yPmiDeA
3L974Jj3w4YtyehldqVEKT6VQvpk17mCU36HbhQhg5WhE0jLZNIgZXMa5dYIG847NQScWAH9c3fC
Er612YJ8pymNKAIyqvy/ITOv5oZeG2v4sRmHERkIGO7wwfLDJH3GIJZyo6KmERscjE7k8VYVK3Z9
90KkDAR5qTpVGcTSfd8/PkyTiQvfHT/41P+qJ1ZqWhAMSDxa7bb+cpehAXOFNwO0vdAAsMHQvQQr
1E6MpCPX+PSak4gR70WY6/rPSYfrC+AMqXmnrnNkoGtSCL/W78G+HW9Xiq4CQ917/YHXsmQpb22L
i87+Hwg9Ck2aVup6B8ndbbuHkWqOFAgLxRW3pw0NZBhCK7hfZ4+Iw0wCJBLraeJa8R7FBuTJjdW9
1k5WMGweBDSQqOH1RA7tdnN4cZl2mrdBrx2x1Ub+hdLNU5YJJrXzYOBfPSz4YQzr7VVPFDGxgEPX
NrsAT3X5EWTk2W3rBEDiyTPHVo8FNdFNyl8awdQQ683aTBt9zbt0rDUTvmtO9Av2R/PpjpmOjnoS
ezxX8KlQuI9bGYzC1gmmMGTwuT1fjFHBmvI87Ah6NZnkWPiU1n0hCeXKKctYcbVUk8jSEbyL33My
h+mHdyTZGI4E6JSX21LzdxBLuK9LzV9+7U477ZKZKZeeMCoiZ22PRZ16HFY+Rapd9zVRQMBSqPQp
PzcniGz/Dv8HRz3JBx+a3L3PhDpfGjE59A0IpAyTW975iP+JgXaSwC+f7sZBPr+plPPUxvfFI5gV
kQpbFV+hs7QBMv0E9GOTckEo1jpGcDB4kOQvlUw2o+qDMYAtCrsv9kQBDVJhHLwo3K/Hdo3wH48x
iYwHg7bEqhDXrzgyUqVNlSQ/bge0rzLAAd8EeXdOshJ5WKkdni9n7RCev2RnB4AajnvWZYtAANpg
M1NLMfta5gewpzhVK73yZFIMHldA9OP8oTB81f8Y30kw9EQ2Jb2oLrovgtzZ+TnhCt6EEh3BTm8t
agncxtAOCLsKNdswBFXE2QY+oDoOm4YcyPwT5udFEvZc34mX/tKtWSAcUgRD7/31ApIBfTZ3RKqW
y3hRltZrvIPc4tWx5wOMaw7j+vSZSpS3a0XAz38X7CNMkeWJ9JyzpREId0gcrV3aFRY0PLVoGZE+
5KOYFPzOmtHG9o5Sensowbbz2YAKwXrlyc1K+/cxeMsZoGh0JWTTq8wiSWN0ttqGi0Cat9UanA8b
2TQ3ImT2RzqFUPhqYDu+CnPsjJOoEOK2bofzJ+5AwCyZBkRdFDyq1ZEgHWIJLCEsEJlV92lsMcwR
FQNEXD1yD/aKdeHxGv70SEt8NXrg1NlHgjYdLkypFCFKtLx2X5VqaPZSmTrz+h38pcLNxvWyZaVQ
LOWglRiH4WeeBHlkglcTJkuI3kOB+uSxRbcu01/K8Qjf3qIa8lUr5zCcKfAic+eayj1i0zFXTq/r
ttlmCOfz+d+/Jh2K+whh2DdXYE2X3ZetMwfw2zp1tEEdE1bJcKtDuy1aCoU3wwdTrtVxPb/XS9C8
m+DO+3+hsV4w/Qy4AHXLKteU9SpGzumsDKpG5KATm/7v4Y0kts4qK3NxMD6cPeq/RKGUxWffZZRI
A89z+MIVxWgw9HHCNlkNa4g7iibtPWRfU+zFiLlxddHPHPIqe9PMiX6xErV5iXQ3DzX39kzMPlBT
InAX097Am+tZqg9xMDstsWABAppIMeDo+HU2OyVGC/QHIlUA9CpJCjU2466FpX8uNTD929cJRFm+
6524upmxhZvNEd40+CFCNHVYIFDFNQby2r2YyG4Kw7CRw+A7xhA9jv3Z9jsf9Sert/gmsRd6EIaE
mdlEDhMEk8Es6UikP5oKckuUWbEiHDslI5RI43UIA+zeA68uzWx58lQPYvK6beogX1cbkRbHvKW3
aFHl4MljZloQTOlNqP4i/gSS5Tm8GaaSudkpnYJh7KeAlfJuTRZ00uFXwQDfBBeWbc9OlMA7SHir
dcm3YCmiIaKqB2tOP/QkSGet6H0c9XELezOdeq7aGDW9io80YID6DUMuHJp7VCWoXcockp8x+ZAX
sq6udAi3jrwb/+bDwHjCQQU3/eQhXnnMcN1EcnkGlVWE9w7+tZIagWTUHzqIcrXKW4zIS9ZrhsDm
KUJmr+AoJ0iljPsFHU72SX8SvI/iF4LCV+Z/56pmodc/98OTGHTaCYR0bIjgKjfXMtTtwyNbb4ec
yI1WJt5zOEzUWAHDcVkp4xSlabK4w1H0BmGRgb1HXIcEHfF6qLfIARIUN300KIfxXjlls5R3DXjJ
6yGKnUVZrgdWwG7q22mcoZB2KkgwzVGucUr+SmBryxTRK7B+8ai8QOB0pH7bkwo+ArGUxLaHvIzC
6/tV0K0476DnT5cNmYgPVq6YZKvDaMPyaTP/UeFa2hUDTRJYOj9pY70nYNtqpGfi3/HrPyQlFYgZ
93NqtnDxKHLVLGSk6xdXrQFgl5+f9jM/EMS0anwuAuPlkSgBpkNVIImWWM9cLIDBX8zixN5QUPH7
RsaJdr59irtGXsqQooi0fnqLaYwDMn/GlTrPIEMuRla2nBHt5QnH2yPkLF+QjHVn+9uEZiqP8ANd
vP/3WfmGNIXTBRwwT72D1oUysME+w0Dml9Ht55z6C/m2a/GcFi3H0tY5QMLVTXLlFGHBOR4A/O2R
txXva8BmuXObk8vf2ZIJLi8a05KH955tGM/1/39oh53dh2Sx5RCh57/Y5AXOe7QZXoxbWI1vjvKF
w7WM56A9Sd6Rk0Jvih4hUqhkGUy887c0IOwkiEWvu2C9YwcqF0BFqdAqxXf4CYxvLPNAtatQjeXr
5HO0v0Z7A/vMQEG321X2v44C57AjF0jmSlBc0yE6cah6m7e29HcPOXmblA/4YTTudB5yIIHauDjJ
zrIJ2A2pBr6YMWbBCahrg0wKicq/8cslRE/TN6gITsvCTO9vVUxfrLJJshjrjT0Zr020jl9Cu3Yd
yUZu5CVqpdWqZUeVyw6Gm3c1DofcpZuvAdw/CW6NXVq6JJs/w13eTww+CHagBEh6JibU5l33fVie
qIIOIxKHaEvbCNRp0SMoENdbeYqB1O57PMqusbX89Uz7lAXVpZWxVgbosvvT0IZCRHGBakhcVFbr
IQLzNnNZBgaXxF6Y9dUQA+Qe/bJ3IOE0UNpvLzqesbXOgNjKRfw9PpOXfy/AT7DPvlFYg8FnS36b
80p5c+53Z1VwmUlNazd/CUpOvwLmr7kVgvcH1G7Ccqr3SRoH1gEmhrT8M0PRsgAoEWBRo6dhzKo3
xcrSOn/A6rKOK7DYTbkzEuoYdyK1rASrk/ZMTODkP7QvGRkwsaeCsV0k1wNCWp9WMhntDP7pcH8h
o/9HEESsyaePOFc0an3lzqWnsdaVCxNz00ltElt184J7zAgG+sD/7+fYwb24Bes9H3YUenLsFJdu
f+11O+nXD7vxw/vgZjXRJaqJ3HQk1lgpd79xY27cV+26pZj6cpdWvpnKe600NZUVnBOo2ug3X5bA
Siom0fa2R/8mGZ1scf32BrmyRcK2fxswJIdJ02UHVjOqt9qhN9EUEzt3BaHQK7t3v57J+5m8j6BG
kWuzzBfPV5I09vWrfNl4biph20NP/7XR/87QcDtMspElX0Wv0HKdeIYGkaXdPOl/ICVuTPdm+PrA
1wobtx4MywNFVH7RLHSv0RAKrvOZ6KafLWHLACHhfwxOXe+TkoZQSb3bDIvMTE3QTvwShW66PEIr
Dd478M6/m5lHsb1h57lGcRXC2mCbWO6KEI0auE3grA1xZXaS6lDEfbWn5FiNbGNvn7nbQL0WfzIG
rNtJOYGogc6OxfHyIceZPUhlMwEkV8W8RX9l7naMWXdWQbQD3GC+TcoUhT+P3Mujk63nLlfKFlSZ
cW+3tELKXB8O/kLO4QcQYGolDEjkdTGak3k283NOcNCPu3XOLFaFP8xlkfwsaa1BLRPcpaMsKLyE
iIB8mJTcfluJKmDWHF52muvH4uLA1kJ7J4dhAbJ0NCUF5i+5Iog0cD3MT4Ne+Eo8kcZCFqDAJt1C
LLxVcr4v7gQ6lmYRmYhCRwoBdXOisUxvIfDWreTG70YIBb8ZjlMfbUAHsZFBfMBEKCqJdMWmLuIO
4fQu6+TQbv6qdEBYWOJZ4peRa7Wj9DqwD1LZQZdSITQhMqoPz2FUhFBvbPfmLBWdYwbhOR4AKajp
2Qbe7SgJjHH7BszTgYhQbLZJGU97aWMJ9e9wE2vyyR0XuJKkzevdGguuFqMSyh4G3F+tNRO3uPlW
98jZZl2tf8m+tDLghW5zuMHFVJ+ZH++5aqud+3hTT3c7Irq7uI7Yp2OFhGub5HIg/tlTtep9Lltx
SQ1H9WSFaiKA8GjA36j2nxgk/KLPEiokH1RlDOVi1MOvtt7aBP+ctaVnl0eAqtZsaOw3Fab/+plR
R1RZbI00511gqGVM7bbFvLoL0ezqWwfysRVJo/1SNW5NfrV8Rp7JA5BMvxTOsrRtV8lMCVKWNe3S
ZK3GqHybqM1OLvNeIeA80BK8pC6NgcXx3W0opHknNGtH7cqUmpQv67xQFpbKQyG0aizu3GF7BN3z
WOX0PCIbvuzw9BUx7/aeR8PACi0RCl30hw+CrCCX/SHXJNR8XLHtuaH5uUSD9d28eV5LbbuIYOPb
vAIIh8oDPkq2NvXY4M873YYzAL/lK8H8fNVxhOC7RvCxFBNgKlOMO/L0LXJbxF2IXjKHODa//Pa6
CeMhLEQaN2rRBzTpHzwVVXnUmtgcnlWF07Mp7Yb29M/5GtrDG/VwpRXiYcAKCDJxCYOc6bS39ypD
WfKhmK++eyFZiVxMoX1CaqpR0Y3XgDfaf3jAWZN48e++ykD0n4p6/WlZHQWXXg9+/HEjK3t236Ov
6MvrmxCWritGkyqpPN7UzocrOVo0uv2X7I24SUTMUyY5ENL1gtohD+1uqKTl77UE3L5wo+UtO+Tz
ii5CAoA7MrSE7h8hE+jEWjEVUdEEmsNwF2B1gfOkdBz/eZTE5LriSiRD/s+va15iem+Gml6UbA9Q
Uv8JsNFzN5i5IrkhuTkpsMTu1YkXTahnQgBXlgdKOR0PVHdZpph7mlZtG3rb0RJMMAqL+iZd3W0R
g/Ijq0T/Uv27OEfWRQ2ttWtIXjo9x7orIoglDZlprZd1tRFO75N1yE+USbIlD34xzPo2VcdNLs5M
LuTowNauAUHor/da/EI540IbfRH7vluEsNr6cddL6WXhQNmrVBQl+avvmbADiTGBaffQeJFWJq61
raGbOfdilLwPGJgo7KZMruBd26sAi4XyF4svXmh34ut2xBMfHpJqXkjRW72nNN2sEDFu8xFmRoBb
pR9BL3mhF1P2m/ND0Psr8U1NnMAtZuxIMcN5xM79dV4LBvM8atWVEclzlxJp0fUirfaakkfn5iVb
GtDv84tt/xYBUhbawPny6BT0FsKHBvIf+gsBH8B5k1Vur9XrO8CaaAWh3lh01uILvilpdgJZx9mC
cevv+xRuuBANPCa3uRdsC38kElmY0GIGDYvuGzKzgpMZffHpsTtlOLWW/r+/8AbhYBA708T4gl7+
wsRZO8LWWZwakfBr6zN4rRzt6U3Xa8dp8CK9lFv6y1QYRF7HSxcSqmyVkCAPDY9rm4n+2DwYeKJl
ix5inmSni10Yo4Fxe4Ku08rjT9kMxcGU/rBIsOc0xJPRXAqdBrc7RcoYcxcXWsEKB22T86LMqEyy
VbVbHToQSIBpMf01P6O030Iup2EJqdpj1j9I80ys7mGk5xURorFTyY2l1rX0DmMZbP4qWS73R2wP
CrT9R/cxdQE/8VgguCbr2NGXFPQA76JTbxAWOi3i6FXjUo5YbyEmpyp87LugBHvB5tSYeUpddIpx
SVzT4M8BZbqsw9a/FZ7vpngZjjeRFicW+Cy7ntGXM/Dai4bYdV6kMPycT1I3fCz1eQJbb3xIpkS6
ZFOgvkvysYa2bB5yc6P4gIt0r5OZa6QJzmKicvunhHdXwhk8lN87yuT0IhrGMkAb2+KAZuVd63sr
nizJZk4m0t718dszlro7FOXSGQHx8Nva6PxC3bOs5zn6LaTZOAo+P3aSuOtGezV/Xu9liIYPnvlr
C+ARnd8s/5fkE2+Ydp5Bk3CCVvYv9pk2dKYPROvyos/uYf0vS23yIB9ajehRPIXgVINqfiIuzKbL
jDKaEXLUiLZIeC/KmrUz890DU2pvB9Fu2N7sp395RwT+U0r7SoBGXuePU34e5hiZVXByF1ykgFt5
WgzYfbJvSz7e//Ytn73EzHmR84zrjbiOYlvyD4XWXhCqPvRHCV2jbSRLJknzfPFIZMcbnFf/VOfA
qBxvdGIGmKGSCXK4BXs6jKtWhZ2Zye4bwZImf2GYkD1qp/xH6IZGaNG8tPsM/mUAL1lztU9Qffe9
RJQ7zmhrkP0iewy4zAdoxkkN/dbn3JVa/eWl5Mn491SAf10hgIH5wHFpTJCYThcNl0pKM5fbm8qW
K7fkcFmdxF9gOrnnQviUKIE7+8XrE3gmCxJ11FjMmh0kH1/jLJrGQZzP/HV9VJvqe7iwO5Dax7qU
v7zJQ3KRw0uKn+2o54K6rIqahW9UWJY1b2l9kkvApFImFkT0a0+cuKXNK0x2PV8QbDxCoWCkWIMT
PyI/kOuu+ZPFtMgCy/byy52FEZndXITA4EatMd50GrggU1/9cQSSE+i7dlZOwGJDnvJfoYppe58q
iMbnmJH6iqIyLAistmJTVxGYT7BJRSQfcOslUCGbanUZEF1zWd3P7UsdRVNUQSi8ags6yJu4Wd+l
FXd52UW9XZvCWflJwv50oas6aQ4YN64D1oHp7ambTcx1fR1vJ4V4PpFQh4ZSNEGGZlxrxElGFN65
F8S/FW9L7oEpUFtPd8ZeKQeXxm/YBT1Wi9oKb0XILFPwjW7KXujEIlRj/hyyO41xYBo1Tsj7cnT8
lckIQm53M6Cwv+zxGzuZbg0a6QGm6lGBoEWSpfBv2A0OzVWAxtHrF04qJk6HCKPjjwFo9b7Ig61t
/AEXStJ0De3z4uB/Q+rhGKJkKba7nM0WuRXvmmhxAlZnDgHzTmZs0Y4fpq8QCBLIIVy35hhcZT4E
0fJcm6RLazOlNqXdopwwBnft3q9gJDDuwoI1sOC/6lniklXf26Mcy1nydN8m38Q76Om3M8egJjmz
Pfi9CaV3xTAm61AB1GLfaoEpmgP5KQ9amwbUme7EDgdADGJM336wdYrgB6Dn9deeA6XXF4c8syn+
jCLOXyy+1DJWQTMZzqNsD9t6KqPOE5QSnLAa2h9FbcKckD40/JbYsEjYaEQcFlB9ZIDcddFUCBsk
yJQlXVV+/hPZPb9QNo+xgi4FstwXWadpkcaHRd7DCElzZAjD3tO9naoouQC8V+y4ZFC1cSzwCjrU
y8CZNG4TWKhLt5YE9zPpn29bQeAK+s2CYJz1tusmDewobk/OtBcFVTf+Z58JHTPPgoY5ruJM1BcI
ojFsTga2Fga88SH/aIxMfRym0NTz75GuZIPbeOMDkIsMiJFOTOubGPQy5BYl9TjahIurAq2yCwz+
vzjwtxmNMvDmG0R2E2uqmqQd3HhaFRnnih89K2EPINkekpG9EP/qXe7JxVLc09zNvJBOAii3EByI
Lgx0I1sEQd8pr08p/ImeYW7eAoEC2yHfFBLaLVycoJSXsRBQe8eIxLvazkYmt8c5GZylk9caaM91
mg02jEs14fdj4mqv91TfuIMb4wBZDYK6Dl7IGUBpzPVwoK63jLY9NnNE3WjlNFMFLTZZB514s+m6
ws9ieLltC1UCWWaUislC2zgODx1bd7s4KVzFGrlvxfgLVV/BLyHeYBNa78ljc7Fp6TBpv3kKggRt
1Jiw1l8MY8+4F8OCiH9oGGY7wVs6Yy724zT89jKEGEaFGOWgFSif6uJSxKg273oNlYUKOdUCKayD
oAiu3D3lAGvxWvguEiJje2hipbrlcaCxCOEMV7CdhgMjR6ZBgOQl2SwHovWpkhAM+27h0L8rYU91
YZ2YUiigv2tXwS/iglCq4eMCVxjMcgWiMesSd7+NZab6UN6r6fTk5Gl5aqZdIvffxtWy8B92KF/h
NxHdhOa+rjqyb0NKhBGDqckUHjl+Z43yKxlY02kEDEC3aRBl8lcd49qxEA7mzJZVbIOMNDcXuGZh
6N0bffDWZGYSdSaV+OxJg0ut27B3Ykl2XFwZlHnoFxui+na7dLHmPZG9WvqAbVfgsu5IiwY/toaI
8wKxY0cqaAB3LgouhxzbFcFU6YoirZjqWB15xTpJaaGl/KzUMRa/XUeTueG61peUAPAHP7CN3MnY
9n5bjKCU4t9e5R5vNhaukdM9F/axhK2nMaYJQA+8ttgJ7lPG2OBidS5fua11yO+TzH0LFhDwZmei
3SQdqpK26ybd9RiXyGViNaJwX4vApheGHJ/Bz1vk6LnTVq4L7avLdThYa2wNc3DoRU1IM6dohB0v
h3EswztAftyXro4i1kId7lXWThoRoG6wntauJ15UC4jIQBnNLCi38gxFetXBzU2+cCUoEvCkMj6q
kUfXhQAyruRpr58DDXFFhukcrZRNa9oVi9Ua2IZOyt8ntfJ7MdbcdFIqLTj6YMmmGf20w3rlcaal
efidy9lB0ioZmoEQkQ5uqy0WTFY7HhuVogfsLR7gX1GiTfFmlXamxqiwfe08PmO92+r054qp4un2
opJuhb9w/zXiaTy7qaPZZYHK/aIi2/94c5nzv/yAE/M9JoCMXV6moUOB65ZCY7q7cTIV+5As0cDq
2GxSYXYiHemkIrlhh6cWzSFZ45O2Jdhzy0/hZjxB17uxVXXIPFPMDROjgF59429PO2YPv+XKD8Gw
O78hLd9vsfLDmdq/IOBCOPRab2U7MQuOucAlMMgGwS2STPQejWgYPrDw9kIZBnIaEiLedS8/XHbw
DdLb1y9pCltOC43psqpK3FBTnc1FCTtLY/Y8meOuLX5XsGDIXdKU6YyImv7HCuNIpYMYL/uGQ70u
GdbTZfGPV+hRGYWlnzTZ76S/lZzIpLWjSm691U+l11183nGui+ViWMXwDMtaW2nU681A/Fiu+rDN
hh5KBXWRHbbgGCwHIP8Vo8mSDJWZGedMJbZ4jy9wGzT1o/s+iUMUM1ZjPT263Kuu/E5AelDFwqxx
3hW9cVgzzpEz8wkqdKbQcmhqHVmljhyvDhLsItnqUlQkloLcvc3a3yxFVucJucRuKpggyMtERDtg
ABIaC+64mUhPbiZ4boCMn6AF3eBDNdX7TtW0i6ZQS7X5SqsxwGQpG0VhY3Bb+MFaPi3ASbipfKyh
KbjqLkuZ96LD+6EAK7eAIk4FEexpNqVhuyaSCgLVyHvwHWYohaF8pJaRpjsXelAARrrbcNp3EKl7
bHJyhsbhbjg7QY/3IsZbpC3NcesIJQrDZFt6h4lQopkXubAMMPLxbQ3SAZzVdQHjhRqRdN/tZUEc
JGVSqS7FcDKWLIOEXIaCFSRW80YawLg5lRqkN9mxKkF9spXOhncZiYOhMnyqIUzJaIkRIeALPNdC
L3vTNaZRlSpDlm3mk529lqPs/TMQtc5Sd6fO84/RO+ObCcBXVgTrClfoCX5gW7MBrdznIDesU2S4
TC4s0xhBvMv6GG8RCNf7e9tzjdDjL3YhGq51+lklQqUGrmT1792w3Y4YiG4Xj3BfBWgKxrlXIIaT
RurZHcWyUTei1eNHfkQYUlK9n6yaFnEqx4EiKPKRlswLpmYXC2QyKXQeqk7gdXPHtqerLIZfkf96
ysn8q6u+qUEShHaRR9NctOHlrtCW4J+EBPRpJFmSXFLISbbboC+xbRzgXvg3I2iYwJtwpW0Xjeow
PrdqMEktQW7+pfr2tVFottwbNJRFgbOPzh5bj7QSAqq6S4T302d/bpfHdFxHe+qTTzSIUqneUky7
NI7c+A9tNpXxk9qE+y0GUh9gAF0AyhNJBKO606Zbjn54WSNkMHlpvuvPZwk/qPaqDJtqfefPUv+Z
5aeOXDVzz0+YWJwLCdbAg6SfFZTeK0fM+scRRuZlJjHFAtB9mTyz1SQKPveaIe2f2uQqpGCaOeba
Q7FQObSNEu5igc/h6RC2TNcJ8nNkbONqjxHqSzrSzMIYMbUnKaFODFZn1aJjSgzEbSGDks+bDmqy
bTJqoh9taVYfGJCdA0Wg3s1mseo4uQAj2gFl2NAA0gkEuobZC5uixuo7+Qx7x+qsb4Sy+W0A6H5K
moT/twEONgDpRdUJ5RLAFg3QiPOQaDWywz3ELvyrxdJXh+WOOHMHl5OB1/pdHTqHbsIqOTWIzlTd
9xVfiVH0yR0x7KN/3oDsd15Cqh/cL9c3adv2q3tvLU8IwzyIU9aww5ksP65t6WWXkwkJHnM7BpEy
ZPOhsljU9hggpQP0uK8FsIJD2zWHCCYNle3XXIV5jyX808ChDXOs3l08Uz1eMX3XFFdrfr506s5c
MZ63w+m01+KZwQVWmpBx9VQ4IbMmLrt6Ynow2BIQuNiONuaV/KtZni8Mdq2yk9an10DO96WrudK4
zFMYB6DmnNSxLmE6/kXPtSvy8xNvXsGUlf4LBr0F+y9yKya6U0SOhc1b455wIEk39VcMT/brUqMD
EYZlT3UHdrWnAu99kRzRnG49NJ/fBddSNMPyTO+QzqkqPxan538zSJCv4Cq/9uCTdmmBmUy7PkJ4
FcBBb4AFio64NWdgMZuABOWD5KObl6Q9UaUDIRWqgmvOUSvsvWJP+kORjZMhrTFzzPUNEJBUoBQJ
ThIQWbPPJJ3tEOqTwPG+dqGqvbwOkX7EBo5i/vMlx06K1TC8CuNB2Dzr07VQzHxwTkFG+3/8noDj
rrBlw6wy4NoW2p7I8aV19uO/SRpd0KNfBIO16fWKIbPxC7Ttb9JHVMgpwqI+hEv74DZjdJ8av4u+
lFukXsV/GkmXYutyyeDQ+3qDbnizFBoISH9tt0zWjU5R+TkdRN3GjC7xUSah6g8zEbUn2Ew5olFR
nbdpDHAz/E99UqQJVXtlqCFYz3iwUcrsj/q+tykRNrbLGNdhHCJRKclItP3EJJY1OiNYZkDssxnZ
/3wwZAATtbi7iqBtgxTPNE1XYq7X76F5kZL8KDUNJLZIRoy6FzQ5koN37KYy8oQJ1aIcr19QI0GA
ZepZR3RVdX2YDvxWxec2jdkFFudWWJ15GqipFfG2irZQG4tAw8AQG7UqSIyBS96xGTIEJyaICKw4
nyG9cZCcpGd9G85W7PuIbjSiFy2UPS6f+vPt7eE++w9FL9eIqBByiNkewWbHy63z5GtIwxlpTADU
zPIY2MiKHWWO+tBsk/yFLuagBm3bHCyv3pFoHsm/2WsxGU5g0vJtS21U65EElBsIvE/78+dbX362
a1oGl2ypFpz+aFo2b7FFAZjThCJgh0Q0WdkyREa6GnLIYtAU51G8mrST+aWnLBYIhZj/f0K/TO1W
b0J/xoV4tv31OfT5EbVFekyaUUplF40qJGrrEcmR5aNwbG65HlH9Y/5b1nYsAgnJD9sEBlUnuqVL
S2t/EW9h97Oy0lG6O8KV8wol89Fs2u8J8aLl9EptOqC7AZo3vNkSmJ8xloG1aI5tlVQUOojfuew+
SRD7SlSRBjBA98K7ADncaecgr5y8jrvyuP0QRX6D0dRs/h75fJip4fLDkddREryw01U/Kv/VEnBM
G6r7EZCq83Kf+lhzD0mr5ARYocmT2WtrcToVOzYJ8uWAfaeVAGwYuz9h+MlQxHsqm3UmYregXC0N
BhG0oKwJICbL1kEXnLsS0CrT6Fd7nKK4DWTMG4oA5hEPRYvAZzOMcGWpJrM8Z9vF+kHGQi3CwwBf
oGWST0xJTRtCj89PJiUqDeVNg2paX2DwC3XGbbBAQrZ/32of8iEb0piS9mC4Os63KQi8nVrHj+Fz
eCRmQUjOyXq/WpB81UKYwymnpduYtlpsjylwMuBvzHHDp+6gQGLevGJcjVxZAze5F5jom3bb3D45
13IDm5gBRbYETWoN1QkPICSYCkMdaXOYF3/G6hCTzwsDt+7QgTCXr2uhM9O+WkbXGUvhwFOTQbsJ
GQtxxKKvOTdIKZmfGk8n6qMdYz9U1z6PPBgmCbKZ+lUv39w/OOptoS+iJq3KO43XEEhoOjalCrxy
kpvYhhGXUeL9Ks3BEhIu3nkCOlEEtggwkx1MAtprnAGbSm3HofhfxG6bqgPFh+Rwg+wF4qdootl4
/Z+HZZkZ8khQMr8y2OrcM2WPOuOFc0nV275yXLW95u3UyUaapB64mMx9BZqRk9FhmssjgwZmw7YW
v1vCTgpvZwkSO3f6BJpBgB58Y5NKbytL3aQ0AiNG56Zni+6jcXIJGo70G/v1X1nf/NFdw+4V6T7B
68g2V3HCI7K/EpCMhEZeA/q6231MDXzuufM2CNjFjvqsdH+F8FAL4rMLWLnk4XBPgTiGmidhdHvR
h1Qkz9I9sTNb8ReFJySehFTEQ3ijNXEOshWm8gEHqZSv3+EPUdA6W5tHAN4nAc+Y4mHFe9lB4odu
pUWsNfgQz6sMKiM+94hAlnWQXkxIt5fh6T/h2Xlqzs5TeETMthqV64heLk+HzOoR5k/tJBQP61uZ
14cUeRoDdtlx42nAWPX+RIt6ElABsZxBdGy28YjurBc27o/Xmdh1ZKNefxZuqgsnNhh0ztDBkWwx
vrP/TqcuGBadZR6xE4gmH6d6vA9MbxfkbbDv9YT+tzgGl2ymsE3iM9bqeiWyVZzblptRQVCw0yze
jyFySP0ukrd4W2PfF6VUkUaeP+ZPbRl7sje6N76E3olnXGtUx4eU0inGQRFEdXJvTAqJhdj3ZUlI
Xu5x1tQdd6Zlj/1osA87SEfOz3Ln8uhXROtnEcKuT6xhbS7qWy/WSZpMTpjaecLdbBGahVlSdGYP
KEJpy4+ZnHV76yK73cHBoLrDUCcRUf6m3r5BYvKENZPqzcsWcyzDWxUCySmWiNtUSI4G/3b9HVUi
CfD9DhRNTgG0icVyDSFUQ1e2l4Rg6FHgYRS0zqbejrnA9suV9KfPCCUXLUG0qN251VUfU0M1dA3o
q5CEzDDV5RZJnCMkCYFzRHMF+FDmzlPc9Y2sQ68bGAiyw5fowkHjKcindTHHkxPkJTsl2tzw3IjU
Mr3g6F73ZIEcCZtVs9Gkz8Viqzv7EbySyUNf46CjKGLzDNecARy//A9gAZzoIXU/uG16KcV9Vxf5
63c6TuWH0b+Dl3HwjEtD+xrQeWH6hXJColrGO3fsvsU/2BA6Nj3JcD7MYn7R0UVMllVrLh6D+EmX
obACGxp2vSDq5SwzCxOlT1lA7JhjyaQVDooDSXly7H6W58zc/ZsrgRrspyIaxZW5cbTH4btfpRjG
c+QptCOd3ydoKCFBhtqL1xbXm++bVHkAHUih4UBdneSw/NJ4WfzHw/gvtza4EJ5FbBEr8yI1dmIT
8I/UDZ1K90EXQbV8cItp1h3DMwnaD5iXYt6ng407qjmDa8Scd7VxG93VxDwCZxABfPj9SB+uASiy
TvTnsHfWnweWT74CExhOZeJ0bFeBP78wEOdXw7AyBdRnXCj3LbacJPFXL6ZhV2g9hvOtUtXa2pUI
uZnukhMevXuabp59PP9a3nj9R1dwzY5Lv6M5ScgM56TlCzKSXwFTrVFYhOv6MAZJEAIoJQZ5RKY9
lgrhu3xIKZ1U0YaiAgumQ+RyWyjpTFP18Yu6WZvbKA6ClqSgan4kauUR6BUmZPWr3it7r+5umrtg
7+HU8KFMkypRp/NiA18yXQt/3c8JysQyvkH5ekJH1ZuAJiqeddFqvZHaetd59eeEbcOBmDw7uLvx
Udfd8cg1iu8YGMt0tcEQJcRDnbnYOwxSJrqGObvk3spGooYSd6NiwJYYC+HhcYdJx4hIwzCVA2dI
+Qfqya99mhBjilJeLR7JlonvdzszRAdxF+WENagdJ/CFBu/Dg5fNDUy4+pQ4Ok/aj7fidhBunkOJ
Z0HM/jT/UJTYNiUis+T1WYqFoJeXGCzr8WJhPvZxPudVzNeBr6XkS2xhhVT4da7ofI2AtxRZ7dz1
mE10mdsfraWXOOCr8QH/fMMFdDpzNk/ErvLmQqFljlVF1mUncUYhsJfks55LxntfYQ0CCvQrl67n
EjapBqiCC6sZKQwQJwAWLRiqQl0sqd4uPGz1Wvb3P7QEUgoOyMtjMmGKNZ+FcNnlLsFjEC0QAzBp
4b+oU+A1hrvVRVXYEMuWHDI4DqVqLGD7mm2ktCNB9REuQQKKW6p2pUDeiathP/KX5EJEGlfWJoAb
V9UtnKCnc0+xcjbRXQxMWUd5YVjLOAntCB9mUb51BjL74Qik0Nc9AAZekP2WJMGTJb/zc7LbDBoU
mOrNarVLL1A8xFzfxwwUMnmyQY4LkF+BzUJAlel2kjWVdZczkST92QVr1F2E664UW/VGE/vTeXEa
7a6Npa3dMSXr8mUyKKKITjShKjiweaRc+pCxiAg5bLB+wFy4vEAxCURR2iD4t/EVb+fMtRRnxfjU
sDz7sdvCNovo6N2k3OHlT89cjGeKluAYI60Zx5fjtzenQTFHMQvfqNMOdvx5G4RYHLXtTwBn35If
Vy9r90KYFtSWT+AHCQBRaC9f9RranP/6SApiTl7ilO7egAELDFQCxGxAMEDkJiq+oAWvSrXFRQay
v5I2TIxhjjDQ2swxhovNL19gosZh3r+KNYZXlDMx6nVQhiZrEp3yko2lImlNt/jCDH4cG/Ba4iX2
BZCEmKNeB4bFVTb3v0lEnM9pC/oKIxPUQ5t3osCauvWDMAg5QQw+5pbwah49oB9tV63wdPz+/VFd
WItS61cDBq1RB6EwCRnnvPbbN/V7m+WcS1kC1TBSXQWKJ/h8wu+zB8DaS7EQp8Q86luEv5wqobll
wbTKrpBHWPxMfgQX+N6cNQB5eCV/6XQHNF8brSICZrlLxv4isFYUyZgEtbmRfPJtzVbyHH1z8svn
zar6uR5Sc5nNdwpTC0j/KV09YfNtmQ8M+XKVEGqU6G7GfEqWvf0HA/3pDCYMeBjehkKxA4EWQaZv
18aMzRKeFh9l3/rJF6GSKchdvz9Rjk0KC2bdlaDO+VbO9FoE9LzZA+uHJPzAapW3c7/7jbPSflgT
gKcQ1aI9NjKDoERosd4aUFXWENhJcG6rmuOeQxaz0L4mchQz3CC6GTq/NIHYvhiYYVIU3b3IpN0u
aKSXVdZZAHuLGtpqjI80Z3T2m+nE14vUQYqPgIJKdIyxoA2PodxHZ61ZnVkZIF7SYHNVeXTx4HpJ
AZJ75vdq6m73uPYtUjuHDj6blgHL3YDf1/jDZwi3G7Nh+098f7iT6gca6fXesKuQsi+reZYcv4PD
qF8uyZ0aOo3UQcinNKZccuRmRIw3SsCniCZSqxVeC9i1Auh7wqe5xWWyuVata/MhBamk0uBcDYaw
RL8vAR4JWgyEVJ94TDjpj/cXzt5qzG9YkV8pqlwGyZT5xJ1HeCvAgnSxHr3+edSaj5LlqTjn0Ch9
IeRqp2zeQHMvu8OO9pwkiR2tH1bV30Y6LqWH3x6hQ6Jz1gmK+RGhK3VdKKY1TYjtDV9sCFMNrh19
thsBAJcruT1ESiOY9HDBvMevY8+vzsH9VxnTioUhu/SoKAbJDPAFMaBOF7KffT9AtlOhNEPclXW0
l/C+AcZIj3POwBysGxTeTjo1sBMYUuQB8WzkRz9ZUTF6uN4y9ZAKIV7iZ2QObZEjuY5ryKdMyLCL
JVkgR2dCtNiJaCKmVN8M9tnwTwp2GFFy2peJ5q//nTuhZpkyifih6oQeSlO/j2E0sNv7m7k0KFO6
jH/MR8jyiXKcUnS1/Z7vI5Par3UU7/Mvo1JNCbV+9SSFK/V5IMnrzFYVwQDlyu9k3zS7dXLtvnqu
zdgeD3QYTUMROD1Jzq4TSzVJH07TqdeLLHRdLNMm9cGmxRuStYuH/oJCG3/LKUbIIWD7Krt6unSc
2tFyjoHJb0aZlA+7rXRac4199n1hbwtaK25WI681Sf5UVmCHSJKXdYYmo+CNABsYkUj04CIfMioP
bb50WrPKfriKIr5HicorH6ju98sw97AHr0Nh6bslE8JUhl4GsBcx+aUXaYvp8BJSFneQbP+WwMyu
doxb+Nj4OGTH3YEyizMJ54OL4A1SvKHRevft4gz7gW7EYMetENLo+FMRvNpFL3HCUlNbEQ4Naavm
xUScvRRnlhZ9PY1Cgv4eZJ6CeN7C4HUsynFTkGmDlpq99FTd9ZOoUWwDZWYgtR5/fA/i0DA8BElr
mgXqJ1PBQBfHz6iQ6XVtqwiosH8bA/+ScS1NUL1X7H0z5rC74qS0+LBxxos6wpoNiZbRuZFscxvT
yx3/L7EyDseSUTfrBacR1oxzZkWQBZpH1cGjsL89tNKI6y+nyfq+T1IfiEma7/oMlAWY590+UfnM
rNdKbGn2WWB/lXNtVtuOFaXoN9/C1L3eKwdo2plB97dmCFnz3GPgSxQP+zFMXmXpRl9m0/96JxTa
Va1XHk+mqncH+9O/s+xyv4gAJl50G+Y4Isx7cSg+tlNxNOfm0uNci5HqeMQOO5pSkhGTNi0EhWhW
iir2B/Iy1SXBFMWVGMBKvUV9pERMoh6cmo+CLSpuqoBNio55FHdYdKiPoGJPUuCxiRo3j77epjUv
cFD4Bmn+xdpeN5243bFhGCGdqvdiMQDnnA5ab7u7hzdjvCNpSChKpHNVSQX7SWMcuwVFNzaKmahA
iXqhEFX8NNS3D1AWGRykTcW/eOvp096Y/CePhgC+LysHolCbCO2Qs0DPP/dNX+RqYisZbhZMRpda
AVQf3wX4RGnWxu8WdEUmkEh9j1/ROQsoOtEHztIkN366edMeLy45WV0e9dgoAiQMLui6podJ3hQv
WmCVNt1vBfkZE/OWA1X89cbOzBNbjsm5BIe64mQJEPgbGdjH7imJiCG7XFGb1zITeUkZp5rsISpT
ZFfvb49yJPMc/AB2vDyPv0efak5FZKflLWokFSnJMAoFAV+X59sOc8sJdyz4ZiolEIRbGrMC3n4u
L/wITL8onqTky4udg+6PI8aSACwtSRgAFyrWwnI2hE2xkPXjgtdGkX6ZEr7c0S8IWc6qH0/oRGBH
GhfddsL3VE9MwKkhHqnk9K81/Al74Op7NTFwTOWhrkQOCQxBk/Gadt65d9GrKIRVaTvQChvUGV5m
5v5PYU99TlMIn35upfJ2PcBWH9Je1kO6Yzs5HgqpJCk75Eq+hO6WuISHa3fRW3nJkGEEIIVsdIOg
ztHmMBtppa3UIiZBO38e6iNAESKUg2I1iwRBh3DTP/Pr6UNPw6YFHP0qWYfYD9lrTaba/Q8zkEbD
HKuf52ie7BU+LUmjAMz1KgW5iSL/MvEkQmwiZyXAACiWWjJsp8COcOeGlii1lEj8pRPnEo6v1Ewo
SIr2/yEYdKoNIy8CybxESP6yf5Pish931t3T0xdblZclau7qgf3M+7FZcZnHyBvReisoC84NJ2qI
e7bUiHPa1R4YFfagS5Xh2BmCK77acHlCJxflWhqIn8nEs4evO0RCFuHhWQW5NI2FvvD0ZwuinvrV
LSgAnzFSwhAU3785JrQPkFOoCsu6JvwDGvnBQk9nXYI7uANZClEtrcWgXlet+0hFYV8Y1McTyQpp
KUtS6taqX7YIZ7PIga8RH94ybf+/m44J4B7V5ynfvzoqwPSGYiHpVRV99QY6somU8aA0JlCsSGbA
K2Nm2uVlkFi1l8uMDkUwi5w1cvHf/nMeIazYc5ctLBnvVcCMq45QGceJH+0Hprx9uNaXSN/rpEu2
3Z8OiFSNM7q+xFO9fsT/hk6NaEZR1RvqAkygl5jIoeOEMGZMyrdXhQe3Gpvb/bHSU8Qk1ICMqtI1
oCzRGM4v3Ngc9YZe8MwbbNAeWWmINJCLEs1wToM2hFlORi9aodvncByjSgys5IVfIASEc0fPafvv
r93ncQMz6rBlGRtVjTPn7Tn7zM3FVPbTS+/QzCfZV/heInm770bwiWEDSWVQRMN20+35fL9WL8+B
Lvi1MTpArOtg2IriFhlg+iIWAJnt/RzAjV504UAQqwYcAl9ofyQ0xTCJeRsz3l7ei8gGn8ZkLSsu
f8+mYA8aUJdOEO0zjFmOoBsw2ZzL0Mz27Hc0NHqdQi09bjM6ubn6yBB6/ESRC5G3zUAUndJKelv9
T7PGSiyoZWJZJ8dFs/XLSDbvQoZxJuG368sJ8v0p/Jqnhm1LHRtBgPscemEV8CdniZVN51ehVzEI
Elz1jn9e2p1/+me9IdLWtRSgZBRIWR4ZrtBrdVkfY+l7QG+udm1OL6nga6PwrZoF9jmAufvj1ZU0
5ZzOM7jV7WatdqEZSNOnnTsUn6C7i4+7tZ8xit2R2BxM4VdkWVYL8e+AzMtLTqLqbGTweUROABsw
IHZJo6YDExmCq7OrwuE8k8NzGOZlPtYWFIPO1TKE8fpf8/qMW6uMOITTPIQ3X34P8xzHEA6ZQHHq
2qwrPjNwnwfBmS4DZWQYiqoEgTgctFqZ6BzeI4awyslLqEx/8r8UhM8Li+7sqz7zc4mu6InYMZ9J
hxx/a4lwRorZzyxA8ds91Gp9rellB52U1IieDt84g8nKs93jXuqJKcpXQB7/JsksXAHJaxyh3VNp
Nmbm1p7SF/3zWaBFz3i2i2t92mWvJ0BOqdRv94syDptWq3HdONcfmbAliKDGlWyidOXutioQBD1P
mjOQLKH8tYYjC7ZeBwgCe09cr7IqfKodUl7eSHcV0+CbzqZJxcHOj9q+ylfD1vZ7LHVw0c9VcRpq
DxhZKIeY2yFyJ/tOl6w7swLap0xykqADI0x8cHQD9pQJ7QOS97LIr9j2Vfj9mkuqdZBCTnp/eKKW
gNOTh4pBMyxnDt6BLbIg0ICpLdyonsdmdu/s1mvXg2aXjfrlE84GEUDToAFh6PJV4asfl/R9sz7k
VfG2LzlvwIX5Hlzl9UQPoaomO6UMYTqEndI5SUA2Y5FXzPsCHxYwE5b+RVVPth6jA2bC1hw0C2UU
lUXoppLTZ3v8JNtTEod/J6wiiKmaF3tZWVvssKZ5dvNQeWzXxoBO4NU0i+xkC2CBPEvlbvtf4iLb
OGmXc0SUgZTLGkiywV2UktfW5Mc4Q3QpEffb2aRsyVl/DrYDovB83Am9wD+IJ/3evq4/Kht9XjYx
TNJiyKyMVvhYnTppA52RqUDMpqkVZwcJjWKaLHmTqjO8vV8kUhNSw65zZ2MrsfKJBIP/SNNLxz5C
Ogkgex9ELKWB88bzqI+snJueGI7AFLebxNt6B7lrEpRgEHo1k1Qp4ryDI+SzMtNor9gpTpI/XAP0
aCvUkoPrq594k4+q/DHwq3e/zgqibbYclVEJqk/QG0r2XQknITEz367lv2vYhf1dr0fXsi96Fr4d
j04kuvATU8TgoYCgr4jKV58iuaCiPAQsttPM/bwask5Ooniru3xSaN9v31bwL2Fh+yq8CCcvS+Oo
SU3n8VfUz5UKcC5ZZrTxIM8VSA280PcERLQ84m4SfnqyPAQQxzj8Xv/pVmjVNZr7e+7nvqf2cZ2b
vRSAytvhwXxrH9jipAgE1nqNy2ZcxRDEYjH3F9OySXrFT7P/1AhguJXyDqJyqoB8YfV5jKxKQDB0
BbS4EEKq/FC/2GgRdMERKdhcsJouzLLIbimWlYO5H1Og0e+qjg07n/XjL+5xexhqfotTjiHNq4ac
SVS0KBFWRqWo0LhuZQGknpSC8PhKKKjHruw0G+DXPyk151m5ljake0VMnWOAOusjKNEZUD356CUX
3Zd3Czd1uZLnLIzpPtZcs+Hqz7Z+FNo8Y3OBRcdvibMFvZY4iArCs8/lGzWQLW2zSsmreX/5trPY
B0P9P2ylEgRxDH1v7eKPYtfVOohujj9RxXiKmAozlDtjcHCPn7gBYSKxOvGF2raCF1chqJkzTJeM
icL0P14A4i/mCChyBV6InGZHF3gL+eavvndg/x4ydXCabhkta6qAcnRO/LrFwKfjCb9hol4jZyzy
sVY8/Lwz2HuMeZRgmjCboYT3rw9qGL2E+2qYbZFBCYIrj2HnyPZP6wIi0r4EWz/UpZTyxX401ujH
X+tffaZOaBcEsMh8tDGdarZX6Wq69brEeoS2xsBum7ulv1Wif091OYnwYYdvx7AwPmfeReI4Xl/4
zZCc/x3hQTn3qRVR2JA8RQFx40K2t0IG1WOO/uCIcEqATmw1sKIn+KUm/hnpn6vG4lIyLlGmEJDX
kwc9GwIg+O3voOVbBgIHI60oO+AW6eJTFTHqRMaOCNYY9wP0CVsF47Ei4Zk3QgLe/P1jIawQRbOO
1Y0P0OCbj+M5vVESOIRaSRV+GgcoxzOZckZIZ6UtcsZY8eUxedajihxNe6Z2GFg0HldKdcUIdbT0
4/+fn4ZFu0EcPg3wjDpcAptoUizP6TPYfSzeUaZ7QSyDpzhwSVg/DOhrl5onZ786c8w3k3WGthfO
k3GDYjNJO39mPbtyrJiD0I/7Gpw5JZbyJK10zLfKDPbDI/A8SSdqf2QQzBkdkjIBts6HcMxuKEkq
JrSV1zFh4uHOGU+AsBu4PvF4WcY4HhkvINsE59fwHG3FqXgGB9nkDDbbgbyrj7YMLtdJSfeQy+Aa
XvvyjBYk2in5nyfzIaJvIrdOhUbpiLsCATo9RV8YZpg1UP55N66dZnA9WM2e+TXBeMT1/MiPwGr8
tJzNiO1DxHxaxdpIoNQtxnCkUCYCjz/lqAFH4mD59iOB5ti0TEr2RxmTKLubhtmbIz/XPFiKxAh7
V8mu6ur+W0lVFcwohWdb7MpWy7Uj5z/nweF2MX1JXBBUxvb2E7EbRTxJdYwZ5QPwyUpeyIgO2muC
wk8cLbGiYFJ73F13jf0Du6Pm2iW3+x9DvHnhQGKG2pKNmaylD6NfHKTxts5vOllZ61qSJ7JpHTU0
8vt/MjQNJqAfHVY5ahlUgfPHnvvvJ1HRK6vOnBLYCc2uyZx1Vo2PKyBpB/peTHM5tmj2qNZxygh9
tiRNA6AQTtEjo4P3le7/i33N1mfdmh4c41266Rql3EenJf6iPUDGOQqLj8jxfcsazcjzn3o8JT/i
bdilTS0/OuwxWRqhyCQf3VT7m0AORkkTYjZyrxJuLArXaeNjw/7wKguO5z7mgzcMU4kveiPL9I4F
R76S8ltKBXosfGNd4piJ8E7CPSviEqRbv9F6B3c3zLgmVmOF4h3hattBrpHEFCNJRKadT94BV1Cg
0xxtZ9CtGVZAE/ttTLrmwzlNG97OJ9fYlAHfo2xth5Ye/HIDXK0GRwfdST2dK7EbRzGUB/YidYBM
hAECUWc/EJz9k0UnH1rmmnJM5lSu7pWyl1I9Z+wsWn1SRsqjhPeJCOU3a8kPcID9q1dLn53uRd3T
S2J40ZHhh3gChrnhnS8FLpCDxEjYgMYOzOROoRo44O1FOsWPGT+JCLJyxxSGGC/P5Q/uxfoGJtd3
/QlYgc7y2AP1NeQ4qzlmeEcQk8/Sk1VC+a7UYNqNiiOH4PxfzlV4M7ag2F3qHqwhCfr2xu4gvKwY
N4zxJkT9dUjneNQ46UKHX432ilIpfMw7+oqZWvlBqNYcIOCEEWJ4+5meW13oBQMmMwg03VL6Q/3f
PTllrl7oe73qzhGx5DuLnOCuMzUdkKVJ9MV+IGKOzddJIGOJy3ITtPzhTT0LcbWcnwZnApo7AO0J
z4DJxsD3dzkc1O8zxJm1vHCdJbqblSM2yWflP+YV5hKn/Tmv4Aoey0y2OxkRTFvboEEjg8d5h2lU
05HvUqRTdgU4quK84C8OGZdxtdtqPPuEXA4h0LwlVN0mkpPdMaDzzsuLnrJUN9XThPgCDFXeDm2E
Mr8pY44Y9cpyqggNwu83SsZAV2gRVNXiYGXhKoGAboWfYsDQgtKe/VdvR0hrJfjyvEK2mfTQi2Pw
Qzv2EVQaAKWt0ZUmCBQkUmMO7ntCzv/BgXMqjFjoJRYfab1MNO08/DVXGhw4S9IK2f/xQjoGnTlH
Kiyd9SkZELjbuprHq8cwmhdmRo08ROg5xOXOWdpIPOZeela05p168dVIFtjUJy+6OOjzjPVewmWd
55T2fV0WnQ6/PXIzWLmywk8OB7blApa9EOaKvudmUNd6mF1QMXToeJuFtE+9pZkkmQ8BNdP8qv6y
ASUvR3uRJW3AXuuZiLrmh/56ZDUYte4pH2DKyUWIES0r3asfNFh361BMMvPgaIWyJlPNZka6LQOO
ityK/nJVg3al0Agg0Tmw54nmRIuyNagzgqVYTAHs755AKlA2hICBmA5Dlgr0hbbY16mINec3T7RV
TqSpyHKraK0neDuWV/4nXskSqpGzHBvNwVRyOdfZe2w7cRDQdutj1vdiS3S0LDpw7mcPN63fDgAY
HlP8bq7JrD57bfbDKae/mJ4G38Srul3m6BgDJoAFLNhKq2pgwCDLGA8V8yWiRUbZzPGzgpl+uZSP
7kBJUgj6gjoNMlmtu2OlFpO0wxv3vEet3LMY1mWtQIL6uSIKAHw0wUvLdn7m3pIRu1dIFMNzmgm6
G2RsMBjNK0yKvarzbUqZNXwUtRhnLpxZLtOLSZGWVepPWy2gFM4d6h5B9Uh2Hsg38FQxwYvRg7fl
ykJDtFZBioFPm5RtcYOoxhJjzy3ugvtMFy1t5dvEoCSmPBzJxQEwEK0xL3qYJwhwid9IJA0Smjzq
Ew/TXfq9SUtWI8HjLaQY2qrztdughIJz6670j6Oh4dbt8e7LFHXEv/PJwEpGUd+aUo/efd3YCgC8
P2lE3T4j6oPOVgZgL5A0y8GM74ozcFm2gKvShpKacMOPRKicScWQRGQ8PCVtYL9Niqi7Hb3YoCQa
s8xeP+j8km3NgeYv1G5zZfgexWgfdifEeZxecnaSz8ULFR1QWRWxiSIA9lmLGzlpWHPkrwFkSV3T
8F0qn9rpe5ViL0TZUIblm/kZZfpaK/HS1ZbHJynckGYjUpc8OvDsn+bzTnn+S3WS6VaI6DhcVY9j
iIe2bwSHY+HZ8Cn/ft5oMPe7UQAykJnVlBClOdDAtH2zqT/uCfon9waDMoOmJ7654QFvWSLB1KoF
wjiSaaVE1lagnfATWPdz6G5Mia5veUMZcJuMEsSqGfda7Gk37vfZOA4YqoqJgdxY4bX4KHrB4kZx
yw6aua5LSEqZFk8JWbW432zI363gWD8TYQ09y1fsb1eDsrri80JTGlnIuHqOiGdDDzAB23N5DOl9
h4C/YofFrehdzUsZQVCRlIyRWopFw/WAVw0DTlOtkVixFCKY2W72bqXPot/BSvSKSoVti3I3pGiC
8PfTprd+DrIoOqxd9DtckVjMfYpFFN8z6FQmkA3CBD085H5Inv+tGlClWh/wnWb6pqnceKoWcySJ
YGqdbS9hvjDBEZsRE7LuoYTqcoEJgPLMyEs0UbJbwMX3NUTaDlT/2FKcskRfLvl2YaFI7e46tMPA
y+lz3uhwiWzg3lO34900UjHbmQtH9RbSWclU/YcqUmE/Ns387o8eLcdMaeab9FLhEXebtDFrXBHF
+xch9/exRVMRbOh4DGFBHJ5ey5jMOfcfvP2Qb3t3EZRUJq0jRzrr7uyQY93o7JY7DOjQZsDCJvQT
/5V0rVgQ51L9M6BRzbDR3snkQ3Iuzre2gz+hj4CVK0GS4C4zMF6g0JrKEqXX16OcZLz6aI5nPSfU
e3h97TgY+X3mJD86GxmFvru6p3cB6weX0qdvMoamfG/nDwpp/Gdg67ly2a2DWEwxgAFAzbDSqa/r
jJqY/PKqzScYL+/UctF/qbzNk9VnFHacBIkEUWtORFRrMljPOD6vrXqnGYXVE6j4CehXNfALHOHL
kYPL5zeNRR6KLmil666RJ/aergDFLFJMA9wVAgLlD8rocQkUN95h46DPEigA/V8523X7pP8lNITy
I8pJvDYdyHBZJJo7Lyiy0dY/vL4Vb6guG7hL6x/nIFdnTwcjQbrgBiEbJUeHwea17KbeERZsi9rZ
5nTiZ7BHk144VVxZLhg4T4hEVyP5s7MGTeC0UoIKXw69TpSGFwGRqEDcRsw+hcY/8Q4zBEK2lmfq
U+3CgO93G86ZVtMNGHcXXN64aNjI5HqSh3R0JfQNgNKWT2Q/T1L90ZOWBLztk5DkTlVQ35dShpb1
AeciAMMu20KqSiJJKS+g6Hmz+su37VKj5zezWIj3YLyLgltc3z+TueksPiG50tqzn93yDKcDZEpB
x0exAmn8IY6jEIxllINjaRY1k6pAe8xKhdIjjCehqjxbMS/Mw88OmvHr7Hvlz2dOt+wACxG27knc
XuueXQb3Y3yAWAvmDVNYy8NqDMRYj7YDv5+ujQyp3ClxgNGBp49jH7Jk7/adpT3IGmemFt1aovlm
e9ek+rB354FaeTSjC+aD0N9uP0ZtC4PAjshBAd8oTlfQrXvIbfIz2TtnpFZSZxpBMx6v27xE6lsI
bgMQLjx4Eq3NT3A0HiiQF6x+kUB6EwTvHcKUVHqerzBArlX0+h/SD2XQWs4oo1jYYhEoTrufMssw
aZhak6U2HDSDbuPoYnCbhIVWIVkzIseYJ3FY2mkx2jzLdZ/gfHwUqLGPhuIn0tu/8ZB7mcusotCg
rxnBTJaGfBH6/xfeRilSjVpIdFaBWgcUxNeP8ddL08NjyJ8EzUvCys68t49JZtz0skhu/IL7ZwuK
RsC4ZAtdd1Ppm9DWvPE8xDqdVRfQyDBVWsI1JC4SaHtJkRntBGdJSzYQbdm5U0J3Bv/yAd0xMkvk
M1fwJ9sNvZ9OtbaXsXQ3zKYShux/AJW7+inhRWTe9Fm/EmA7crbRElNftym0tZzImXKlgGT1Dsv3
TcyUENOIr3Ng/tQTIlJkDAymeFFl73ZxiIeC3fTPhxIQWrpHqn+K6BmOy63843wAayObe2NKrf1B
33RC1ogaayZiuYjcAh7aodIvins3gHJxg1CTZian5vRlWaOqG0vK6t8V6qnedLMQdQv738ksSlcE
iQh/wmqNWBU5GmeE77bCdQLODuN7OFh22QutY2/Id5jw84HpCh6IdSgTKc0j/6pr6frfFFmYuVC9
Z+IaigwdoeAA1/sfIkodiceHal3EDSKIc8C0pHrRJSDaix/PN61gBpGmf+f9UbCKUYRtea4vlfgo
TgXnTiTIKI+04XBB6TD1oplVLfJX23V6qSSUg9LqB03bbZwJoBS2Ahednhv2dHp4wx4pTAoO1w9C
4dSK2H1p2ywqr9FTInnKnJLNtO1Ysl4DOXKYm9GjFuzVsC9eH0Y7g5uMYiALsZGTD2miFt4GeUog
126ygwz5r96EmkNfanBcyQHsz03yvBdNLfzKKxjjx9qwZPaSK1lROUt5oYQF/H1pnCqTM+VJCPR/
8S0HVWATsSul03EB+1yZXXzBzKsQmosT8Zywu6kKtKVlD35bQtX5ITFh4lc4BUf4Gbc861iIogx2
fhZ+XdXx2Q3/57UK+vifoJtSft0bJGuT2VHdmjOm8GIYqSlm+z2OyGTCHEMfEThsMxBEO+IkbYTm
di2B0Zk+adPd+bx2nbkz04vgfly5kkfPNvGaCk4PIZmSAfCs5zM08bPMzPozLCOrHgKKzbcWbR9x
eXdfA6z9u32rp2F7RH2r5qhovM468spTQ0R13DYkt/yVYd5nOvtKx/ImvLDD1ZJTsORX/ibZ3iAj
ni8pIip5oiLuotoJjhcbzpqKVnX52/rDZI9O3yCY1yXjtCoL3Jjxm3gP7TgROK88gmfIOuPVuzNQ
ogAYpgpBzPmAcaI1ykXyGXx3IYRO5CIxWM6Q7xx2oZYrWjVVeynh+7iJ88WkxdTuxW/eRqgZhvbn
xwRI9lkqQniEmE1amiMDBnaZwxfoXD9+pdTfiT7HfyafKaPHk4U5uY+yt/nNmt/K1yFfnIT0Ff1E
DIx7IJboGrRK51143o+z6Pk8Ot0a8LIqYiOepP0Lsc8vmfHWUVt5/LC/307OQwUd8lIxNg8ivojV
DyHOFuHQkqLB2Pa0hT4daUzR2+oztPyWY9QeQVobBzPrDEUYp2zEyYhsN0fGUKMh6IOr3iXXnarF
jZIwpYdfSuk6i/SJRCpxQ0kC4oLb2mtTQwZlC9UZwKkjtYlplCsEj1lBEXMhHXiVsvFowiGpwPY2
jW9BziSfuj7mcKQtUZEfge/c7Aosn85gNLtCWHvxYIoYnx8cJU4AodDCeb38lAVDC4g9Tkjf9BGi
N0LHcF6ml9Q9q0xpQCM0wG0iIwk/5IrAIQpHdO9lPyn/6vIDDR7qaHV4Z4uNfNmBlvwbJqULxWG+
0uOUYZArt5c+SRn/V9MtahAUYo42q34mcr4jnTSz0Eno8VN8dZpy0ZBvUX6RlxVWJyhEIKDX2odZ
7jC/CNKQ1yeZsOLSI90zQHBQCHNfH5G7goibJ2wciHB1yOGp3yoPQmGHgQ8yJ+SbwmLBYO8+mtzz
Zj3XvhCO98Ug473CfM6w7v4xhrfE8jdVVJcb4GwiJ222iLwbVKyDIX4PbD6j15bndx+Q7tnys/45
B75hF1qiXirIMvqZZY+fMH/e7fLPAgCLebJVAj7dhBfd5Qfb2rFxjx1mCAfljh82l8gmm9E/ZqbJ
xlPHeeorhjjx9hmcWH980yR4zX1t1uh+zwV6F1IRwNxhH2437aBoalwN32uA0xCZ7nMwzvcK91MK
vznyKJ+ey/xbJoJ5tl98dsXhrWYjTscJcy6p3gLZH9D6yMXECgO1BQL5Oe5u0QIx2RnxCGtAzEVI
QmBYA/T3I58zJvvr/8R2lPzlZ79oQf0yR8M9P3JvU3tGlxAW5FTDMFnnt8vCcfSm6XY8SnUKVdGg
E+wrNHRtR5aiYsAixeEW+2FSPfsBQHd8BYfpy3KzkAcghk9UUpkE6j/QOv+RN/vBTEqDEQqQigDv
YdDepd0cE4BUmqkYzR9Ypu7l2I/7TiFcAXFadT3RxM89cCHN5EuZaXVLh79+OsCnrpyFBTbmXfl8
R+nuJle+vh/cLKDnlOIs+ucjmSuK1T8V+RlFVZn6kZO1QSYvfiwjtIzDpRagYEEekL36eiom1m5h
dB5jyWZO5A9odRFep7s3twtGWEv71rOfGXThtphslwWfNVx66fYN+OaH5bKlvpuZLBxKiYm4t9zR
N2J6R5hoFENClQstguxvrMiQrtwsLvIc0H0mtdlTqQoj57Bryv2PAEs6zSo8NQMXpbkGpt1k3C3m
ZOuWL8dFGs8WbpHWR3ohh3C7eEha+G4L7UzWcM2ZceANB/WpW3xtCAFAoJFWorRb3L5eUiceUt/a
4D2S1a8d8kUf1d/5cNUchE+7oHnX9a8jTVbRcuopyCCSa0r5GjKM8vNJ/SX5ib1WwVeg+ro87Mjn
KLPUBhdqtBgeBJaiW79m3APf//cjfbluImcKjD8s1HmENtMjnJfyBzPQowvlt5BwxjxtYc4pARpu
X2NSY/ofpPB6OTejc45qQM5e4vbvU32wzj6UF/43yWFL6SS45bRBoNA2kKiW06xlgaMN1kwOHnA7
7oBddRbCjiLkknOcv0P11zLQia7SlcZplA2QTX819zjtvh4frZlTvc/3+G48pMHuCTf/XzcUJxLr
fJ6wnHIZExjx5oZxUyH5aZ+MBE07rhw9wN5aaH6UeT7GOU5kumu+JwmMNDBAEx30b3StBkvhG4lZ
J0G4rnmuUl+kSRpRXGcPmmZ6zAyuOB5Os6pvK4zgydzsU4TH0lr1EyxxhETj1aMt41RyM4SG/b+C
pxquhCn1/Ha/OohZZL/FkUCWlwXG/ZFIADkONfHR3NSNkWRxKBvrLpWDbJPlrgBG2BPah5QeSQmD
y7nvb2oIS7lQWGZh0Z99/UrWnWeBZcCdSFB0bIjMQviek92mMYZGKbyn3WyJY8VaDZkk+QZJQZIl
PCn3mpPfXBYQdAQWqnUqz/KQXa6b6nXdF4OXZNuNwUwZz0i77ILYahwJzKQqlIfKgLrM0O1Adj/E
XsE4nItdCc96xbNlSczeeMWdjzQp+zsWjp+DbsuOegj4sRQzMb4+rh3RjRaKoCQIL8fDKRxO1fU+
HHv6jkrYQckiqDL0iUdqtjSvFJaUkkkFk8yIsLWqXiaQvxXzvTtYhnqpB/VrS8zmtTE1KT7qjC3b
66443TdccQJ9MtHZIQsbrS35eUnynlaKlTSvyx6TAPLp8peCxQr4DrEU9RrDEIQCEZPWlZWaUSYg
Uh5N8S42H6iI6bjgrqN8giLhEb7YsA609s2syJPx/XeOqQEBD5nymm13dvFCKSK9oHVn43bJA8wE
tgnUkyxvMNr74LzMVWAiqFZFspAxKZCxYuD4KIy8wUCJZcIdRD7C6PaNZtU2MO8pvC7nuxhA00qX
sFkMbXB5ptXVOQbrRubEHi4wZZhJ43hT9HQtGagm9N16r6evgSeQqPzTD4y3oxqqccQnelUgFJha
M4vPMi7aKdS3qsjgeDHAwqhG4wjeOK0O61oNUussJ8k2KlTWS7OdP2WLANkjKT9U+EoUqgDZZw4z
A4+W3rHG3liX52n26ckSsUhxLmmfG6GtQDC53E3LphGPRDjQE8SEElc2GuwoDaoYmDBstnOf2Riy
p8YiDu00Kch5yRrnyUmMlNX3ozRqGrHB50A6PkTdLt/dZKrZyQ+LoswCC1n9vbgKK9lVcmM7ASUo
1Qacsi1MIWp82K8AfhkWcPNL8SbvKA2VgVQw62FVon7HrMnlZ95pMcI3tQM+Gmju2FAUa318Ndvs
WAr8Q03pK0UwNKC6RNZsbhyaZo2WnrqW3hl4NPglmHNdHEAzvBLnr6gXIER+PHZJq5E7op4AFHji
QwPlNH/r6BxIDl6bhnJowKzxXQB8nCf2WEaVTbLPhXfv/KjMFrfftEaTytlkmUb7W+EEwryipqkB
+27RplzQ1Jj6Ud3kA/AU2/W+Jvtg5nRZVXZI2SZG5LWP7LujR8vyjAxnEn6c7JZTC7LxELh8lbkI
KFbVpiyiQ4BF9OQSRYDMIbsddErLwHMTzJvuirv7wh6pOUMfvALeogjwi6QXDmIYVKI1kMKydb6V
4BdbHxZ6gmNGM2wTfS+xKDzYwWS5uWpJ5jbSSON56I8to3UAY426h5pfEou5sf3hiqXxp0Bis1yl
o1xxoRr+/m5tJFDOlCCfZLK6BvluOhyA1SRjvDx648U9WdgemjDFAMVkhN5NwWdgekGAabECPBRz
wqqqAXvBVofmeegcXugBY118UiSkauuIbwSarhTDLAOIJWSQoMSB5QgVNSkRZiMo722UVIH3crHU
JduISN0SFxZ/Qac6EQatoeFq17SLFYwtgAY9GFmH4q/SEJSEanCnLkZWecBO0/z5EOB7940ba31d
OOL5Xl168ziD/TuPUTTanfKVUVP84RMEXZblywdstHbUHkCH9sxdUAwly0BMkL2imVvah2B3A4mW
Cw3BgoFpyMuLSurJT4SZd/FmRlWjUV8Npz2kD5+sTScbFoC8ZqncSPexiruEJCLYIqLTDBYcW1JG
hwKbp7mnQPnq8tTobh9DTdxtc2i8o9j4ay07sd0t6X3hQv2ymI0h5GDYhITb3KIZ2n+YkNB/DDM2
feRhs+RYU/AM4S4CvQPNgOMGOdf3rfLa4GAd3BNSRN+ouokMCxVV2JK2V5vnKWjwO/VkdJ0JyRw+
cAoGwmHBoFAx6r3qkSMJR8W/BM+d0aWHbmkUMfQauMUkkKHyVWBVoF61+KjOHtC73P5gEGKDyVK+
VzsAD4BUqGLV1jRYUaVhNhQJq6Rgax1mGSd8cz2OnW+l3Oc4z6Wmz6L7FEp1Ycp+yhxBA51ffmVV
T4k40XBIFgt0cUK/8UIjbB6pXTXEuk19TUX2KZfGIEJa48v1LbMjV+akbr0onMUAK18nt7q+X3Tk
tbUgUHkRf6ZHVNKZKLWHFV9L8tRl/CRSNPqE5c0yn8btN5HV+xmaqo7vFof1OpuymvNBsRiJy1rW
vN2P11y8Y0L0PSF3AXlBvPKIZxkj6p4EblamjnilvlaQZZrYI/kU9/MQ1apOLg4L3fHVfNgGwI91
2Uzd7ry8hYlJBreShYxSbNGYIsyN2/88K4gs4bRRITNxmLubxzovVikbWLYqqh6xxAYZehy9klKO
Qj8tjlJlJANS8PHBEy/L0krfNVmXzPF/sZb2C9wyBr5kB1Ry24u+HBE22UHwjV/Zwn7pmas6Y1zH
wVZJVGzjlSP0Pq2Hq+JJ7FDN5GDErEsu0kdh9UUuYZp8pqwi1wnKBFbPok03Z1mZTcAz6stBqort
TAydmyq8DHLpEIdpy7OHqGJet7VQmux29FGWIDMT/m0oboSN/u3vs0VCLzv06MVbQPhxfH3rkFVP
0xxRy/lpTbW57Yxr9RrNTvrlqf+R8Wy3yACQQr4Jgn/VS50CEvNmv4rRb/PUxYHkwzMn+l6cIYNt
EkG8vG6FP+ZEkRYQAMnUWttK16Xf7Ayat58bXUxaVQcW4v3UGC9dXeqOPD5Nhj1/4gJPZ80he+k5
iAmlUuIfpdETGPN8xzuibb5NTk1s+XTdePRpP5calP69vOf21GP2LVNBYQ+oZ8AYURq3ssePPV4n
CXSieFanAhnFepS/qerrOlxlxynmEuwUpTKjPpU24PgM45iYauB8z/Q27aTfkgvLx+vyaqJwsoGN
fXBQvSumaAuAy7xc1KJDrWi76XNFavuphlb7ZUcs9yj6WS1iJ3duNh8bpV7Oj5VHXjrgQ1Bf61eE
j4B00P2QriQX0dEp7Qqmfq10z94Wxep+GESZpcWZoPIJMcM62EepPyocRYx2Thm8gtLCMEkg4u+k
uAjf8qi0GobaQqSWQg1solvcYLznoQejyqtEXdxuwPuGoad4zv6fdtq7Nk36SBXH+5pZllh0bgQz
rqAQqK+cklwVfl9pmrr3aCZV7N7vUCyK26j4GOd4nV4CheBmMuiZCwpVoJ5eQzc+8oQWtkRKe8D/
kOsn4KBMIMxB9OS9pqIp+dBrVJcWIY5M2NwnXby3KXl9ycSD23V6p4+Lc5sirSMDJ57uRMIJeDEg
XJHxli4+Jw0c6N/Pftp4Ekk8RPJbG1jTqGO3jm2dUHYW1uHLTp6HOykdHEVuZVbBLy8LaeLY8K8O
vw6QJJOAt1TFPEm3xIwu67rKZE86rAXrZWF1XWEwgtGoCAdBKOdYgB1yguiHlme0wTzblghnIZ8s
krWBfgeo4SqpChWExDdcOUdD1aO2ek+dmYci3Kw3CgoqgJt5vKMxOJMs6mZQictmoEsUtUaSbk66
Mq5xpoBW1R/CYv4bKTjsOL9OlN052r9iXOldmJlErnaITv/3fLbWuiGPeUwkky1SHeNNEKFUqutq
2CwuSMJVRoQKZoRFP30cIuOc3twC3wEOX2pLp3Gl5mVAChempRapT92f/pJE76ElCEf0SKnZJOi0
VCXgKicp4g37HdJMbxsv7hXfUqIoCa7av93/WshkFMtWEmpvYDDBOAVyKP7rvrZoNEtwZi+r5SpH
6jvn9G9W8ggcWykpiJIQoHFy0WFGEG+BAk/9LyiOjqL3PXxsGuFyEbXvIABvctlx+eJ1zgy6c/eR
bYIAigJX4uZ5VmshcZvNE9rtt2ZH7YvZiHsYYlFsVU4wpG9n+koZE3GzWmrwWPkAlFNatH9Al2uJ
AVWWze7idLKO0/oLqLafdvJ/3Q1f2aQKB5Yls2b5xLw90BxxZR5RKqNfOd8ZwnZmx114zErgQCCh
rhJXDjp35t1VwIJmbtuh3Sq9V3n7SPigf2J2T+zZPfszNARuBWBPj1Z84TAnt4oio+CZQC9t7UWO
RAYG1k+h3+F/sguPzg4nm6+4y1FfQkDcxNn3jS/DMR5+F297eN9bM0rc7OvqWQjNAO8J+e20cpjD
2/WScUzFQ0imsmw2TsWAlpx4+s0L/yDhAsG1bDDqkgo8tgqZy4D7p4vXCWu9ig6kNKGLB+7OrpEk
dG9J8AmiANW6AgXb92koy0A/2G5mQQbBK8+LOSwRkh9RwPhmNW7tBIKdHBPAVoSLYCaMH/73cLZa
SDrWtcUVhrhNFAnfwg9/BkuoYprpqAJvIc3xZt4qhJuyFWD+K4sb+O/VQJQwd16FCKlhZl8nnjEK
zsTrPfg3Nw8e9OOZbHjnj+43H4ejHasz9a5BcQeqM/dvkl0cTbFFQWEjSaLSH8Oe3ezvJQbdJd2P
qEvNwXj8IEgARZHP4MptFSmuRNr4WJ+imNIXMvS3k0WgNWGa8/Qlzvuv3ZqGf/F9nOHACkhXyCIP
hi278scwADM5gaIMDRjY6HTOv38AY0p/u8Vls/lJj+LfUGgHmLPB6vHNQJ23ij9VSXcuuLMS9+mo
6vZZa3WUxsdcHU3e4IdcdkaUc5jrwADKXTVS7Z1YIVtmH5c+xUFFyF3gyRSSc1BwDOR21ITht5lB
dYkFl0nGVtOHBm/2wEdwf27s5c7mHmjpnOQY77mqG7ra+Zy3gcNxqs/IPH1CZuU+VM4Jeq//QoMi
QawWBcv8e8f0fnOZWB0KWo8d8Ln2rift+yP6ccDy9Ho2+fIedLTJVi8G4uRbi6ZltSSTeNljeYtK
uhCpcI4Tg9ccAOc6W4gCPKxVhPn6g0N/oP6eGgLNHoyAoPIT13HLT4ra5ZQpmPQuFRy8JBnrLrvT
BT4s8GBvdhrI0j1ZofXz12tSiHcRA39Qs3u5z7v44Fn8c4CiBfbtdM6DcRnfn20dMXadmURzjgPi
UENLS5GMwvXue6sYfP4M7VWPlE52G6c386iub2YB7INOT8RFlBLnE+0UnvhaXIVPhu0x9dHjVrv4
t5RJMN62hXPWZEh4JLEp4o2T23tVE/oAdyiBsKLyJ6kycwWp8B+tIdSisZ1tuCtwhdpTnxsmzKBL
nH0BjidkPHbBVv7DH4aa7vyFrMjfqngY6zHgoZACqDyq1z9uVIgbg0fFLPtRsBzPOGj4/A4sHakP
dXfUIXueLsXVMkHTPLjzKdBr9YvPwm3DzGVKFE9cLIw0CFo0tKe0ylUKLtdHhW2hhmmhqL63sFyM
AXsRv3e2tgqxOjW0JBVDhn0eWa1z0OwOTZBeRXkXaewyLgWZZt/CkOOUEc6Cp78XvPlQeaAa+LJF
/sXCXOd04mMe5N6D85KS1M1FIe1QwPvafI401+68yhGwr3c4rkZKC+dFdk+dJg/h/zyENx/h3ly4
N5EicRQ2sDEG3IfJ1iZfEw5QbwGNtFOGU/EKdPKst8e0N09NN02NyVMnJX9Ebp+brcLy27lwmUz9
cEosvydL+an/zAhHAd4O+B/a1o1kAN5oUB6w27XO/2Bz6T9SANSzDFeIYxB4H7Eww81RSFbF7SXZ
z8Mj0dmEKXjqpYp1bkeSVhkNcB5csN72lKckUfQnfNRcCgJuiZQl1ahzMVouJaBwF8VuU5HsaVTS
4ImqKqjav39zV0QswRWgNREfrk7VegQ3brgCZhz5SchDjHS7Cv1d6XI4f9eokWseRLEgWVfkYNax
U7oqJhEwFmDRKZPkp1udZq5aSii1WIUzz5u8USwpAWXb0tR0ITZtvzZnIkDEdzaBi1m7CjoDgocQ
XwFAeMRSbaHUXLANegNVwCs62KScz5li6Eg9jbEXxDG1qVrpdIeAuOuOj3zS7QBOb6gVQavKdnpt
d25JMGm0OsxlWrht9VzsUy/YAFrl7cJOxGUpZ01F5PPNiwSECYS7uuTxecwfvX6e17+Crtn5EFVY
BTO9I+mfJEq6FflN9tFa7sLdv5IqGhYCuy5TAchWZQeh3qdYXXnisg6wgaAnqPfALcETNAeVat8x
cy/jDdKWOI3lu4f4W+dazwAoWRA9FmbdXpdYho++h7nLe9qMbie1yp9wR4ex6INb1sYJeidGcX0h
I+y0IkKnb4jcbS/0moVXJamDbMyWv5uDEd6LI+XhONF+MbaICuIzWg0lRkBgRErBCOgjAnnpjtCo
FyAy+Jc+rkZoiHHVysemlizFjyFi6GAjG2j1UmKe6VPhWA22AJE5eNio2f2+ZmDbbV14wlJrDolB
BgrdLeH7vsLI36P4h5TngyZyppb1KEHdrrowQFhyZ3lCYDowX+ogBom81ILGAAJB6k2x1CyHZQ9C
XfvLqEgQ35I7xlsTIfpcJxd9bgZGU1GytdcDaJWPD9gFrOEcLwFy/WVDD1Jz+pZwsCpSTjrBqSuD
CpVqczTP1j2615jyRnoDbgJrCZ6cmKJ/bEFE3pXHOWtqfGPewBW6RfK6dwKI6f6/OCm/O5xXDxCW
+Y6pDgHe4SPH7EL+rJJyAu4GQ6KyiHycOLd+RWxtFUjmqhfdocSONbTQ9Fjlqe+pIld6NjMDQzcf
xvRh8fhZV7KpYw0j+LXMoHXdlKTdw/+VPO1eR7tLj9SrrCxZ11foVEE/sOrXNdsklTokrycQTV0b
0pBodJHMU1ooQ+NPb3JHagdBhU6M+naClkNHbziKaMf9sL8A84T42pneLomGY1og58Jj47wASqPv
Zx5kgiz5qPWIFg4WHozfZdVZFFn8/O/G5zB4JD5S1Y6ADU0v4JAcfjj1hLfDzmPCy5Tz0SL0D4Zx
fZbftDqo+ogm5vdo6GVD2eXXeUtssTB+AXZJhKWsT4fyB/+smpXixLZmoBkExPgcJ9PRetveXo0h
bZLzLbYaQ/KR8Ml4VOAiwYzpsQCTM+dsWYFDumWhxql5AjO4/cMGyBoVnRP2GVmetuaTeuw2KkYz
kwwgJtLnXmbFCB9/ek9ubgLgivcXhZeIQEdUcbvUWYK02fCf1bSRvYE+ysjtItEXO6Zz98IFUstN
qnJhwcwXoVN8oIU74a5lxMJTnSmnqibN9NskUKyVvxO0DAZRVi0Jr4x8F/o//BdKXcY+fTfJmzYz
FnCvK07FfoNOvfUu0adXmv/FNCw6AOIkKQc+PZanpNFs4mF5ETA/Lv3Xf/Amm97P2WbtVPeeuQwE
Cb/D/P91mNE3KOA0H719GMkQ6VzUV2+tlcDnEUybrNTpSEwP9gBiqZF+6ZN6k6vHDc2A3JlP1nAA
ip6H0+41AtAt2H1ioEVDgFoDAgGaoPkjmkUCNJZvthK4eq2qr4o74ffH9Uj1nHufBpOlqAtkhEW8
5uQt2SCwMSd0kV2D7t/oJ1f7AU/7e1Uz1plRvmzChKCT1wNPYDVnnNCiA4NWJuyDxL2igSNGjkAX
d77USQGccTutdBfNrUE4fNumuYIGoGHU15VqBx+FosOt7oTSkm83ITlXuJwpINo52Eiygsz1fOao
k8nDc1Ts5jwFUBufWEqxIdAep23ZCd95GOU0nDi+QvPQThxnHn+4Kj6NQ/kIrmcYUPvVB22GMQg7
N2aet1MFsHx4sHpQ4qIIWYn+uO8HU+h8Hln/j7Ce0cz43N+qw7e7Gm2ss7WyvNUcvfZoLRMCVkO2
1cv+YnlgtDZOY6w6VYtSzXhvmGJKHMmFiBLOc8OkaEjQs3VkvJ+ipIqRbo0PH1silVhpb8+xH9A7
pFW4PSphCJEJBn7++duQRULJnBSHIfNrdD33AsvpgpFjnphSNaxUSC23knKW5wwZDuC6TaDye0GN
ESLoW/KEFFqFnsIEJg/e/2wVs6EeL5K1hKtRT4fIEDEPYXjw+0KY/a9Del2GgMskfLNtYSLEojUj
J1RSbDaH73xw73uycZE/8Mp7rG8reUPBCSmf5QDvcRhEx2CUcYqcbdfDUhfBJDk1HHWuKaOWc3TG
wkqTlkj0qTK42Qb/F9addYCvXFQTJcuqyHiOQNbAnOMS+0zXll9ROYSUaNGN9POtDVlflPE9tcZp
YVtZZXifBz30vSNIihU4wZ9Jpo1CLJZvudyWLCGp9ELzH8uSi7VZyXl3u+YNaYyUmojBqqebb8Pw
ZYwHmwnN6VuC22AxocBHG0AicsawZlzRvsPZ2/UixXwHqTm+QBFNofFlOKVxxR7HIob28EOfaFFt
hGR6ElpI5iq7W8Qz6YyY7VX0J+E0XSlEmMgtjozUaHok1AZY65xRcoefqVNWo7CVZzQMjI5NY7Q+
GMEwoQALXHy3PUSD3jTl3R+x9UkYdFPqsKK0vE00dkw9MCjTlg56oYo3CBe3uNLnclpF+IrtAcvX
0l3sr8lyWVIl4lwQMAHa+vmPCBrNF48p/lAztCzxgjQ0REeitNp8zEh7rnnoKwL0SjxBDJyC+/5Y
bA1IOZhJSpvQnJw8zmpTMdtzXNlzuznXTICMBE3io46jb+KMduJu3f/1IN8iRczQHE5Z9RLILjh0
P0dB8gXWD9MPAQLokqeMXwWQeeg78H9nXOwdIhv4sw3QsvfDtQTJw0G+MkRMyjLBnX9PBmANL2rM
A5J2TL/RT63dvcljL/zKGtBzBYiC8BHhkIKhSJuPclgnO6cZp6zCkCwMonzuh8qyOoZs7PiYusiu
a5i+dg/6ThiIOkWWnpgcTwXluQkuEbHzGODcpkrKRP9i6A9hid2gFP6hk/RUXo1OCZkP5yVSFWn6
uzqxMEzZkckQKs4+Dy5XymVPjZ+jpBe7QBsrPw8wRVGV1uc9koFMOB+T+jfFEzTvq84J1hdY0KzS
qpZZ8PtKVoDdKEtuMj1+vqap9fXjzry7sxNGufDn35ZWP7wcGly8pv2ArMwNZzwxAaWLY952MALo
Lgh645g/uJrUGoXjfZFLjLDGg5j0vl8EpA4AjrC6wIkNMx4Rp7QZ+4S+po6GEiZ0C8QH/D9pYngS
H/RTEfLDbAT9vN36SDdZ01xLkmkY8nJzxwl0DlnsVhzRpdpMn09pxDh9tb6wNaYVoNBVLTukkBlN
7rV6b+KNUuvP2uEEX/KploxL4X5uK5qN/LItJ+Ny9sy9RfIYFaGwUE2AFRtKRIEGvy5FAUXafDCu
SV8CH9LJljuzInhrNLCyjfs+Zv0sw7pQhiQZp9n+GCmsKY7BGODUvH66bGn9nEbUNeubBBy0uodJ
32iSbgees1+XeJuQTglZ7+1n6Cxf4jPmHPw0FjrPXD/G3BrRalr/96oxMC+0Z6B+VK4HM4JLmikb
AHKoY5DqbG4+FJnp3tWeinsZfruoasdlgXtGgmIn3ErNgSSf0xyKcjFLAhzI1cJ/8ctTNRMYP3kR
VKmOzQilxUUUf3335Z4eukQDlSYsZNntbimiyZkP2CFVf9RYzfdpIXCteFhs1r7UI3UDW3cz64jp
VIfvT+FJPg4vZ3hs1Dva/Jq7N5ptsaQUbRcG/YxutJ03/toSKdMU2TYlsvrsOapbuIV18hcici2K
g5DL6mDI38T7ko82Wd+UK8rBRstVrlKt51LReQenh3p/QDW/ibPebNFXgZvKL+Y0jXN4bkMfytqQ
rANV2VIVDRajkpmHIqwpDzB3mPQtHSmtOJLxQzOswjjPGJdagOEgWsEDSl/S/lNXswUlWqPj9OIe
XUvhp+36eZGFJgpFslGbmjJ0LsOvbmac1rb3aZRrFZo1TAm3zrVE3goYuBODGtzqhKQwZIqW42dt
JM96oViK6vi8BrMs8rNY3VIL3rob3ye7hszGJB8UD3NkKpS8sFaptZVV9nNfNYSr9ial/6MWh2PB
WB36vMUsfDJgp7Hmjs3Fiqwda9EIMb9cKqF1HkKaKzVaiJFAd5nxgNtwDCpes39jDZHusLZQ1+A1
z5/nsUwo4jmP0kPOED4GLJgN7iqllafPUgK/mAolqp4Pufz7YijG3odWaZC6PcDCC3rgkQxAs9D3
eVLM69e7g1zoSWGjzk8BMnkudynnlIiIQD2O/LuV/UlUs9q9t8Ho6lEONfM4QgVi2Ozv8zT4M7jx
uH37rQ03WRo/2iU0mQeHiVQX7MZvu4373PgJ9uL/DTIg+w4qZ9LpkxoHmKwrrr3oG8dRpmoXmccF
EcXs+piqB7/lW1Lej4OvftGrIuVBkNqLvbfRnvZ3njl4/eaOxrjNnbZ4adUh8oBPdS/+T2COcqeI
eE4zB5AwNgftW5DHvUIek1w6GKHgAiPjI+B0QWmE2VZAUYYHBT6RI67jg2wIvEfA0t+2V7MeP6UZ
wNW+sgrTRsrPHWvvkB2ZUIskcxqDFA6XoKWqBx22eahfCXcwSceoFPToTUtap8oe16pgJyPExwHD
s7rlLjc8DEg8hDuQVfji9Z9eUVJoBSb1UDT2rz33nD0kno+Oz6YyrVONYi4NGCYfZH1JweHNhuRA
JP4bOysQ6mcsEP/s03TI4KlSPb4Mpgae0lRukV5tdKMCC6PGW+HMZQ8ebfquo7AYE4avM3/kGoTe
3Ku01JoH55Jhkg4777W9Bz1LPW+4wpOYCK1ksKyiQ1cUsUa0oZXJPNdwIJZopapDx4fgez/bq5Bh
1El3CyofRt3f3UdTuURR2H4TRrRiwxmyJ0dZV0FPispFgm/Qqf5ymTuszj1fzhNhd0jEbazIr+HD
p0Va5V2/dG1VtRXXXeDAc39eag9YGq8IJZUAxIF+pDjASHFOImd20ByetvT51CFfCMqGuEBb4ynw
OO8l2zlbvzRi2EhgXuuzfo6xyBEj2Jdv1hQUHGW54evDCfO1Jzceeg9mZWT/481J7jUAux2o1Gqd
wyrrV86eAtnyGH39xBNGZpNPuSf22EYDqGeAZ/e8LBw4sx2OxfN5TM5DBhT7bwg7QMCd4CohCyDU
MCpfHknSdR1A7drx9JHVZPNoIHkHGI1iXw7FvoUYmWW/Kl70kdx3qokKUeSaBa43m4LlDFXtDZll
9p4PrCbmR3vKZ51814DscxiOTk9BTtUgEhsdlyNvMzfke0xnwBmNQPOivxAe3vW0iopSk4Z4TZDF
/B25ejH8rYbQKEN5XmtNXqprPHa3SH4U2p3IPVeX92mLkBFn/4GjfLggUvkfDKWkmZ5E9iMHAkOc
1JNtXUAMlpltoC+I6AVPFsn4TrR0xBq08WzwbEO6XSIAqEnsoGOxOgp+zuqFxtnhaHNgo+LTGnBL
XoMqU8saGcggdeoYpYhgVBlEBkXjEKOAChFhxlhDrERbpBv5LJNaA8VmZsq9ySZsE9L6P0nPgUFz
MTNcy6apmlCICo1BwpbWhHqTqOuEBT2KjUdc07dfqCMggfwwbusSR0c7WQ8Ue07AUJ9rLmIxeCgR
4IYWDZRR0DBpOpmFQTlES6z2wrcCvppTP9/d3TQeTsZC9FVF02hbAM94ZbnM5DYSt6XjsasRYZei
85nchy//lGOlSAN4/7Huu1gK9J2ojkvTAsK3y0we+wjsZH9B2XMKhzGj+GIafA4D39OFMQKg8LOL
h4rqlF5JzVC63bazfDLfUD0kjupXa4qi0GFEaaBtPWuX91B2aemm/F7sZ/3nSn6UN+onc1aY93CG
INXQhj3dytBRYkBj4y/xMzKZeKom1BKKQTkkkbaFmNwS1GptKKjjZZoTj0COokUvJT6RQJmgqPTr
1r+3wXfJjwTwVVqn0jN6pZc7hZq1yLrw/9+6QQw/yfE7h+M0PYdOo/mi81wD4uewEkvCD1ySSbPt
DeH6CEPHJHi2yV46QFcK4N622MugonR0JXnCt+DetQqmUq987Yy2V75yWrtVyiOvQYUCeJ6aFWX0
f+nOc08xM8ISmrVSGzoip3c1BI8qmpqHa/I1XAxrRgN+dsdp984/KoY2qRwmFyCA04xm+4BM2kj5
FqnjgxRTnJRd1PBhzZb66J1gqIJcqcPfkJKttbeycXTbka64Z+5BqDaVFoQn9DCxWFDTXG9Zikdm
qdjhU1QOOhtBPF1/FWzmazNJpgfE8GbR0mnL1mwtMvI8cfJlhGLKNWb90k5ZsUaMZ2uJ/UTfVqgw
O7fCcYKCxMk1TDTRndoMQ3qSnzIpJnT2j47J1EoMj5ibh6KIgHiEli1SBXhn2cJa9D27dnoZ/QMC
u59rIzPQcMfUNSHM9Gqtaqif3U8lYf1/Tnbhc9w+5EbkewzXVlzTAb8K+3V4V1kVgzuYA5dRMZD/
jQ3rIrEqiK9qlj15xt78K1iSWshCFTv6lNPlBDWys+1j5ZoxY+YfzFxU4+r8Pqq1hj/rOyFmCEGa
OknFqRI388mz9cA6nPZSpmgMT29bYMC15W4kBOkqa5adRrZVkOoobTc37p9TCuPBP0ZmCSuBKcrx
fbh+o64ydlYjwuCotOp+8hoA3r7EfV1BgyOy+Kmp522M5Pu1REG/8f6rraFPI6pfukoeEyn6h2g2
nNtfHOjcEPCDKh6C4hwbQPcQ7GA+Z/IZk8NJ8bppgJquiUK1jZ6AJnVoyXT1fVUirTNJ1uz1bfdn
61gMXzxwDDvLbA2eK9GZkLOEGHhgY//GB9zjNV/1ZS8twT45t/CYzEEddZV5uD2qV0sqhYNqGTaN
zFSCcGbIH5YPqYGU7B2GcX+Ze40sl2Bznxpp6fI9cnRUzrRMFCRUm08PvZ5IlYsvp4tGBgq9RrbR
/Wg3SPArOji+ODqtTWWfrLnauzdQ8BLD2kQJ0OdBtlOWQdA0eiU03bshQnj+h1JOmrstAKYKqjIs
rFbDJeZjCEAVM3DyPNI5KVaMtMZfT4nGLBze8wLd611QfmmYOZ9r2z47xVsv3bPkWk8hegnpxUsR
tNk1NhU6INVBB74JlNtd04Gafm8AbQvxnEYRin6MxvylQDgeBvx2B8tmzQjX8RknpZ7ApHbueq0Q
hnd/pILS71Jj+sXVylgD5Ow4J18dnUnYGc0eLe9ytX193d3CjJeLDEHEZXqKVSdDuHjimBktttIa
Aoka3BgHPZNMR4RS/+CPb1d+kfPCUa0dQN32MbQqe8pP32OYJw3Eh+EKs4x34nQFHBL0l5u2dcPE
3N+I+Mase9VGuho7bWEurCJGSK/zLVGTxrWMHFG3lRsfZVhDSn6TeB1R0dkIiVTe6hHC9PV+txcI
hy4YocE1LVY44Owy8SmM22/3A7NIcuuz/lbk3rIMWq3V2rdCQIbZ3dgjVgUo4LHxLcE4Xm2B6N7A
24fmQP7Yo2Daw0FmtGOqrOIEvxnK26It+AomF+JhcTp5IB9pnPh9YJ1TabETjVuLBp7OYgit6oCZ
QijRX6H/jOzrK7i7SKg4BMx2U2SPg8SWnJ/jHRC0FCvghQPy2cjIQOrlnJfIC64JOOJiZVyZ1AEA
n7NgVJqgbIgAuy82HYdYojSGiVWu1w1vWdPrDfoPDu6BF+zRYAahZgkXNUhHdPn66iCuBNDnB1UN
otNk9iUX40w/RJ2QBCRUBDQhnChf+H6ajwVfMbwir5AhboQLV1x+9bCDYPAlx0ZJIEVz7E/NbqDg
oKPykHPuiym8FZ/u3PbIv1YDshM+rL1IvlAQXifxVGI27tcgjWy6WCkefqYPaFqVhjabmCnhsjdK
lOt5fM3gmFaVIFsJ0upkBRNs9jddWkivGWeWUnrduRvi4EGFHxhkvCx0zgokIzgEXQbcY8O3+iah
tNHzvYxR1qODZMOyjlwLmPil5Jn6R8fMyj4a9sd0I1cSHoJ7WVztrsnoUIdTg95S+6oo+1SQTl+y
o0yui++XJizxkcfN0PBlIPChMpwrntWYAMmGLevaKwQJhETCBUslT311eEIFenpL8zCcIqRJgeED
9oe0l/Q6UMjuyxJ650wwF3qQ7rLn9vUAtU23DomWFgJzpEFw+820r3God9M3HiIap+aQn+kaywr4
NGdo+z0B4tRNYOQVf5ZHY+0IyzYoDabIZupsGxrfH4uy73yvzsp6NaWuKlpqCZLL6PQ9U918AZEP
CXsdBD5cTKdD9H5eK21ZxXbt4PnlePUFLqROjIM5iwCLAxAflcUOsXxO4hdytfTZp0szrE7ahYHV
uHp1Pcj9WXSspBhlq/Mxa3ufj2u1w4/3OTNZGVE0EVBrhBVJSbB0OPT5HzcuHprAqHj/yHijIhAo
Am3DMbYnWvaAN9u5naJirT6qBNdQjfC4AoELM0dXeNi62vPTwp0uEJO2ns3Y2ZZnXuK+sfbl7iC1
I0sa5JpSxSdHjcHzAKaXykB7zZmDAIdSjfp3VdOwiL3y+SBB6TLWi/z/lZepZ1bsT+e7M+xpo+2w
LVraJmsGewVpBENlQb+PXBZIXV/ybZdc5XmV0+qjlHXXsYGhzUKHOYUbnIc5j/vgRMbrES6tGpxM
Ju5uesqKQWJCkroMjPmw2+bR6/Hf1ZEazB0NkqiqFHK9PmIrjLpRlXLxW3HlAm63P51FoJb/4xWE
9YB3f818sfNEy3EXPf/9CGOT+ge7JI+0dGc/+TiTW1sX6bRcW5wSpTpvxq+1xxjcKIYNd61TptkY
Zeum4ZK20PsUWDVK2JKhn6ka4KrzcolpKcJ0z89gXKUTlowPApeYbVkZXVYmtPfWEKsO8BpcNjr2
41m+POP/pbY8ITmOxNEDKrhXRfKBgYf8Bxele0gf97rhFWSJIr0v8UoWOxOVdqoSK3O4s6BvGkgz
DgqJH7LAAw7gC3LY4b/29TohyHBsOI2VwOWhpgRWaOoBZECLfYy/mhfnKZZkREj0nwUZ3/I1ueS2
9DH+JSMTW9Te1l4PTPJ51VEbk4duTN+NpfQ40pvMLKw7iv71i8EoQfEgM0jQ4Zpk1MdA3PmJCnho
2J2LNAzmrGADr87ss81FGIaSn07fic+YYVFTGpt3s0tGPTmdqsNp7Zn2P/nJ3zsL23BKFsgg+0en
S7T+y49AsVSAY3AjGuZ8GytIk3dlV9SOxNSe51Xjt0aDnKZ3N6pSL+6KAflvyg7XrUudiuqIg6SB
vbOKpHeUAZNiNK/fHQ6ly7hvAAEPP4+CMEceBP9PVuhXHxmmamDBsla79dib5AF9H5ZyQqPUWaQn
vLVNKIJx3MJmCMF9iDDjZDf+Ui8vIf2fBVVfpa19J/VbflnCEaYX/fFbItJRB6j+lEN6CBD3Ky+z
kA9MJLBAClG97Ay7/+hhLFL72SOYrGx8tsHOPTvE3UCncxP4Yz1q8HnxVxXPIQ3O+TaKl3QJQ0qR
p5aP0q1DYbtZUzvgzwmxAwnaGcyhSEW/9kHgIaJHe9fHSjOJYH77F8pHtIsbTdQ/b/gSFPOj5hFz
IU3V6CyxQR1mwBSo0HYnaeqEg7ZfT8I+J8Vcj63+i+1O5TIR+rU4YVyLUdPnf0iBNhkuqwqt8PNq
PRPfPXuK0kUFZ9hduJdrgX1YG8paQhS3x0Att3dQBqIORY7YCLUswRYDyuilEAolmZtiD6z2VpLI
hReaLAJJ2KlZwG/sp6DtUq1+c1D+fsdyF7ub4arVqve5To3IM487zCmcjG+sK+GN7fMuqYSelf05
UETIwyv6ByPu8AP+9v0t1tYDKm28KHWtedjWNAHTV6fDaPeKv+9xQnY9TdFLbh6JlyJ/GgB3yNEM
Bz7vQ03ZUF2Bl0sp1ZxIiI2YbI5piWTnyGmpfS9EprsvGgiZ3Vw5LrBUeFkqUparjhfp+0cVYeOt
y3G0u7DGwU1BLGCYkmyIj4w1C/71q8pOjKT09VSzMeYiJdAQe5Ykr2s1Sy+5H809aOJKhrlyqV09
xajuVM0lN2KKg19iULna0pKpK0/H7kE1gQxrb8I+LSZUnM3h6GhV+Z3QrUiJaTVGZ7H6g/Ip2RSF
31jrIPQJrfk+rra18VQOIkzJyjgPBzvRyx4KZCuOmSU4x5GlfLy3LchMrphSdPgNXMbAHwYsEsgZ
MiBD7SDaKNI/zBow+mDNjcy6za81Lyb3BPxraSpq8jlAsExy9w4YwZPfqvpfsX6CBLtU/NhrGnnw
fvtNDZV9U5kJm/SMo1OpAOhZpzIQ7WH9itKROduWtCkV4Sl5IC4jTdwkX3BR5BAAWwaldmDL1Z/F
WPzeygGKe82vVZ+yy+3zq6RgZK3BisSk/iDkjHfdo7bzGF/VgZSpEyUKCYi1sIctPYL2h+buedlp
BHSqV2C9eG8dq87JYn/HwsaRg+BYS6WMwQZQFIrzT0S8DJaSeEMxDrEK2BVNaR/vut7T2zEnEB9P
ZmE5uie9rxGBOS/9QhKt1DR3BWgQLGXfbgUBe+xQ+EWbcS+wLluzHEro1XUuXlTAa61HPYlzlwgT
iiSuWK/g499WoFlEV7s1WGeXHYweR9yKgyrKO8ZXxKmTzU1hUBQcsnXW3KsDWiy5PIuKTx0zJ1eY
3vukkA5EI0wizcWf2RVMY6j1thtTvvK1m7uQ+4hLCFF7P1L8upLcsfonxYCimGY4MGCSPWOrKC5+
siy52tqQeGMcRPxywueOqyKL4jw3KLOaxN5x4XE2jM/C8oRkdZy7kkaHJ8A4Ynu7afYFB6uSPpFj
dksSjGyB2DgBZSb0CNs79SyoVksOnhaUwkNqaZRmZyyyuioYn0et+L4Po/qmtz2wKZgjKygVcubR
oYycJDd3Ft4T1V6/nrTt4XFzgTn9eTMLNPrz+2HhfrOEqpy9smQncNPMC2Wxt7tb0OLnJEodAOKl
o8Jn3Gs0SseiU2cRDiCYDXDlBRq7QuKJUzNlnf21rq0ypI/XMNxuRTJt1nWw4ET0S9kabCr4epf2
P5Y8PIk+3N5fab8Ku13TwFh/0LaAiXKt/vilAQ3///g+jGL7LFofUfQwVIVf4nACix3FcFcEWt0/
IZnRjEc18bwlU4eKc9EdX8/kWA20E+KruW6Ws40uydfe8iqjLgozuA3gtAwQRiaE4nLc2QeFX/cl
ad6neTUG99BpinTCg/LWyXiY/Xk0YTU+neadekk93C8aLrLRdE+rmEAXv0Qz+cYLbd1FihQaTEQ0
vAe4rb45kIN/133Fbog1djfZIjmwXM2Xawmy9TjUpiYIi0hoix5cCpiq9LZrfsELESTxgixTuYR+
sROtM6egXvamOKhK0VEoOLca7e6Rmen+Sjp2CaQyVJnAQQ1p3pzjeIt/ebpVoRlDibm9yatXvsh/
MbKvdt0GbM1MSG72V0QEU09AeTKBgwiBIDdONMkEK1jpAO0tgZ/ipKunwlnOvaljBW4A8qvrrIXO
+uf44xfG+X7Yl1f/t5l6alZCCF1/A/2/HJTHod2+7uUCbimgpdSmexqrhjcnWM7e7abuGUBoEJHi
nZrkipomUVpVeU3uv1pDrht6j7mCbVnCSz2N1tDYEDBg088lYMODFks+FfIb+i2F9soOW+duWiUN
OTdZydneqb9i8V5Kh6cTIosuIW7mVYMsdCIBbE/6/ESKYSCqaa/vM4SYpY89nEMsYd8gZm4FBOzE
sZwr7Y93MS8YLBMLpIHhlMcuCtliTtnZ6DHL0d5pJr3I9FyIZ+vYfNPpJALAlCfQm4onIS8QKBpj
8oVL8o9sF3HtCA0Co3l7+nfpZajaOFSq6KtTX2PyQtSQ8o0v+oI8UDNMSJPISyFR1MchhG4Ptedr
zojXXJX1JQWPuVA6elTzvQkWYGQCLh3pGSbxRiNM8D4tMuIQWoLoyh0TgFlKsa+zKQ8atcQR8nyG
4KJR86jyaxiFmDQSeykCnsrZFD9OkjGNrI9HG7qjr2L9+cddmPTfAU/asL27o+pvb4XhN4BQF5n6
s96gB+AjwdUZ2A+Y5Mm8UCwJsrrZsOSxV1AgzXtV4x7Dp6sNcZWL9BTRRC84oCCfYCK4pTku+Fus
mBnlnv61ZyoBjXKhl4IFNBegDsukwZ081Tb9gySMRtKJ0MYv7ZGMPPDUhidEu4N2iLsm0xUZ7vHT
RVYwexf60n0nMLZ7WVS399kqXmOaxNA9A5jZipXKGZ4iJ6wX7FhzRxqkTbgjw0VjrGMZ98HMX847
QUqpd5hGbiMGEkodjizxaOp9aDPbuUAO4N8Jvzo/AiGtqbV2IKziLmFUYXPFqJbU5HUWhX2lEp7n
12x+srJOIrSz+W5bHzTtVGnPRm/gnbBL3OhS6Iytcftn5ljDbpTc1pJufde1hvLqx0sz7Ih59kGU
j1gECYSQO+yR1zsDnq29Mx5Tvo+wOKTrS/9owLnX4GNFToya69V6KajLsWt2KpGiAmy5FIz0g9Rs
Q9liaeCiFojC7yx2uf6xT6xT9tAJQu1f6lschpTUeFjaV0fpjNKRMVsJQP0qd0kDGAPntdiJeEq/
/BO1C3n+6RsADdu8kl/vt+4ikbgsQFVipkUEPea1sdP1uJLoXaELHzGWdUqN04uXjzHanLurv5cg
WfXIcG7K8/CKzNkNLbBB2V3bjQHTlzUdEz24GQ/v3NIYRRPpraKZQhzBtJ848BbRwcLA/tSv5VkN
FwcX+p1mLBtMsj/q6thma+PP7uHw/LClEh5uk9zV16GIISY6zIGU3u3ffvweiKWvqPhssV6EdqBm
FYfYY5okeHBmZnCgJxxAMzScsW/UUXu6mMJOryIh2OE6ICX98bNwnSOANmSsL8iay19BVGKqACoF
zc2kcs8ikjlYVAf+G9G04jVZrSP1jLn3kkndHdSHu4gfWOcyx5ZRawoKtyFJckMcXBTXe8R++4fF
JaTnidMeKngGM3QcxS2eW4IjG9lx91fkmoD5vl5U1Dt9m6n/kjOIJuqMpAD6n1eRVyji81DyDHgB
miFoP6ZJOUu2ohWU5EWmro5Pb3RsaFXbXI9rtIwVR0k7rAt76AXwqyOoJTgw0pYIEeMWHTQGb3rA
vQaNLUEkwSMj9WCz/y6dPtnbok2Nfho1GvAv+nGwZTBL/v6WkWnfnkmiIvM39dU4m4WReyJO2z5V
bWL261RdG/u+bX82D5a6Uvq+VP0ePQ65AyUjmMKSt5OfppEZHr23GXZMOOL6R6WqR7Y0LVdR6cl0
tlVOE41RcHezPj6j3qW8O9jECUluZDztEf6gpQxPkAAh4dAx6a94Ba5bQ78vJFJDYF9ECLobnFe2
dm1sG3uHinWQpiznKMwNuuQN3LEchesDKXez63ukhct2ajHz8ZamIeMYFbufr1KDFM9D5eaeinFc
kFbSnKtptkpv7BTh6U4tffXJCm8kn0owIm47neNiVO0N11JqKjZiMQYszMZJ7XwCD2hwYmIdYmtw
7pNrvSLe827AJcKNj6qCggs80ugoFaWzK/7DTdaxxDnGKaYVc2XdsP9BibLIIWOIUD8fGT7wvjzI
9MyaPyrIDbv5h7S0MgXuEkYPy5gk+9OzA/0qEkWdz08HKj61S0q/fgoPb6swGaeC0kMA3rLMKlW7
8QFqpaH1koutN8f1eb+vpv91nNRWZIjvlvw0A2SfcbdZHLBmcbIuMMm7kK40pY2jsS3vfwExd++I
dRnHwauY9VTZNvk2S50baxKPU0Lx8lPpgCVcWtetd52ihH/PMbMwhSL7j2pwYowhsNZzwy9X13NZ
Wdz2ZgZmYMKHLnLGKqTNQSuhWTx9WTRmKY7HGg3SZJCYPzAfJ6nGf0Lmd6NLPg7FMtkq4GzmZ5BN
2mUJmdtiG/fb+nfj6MVon+zC3HLX2LYtq5MEnUpycrAsHjB9BY8nz6MlLn0b+2jPE9bOOstVzMYs
64+ovOT28kQTRO2J6KDZqIsOQVwCANcYkxQgo4tp2uxGW5HLyqDr/e/V5ED44J5l/NMfYJAJ11fq
O+NKdnF7Noi5fzLUoBiBVHBC7SXKztHhCTWf2DFcq22tPSHRnPtuCSbpXS4xNcP9niPkbZJhVU/8
uKYgIRP2lvEqfKJnIKxZVevlqmYOGykrndXO+0nXQI9t3nI+m21AERJ0Tg4EBVGW5BBPl0hmnsew
PX4ypcvDyZR3E3Bu8x3sOq2P775l1wAlYs6TEhowj9URKgOb09/3pjrrpodTXdbl/xP86E696Si1
kTZm41j9+d+3UFkEDJ0NaJPLFEEKiVtJ81jluIb6Y9DagjNaKMoA+Rj6b1nJq4Fg6hm9HbuVjBzz
ndfUbUS3eCuu1SNMyniv+ks/YSjvScbjjwtC+SUoFKpsF4LDyL9Az6k7egG1S5fC7exuUtmD/t54
uj9hNZsKMaM2n/HMQaNqpHAovrXInIiQoQHyc1ilCl/sb3lvaxJ5GCqC9BUQmiglqu78LN9NAUna
oOgeDdaPqPliFP01T0Ie0GApoL4X71Z6/Zxq8SDdeOKoTld9a+9iuQA/geTj71X3J2HeijeByMBP
K07sPOUVb6i+/YRG6u824Pi0FvrZvMOFanQvHQtiUucWJ/bo5VUoeLZyRHoP0iZJkcA5wY6s521R
QQWyuCjFvDka7MvdJ8l89o4KLt6b81sDj+Ni298tkt0c9lB3Cl2ceg0R3YudWuT4HRfWYuBMSw7X
K4TZyy7CLctOUdAkJ9/mceCRnT1vJIEv8GMfQP7lFv6qN+iy/dgx/IR7oFPweJEH0EqfhXNzzlKk
1ms0E3NCjV08esBMY/V0/XGJRxRZqTgYJaN0CVRvaLX3nBZQcWchDksdBjO8Ou4pzzcICbCRr1Gs
BGuWresnmCLro3o4n9cr4yzIfnuFVDArYO92a5hEnW2AQwNX6ij7JkeSHoASxYVggyCpXme9StWZ
znB8EMjumpKoL0YyTNF8H7W3d8yunZs356pg6T7KdFk8ZTM6ryWZ/8iBmvJVQr8zykCiDZn3a14h
tC6Q+vbXojKNpJoz9hhevPJu9ttUzpTgsZohOXyMGqIT7hlcqbGqr8aDPSGYZ2113KnvdAjDkkmW
k7VyYSn1Rg1zdb5OoCaWAR5pkNKxJOHvcgWv3lMw8jKqzrUyC/ezjqJXNVGeinY2Y4nSgtkXUjrX
+UTA+//saGznxN+Bw1OuK31iXpnVaiAxodgWhCdP3SdcDGyCTP8qsJnIMdSm+ujYgvJh1Y8jGRc2
o6LUTktL5SBAft2wgmCF7Vqi2of8uoc8d791oSsT3tpR2WoYmaysvsf33xfxz+2SH3Awsf9P2zhU
a0WIQQknyL8Mlzy1sE2PjcZZS3rvzXi/L5mjv/Ie16TOrU1WbBDc/dicjNZ5NSMFeC8mF4xputFh
1F5e2WyCgdQhMVeKE13Hwt3PKmZ5h7yAUjwdKCvsElRa5TlZ6Jm+5w1z21PQtIBJaFhYjUO75i+H
AeOXp6lqpmG6qUvCV2G7meB1Z0SW/m2GVPBfrVzdxQofW0pK6CB+YOm25Vvut0fpBXU3zJ9AQFsi
X/WGPb8BUfTQoGhhNINxstxDWUUMEh/fMgH7BowEOFQY1ukHC/vyUUvf3T04DIoaf2MQNhZcYYbp
s+ZDFo4BizcbTAaFTd/4H85fbI1g7kEGxS3Znyew+E08WdAp5CjpDR8eab+s1SvOymCt7xRijE+k
cNa+T5hkMearp7dg2yBO8fovZxIkfnSe5nJDdnvAJhunofyvojFBeGaPHjf+VRL37LQqp0mvSIH8
jMh+YCiSs24Gt3JjXI8W2VAPTF5d0uQfQf6eRx6CeDcfOsqEstQyRE5JESwdUl7M/RMp/spkWBAV
8WSPXb4Sw2yeBm6XfNLWCXHVeVGb15puZrgXbgO0PhH1c4me/cxrnYG/waw0adspu+sazleTbtM1
PYaAzRNFEzdsdfUOu5HDDcEl9hwnektmzA/ruGDSMBI+qaZ9/cWaOMgzBZG4ZtS1gqIR9oPBvGlM
w4bpSofLWxvYbr4NQHRf3lZnFFEIJA77T1aOEjzaDjVvUIlLu+hGFwCKDfbad+udk/AQj5YGyLbi
mP3MQudh9WIeoDBxqfNFPUiq/eyWBDut2oCjA1dPECtKRFjA1bDY30aaX+YePRUWZjJxeOsaZhda
UOHSzo7fxW9jTcF1ahnoRYow3H49CU/mVwb8dqs5vNRo+7mW8/djqrT0Fm1JgjOIVNKQDYoyjjxM
tY6pcfl9D/x7c5/FHdyS4Ls8ro2LOx6cSGQn9gU+P9mN8tkgYpT51BO55IjQaX6Qyq5VD6mcmYti
9GuOTsHI6tUm/DiVmeXt04cvxkXua37cP5SmtAWW2z8JZRcJxZWREdtTO+OS+fMazTZ5T0ZLTo5i
DxLN6u4G1i0fh9G80cYTnOV0rkfEvMVqV6LEIb73GmosFLWZAcLWOBH7cP9OmuvRuBun6TQuuNxG
TM8Q9gBFVVlA5Dmf7Atlb/Vp2ydJ+ITZ1mBOEjD3XDeCw9NtSAnH0bJq3ezYxHNuL9Xbbhgjuy4A
0VyQ0z36C/91BZlNnPIzwhZocO2mwHYEeikveWx4Rk5tWQ7Xhk6mwo6s2eiIc2xwVgcwevbivgEg
OCHGpnr/vFIH317s12aSzcD+KqM8oOzQtoF9n/zBflg4FuopqIu6niyQeBCm3uWVQrxA5ghKxpjq
kebNg+Rmbh+6kXDoO3hCd/oLCgqPxcMb5UXFVqKPHRErUfcshhpDA0ATP77asILnp09DTXq8FiyN
pn8nM0f7U/AcEnW6r0KoukEHlQS03flKLMmbktMCwppj9+vFmeKtcZiKNm/91AdGhTSHLBoWxk0L
xDvw8EsYp+PqmgN6MoAsxjX8utyU36pDtAAC6pEL3qMXVwF7SPFTlvDZFuH/axwuJx0CDxyxeQOZ
fF68HXZQra/raDfzyUbdfGjKLUzrVBid55Witv/uN758618DiOpCnINQGfENaTpvBV2DlA4EKbja
+qKzQ5OBSvsfu5WBjcYdDpXq0YtvitVLOZXTueFeM48Nbuzl7dC1RyFv/CyU4WcfortHfgwAhmrJ
jNvVVjrt4eQWTWYwDE8R0FcPk9+slTBv0fNM0xxnKUir9upPUQ79kiRl8tlkyI4rolJlQhbo0W4b
vF1qdMBsIJvgwThDYvnu3Iig1+mm5Z+sfgbpG0++3UgGyoBJIlIlHX4I6pb0OAfv0De4cXTLvUBz
rRdj+VbxuucleFlUaanWqcXM2wbMkWYIHLqP+/gxMAzfilbnzPP3MVtTLk0y0akIKeONfaUD+Vy9
/roIvFhwBFTgYxo9aEJrmZlyqWEMMnEAcatkyTDIYWuSUT9S6AGQbXOhz0vrWLdeMTMmDzPIqBYQ
62dK/F3AGVDlWINCZ0Xg5Caa9YDk6rGnHaBHBU0C9AYNcluOg/pIG5/yHfQUWdSOsBM8HKgE8BSg
E7nsu5pI0sEA/EQZ3ZonZ2w2UbiGA4+nxpsmt8ICN45idaM0j9jGHA6rxk9IMWoJaEN09p192+np
DifFffwuYga/UpCkd8ByFA4HWEW3G4EUQ9LipGAkSDLfgK8ou5GQmKV5+WwVLaivW7VuPqrYneLC
z2wc8IIGfmRBBo805kcISov55SJxOcdP7Bw1j3RuQcmBfkuUPb3s5+Bj/x7UY3dG+VJMUyRgW7VS
vdXzLFGlsyzwnZSovaLGmoMF8b2HvncOLAFVfkP/VMxgQWB5p48Er4/ezYGXYcNoOyuNnrHnPm3t
vrQ5HpWG+h/MS/Ru5DurIC0JwF0Z129tOYCNsoPGixJsNSZ8URLLhnWbAVITjyg5+VdZWqzoRJbw
XOXWeaQmOuooN4UXB+gPrKLeF0OgExzz96UJ7rKWgiIS7aTPaKtzBdzhZbbgWELvxEzFBKEVFzKb
2MULfeZqlTHNf2NPJOlLQHB4/l7hhQxLbXw/qiABJHZD6TGiK7sBlFQ7kJTsQUZWz9vTZdnRnkMO
AGDC+OPWXoSYaGNhlrW7w1JqOMQDLAmYRRJfJKmR0Blh15VPtnxaGeU/aiwbt0VQ5hmEtaMVLjmu
kpoA6DL2JrSD43/swCUlTSdBPpe3ot19wE91T6dBRV7bOYkg4aytBTj2vmIvEuH2VLLQ9aJoA4th
sHcXk9dHV09Xz/LZ58hv/RtWuois245/KkrFJ5P+lxXUTdh2LCVwIFLt+jlSn6+1paolBWh/NIRE
zcf5i2dnxSjytPj+RI3ZheR5Y/KapjB8luLnuPvWr3MjHah8MKlyfSODFWTYv44mZjDSESOu6ix9
Mo1VgDheCvftX4lcjVRjtbTzzo+upxiJfyCRQR1wgj9wYr/wzMnYBC0pBiZu4Ff3xugx6OPfh5bK
H8mZfkWdHwmkKDBUqfQo+vbh8EJA+SP8srmPIP0/RDDeklOwM8Q8q6Iy1ylhF2q5JbrCLeCBG6Ha
i9lL5XvgHC168wZ5ybgt9b+aq0uL2LTOvWnL2PqPvySZjalREevvE9MxdGF3usBo1p+2POowHZNf
sTTaKhpLE+hE2wg9hS6hDLCmamGZyUuY3v64by2CJMbh2xIzDlXyqXsZD1g8XvamjNSRduWcvAFv
NfDxXmLyd2UBpamqDzfJuXftrroF2+/Y6yIkmzhQLm/oqqdqvZKIhthu8Ka5P7gLMUuSs6GC8Ofj
M6fH2L9YV/kvXlOg5ILstfQKoFAwOfhNtf76t86VuVLNFnk9hWwfdtPQHkVqoBskPgC0Ovml1spv
DLIYmhXV0wGQUDdhL2/i/WTnQrtDD6EAk8uP/fOPwlyv6agx7cqu6c08mxQzjrRO7uRomUx2fZdr
wq4jXN99ERh2lkIbbky53sf4+2Dq0TYWoXAbuMfG4OepzfwWT3Jgx3KaNV5SU7hvXrDpt5d6H8Xg
U9RzxnNecTKijWx8NMmqtH068nkK6P4d9423+zs0mrDm2B0csm2VtClwKRKgqEnys3qoG6Lp1I4t
wuVV4LBe8iBbTnNReGnh+RyNNYJysi9q+r3Pc7Xq5imNXQAdB4x4yWijT65+1nqwJO8jnByf4df1
kRuc3r11+L/8CR2e2/PuBW8k6kJAVTuynNj2HzzH5GQ1BCTQGLeb0ivZvXmwxwgA0mR/uCHZmNJV
pKK9dEVNo8QFq4dL4yuEVM9VC1oAskt++p+xnhIwY5ebt5kTLwdWdkoS+3VN4xPDDBkNLTZmcRkk
cj/M40MtWZf6nWFc7gug5v+b95I3J2Hwqg+jAL1e8wCRzOTwgGCuq2fdUFf+HQrGv5ZQyscSsGU4
J98ynbtI88jLWE+dNYE8w2DnWM86l/4YTdYSHQ5ROIYC2sa8jJ1ircaBtlHFy9rR0jYo6eXvGqrf
UCh05L6OlqjKc+2goDbRtNwuLS48Gi/mg61w1+nVCTSri+e5Yy3Ue0uD5PFwV8e5NPUJmoNNh7JU
DsVYEYdXBjiB8beuZWlSHdafu8VUktnFvzHkuX02qSY44WoLjCmbb3h7re0/x4e/jDUxmAHFg1qs
OdS9eCJhDuiktIRgNMT/ioC5sO2hZ40iyOPEhC7g0CEMDNpvuDXTSmVYGG2F+qVlKRIkWzffygZA
emg80AUbpILX5IFTmxMF7KRr0K+E2FgCQoE+MR6GsO5ef3wt5vnxKjUG8GO4n5KU+713dXFIAPob
wQwTxH9fBJ/VlhughnSJhO+/Unkk2BoJdCNjakPtwxuKl5Fjy6DzLdp7cCxI9SI40AshGbR3LOh8
Sh007CzVSb7PBCahQsJNfFXcP++T6axjLTpMmru6wwoBDI2U9FdDt9Nz+fke4M71LvX5Y0keFxLs
wjkQWT8Jebh3AKS7jvNVotBwpexe7YSKYcuOSAqy8UWhxRLAKsDeSYUk4FbO1HatEq6kvY0nu7bZ
/QqiAqD7Q72S7hE8yFqzn3V+YqSe2kc/WuUgkk25phDs/1voH//u0bSJ8VY19+QFeg8d1jj4722c
muE/9YjJO7fwk+ZVe0SaPrxjr3+Zsc4es1kSGbukAzak76YT1GeHwc6pW0f3JXNK+TfT19CcjnaJ
hKu8+eJCxeS5dDz3NRSb+O+AStALajw9Rn40oRjNQjZwJa+inJxq1Yh38WMuVesmcYS1p4114I9+
ki3ti9zTRpgZh52g3IGqqQIrNJhHqIrVgoR9d9r1EIEYk0HKyi3rGXbo/YmjRAT4U2l+t1qchWbB
srHIIDfEt546b6wtHk8n7aMmc2TZfaeI62i5qaN4BcdamDtv5FBox5xyvLyyPfQ1Cuf2W6eRHe7t
YRMX4yoCpILGjHn2C0Sli6WG1kBQNXGq3coeYZCtEIgipUcrNOZrYXM3Nm3caQOsaMm35sr3PLFp
TuRxiI639HngkKDFguOBVTICuz5i4C9Lo7a2awfGLbb/fpiXNXfE5BqZwV/q6q9MtEVhgIYoq4AM
lySslq5wxLmK6OnCJc4dE7nwAv2pIrSTJMl/7jUMR0T0wxK7pAuyoMVN5cHxyTSntrjgE4+EJwCO
XwFd0UnUL90f2Y9U09tckjgbJFtiaG/pREThZcv32DCvMA7QZQHuOldIVL3nJO+ZeJlqsevxac10
5hdNVuT61cocY23iev/O1EAuqo6Wi6dtuKE1FOVGwVNnSkSBaELPlvIGbnB6ADrOfDYC8+bEJ1Qx
7iN2vvWGRwH9ieQl0rRyncMiqObTWrBS5oWEsSU5OH/RuSxj8NvsNSeazqqGMRRoKrGz3/SOxUch
t6158qi1VL2+5FUtRi/0MejsaSr7FQu7K0AEAFwuiE6hPR6kaJQOuPsY25aBCJvDUgTwYd9OhhMe
oE6gZ+KfGuDI/JYVHOl386fZwb/Poe1Xog8hwOUlh1DUomD2mThPERYUgklBNZ7Fuz2If0gXW016
c+vF5+lrR2BNXP9dc0YJeH/2nCg4HKylWZ65JeUgjPBLBswm9MHBI6BCUQfHzEScVC+laG7XL7o8
bx5WQXsnVrHaZcgiCi47ucYUKGors58d44YetF84ln6RCXvKa7Y07E+OrSeARAHngLADS+SiRRsj
GdwQhYg5m0CmxjqqL8aJ+h7xB0nxtGCXh2WQ0rVW/HgQx87fwvmTaXndNlzoI5F0Lr+UYf8qXbj5
sCYvfNSH/decVV94xdvDvMuMfcCEOPg5cEH87E+KBRoIsUBHmlvugWSQK4UXmwY7jW5YEbtYP+AU
tYoE/yFtJ+dDp0SkfOVRhyYbnN9CcuzsrIHDEAaAsTNcvdCNPPWPwPzVsRpzE6y8sK9132O06Zrk
JD6+Upc8jW8Tyl5fAh7rpL0MSkT03T3qWnCuXWevkiF+VQtvhHkSeDwUh2SRmBg8CEPDrB4mR7zo
+Rrewlx+H6nJVnRskrzm5szqh03HjF1f9wIW5YHQp82F9Y82RIvZRGDTnyK2bDgnebhZ1BOKDA2K
Zfq87kSe7TWAGdXLKJjkhzj0Tj8As6vvUbbtIoQl6f8WOdYyanjzNBhvPFzIZapynMBtkNQnYkjc
PrMeqxRfcM8E7spYkJlGaQV0r4VsPT8QwmWxtN/kOTSrtpwdWAlUzMI+QPvmsVnBn2XffZM9QUtm
ATMk8bH/I1huapunjVABgHJstL1xlpaZRsqMiuVyEU/UXjsjYr9l54yZMBVAeAGsuI3NUkLycKuy
nviA7KS+aywJpaAaWKesTtmbATZkke0uAcbPuPgxSv8ItS+2a1y4DeaNNIGbAdfhbrTWl9ZM8/Mp
/L3i35l3JLgvy9U/VH2/9qc8BVjxlMbUKrNzmIxZn1akRnzmpn1lH0zdqO1oeOvgikhonHD9f/qS
9MW3oLCsgiCGcrgOzvkFcK116kX1sri8gcg4rF0J5c+ne9ydntyiAtaunE26b/OBsZX1wDWL3S3G
0oS87TVuF20zGv+NYpcki5/cIR+kpHr0xXPKZB+ZugQaHVd7qhcnFSZnXuXWHxeyCDhREq8lPY5f
BTKZNTyhNr0Tg903YHMRlXG4uGNpZTyeV2UUf+otST/pe633dPv+3aJbb38QCZEQqFmvV5XQfhZn
YQHQZD4cPGcT9i57KvHA3PrkJCIy97cVh4i24gyf+yITfCQlBoniSpLh82CDLTnwPkkC/r8xG80b
9ff8Bp4fd1NW4hd5iq+h0ceTl5syq6XGluIj8NgTsiZnpK7T2WGHHDti25bOjw8uNtVi5Hx3Z16p
jlsaQjOlIQQl87SpUp9Mm5QshX9Oppug0VafP9Kc0GFDIqwc9OdA6QwoZ+A36wEoe+6QqNcy1Zd0
yWgtwlUMrH8aDU4X9YNiB2Ikl0/UGZLlAOXgEaxij1nCK/3NuNiJ5jQ74tv649bo+TMKRybjVbJl
isDgeR6qq4fpjGE2sZNnV5qCHZyuLmKeGlJKMkq3kjZ5VxoQG2MnaoRvEEqtYpMldE+hleiFNxaU
6xKTLrC96/HPIUDkLyWEXz+7AyOXW9POhyNCnNchmqruNHmWisHMRYinG4cCOwOmqoaJDSKPX1lO
BAcCxIixXBEdzO/3XbFXa82jVSzOjXyLDGW+7vs5HSAkDZpzBwF177b5HrbAsipyee2RNMJDLeL8
QdDyLVF0+1Nxhi6UesGeDncZUOCnZ6Xhi5Gj2KAKrWRepIv+fNO0xNn7okyDTcNnekWj0RMfYU81
GFL9p8gQZzba1WOCNVccAIfs2yxtO9EXMHh9fzwRlJtmShVZGo9Eeb1l6OItIqBtd5ZYdmiDacCg
zIwWJsLDxdLt/Yn7XuWNGkj0MieeH0MJerLYatGgGntnRnmUyjB2TufxMI0DN/rqKFiHQiqVJFqi
EXNbMXmy82wO/QFMMrXU5A0zb30JFPLo0erWPckSnDr47/cjfGSh7GEKaa67NReisBSc+4UuQy91
px6LpBsQtjcevPfnDbrPxH3Gb/BUZdyfnLMbe39Uy8tCX12Ixt58tQQvVLkjfuR9ydWLREAdemRb
E6Ca+oiDa4G7fLKvn5qFS4goaffEksCyfptsa5MxAdO/VGAWY6lnI1vAMtMZSEIJgJtWjy8MKu0Y
dtuIpmtYJT2FDx6OKCCKTGXYxYWBTXPa6isafRWq931+FzvmRiS4Q3VNPTerURxYPtVOtajMjXMA
vFf+JG1A+Qg+VzjYVhcEwq+i1UAC3rGelyylP6hI8x+ntoOD9eO7EuOClJjg80zhqgbEGz/iTk+Y
WisgaPOZv41y4LtWno+NFqfpDiGCXbDZJxEF+Alx44l+xSRyvx4XdTvesuaym+t+DGwGMZJwya5N
TQzMv6LmVpbqo9XxZqc8h6dsonfGHQ7jL4qROgKdw86nPSFiAKqNEQoRxldXpVNEKPujam4Y3cnb
d/4224EwQOPeioa5L9pEX6LGTsq4UnduWBlPN+U4H1VP+hpeuFMD57Xk1J7lmQnPSo/HiHSwRUz6
EPdtBA13/sVoEZHg40ZXsk4tawBQpLJT5RkO4jSVSk+8liugKo5Pq5bBaOcP8qw5ULVCvYdt/s7o
GMGKVCvOJaQAvlRQ6xQe/oMB+ecqsOd32i23n5J6x/VoaivutLW12USUJ7mFtjsLk4mYZAPd4rm+
T4A2llxefMCoOoeTqtaImBqx8N1/7fPmrZj91DAJSth7IX+BdNf5r+3wTnZ1Ztfz9Lf6kHd1mjjt
aKc9o7UIImyNYBczx99jqSXLeNCdO2ETXmaRaALpViS8TRVvDIvXIlhqvaON993jToRjCtpIT1IW
BbhvkoL64hfDEJ+v+ccN1WGUPAsKQpJjrmdBlSMPybP2KYlcbyEZnwUzoHQm5kdDgZDWgUwkLU2R
FtrGQgbonlZB8c2Kg/1VOqs1EEFtmhyUN/1AllEEvUqSnFnaDpKxuWs6fm0paIeJCs0LpsYi4LL6
P2y3JTDodVeLTNRQdOwDtvklgf7D8dhPZ6Kix6JlFffOttvtHiv86iHaV614STuxOl8lovu/P5X9
rGi4P0MtAZuIixrZaKvwmZIr1Lgn0Oekd1/ij9sHFa3drID0EYwN9G1+MpPyw67D2JWPEe+ngZcP
1kv2fFNDqFul7cyPxRnqr/0B0R4uS+awBWYzAqJtn4w0Hm8yo/ul6AGsJk9UqPQbx/T7cbg8h9fV
PKwSC0OTvQiDVcskZd/135nqqbn7CpzkMjFOV40aF7bsPoWHp4LLUFG6ayUnz0eW6OvLNu648v5m
yqDISN6/sJ2MSBHPVUsXraJn+yT4XbnozL3972cJrdKrZhcs2GX11wuY+Ls0/OrPmxgHB85Ya/gF
yPUlaifRyrxhztrI4xJnO+i6RAvv8iq/80ufNuADgGV1036zZ0awNaRJr7qCudaNb1rkLdj/Hp+z
y3G8ggR7AYxsnXye2/9ltR4TSdDe9vq4QLFN0QhpAZEOLxqmU06gbsuhegGp0CrgpPeb7MQgjAq9
gXm5JLl6XBkzBRkjGmIAR+yiDc1A56JoTcSfS4RdAEEcroUiLtTqRVbo7miIRfCrBlooVGdsoNIt
Y4u0ZAp9DV4SK1xpb7ZZGW1xBQpNCw81vZzyakoakorrOJM6l4DSHfmUSA36sUGKLRkEW7uqSign
ornxP5jd0rihxu3xzz7T1Do6P0Lu/O9dlmoaZtO7EiLw3mLWs6d47mzxsDCu6ym42YiFEpjCdDTn
3gDQ00nKc4ysmx+ap/RhZZImdxpGpuoqcA8xqMmfzhRs/8ixGSrjUIiX/+Ux6fXZZQyx0eye5z5y
Vp1kDrCZplb4MCmosQIOnVY8iKMqdSczLm96FBG5QD3oL7TcjYFgKH1jZsGHJSzhGLZc5y987xjm
7v8E7QNUvEHJbO3e4dqRRI/ce62jXPLzWkPzd7jyMdAB9JJmIUtponMBy9R+lM0rLW0YmUEmrDDK
mv1L/X/VqpxDOFsj51Ud6/ZcRzWpyYsjNzVQ79xfGo7hp5G8jJYvuAa7WCX96lw7yrUgKWWk01vh
NgNtrNyOtXgTnmHIbLvZt59B4rAlq53DDFFajCgt0z/Pri/1s3OBBpdjZSuyjHRLzhKXxbXelm8h
5x2yrmPLroYKGCxnJp76VNBo1B8r0j+K+70RBlolej6oGWRs/IZTYONm+n2X7DD+vjQZM8l6ySUH
7RWFCEUDbPrgR0NoGFo4/o0ZPDG/fCruOkNRk1J9jKTSl1S36HnvnP2ZELiIwpSCUMDET/52qP/l
RUeeBXIhkzBh6yNhINhZgnSfeTxqEQNWlRoduwsJtFw0tlPvvNEjFEZRTzhpTdNxUD9QX2wR81Jw
6b7a7JR8rtKhT+YvcJHlBcQwYP9pC59uL5wtAZyokKUuqrzlaPU1TBbkPJbC4qoR2umfzWOPdj5Y
jnAo1jLo9YJ5sKhzhHNdbq3wRcAIlpLaG8qOZLCq3sosUbI/a45NMgNy+Z0e5z4WwXsyAID/Va5V
0SUBEVmNlteI7njk4I5bk3jbZUlKRBlDUIyMYlzODoFmcwetrb+Nzfd5MZgO0SUxnEzDSXJLw2bH
YI8WMQiJwC+NhxjVKEBSkg7pADkl3VCcrxxMzkSAQQX8VUPM2CaQ01UcTaewXdqdfiTrRuDvdOH+
PUHLb31X1ryIgFxg6p9H3yf1EH6exGO9fvBZXBL+xVdD82tOWf2VLys+7Lb1fyEFKNW1AEFp6GSv
1zCxKsUo8IVzbN2vZQmHzeFsS/oIYf3pbevsJVecAgiqIg/hyEEEod9ZWek77Y6jlUvVfJvX8Ouh
11/MRTNKXQeRVQWEHsg7qNvja7cyUFQWD9T2qrm4h78OyRC+ZwfXpMBZzhpLU6VwP7efxTJ2LbBa
P4qZ8hjy0miB5/TJ2464rYzKDWvCWR1MvgCB6IeF51RWyzlgoM5Pyt+egh0gnKPUBBccSWy8zk/F
+haQRv4TmPXEskpS91Vq9q7mT0nEYd6deya8tI5MGo2nlGw1XxWIjsmUTgxYDOSKsKs+eizDlske
hJj308S6EgsvuMd8u9R3BgZ70dJlAbNlMIjgtPq6eHaoIcNrHevGWnjyr9elmLyLbBtyaaempXwD
x3UfJvjkPWv7GReiPeOX0/TEa+O5+RndNxFLgYt6CoTnSRSs4Bszfb1uW8G50+ABcUVOqyM+1QWy
uA6jP9Zya2dnN6KvzEw433AYBR0lK3VgpxLoLE3lqqpZ4iuv71zbG7WaUX41Xeps5ActPm/sF9VK
1pGOLsziCJBPD7qBnjVX4LvBnaxgWccDV4MZNCUdRWIShy6oITPmu6J4J/HeN5cAJ+x3ID6HvM5V
Po0l9uAuobm+XE5S1j269cN5woX9Rkt8/0KJj3+Pbe/SlWbPPiDcYqZBv9z4KlmT+nh7jiYmHBzf
I4huSi3dw9flwNa2A6xhdmjWLz5ApMmwQzIlLWe1DeKHMbW4vsjf01vpP6lASSmMMx/YkoRXGpAL
vimgn2p3Bu4/KVrG1rUaCTJJdixcc+UXmjo7Kp8Pm1aCyU0EdBNsZvkR/1MODKGa9nXxLW6HrqA2
K3mGEHyq4sS0DWwmIb1RrW8UQM1KvkrW0HOla7RwGyAcR/m90b1mTVFitvxsIzHHKsXKZ7unT+mB
IocHf+88r1r4xTl/WOaAS3gQ1KGJMiXeeDSTytJH0S9Bpm5jo8lUdgP8qhylweX6QffJDjHmfc1F
P8/Sz7YfrtEYY4kxHHvxVZx77owA0nDN3Y6/D5+gB1i0NqIPTh7/730bdyataAeKs9XyxcA1oTpy
9jzWTp8APFJuhF01a1+G3RNe7+JWdoqs3+w72jy/ILAtsCurjvBpRYLfGUpuE6sofucSEbfm0V+L
8cnu2wyOqRBoZfhLnRfzAOKj54O15R0pzKbH8Zh8SfNppl0sLIlvz4G2xT6P1HVR6Px+jimguYpo
4k+N4e8ooYhbnAwIJPvsTNRlo9n5BmEHJ3bgNxRokM3lDqXQ9Grf5Fhi5LvDhWDMrnMEIPXfEyYP
JD4y99zOi7wIxU07W5i3ZyPdovW1Xduz22t8JVYuN87LIHvM1wVu72ulSKeTckqO3D/ZmHYSAAGE
yEld9iFE5edfYjS92qSfuZCYVJJA0qSMHMLrMhcHbAlq7IMBpsCaemyH2uPQrN6tWvQ72z9SAZG7
KaaebbKdBp59OpfoCRXQYKNxPd1hmowdCmA+uZka4iiYyl5qyruqNRP8251ytpXmBKl0oqn2Hmow
7ssNyMUjbTFTn3mbw4lmdzSsr3U/i6/iWgKCSaoU0eRz6DItGIZ+xaz7hgcqNIN+C5A0ly61romu
TRH9lVgOIcS531H/2SvICo0eNOjx/6b8ynSGeT6DGLvgWSm1CQLL+d0flnAKgCKWdrYmW2RTVQL6
AiuMn+tdbdE7tVqDs0WI/zkHMpaiQP0P/I8mZxkO8U68PWjKADj6riChTH7mC4fT0eX4nPuzDzxp
5ER9PqX+2fJY+tsJSLIuQS5Uz0aLYDWs5MBDag0Wbmp9oShN8snSSKRZw5QvWlGnyt41SWyW5FSM
6hRiuA245BCfkzCV2CMxM9v8OsKDG1HqGYVhNiWXxA105KGji+tc+AzgkqBlXe3kaTyVJBGBIcSS
U1JezcigbCpyWF+BMJ4m1OdbZgz74ra8b6wpl2f+zelmunBSwAB6egfbpfp7QsTCY/8eKrXwjzAO
uHnN6pO2VZS3l6dRVQ5TxxvTy5YoMRYGUh90bsSHoCttImWZbj0yDFc2epFXGF2Nv5cgIwyRZqMz
+O0H2r/Zx2sNnhs318Yg93IA6vqO8bcSf1I8QAevT3fkEwnbf3K3omc+uSh+lR3USOQMoOXRJSC0
z8nqV9qm5kaJgL0PawOinklF4Tmi9MGK/lU5vFUZ99/7aRIYovPVOXTwJUz/un6gEB4x9D2uLkEe
V4SHUkISc2TEHSSn8hlXu9ZSMH8eOoRgP4spsLr8UyC7p9nCA61NynPf5koUXL70LC3dlrZASPVE
u7aODHRQzIowf1NFqqCJcE+t4t7/QH2L/BtBmPpIji+Jpw/CkLY53FXO2mWNrorfL8bMvVc+FiTR
n8mmAVQA4+5AHIf5dCRMYopAXf4wvbOIBgnbwqgr/4C3slMASzq7aGzbTaEJBsDRyStz31QTqtAy
nftKr6bMnfSgWufxYwPjXuvUE0pOM86mOWuvEpcIY7myNcngFfP9YAjufNxup07BHI5ySvY8OQAh
XOngrPIs4uOe+CvAr8InbwGFFDnv3j9XhsswsrpqGOme4LX3ZZ7ZPBV0h6lPaWGabhkNZsUgEyNn
xeNAQsWnGrAR26eTdrun64IyKoJEcrjFqNaOP3pisvlRSZOEUCt4cnhqsuvjF3dnwXRBKLdpsQ2q
rqDc2bv6BopbpEC9dJy/gWNZYEs2lWP+MeH7hVRK3xbAQpkUsKd9ZWW/ygFyvpHqGHKpo7GnFu0S
q79/f+xVx6NPVtQ+XQEhWNjwASM2IfO+Bv4PfNFWHbTeOjJXiMvdvV3ehAaISToIOpoYIFSkFJdY
+jE3REuXlsDiXt+8t0WZFAKwmTMLFB2sbikdRFl1NTUBTg1Dw2Yhmj92mTu11k6DRyqAjQiTdCGu
Pk4EbOEfASOBohI7tFTfQSDCFVdxDe53RfctLtThre9M/aoYn4zHOn63T25CzYub74KY+L+9P3H3
ZMcKcTLXgk/L0avHfETAkwP9iJ+/O8RlB1uqrIfw9W99zI1Hefqvj6E0KuFpA2tuRIfIAzlibZrP
0tSmrOOPs2huIGN6yefSA0p3gji7G9CW6wxY7aYGpGKRTe/dWeitEkTmuoxmTXVUPYB9vT+7L/sp
LIvOi4CFZPb9g2dSIP9SI5aO9kPuoN4J25UMlhjlGgrHm3470buqXXF8PxcRQyhlTabYCVhwgzX8
bJH2rG8DMglcV5QqR+yVFIJdLe766CA3jKxu1PInORH39ogGp6/jAyLur837lBLSoC0EkhHE8WIz
VqU0BUEZRq9V/F1H/M4J9TgfLmgq9SwueYwF4T3QNTg04vPvz+xzajZgsIGVI5A17qeoQl4wdOSR
55qcQTSV3nVkFZy9OOuz5gXlWPBDsfjASTt2IFx0eQzsJQmAuZAWwz5sKcAWuR5oMMLScqywEqMi
epwYBzU3T6npSSDCodEe6wIiSlPc49Lv1AFMrAkBWOJ9C6Pnfv2tnJVaeXn8LcGT25ul6lMZBgcd
wPTkS4WXhBIlX5eyKI+uhP6/4G28xadZsVwv/UgoNVLyzTk9nAcvEdZZRZ0r2q1dtayx4gDpbWUE
06l0DHcwyLZmRj0K5uCh7DV7CniZw1CjDIXrlZu/XYOF4qG//CYYkZta/7f//8+uFpxtD+SUYTrX
MtKxjfSNf/T/jQv4ScrxogR/4K+gdgVBmLdxBjF6HFXbI2Vj9jsXR1QG/G4TCOs2l3GcqL6DjE3r
Vd5xiBcZRNvl7kZ1kmsmnJBfkdvhlQn/bmgHabxVFKx98UJDbQ7InHebinyNShLDmbh+T3RZd7lk
7ISXSsXP3AdXOQQUFTyXrt0H+dOsOLqhGkrbfvmxPKT8f0E4FdLklyzPAY601fh0bM6blaZIs8+j
voxnvg1jFhTY75TUa3dl/f8O6pxhxgW1kliNi21P/XXsCmP9Rz3Lmvze0i4UMmZsSgh4W2DvX/Kc
OmUvp2qz+fcJzu6dFbU5LMjTQjFEVKv2RopqevirZFeOxJEm0X9ECWzcf8TPzeDyOFGiN3S6d3qv
ZEnRd6gOcLGcyYUsRmQUP0cZaBmELqm7xTyGkuxlLYK0gd9wb4900N/FnjqAMNoGOmUjelFMCqbZ
OEWb/VOpTwSv+Y93BsbEV27OqVAFt2zIjBJ3j1XryjH6PdK9B/fQxAHDL9iQ1wZZCLdg8YPDkOLX
56JKoxRGa4M4CVgl506Uik26EysUHN3SKdmH/44N0ll2zd4r4J3S5nXIG1In45w+/1PuK/NQc6xY
q/qiYrgJFBF1BTEsFQmDnz0od28DEqd+JuXJe05hBGVKP/W8N6O9/1eYA08GNhB/o9s7ZaQzK9sp
k63V+pwqkTVU5LHYHx4zRfv3OJSdKMSfDZxCIbGTc2hY+Ny4j7KsA6iWlSlWo+dHb0jb2IoE9yr4
hXUBHSaUg1UjPVzHL7mIHnAwl5ckk31BdQATgjrpjoEJhUK2GrMbXwK/xvnfGFRJCED7O5PusPiM
69h4Zx6vj4QwLW3PA1fdH9Ocn8gBeJJhJr02xXLsMDDJ9KjAU+q213y++625B0BkPunpUIDcuEKy
eAemPIqcJ9I/q7kQS+lvN/7behsfXapY9WtAtz/K7M28T/pr56jEj1xCav99ALHrvPOYO5lXso+Z
dSUcBfZRytNvOvj4Ho2UFwOtjMP8NPvnul3gKAF3G4WDgxKG9KyAOYBkHVBcaYmZQA+Oc37E8QvH
Eo+wS1aUk69obiebTvWd2XZzgooW79oPYcFTqAkIylpN8vSBbpQF9k2yDi/as4QK1ihl/8E4VV+r
7YlPtRK5MbTRyJ8VGxRGrXNj1PLzlvMJLu4yIHsAEbIgc416AfQhHMgObBde1W8cN8up28+23aV5
C7NqEBdKQhIxF8Vdx1pbyZH4yrTXe9RBVTbJxsYywG25VMEPPkZNLC1C4sOTA7vcA68ssdmvpKYW
4vmSDPGVYnxg4HZqv7LjgUYB55oH80tfeeT9PsRfXvi4R9zP3w5BqopAph0FJ4SGDvySpocTl6oI
ksNWwkIHhUd94/SdUznSVEYqRijfjTcmI91t7z3Z8fgQKwqvfA5gB2cJDLHLRdIcgk8ZDowk95WD
aVhKDxG2yg6mWqD1M0ldwuDv/PLhKIBEj5bCkmIrik0QRzqNNu4B8/m5Y0MaonNA19yEAqjx32LV
kfJLtBhn5n5fpaJxU0+sNUeYGYfijxrcRPIGhNxGK1mxoIBvRf+3BwKTHcWgwIvQYIJ1aVjXCxf3
maBzumwGm6b9SICncW0UC30GvelM8mhXYcTny0MLUI+1cYg4+hmd4HZYjT8Ynx+MRVAU6Zm4JSTL
mJ/g3WgrtkqcQODZ+lXPrdVCJ2gsqQVaxXKodhaSp7SfR+8/QGDU4PuhfXUqS0mXIdyicb9z4vVm
X3hVHIu6s7tdvvbgKiHwsCd42v10YKapM8pmHEFDyPkqROrkqoiPdyaHfvvxxyvFeP1gZ3iOvuPV
RVWZhUMC1g1RQL6zdeK+nsUia+vMxPqODTJkEFFQZWY4SKSNZlSiBzZB7ABp5Rd7dRXwrVW6K2ZT
sv+olioLFfCAt4ciVyd++MCJAgIE0X9+5paMSuPPciQEzQInR2NTMBSa/vMJ/2dA2RSPx3xiYdlC
mbn6/H5mQqmO25h7A6OW8KeIk2NiAE2Vr2WwBx76iL8qgfOfqtRt9UoQYbghlLYRkWPAdtik5YXZ
F+8BtCeyeWthtj/6RZdzlE5yKaZiXUIsVCOHSdtgWytN2IdAZzyfNY4Wf51YhPEN9HNS39ktJbCJ
phCrpP9injb72H2nNVGo6nUw5JdIT2YQ8AewLP1UZZtYkz4XzU4i0LJhVHpHEJReTPffGBnjTPyH
Ih+DHYRUV6ClkBVTQw1eYNvyWXBdjAineJLZkjo8owbG9CJhs5tJA1VjB+aH8PbJzJL0eDz0tZuX
mdYerEHhd+wb9OfhNzZ4zkkQJT3x3uSUwcFpJQKmtTIJ6rhkNtzs9i9SiD6Q5L+9mg8tMVKyd1Jk
L/FDfHkM73ztDdHw/nldtg1RcYToJSxGCmqkhBQq4RK/zC7sE9zGFQT27bnZht5/aXggycWQHuv+
KSZmVmeOfaZsgsW9j8oHlhBnxPW7OMJnr4SQ/zrpvGjRkzGafVqY2Z5f33/Im+MAc5F0Hi/OXgBP
XW9uhl9IkEBvVZb/vqKQTyalZ6q8vXhDMENxOp2Etz8j9bZW540jU6LsdDKVmF+W/hRXKo4qf2Jm
YNuwm/c5R01M08Bd+8d/7nZb0VqQrYYVVLH5Z9yaWXk0TS9a13wPXJ/KblwipnP9Jyx+2fVM9Haf
NfItJqjJAR4MedUiY00hg0OEsyScLqXINFSEKPFPykzCO90cJdMKV0+Sd1LHK+fLilayc12uaFMR
rcskae5Tu53NggXvY25vMZ+oSGYtuUQJghiSNJeT/PVi2RQBuBYgT/aUnEwNPiH8AIzGRqfRnMIL
dp+Smaje8EyOj7tRAPMZ4ZmiH0Zvjv21qCCgtyiL3h4ZljioEILJ2dR/gHVcpU10JEVTBrCQQRle
lRR7SegqVvbioynjO4tEGb5ooLtzQt/3swCj9aQyFf3eQdrZLmnhVAC0bo5ZWGOXpNEXa66QfKXY
AZxhPhIvku0Zmm9CPZoVpOpsrNME2Vjr0IQymjVWU5999PW4LmLOO8VV+YF9tVDF3hr2actdLbCz
AVmsD3NaXRazY/TAT6x75TPNeE4UHLKRpKjb/29TZZ9ID4DCK7WzV+mcBxpVMeiKs4whLk7vZrIl
LWByPLvZX9nMyTUmC0Xykg1wSrJ1LESFwg36FAht2pyk3p4qBa864hKtmzY3lRT5jLoTRHQvRPjQ
TbC0DTotyq/HhjBIBToEvAzAchQAd2Mh4vPncIhROcVIphj4KNFwHFjZln1LBxARHOvH09+a3IEE
Kq/WbB1xKtzV6yrW97Md5AATF7w4RAt4XqORk6T9uE3HGCQyTUYYzCrFdNSSleOljjY3rmisogmK
2OCA6pQ4u1CKrr7SxDkwm1LlUGs/gBWvetBGaxOasrAhHSHcvNa2gpljUZb24tWu7s76TBjZxGvi
rivScXhCCvUP1JakqceDgM/OGn3NZwH4a2kodLFdBJ1HlJn+Tk1eNcUYlGxAdTviSf7SQ5LbwGdM
V0SxJywHZ9LsYVy4pBBtCN4n5Wmfap6s67WLhekTYIE2iCQvA4oe2kkYbeapy7IqoT7+rAY8voCJ
l0eDShKh1B8H+FubgJgCoFRXCTaGi0j+DiqeBwAGUkrQHkfD9V3MIBqpNaWgbz4ttooaXVup/tOf
gqOAQiziCFqlyXq8lKFCeUYjtCW34LZs9igwAh7lhmN11yLRLrYKNubfdt8cK+nMzSPwSIywygCa
TocdJZT4mmfDPdFq1fswstqgl4Ua30Fk+hSWZEwIqaNjRHP28W2UJg8Xs6/2g5Fw5ujpDVySemAv
E65WvRMBfpHk16CGuuWBXb0h8+P8JQvWpXxZLcIyiPFSnr22mEy/Jgl2Yww0Z/thL9iYBPHanA7V
3D5sldr3EfJluv/xIBOzB2DhMv/NlUwMWXVgRIWcGn0ZzE31dtfSgm44kJhpwA6ZDHlPAqFwzFTt
TfJa9Z7yCanas/1ePUU4HERQj5VoE38CSsTE8l1yF8J0bHn3jkA8KV12a9+6G6lTyEbQAQ6u7cuI
xYg7mpzwk4PDNhh6BOdjP4Lm45LhRuurZjjAlbOp9yxX4Q5bk0JdWnlardU0nspBoNXzhlovZeTT
DEfxXvccY1v/ZVb6s6ydVTsu0DlzmsuLkXUMPAEf/1ijjHQ0QKv+vubeO/703ToLKJTTkeqZpY5D
G9c0R0PsgDor0iPWF7vaoZBeepHbXqp34Jh5OvoUJPvf89hz2sYT3X4n2AukkwQdfRIlai/iD+2F
30pr2W+qG0VBSoFKOwM2wIaoiBCjn5H29FtVAC3CJfqZlQ7F65LdhkZ6vAyt9KAY+ETmg6Phbe3z
g+8DXF7Sfu4dmitwsvsnM85YPhRTzfoQHjaosSi+fsBggT9DvDiCV1ar7XRk8Cfxucn6ezXrEyP6
s+oo4bYiE2SBMNFo1rmJYtjNMqlWRuvGxLw4fp0Gjunk3vwqgYWY/Y2jvXaR9DSJL4tQJW6MvvUt
bD0+KRnAsh9qwOwcKNTp+nMDCLJM47XsDf6D3UWzDWA+hFZx8bcwlLS36BI8gYmQDYCuN/QarNSv
IE8/fnbr1AKH9p77vYHN8DYyXweE3USLf9T1tvV2wjy8x8TJpk18Jtc8cDTazgfKCuMKXoR2HzKL
auprmLr3KRtBeKe4AJSUbgcHh/RC51mjMOUDkDNUQhS4CSpmE/6FO3g9rwI0vPZDd6bn1Ef0ONcV
wv7GD20kVlwxCVY5UOk0rJtD+aacmUWqap3T7V751/Wn+K+NPX1RYnYfbkJTzwwS1EpOdRAMotl1
wWecF5HL+2Np9VbYIRPUtGD3+myEKUqKmWuXhs8eImMM/pvq2zm4HWU5IrZ5twvdqfZqWBzdzJNH
dJu7FMxAZ9gqw1y8oeyhjA14XWi8DYjOuiB8cGSA2+Ios7aQFJzS7KVTo4/InE5Lra/Q/DE7sXQu
zmtP0mGXDEUReSmWOEoI1f3L76ZQeGSu5BdoDThbcgAA5nDK6mLDZ8sTF4RpMIQ7PKVhEQHcvwsW
/Jju1NSukLM+uHveKu6C51u77cOshRE0y2mibKXWXVUItCu8FK+N8xBxmuxyi5kVvPh0g0qHQBt+
Q+aTHBx0C5aCtd9H1Sy0fZhgbQoRG+O1YYB+T7JDu2q2xeIz+Z0MWfBruXGYDbpv/vuYaRVTb0gw
oTddsUzuqclEA2mJ3aGNuwt+xgUT6TVAKDNmrIkgKLcLZCWImiWLe2gcOaII+tkxuHm+d963c81H
JHr4lxCAfjLk/wAGw1tRAGkxnCsEEKmreH/IkBFaW4j4Ck5Mhv/tj4bqp1ZMgW8tdtfjtkuUkVYw
Cuds5Kgw+Uwb0+PsUMsQ2PfOGtsY3Yqo/+astFkLer/EbSjZH30Y08JVzdrOhQr9ZvIIzg0fBN9l
/1jSoys/1ixwrEE49XDGMyt4UhOfAr1lmV3yJ9hOj8atDWkMm0SMOy4IBhPzmd2ZnY3C+M2j3qX9
rnZ2AThphLuP9MMeZ/ZYaqFdGCHTb9rVQjdlMiG/prgOG//0orCIpM/8ViMrjHwB0y7eYXOBEDW7
PgY+/XZVUowBXIGBZfpLdofMBKpev8IVC5wGFKCnXx9xPbvySUBi1Wv5TufOp/ZIhOYF9hgcrgXQ
1I9bOnzoY1pZ6fMOZuKZFREaj1C6SKonj8gSf6OIpgD7f8x1oPq2pYH6UuVkhJTahttfpvPi+GPt
iWJmD1UzXSuO9ZiZTEtJ+NNAkYWguZFPbo0tHmCQD3HMqw28luKelPOlgar407srXJTmNLFGSFMz
G2maeavq7bXjlrFCF3Cb67bGbdIyPRgCGMR/QAOG8S/Z8CBr7FPMTJsmnkap071xlrUwCusCd8Xg
ZiLrEXww3MOkuJFXCz+d/L4I+qr/VupwuypsWiSqNAdAX58aZnstUdZWPUpJkn26jNH+F21Y5UnE
T3zoVPU/tyU/1roNe2En2HNK0eRIm+/6HA3jHk+FFBXsxbOcyecdjFu3q70wWgcZOIIUiZMUqeOB
BiE8vkR62mA2fmWNadF8Z307flZDGIx11YyIOZdxxMOWuNqsvQmUraU/8J9RoTYo5ccWeI2rTox3
S5kdxwrQ8r//ie/cEqbszTN8l4fk7zx+3vsXr91B80wouyb+4O1IozvQmII5UQv26gUs+qXRyDi8
/100BBIWXS0np/zACsgrZULwiIgVDRQ4Be999GtDH9eqY3OoOqPtc9Aprh3MDK7h4iuFQkYsi+u6
2WhihcIZbafcUYyl8Ik2G6RQkzvneIZSLmneidUrAPRCXSsonXVn21Mt2dovxvQahP1yiY4bXU/P
9M8/+8j1+C6HaWBKVTa1bLlrXilUzlJ5+NCZ/08VYmW3Ej+vCtgcgYw+GiO+0g4MibjssCPyNJVD
xJ+iIP2q+kzLXV5lD/+VTRG4BBdBOYJhZEziG+Stufsc3nQ+LmZD308GFbwcW3eJgKwYW9Fmvsyp
wBtVbnh9ZA6dB8W2uM5aEKFAkqZAlgQx0hTlGLKredbJOOsyWE94BX0HqmVluC1XMnGNtqwpIKf1
SZThClZOvpQW/DUq/nTNUavxc3+nZQBbEMgwcMTePFI3tu/yvEbzPNYbwt8uY+K/BLyvMnSBdDbr
n+vqp2dmC6ZBr5gRkk4tiDKcvSrw/MjkQzKgyIW3l/bWU3SalGhR0U2nNtBkfcWfKX0wTdvnACjc
ws0Z/SdeJGqtA2tTzE42gSFeo8Y+rW1oObTznHWbcyVffAg0NAHpTD7S6rEb+hmZvCGgCZtDGRYE
twJ5JGC7xZ7PS9l1ImnGZ5xrtlidlKNRmAF77NjaAaZbTUVDmbfsk2hokn7dyGNl+siBoNiOkXKk
XUqxNPj/eDsmSWIQDq0FFYBwSq65vnKyI1VI7aJCH0XPbGLHEynA1sBl74v5iurWzouCC0hJBmQo
3sNlsfaJ6a87Z7GFefMtn57GHqQ4npUdQ5AnmlQ8SpqNmQU8ayxJR2WeoXwk8K0v8qg2ZrO4tz3t
3cpS1x3LoCCUzjgp/alj5hlxHIt0L9y+C3EJxfka8SYuublSfvppUejE+OL1BSR4tcSloLttiLs+
gjVYqLthZGrTi257fTsaWvSpX7PjI2X5c83o8mNil4LszLPsGQpzIaRht7zT+sRBS0YS5/jc7gk4
uuRKIGNhQz/EKPSlIVZpeJf/0Nfpp/AT6nnKET1g9fqSoTnhcLQ0DrZ6eDI1eqgjHvM0jHh/riut
2FLySft9aZxnP347o9MGKlhidHoYmlOJw5ColC+SAfD/uU66+v2lP3zFPXf4dig5MNsNgXhgPoYb
xqZV+kUAmo8rzcfD1muD/W7ICSxbxmBldbEbNeiLXa4sACZIDjfD50xERnhCLw99z2U1VzeeB4Q2
FSl7cnGtROh9NwigJC5ApF8VozGLRFIFgUMzhZW5qOb/n1a52KGzMIuami4f8NY+ts100UoRx8ms
Xe+vfm3NeHY4dTb2WJKHjwaTKsqUvhDWqxQ/Nv4vU/K1aivLSXgMGP5EHUhnPWzVEFF6q8PfrKyZ
YxQWwVk6pTfjbpbcXOclsFjRETx6dWuskqrXhsJOLAqPQUqkp/WR8PdJ/+W4xeM+LG+1b0V8cfbf
c0H50hbTKoboW3W9QuGUvU7KO9ptBMBPeJ4R7HVCpA0Xdrl0E+GNM43699AXkVgdUATvWKagi2Vt
MEo/MhEg4VBumC5jhMZ3i1ksBQ5GXoVmpXONNaLZV+Brt/xUqKyXNcgNQOhOI6ypgcYrwtcSKEim
u+igElovee/P0x+/R+LDH8Iuxepcr2czhAVNgGPsIGJNzMtPbpC1RDA6g+spdlcDbpQZCRR+FfOB
2jRud3dIGfmmnBzh7bmBaGZqB/FJoLAThtb+5B6cohF5t5+eLfwsMHK/MtvrypbW2FyxDXFzWgGr
LbVlI1aE7IOYeAyQM011b23gUba3b8CusR8NaI/Cx0XHdAUR7/cdeftbn7vf0iT89CsLWUL/L3Wg
LuBFZXAL2TvI301G5BUNlAZJQ7uNqw+bY2nDW5/d3d5iNRqs+N0sruN8uHJ1QfIraw3kixQEZ1qg
0dDhZT0xx9Ma7k4j5UpD4o0uuQYPaj/9NLY75ZeKI9ogHNKrL+9Ps0K2qKPmTxdoCNlqEE1UzMHd
V3yggL1SRNrQhqhBl2bslm+LbL9N0vdJI/7quMkVE1NyzdBEfVI3WGPqiec2EyGRsoVT+iyeaEWi
0+RNKMicsG0w4dpk3L2WbFOePE6Z3Bpg5f0PW1esyDbdU12Bm5ei/XdqMRsP/pk2jFyOEO5IwWTj
nJ/yw2ZRIg3FrInh+SeuyMrB3o368EfOvCfAmhM3QdtF5xZT2veeYZ7jVw02NhhW2JNQ8dpSEQ2Y
2OCPjb36YKvhjVE6HmarleIcKwNqUOao6wmotPervlscEEZtcBsT1v2CL4oyyl2LGQwpWG3+fdn/
5jhKj0oJC9f/HmgINS2WOrJbkgKN68zWVOBNjp6H1195oDhuGGL+eHiIXMaTTRXk3zQ1nswwr37a
HX50RlmZ/+IlEP6A61zKFWuMB7C+mwbrHZTqn6x4lLuNxIHPROBKQrzLFylNs9Y76tQ2qjKFi12y
VljaIfYy4vlYm8YH4ACO9kK0/ZtSC3dgMvNc1xmStoEMGXAR8tzrux9fhLbktcFyCVcHCIITIk8+
MmcXznyBhjcCO4f28wbdP66fRB9MQ0ch2e0amy3iiQgj0TcxKAifrVVt9Jzll0lTYqu1wU5/qT2u
UVsTkny5egXlJVQq/Fpo9BrNVlxoa8a+eoS+SV1lwVSyDc49GPzB72y6zOq9Ji2h7tD/2VymCh00
q3dwgmjH7CtUDNgR+iL/oQwgAMtcDVgCWTs/0vyPJPiOTq0Hkz3yoY8WY9YAxDvjmLk5n3GelnSK
1PqjIe7La9qZg2g7Wqy+KIr42+LCFkXHaILPnt8Qq/c/W3T24FF3RyXTTkqYhYF/ktgJLPjnVGlY
dte599FETkGUxXaHi93LdbkgWvl9q918zWJVXT6DYQ8XwkDI+fit/BgjobfPRfJajy9YIsp0LvTZ
12WiwRfHhj0XxiZUl3FrMFd5nEXoXlxsXR7rrob8zdKMpHBNohXMPijkDyggj5BB1itU7c8BV62u
TS6QH667tPu6JdLyvUjLStGWqqjyIfFemQ4taWDFk/4aBcuVXefx04K6jwmYsdT+sXJE4w2ccifH
zAY1saN1LdKCjHvHhQbcsnfa0gZ1AV0/idzjQqIU7nQGRNjdheRtIE02qtO/MgzsMVqj3sM/7c6D
mrIUF7xP81ohmJBG9N6Cz+gJ3lgNr4Nd93TBfoZakMK+QtKGexVPC9o3Hl1Kfsp1J3tOadR3QPd3
GDaAVKuLqApduh/pw8b10Hx9kRZLEFy7O3LMet/voOzOHQAiSOhKFGYjsJqJL4MtF9sf5UlOzuqv
TmDZwFF+p+nqrHjo/8+iCDjJr+LNIIPrYttfDSe9QltkyRPwrLjYijlqzD47ySGu5pqfGF7kSZ98
2zlF88dzfAoYzahbqoqfMyLnn2bt+uncHyAeGv5WGXkwV3ll4FQMUfZgUZg6E2qlDjiUiec/6dbD
J/Ie6H88XBv1AwrVCwcwJ2orR+AoikSuQHks0Z6YzhzrTy27RLJW7/yDdqTLh1cEeVwEpeyoXGUS
PrJEimeB5in3kZ+PeL6KsNUP4GlxGNWC7fDmFn4EFkPWqUN/1VanW3Mto12dPjbBwjRoy2uuiM5n
yWe8C9vZRzBDROxzDNsQgqYcVIkKgXU3moMCDXIvDNb/m4RTOr4IOQ44bR3o3a4ZH63kL2v5VuIq
xnRHZtEYYEorBkBfPHgxCJ6h9Z/tDhfzt8KsnnNj2WQENRSaLmFJFzbJQnCvUihTujasH/kCFnH/
2R703+KXHqSUcAmSaaoUC/6Sm50PIkZJOHIAjpNxRQiN2a0rBdaU3/9p9vpGm5xlF4cBH6EKks4N
SAKrcEIDapxeugr4xTaJ4llYGcc2L/9FV1DhevJ9Ya7oTFV+AWYlzJ+01a8t8h/cQR10d4mfcm+J
ly8mc3K8bxHkBlDyNdmEhclJ+XdqcuKUSh/zB5Igp5/KW0hz6lByfLnStxD3CF+1V3E2j4rHGE6y
CsQtg8etBCW6hPL3CvwN+6LaxHv6kI3x0/ERq4KZKVHwt2WvSV9Spgg+fRT2aO+MoH8yuM9jt08L
o1NyLcIL9nt0JOB85IHbexaFvCsjw0FGbMbuHZtpA1rgrlQy07OPoAtOMgUHcu0QVAiLf9xmGQPQ
Jx8EJuljMxaty6qKXS8c+TsrMGbwBpLS/kdV52IQ2vVAJpbXmHnbzhCErg9ZW9Q14oZCNNkvxtxi
ZUTXAqPaS4ysHkMek6vE9A2FmY/EUBetjAbuNzJ2arcgF+GeGQZnUK0L9wJbRMaIm4oOJOpH0MPV
5YbEzr1wrhD+ovgplCvhRDp3o7FV9kv8r33hujLXMw+jfOGaYjEKFwn6YUXydcdrqa7fOLa7kbk7
vY3RAZ6ry/zYeK8UvboMHLN3DgRggR9LV2VrvhxlXQrRYL6BHHY17dDcCmU2Xrvi4jmB31ieExL+
T/j+oOO7o52FpORnhpXOzrpyC+YWp/5N0WJgnxsFZQSy2UOJFwkmGB1ry8BQTJZoqDKMI8hxVkLQ
kif62pmSGLPrhr31x8GzDp5SUR5Cho8ribiuZs26Mt9VizAFs9qm/jILD9PmFK7HX3TZjegreuvE
rbhqIKGxaRfBflBww1843mNRlOPStLFR6mqMGjJE59jSU6aRVxz6LClth/taDMgiOfpfeGPLOXfW
D8CE5E0i3lLJljKddrde2g7e6s/SUhzfeNy9vGHt4QXwwNqTqNd1HMa8cHm0DJ1HRQCELZT75GAS
VfVbyiD9dQoKpMKJ0+j06Yh/dhc8ODTb341ZjmFf10Vs4Lsku9a5m9QbW3s7ehCVd5642M0RgT6O
79Xh7I4AS6rylY1Rg+COAglLN4yBoZkJQRdSMOz+GW9QOHfN0lnIAS4zaq/sXSbs0ZLG6iR7Y1/l
jVQeHJn7xh8W8k7k4ApWqJ4hMxAjvwy/uo0NvjhSwlq3elVgV894OB3nbNJysXybLcxjyy0zSSki
fihDISKV77GMggP24aR7QazaA17hVffVyNJB6TueW47DzwLV9XRRYMKQTUceIZ3riHdYrrzJIFGZ
mtYMTfDTbq7YU2STP9iDroxP3ZXNEQG3NSSig9Z38tZYjrkIqUBkAVJYqMPF78CJr+cZEmF8ps60
dKTe/inxUNul5mJU4w0Q1/VIfDeBiw2px2G9irX9SS8eZJER9NmZgeQfsEhmlywHJ3PuBpy+0TAM
HsC/X33mKqTV4d/dtzk3o3eV7ZbBeAJKh+o6SqcHqwYviNb+zDhIzmUq44TaCpB/dke2OFxfMbUH
awKXyYy7N/A3Nqo0lIiO0KM7KNLxslmZA8qUZIPqATn819GiW6vL1I2rt3WSluV887O9nalf8khK
OmEHPzKNYzzcGjN0x5or17L71uzWVAUoi8MUyC7jVk8hQBh4suvXZDUn2X9DB/ZM7PdsSXWEhwY+
6j7EyIwWLvbAUEcHcPIofiH8GFTkXhQ9gOFlPBbBPpioZ4pza0g8Bq58Ma0j9b0ToKRNJcvSLrz3
5sfGY030s8ANuF4UwxFhV8lP6G2AX2IaOlDRBdwJ4i8o6I67FK6xThBisE0/ZClA2W4l4CfRcWo3
hZnLXFHzxv0FcW7keKQeZMya0Iq6UTSahYGenFDFIwSKsSz11TRhBeAcjaodQ+d3oIidfVMVLX9I
1h1CJ9iJa7vlgiJ/6nc5hA6nbmzWliVAiNBFvehPy0MP0Dzenr97W3hO2n79Ra0LLYWAuQexEgA1
dOQYAe/HwHXWOAsyWAAy6pubtRNK2sZMi+m6qTY6b4UO4lXBKjndWm6ou4ej8NSFN/cU4jahHynT
iasx1F2Zz/yeYiFc9CQ1TU5tvNicP/XcT/zQRX4RFoC3opKzXAc91jSEAcPtLLMJH+Cee8RGWnTB
RFNN8uGWz8PXDzV5KQXyX9USaAilr8Hixo9xMLS2a/2+UdNjFqjKJVm0cGdVFgGZdhWdzovnMNJK
ZLJd/X6/EQYe9u4baHUNqnzBj7rVF7lumuzuWaCWJGhZrqnJotrfaOZLG5kvFHl5EtfSFx/V1W9F
gYEIzAYlLLWUaDmJJRR6fUoqOeQ75qqKhLjkRXkqH/tYWGWgUw27BA4zxtmPIXEC8hd3bENLDlYE
vaAbUaTo+Qe7qFIfWcHff3RW/0AjCUrwg01Z+SgrJ7LlYSt1+OOaDMqHnE57NO65xozTBcvgWqWC
A0YdNdXDRi3NvTQ0iCin+YBbjkawwn/6g8huvG83DgxxaWn4/Wqqj5VyBNtmp2LY8pT4hKf8CL/B
3mmX/NSywsfWbrsD7yQnA/8OcfJa02qskf+0ZkYyfhg3pLI88togqNEEJMZGWYX7n4jXYXPbZswM
2fQM2Z34JNtByW84pdQhofqorz3yMC2IBb3RqJ9RDcbMsx0Z+p+Xqj1dCKOXiZUM47v6wK8ETjtU
lhs25DG0syU1PjZOqcO+A57pVeW+J/bEyv9J52EC33zK8kuY+KRj6imthXsQKJWDAdUnDYUFjUeC
QHj/fjOBMJ8PEoFtrF1VFcrv7zOPPBiRlU+Pf2FIeGDt8/fCDa/lZqUsbOo858b3J2mb6xESkaGS
areBtkOESU6Yg7cyOCl6zXaZ6a1So5FJ4KsvsA6wPQH60NJUcWxyvlaskYBu6OS4VdXmas8fonSY
2CWNrHWJ/wEUbf33NFbV9GMtFgBgLbnNLKh24i/6cMZ9CUAwG/SupVJdMZjZZH7e+vpwX/MxGMvD
kfDL9tbVhyPPw03Y44ObkhL8fTYBT9nK2gFMZv/0PdFWKcd1YezFKK44NFASvcCSdLtd5sitK1nj
1bB44NnvlNERZHOsN5dKE1EN/5i4sZXaU1TzJlhwxhOoGX1sUc2SVB8H8eYb2wo3KualNso6xZRf
PIeAIBsPpixhPZQEvvhd5YkvoDMe7P1pHF0HDT8IOuqzFtjhwUcmBmCG/gGNtAI/KcyZ8odNjfHW
hZxCb512ytRtELHZMe/DQb0Hxcpjzub2g58RxZmSajR8X8PWyAWKP6SDv3jBzf/iQxGBLvIG2VcC
nXZpj3Uo/+j7jXLvjqvE/5y88snPnb3oXufAmQWsEmLr37WeQDUCT7WI3T19YiXN2xuyAHxoa3S3
O/O7gQmD5gF9ZqK4WhUEeLQ3cNeTolIrZsJyN5fyguyam32p7J82a/b6r3JeG7tFojWUkycZmGg5
CDzbTsrFo+jwugS/OIAh/XTXZnMUUSiqOJBXWKOFCsArRrh9RYMOZuO1Lms4CC44qy8MtkextR7S
7jsH6DarCDT/T+CVmCWLH54QS7WeGIQZBweqNlt0gk1N8CZ0cg7KV1giGEf4KNO1FZe82LbaeONJ
wd+knQsAwQvWItoc18QHdVkSAkHyxHoNVwI+J7XM0zDhpX1YJ7kpu+IIrhOeSvcix3HvlusEkGza
dMzsW1z1xCe2K2NU9Yrp7jIXrud4KQFv4OTWFQDMVoVK1esbDuxe5DcsEmu5vp9zLbn8umWbvXoz
7fzpG2C7ob+6SNroSpSMgTuURk7vJx8U6JKamU/zll9xf/tCtP6aTmhuXDbS6sjGG67pZrhm73hZ
34b9KCSySkI6sp4jm2hi1EHrAFH+vAWyIzDFq0waJv9Kb+OcdxJX4fuZoOB5vmCHxj0DiqA0yAwb
982wh7X/tMyIhp39ne7WX1g+TxrLGj+99u7/JGnPtijmMtjP7JNSi78lbIuWhmb+VJWnQX4meuFa
miiBvpXEzXb69b6Cmuf/St/c7J2KzSgYvfCq5yFUFrkkZTso0b4n3qF+RAd8jgvkDJ+mggllLLoM
7B7bN9ZwheVzwwgXiY1Ysbx0l3weAls3RAhOYMna2HUCbClYR2y0gsBjgkicn2TxjD1mpF6af7LN
VpPCSAzSd+xi+n0TEx3Bltk1HfF9yap9MCVl5TMGxXWYwvElRda0bfPax485xTHWVIt6Au6aytH3
llpc1NhPX+pZToUaCFy5DejrNhT2v1kL2ByDpmFztOZZqwoPWz7UUaS35o3yfwCF9lOmp12ieW7U
epy43iKtB8uO1OJ3sloifGCFxGK7VyqrEu9j3V+Pw9LFa20MPcS7w3noMi2mV8xYENqfB3buPjVe
oD2sJRRUqcQCJiu8mxST/UaHqcgkuPuT/ZfCiyZrLEP0UYbj3Q40Z+9HpBYtECwyWz6U1qOO0ah5
mM2HqZBDu15/9wKNh3UTmW66cghMMuf5H/dm709IBiKPhkNHwtsKLekmlsZKAs1GOWPWKsPmIN6m
MIbZZ18JKmZDMqZqVoiokvpn6KG6E1WWyS9v21UxpcTjbncotZb6zExRZ1yKXuxn3qVQLXdTsPxe
i5OmtvyIKFqpmMxJuu1s+jKxpUioEVTdjkGG+f8/c6lK6/1gfWm1bjzc6CdyKupFPfb6mF0IONqm
ExaxT+BuldJP2+BE20Epc+pMogOlxkuH4UlyQkDd+Wi20QUsNLwZ/9JoQ8vEH/UdeKx34orIQ3k3
ODGM8PGPyfubYPB/K6t2mELRPalfSvebLcE4zRoRRu2Vc99aqaogBhOppc2ObgxGPP5+EPefNvqU
ydDvtoMzXoH9sAOcmOeQbWFx4J03UkSSPBQ/xGcaLFx8i0uMa05YRIdAySFTG4LEusQbYxKjsU/H
BsvE7Qv4vN0+jy1dc1o+JkLUVg0OI2GY0pL104rrkzeK0TPCzQ1C01xJZhPTLzDdtEB6bu/1ss5L
7UI2uPF7gMXpf87wfWqtdrwQ8q8hwm2JfqcwLPM1HC9lYX0Do1eio4LQ0MYLOuJK1lTbz2gyP0Ut
MceG2zCo9b50YsZRhhFSKToTh53mowZyAzpkUTGVvALhQvZtp4VC8qA6UPdmQRC6IO6XuSJm9a1q
9s1GWpeDpmXMIvL8stswbgCXWpx9UoFWAlnF8/IPsMVPWyljpzqWffDbwH+PqQ3mF6pLxM3ul2Bh
gctUEMe0ezvQfDq6tkM6A1Kw+OykpnOTmR7CeVVMmjl17Vyg3s4qHBlwsWwvP8RL15A42i+2JzdG
VaiLcKMtLETjiDdKl7b5ML15iNpIahWqV//tSYPpNs2p0ekPa42rbBgSJvO2Vtl/D6yeYLb4tVC2
CY/1XQAYnyDOjMWW0HVY4SKMg75cVZNFkZeWtMLRtMtTc2ztf+FoMjRN53jNKyqpzvDRqal4Zn0g
L2zvH2qUnW9ojpTrUG0jlMTGvjj9l3EvtMvK+aGT+UjnW2ASlZY6ZuaVJu9IY637IS81z+qNgQal
bMhzwiXqoph6xVa8cGrJoIW+hCgnDhLDDwddflHzfATobHzMOtfF1KwLLklhUbq9sbaAMxeXbzYE
l6I/WAoi70oiHp7xAMlH3PsxtgWy/871hnPDVNlvqruhwmQEkdsHtFZWCJVJE5frm/ZXep/aGRF7
OdeCbADDPIcpKLsuKXqYWWenHT7/H/eIV9m0qraDbwnYzmDltwXSjq3kh3SxBnqokdkDnrK8TIxE
vpDBGJXYU2N1uNN8xQ3ew1Zlut7T9OehmOy9N9Dn3SjtKDiFBbXVq/2bnY2uSaFWYmq7+wL76VFJ
f0piQ+UjAz32ZjeUhOchmgTck0qr6OYtrKE34mbBO0NqSRMMHQs8OmbpGKbLRgXllkf6eHQiicmK
0QC2WbctjjHtUWLF8Z6ZCnZCRhVpJ+tx4kEVyYTzPRFOhVwQ4n3Qvd67kKrfRLgn3omr8ujkrsPG
+/ppKOVREL58ZUyo5z6azi0kwyKX2Pad1sinh6GQTytKzki8neFGpw1aNqrwz9nuQRQfEreF2wao
8Sm7LHiRnAmZYc6K3i/Ttyi/wawVA3HbUg+297JWdLkOoUedDdsw/mw5U1GEdJjkqZsO/yuaWVy7
dfSeQxHFeFPok/sVcZ5gFJeYXDeiPG8VIc+mS8qKDEJTlJ7G7dfIHLMi/VzTsb7sXfwgTns8CWXc
VGn4bRWqaVrGrYDgB1ADzXFETBYOQMgOLy288//E1ni7hI2Xrim5Lj+LBCk6u0VeQa+QRYXnlBW3
iFdKBfOWgQ+twHOoyTTHxCNHBYuzVghZJsnD2sGAOq49i3vXO4d9EPPl+iNWX2X1XlzbIlnWb+D+
GeV8JRyD2AYDkfFfC7a6OspiL6h/vHOYq8kRdJNhpevyQC3PAv//b7/1q60/dkRsZ3d/7GXyH+XU
SDNKha2c24qfxMD4PA5os7Ed/kbqXxGdq8/dboQmteK9Nvag57aAYwPmPSEcKm14lZ6YdFLTZE6l
4r26nCgA5grCGcfHKqs1owVGB3MYelSI0kSlGkx8kcYgNcBu+4CYoKqrS4j6wMBexcCusmHUd1u5
5g9TdwvNKJnVuUzXx5S3Xn964LpTKV0KCr1W7vlMBQ8nZ2037CGbu/IbC+2wFKkcS9Ba+dneo5O8
hBysFNjQX1QF1AB+S68IEqPuVpqV4dkhZHSft6kXq32+NrHARlcU9ZAfSgHiTm+7E6weX2ujU8h4
h7NFnvju5outu7N/RFac8Sz5mSgXAC6vBeqAmXPyGpT5IBJIOK/TRqtAPv0EzF9f0C/F5U2z1ido
AToRDxxUTXWPWJMyff2B0aaTzF6aNfGFRglsEcbPyiYLFYpXsf+3n5JyOp/ACznWiRqk375aukZC
KDln6cnRxGAeFvP0jW6M6oKihqQV1Ls8RdPXAxGykEyG+wbrf0jJaFPqu/hzH7bjUmdtPezmEslm
K/wY0uY007PF4U1dx8OZ+0VDwSekWl6BT2SKQJc6e722EJzKqe8/i8gltUiHKCa/MVqiUeB4ZzFs
1h0n4ZU2v6KulySvRhqqcBncvyIllHWzrfZ7uvwuZz2hcXDfRw/awAa6E8Bzzf/9JZGyfHaF9Mpw
W2TjfeQuhPRqcxhP3qUigwpZTqLrBBznIrkK9hAOIXw5VHDSlJM1SEVakx7e5yC7slGJm5h8NF8F
eE4TgwLFPBunmIScI045PhX5SF66u2bAAGHK/a9lT6fmxDXeoaMNyaRpJpUi6lQcaVZfPywqr9/a
7kpH+d4s2krv4ZK7JHW+wPARI0tYXrhhVupCH1uROz3zrInPs17p7GopKbKICF6PGmE/E2YOSaIU
mbtm9fqwlclbOFNLwa8qeinxuXULUOvKq27th6xkS1HqYBSRnl1/5Ag12qI6WqPxTB0/ajHB8Y69
l8cmljY4xyTY/abLeVXqm6oJ8JhBDZhfZinUNKa5B+4l0nPjJySRU5kZsz3T/hjDxyPIckJ80Zsx
AAugsNh9Iciy252aXGls938qT9HaatZC6jjcnIunTg3mbvrcwqFXDN3kPWD0+Z0nZnf9dAM2Q8Rc
5t3cU+70ZhNLhjwO9h3HMdueQ7iZGcKXWT7v4X/2znUBPEG0wCX1gYAFAkmreBZP4NM6BfXa77wE
BS1/xkCP9XO4OvRq8DM297Xc5sq1qBS3sydRh2LMRycSrP0MTcGdRhVHjVugJvNFMoeQxCbXMAtS
iZc85/0TQ8PXute4degnJOrBmvhDzCoujQ7ZzmBy79ixf2UI/e27wx6v3WSK/YGOlxH2rJjbY7Ej
Mvry5TY62yYKSI3MDF9LV9H/Q9T7IyHu6mgHlTH/wodXwLSfruYxi7vyAQf9LmiJPk9L9+LXW/91
o087fRRP+18Azox6oZoiQzjMEKf9T0yQS4/zFt6K4reUoZco1FzOziPOfm2gof0VvEMaz3y+H0jZ
4MQCTAtux5j86Fcqy37fmc8F28PSbMYveBGU99BhQmqyH4QuWJPflC64HYUv1E5BkRbIUFVUGvLc
jIsHvYyzLeRT1YfSJdgd0u8gKqyswA1bAV+uvrazjtBiG9dtMZ2qv+k67DRMCzag08d/9uHb0rcY
y2hJTOlLsEJiU/ZiZ5dejBxbPZjY5Kit0EcNgFiTLcvw9mrHVjEfCO91x1pKBlOxs1C6+YRGWl1l
kk+Zj6llreKkNc3gyoGzTezFKiD6hRhb4v2BmyKzUGBc/FfblDY1ATCzLgh5NkcN1xAFUCI6kX8O
vqMDk3Y18JzUkLVFTddkb6c70PI4830Dk437Lhj0cXt8aubnQkYXOI/ZKep2S8LremMVXkZKS5Xh
eidRvHHaBH5PVqO4rF/mF/L0Fi4YlkCPKmtcqWgxcj11jr9UHOgFOe1OWxJThyUFDnaLEB/nAH+P
eZtjWu9dNIv/u+EYhjyLogm3RZV+1ogZrkpZvbJh2/uiyrr+aEUDm5phuyVtZU7Co7cOwVryMxvd
shCaLs7/Ayli9RNq7We9mwSxtucfpIuyK/31OzmXOtSk41xOGD3TlAusEPrnPq2hWMGxvEmfWjMt
AyRVqxarjFfbcXOZVSlvwHhSloGwmDQdkqavsHuXqM4etoqIPJ9TznOKxdHgKpzQbcYnob28F8vm
IZmVFAMcI+s7oA3o8KLvsY2EOsLdu2Z1+IpXHmn7w3XFNrCtTdY832gtEdAT+9XtxDch0oVXzORf
llrugY65Li8usJ/xjJRUGv2MPgNNGeO0lhFEsiH/NEu/uTV+onxG30u+qOGWYjMlRFvVdWVIHQEv
msKVhQAsGI7yrQarnOAwUzRLZ8YihdQL/v8GXBBTjOi9E625JHp4hqS5JNY4SFDDMPoBFH+qQMCY
ylW5Q4BgypYzvcj3f8g5Qgln9oOqxjBm7phL0aEnEPAT0UpOnzjTNRyhmfdTbSZq3Q+FkvW+jUVB
3LbwBBaVkgtY8c5ab6nM97S3E4TQO5JzCfpu+CzIkc4gn/Vp6fKyz9eEGhuBvLbegMR05H4YeV9C
ce7jMQCzBU70RnvDrpodf6dueP+pR8EFtd0aKK47rqcc15TWBPgf4XevZyFfuvPTXxRRTzBTrJRQ
wVIgUTBQqSqQHXfbRr3A9mBaXVwbdwtzIjAu37nD0e8u3QSRDIkqnmS1TyHbkzYfvZTr43R1dWOB
4+xo8yJGi0CYq618aCZC3XsrD56orfH+piI+DVFGWnVxmKJpke0uCgWTD5llyo+2MsA2b/QI3SoP
29BMtSoxuvR8mUXExD8iyf/51mEsC+UbEpjAgitI1aBbRodoSWHXkaWzhOEMA9x2giGVP2jb55IO
1Nn4qgeIy3AytwH9tJCpz0uoV5g+DOShrv5ZaieLBTGr5RjocLsFUKX6e4iYcWURf46k6iTanWow
1+w3PgH3H+tjYWlS93gCGX6zCGw2fImW6RWeNbMd8FuS62fXleoHtJAAXfHzSTlRLx4z0CPkcpMh
VwbXx7fWyhaQzw1gjSVccJZGqmDtc0HOU3z8ilFD16D2mht0GZHkl8LbETyO7+F314IhFv0Zy20w
m7z+4KxWHnrsxFfGCcR73eERh1q0f02BMQPga1gfqA1mgB322gbOpIOupCX4jCzaBwHh2gxLutMi
IiYhFSCCO1iJUMbGsmkSe3iJFUihasKhfEwmnh8Fp0zdjGL/DJDfYutKySt8pwcSOoVQ8D7eHVD7
zhuIUsAebCsayQkMiZJaFBxn3OtQiikqeP+MF+9blnL35MV3O7XaA6d2xaGmNsCwUoCRgvVycAyv
FPH2v2lho3tewc0hXppYLIBHOwr49uwcFhB/BtBmYwaUcySBwZGLKEPrPz5h/MMX+kKwi/Dr4KzL
LSDF3CbNGCP4DrCF8tDX73lm7OQDLrYC7XGGHxthY3Apifa7ceeXG4wr2OgdgDKn+yFxUG8taiHy
QjC2LB0ZtGri+pirnNR/gQT1Oq++KhHVov5XPtAdzbzS+prSxAMgEl8aOVSchcxXRJKuadINlmur
3OGisHugMCAK+/c6KXOvrsNW+qY5GHeAlNWVBOM/cTIlCLDmi75mNDA4MIwtSzuQWOyc/0Ni7wzq
DtNv3F14d82UEfmhYYHqQXl2M43WduOHPfoCOdHfhWK74x94pMbMGB3E0MPbvYgC32VGwsTdzvyg
PwOMPx47D6kVBl0e+X8WZnQ8otjIAv4CmCUtO+0HLrLMCrge0UZnPkkEfa+gN5mqUcuZxYY5bg8B
RNJntytW4bH+3BsRdWRSYPvL5ePxP1xzg71eNoApY8UwNqER8xtgbGrPdV8zchp/RGYl+bqVWZY2
OSrvOBSXd30Np6vPSUOjS4wxc96tH6Ahxu94ov+kEulULYc2qWWZKP2w/ZTfEtDRlNKUHjOnx7IN
9j/eaoVnVN/mWldHVTk/EMCYoE9fYArMOX6IEeap7QX4D7Ejt7k5AsJIlZiNXjN1Ea9LEXyTSjL1
0AdGh2Bzqdh84hGWzOfEi/vcg1eOnk5BjV8ZZwrEtDw93JUh6E1gdBAncCxbS/kxvp5vVU3bxBxo
w6yqr3IKCqNQvIWeG6CF61iOkedZsrELy9o2EvBEyiEo0GU3wkCdgMiGCFSf+Na6/e17jQu2B5CS
Vy0NME2xKYyTY4f8ll1URD4g0ea69K0GKXF5PuBrKNZjZ67S2KV68NfuHmsD/ngH1XzlQATxYf8a
fDpwxr5r1XqorpSuNQ5PqWqFPftH4OZMi++GpWNDHDD9BK71QcE2d/blhAlJQSWCUL649WTcc1o0
zh/GOv890KDN1OGFK/wnoYFfoCCLspn7V0reMDh4fTTEIODqqiFH91HoN6qYy9r3OK1o6ZTtprlG
HbwQlNhIPggz5RgGOoJ+tpoyku2HVwBzSTHhaBICnBmW9jggXvPIsJaucS1WLQvFoyO0i7jNAOYh
KQAeDxjasKuu9/zqTOCYlzMx9znYkl8IZTs1rB4MPmM8noMaJCAPCOiK/ptHLBHznLEnEwrq2sFw
SvGHFa4HZNNKkak7MlWtjPRbDttwf+o8UKNA6SeVqhr2VAOV1YlQXapKrxXCjVZpkdp3KYUwB/z5
6U8q9I6fq7f8RCb5no0P0q1iFFw5ikfGv1rDDkTyB+Nh/QQGsPwyESWMnVEwvu96N5VKbL8AugRD
du73YcpQdBJw8upLcrElSJMz+WT2iGGg1ouYP0wtuOhARylPZL6QEBBmOqrJ7nQzOKTsTXCTH+kH
5KysTewl4uW41y2OyxsVyGe4Id4H4ebYoBnWxLJPaD7nIojJqySQJSrj1kFWl3ke3+gnQosD02ij
ZC2KVcZ+bvWrR9WF/h9czjthLm++5axyvv7qvy27Qg9PNDLCLg7/WJTjFH5Q/4WDkQnhG9ApzJut
3HWpTfqc3XFA+SW/NQ1+y1UqTSneBcnCwP+/8S5OFAvXskPnx6Pa3UuwmSbvvAVL+PlCpaaU2MTA
7BUJO1LqnXRAnkQIQjgDv+k4nZBfZJ31vn/REroO0YKYrNGC72MW9Rh5R75ZXslkKoVtMvGlUrWi
rkhw6J7Oc5IdWnRhKrbgJC/6bBpV3b0gLgjK4+IBwG6PsT/S3z9HMhIV8B98htvN1fNDIw8ZNzMs
jJEehrBKODywPevO5/6HCxPGR9jqv2VVGIVBnyg/Gu55P+AikfwO5D1gjQfNJcFJmsNnR+gqhyOI
qKHGOjoTrjNqLubkUckj+6Leww2k/NuYI+BZ7rNmBDMJOt9s8dg4GOC7+qGJITnl7DwFxj9/KPHK
5YPiF5h8kmXOfZR8V15TddgL+ds+WHabVc6seh45c/wGtywnp0kCoMldee79nw+ilIY/sNX8l7+O
/unKCazJX74MpHnTy3FgvQKi2Sg/O+OT5vxpHDxvw35yNpL854lKZdLpJq6MjD+LMPMrzAgDL0iz
CKhbVd2tgC7YJHo4CUU6JSYV4rmhLrWMssCi6vQ2Z20WyP5Jv6N/c9j3vgIkj4NT0ifdYVXNADF8
UIrPzKvLswiJX9As9aDx+4ozxs0YH0VqauQaFTyM0AqAVOHquE1/t/0AX0Fg57t9FIvrIHwfqi13
6PnOftodNw4y8oaAg/ni0N9rWU3843lJK2n/+H2cjjrIVYc4idkqWPr1svPnMDXk69Srf2/Rs8Fg
K3EiPqA5MblV9ky4+D/xTBfCl7p0S/g036RWrhYQ84YF8bu2AxNkmPx0VkemONKLRv9oW2U+TAqr
j1CK1/BcDAcQ2JUKIQ8tDQ/e+0mKG5AH3V7pgQE1cPBaIec1SFVkpkOEEijSUgKP0zd3QHtT2EN+
OdLW8yiqk+EoGFekCKS4CTbUj2EOm9odPv1QVIf3ONV4fn4A//lqOz0gTxO3UU4T7TTV44ZYxxXb
otn7vqqTBDE9/qhkkZz3MuwiMQdYp4oxsdCej1hZsRA6R5gcjYE+h4f8kxAdI/q2M2AiWFa8wCD5
fOaAf4oINGiKBPHGFfw3Xiye5qbm9WJYaRF5XsJjNclmkAqMniaDMMgaNeYXWwKvem7Pbc5MHVPw
xSO5V+3ydHFVRBO+zmSWy9FEZzIVA6vNl/V6/u69Ffq6LDOHvSR8E0vOLXY0iIdWAO7/3bU0onzV
XKliUydMGX9fASOMFAvqK5j3fKvZI7EKCtaKvouqsUHldyDWgpLf9lvAy3ZAzOUZVv9TuqOzfep9
HXogC96HuEjqdtxRTNJK0CMQn2JhM+NaaqgsDW6ekb5WTS7a2MadBjO1vb+xMzFSbr1Zl9sxwSrw
+JxgdK8zOx+I7901y/AJcfITSpvIJkk1zwcM5rEiFMiHhhLHz/D6KQEg+ZjfZIsVm1SU+NsuZqgW
GqOl+BpAtcccv6e0FpxTLuEDdL8lRFrB9MMhwYFaIj9GUvFNhkfFEue3gjNuyaObzp3YCzkY9CUr
ATopTh0G2+yEq9ajwYkfZwYbtOcv0mokgwS3qI2frMDO7j18U/fHNnHQBpDCAN4qITPlkVb4Rhx4
e2etnlSTQ0Wa7tz/rCwtMUYdBfbb9GFRwDPibSb0RU6UmNn1YPZeEIgxcmTEnwovgbiYmddb/C3n
j6BYuEiyAjGFdEEqcIEnCaClcNDb8aGh5MSYZCqYgSm4w1rgm6QYwY3JB8R/h9ftsi3USSBaWpW/
6N3R9U57Y72oxoir+SrMivn9ZL5wLU9SLLsuP57Gpn3Du23E4griBWWyI2fzIa7zB4eoVfi3GG1m
nQiCHwC7e6WKSQIAGiF/AmkmTFYGZokxaRxa3WAKxIEABn2fXBfx8YfxFoZpL+lGgNPxlRKyTT9d
Y6mVOqcO22wqPFNozLUhvVVHpmSVl3bkPJ5+hNcj3fWXlniyXVxvZEgv4vaE2gqRpiVppv3Hmtp7
vGRlESqE5y+Rlngs1QcetkUdYuFRDe6AXQmDHyAu5hhzRoaux7qaw3aRGfw9gaN275vo65O1BL/E
KiR8FtNGPs1bOyYS/hLEHjatuwYVKScGI4RuLfnoU1msP4QtVvewSIOTEIa5DDx98tU2JX1WE0AD
Oq0nf6gDcvtnQsHAbJKf5AjjlnRTvSNutn3w+McO2XJdiEo4BA36gBAyuXSSHOeK+CNg/Aff4+21
OJq5RXCfKFkazZKa2bNnC8+9qAPK/qYZEm5QXocK7+/LSZbYzkxiMrHq0LTPg518irPAGI3fIRkd
qFxn9cpg29vS/lM8MB70+0+nekKmKl1axUfiEbtIasuj12Q8qdHROfABSG3wDsx/9L/kmTMQj53r
2Cb/+tR+C70+G0SK7t9nIGSU2mNjF7v0CS4hkAKMnSb9HbXkvqdpCXSNGwMNzPJjmvPE8HBbLrgM
Bmb72AwhrcHyMuhxzyMbVDVJoAO5wLJ9RrqFCDw+SrxIewBWLpvFHLUsqrWSNsohknUpNqOYDLIQ
onNx0mlwgdsIEdRU+PbOWKNsn+rHB2hmDa4Dawq9U1DkCdcZDcKhBfxNQ/ld7Z7LH2dknw0Iq6ah
iW0+sJ4JHzWvI3Rdsxus9FIgLR5GA5Yd4YGUR73WAG8FLIRG/XqKTCsSkVAksGXUFq/zxr7K+Knu
dxA1idZ9u3elwym3dKQF3fzNekOQ9/Invu9Dvgc5V92g9V3FiTkdIdZxFhOLkl3dRZ8l7huYNgFD
5DOD5RWeof+nEXAs3SsyvQtc9qddrhAAGBWfIgsc31Mf1pWKPfawfVISwjZxndTDXmM6SFAiyHn9
36SoqNxFnmA85UfeYMPcAxr45G0nrOpI+7+F8MDvj/sEoMjB1Hx2YB/nm6t6zZz6ReYTxbER2XyK
TgPdZoKlBSkX4c0BLMQzKHaM0KhQUtEPWPapZ1TKKneApuMqWFXKvylPTMMeY2SbcZTWl9ROS8ff
hoAy1qQaf0emiiMNgtzLFimLsQ5J0Nl9JO7ocBRdMTJvJJaoVrpy5fv662NfIOyDcNsu1PaJ3uyr
FI1/jdSJ38SxAB5sYAG9BzNX9THNGkV5dH6++PChtwS/WIFzUDYqfi1fk9yfdY1udZzl1EyIrahM
1QEdo/uvC3dRmNWLnKhSXf4XZ1kfuSJIOBWIoWLo2xz5aFdCvzpbhdCmx77gRtKd4Jo3CXoN+maA
2n/4Hce8Lv8KDKsLnjuhhOCVzbsy89RqEFHlxgrt7bSPRIJXESPuH1t4JDU1uMSn9FCDIx51O/G5
agQu9OUgB13ZY5J4fVZ6oSCkP3q4zN/pR/uETY0nJnJe9/aFgH81YabWIj3w8aW28jpl6wgiGd/R
m4D8te4iLahzMTFbkn+DhXzKVvNcEB4QlpAWygYnaqmwe1EBUhJdPuhT/F51OzIIqKfao0eoo7Sq
tJcp43NiZASf9jo2tFfzOweknkrbaHCek19G+X2DevQZ4DNTvrjkXYzHnNsLvJvUQ3TpwpRhJEOz
FosMiU0+Zr2yjYQbaHCAFL7qgD11KJINvqlyJ0zvLQL6ZwX4dLF/TOa27f8zgMSFSNbzksIknnwN
qQq6E91ndIc0eb/OAduj5r8CsO3JwJqjo6hFsYuGG/kQ8ByB5710d4lni3ibGT9JwC974aFGq1oa
MDnkqayup7DeL+RENAUB/XEolEdPeGYmjJAeRaOajnmD3vrkzBjQKwoP715nQGj/sSv/nQGiApmo
2xsQNWlP1TqjAxXIfxPx3+7e33zsc8ySEvLNYq7//ZL5Bx/5HQKEEeyibwU8Vgx2FYEzOeYzW6PP
yqgBc7FHu8NWkMTggG6eo3WdebcZRkcYFNYU+wIkRYahzobb4kJnuQpgSP/wsV7KfCbxWTtAYpWh
TMZrXUUEP6ucccv8LmAIF00jvIJ5qVV8xCt5jdomAPcJcu5tnr3pxoQqIEabiVqBp5TlTsGGVPVO
lri/ypBpR4DknflxfRSyRceVMunvBUgeN2mzjVMw5eKb0VqdfBnil00UOF92AJrdWNCl0pgUbGam
yXxAeQDnLrkY0pQKyvWr/jaE3hnBt4IGaaBnh1NUwNh8FM8Mjwzz7LmzzLjBFE7+DuyTUcVLA7rM
DV6hAFWLyGA6X6j16x/ub2JYjDW1RZK6dPQdMlR6l01Gs/y019DwGz6t1ulWtWMzJs7iS9Hunbe5
DO59JabO7OaQk3O8MbpJ8ti2TynOOZYiu/8ybHOAK61WUrvN4z/2/QCBd67GjIAs+DfHMC+9GWhb
bf2g2mxWkAtki8M9C9mIX9RU4meoadXn92C6IBT75AfJxRgTq6G4ptM6Ad6sPqhQfCkV2BPstrzb
STL/IY0L9Cro77CjTeYwPtiuDdtGDS62TyBzex6zDrtGt+EWYDe/onT5ioZC3kDhloD9s8VVcVrY
I56xSJn0HQtUEfn0UiXgVyazAaVCmcN/+zkh2e7qHKg8QyYDCWA3lx8G5I3vMq70QpVZ+244fZ/k
rSgnDXj98iGknguHJtqeH52EHpFRfRs65S2ViPvAkJvRu7WUiEniCNHXF9KsRtXEX3LGH2zZwHUy
QRr7kiWJTazq9viFs47cx8K4D510+VxX+8Lt0zHbJ481ObgXe6FZevR+0tlFPaYtsKFZwXHGCBLJ
YkDPrRnUhRPweBD2Ox8sxsID5Mlph5hjE6XMtJMPQ2BcNhjGw6OWbhXr+3It3R6Qs+JnNPNc6xm6
ih7UQw018JElZ86X711TehL/7cy97n17IeWbBOSk8KAU0YL7kZ7f/LUrNnsBrAgfzdiemo3qMRBY
jhowygviSfJQs9EyXC6DZUKkvKioXQZkb7ZotZEC/5jOh7ziv8FBmp4O9waKYr2rEDhlQE1qptK0
d//jZwheX1HQqoleZn50K9DX7POfvAGgcO9wJoV6xhJCPmtuECpMCHXtEfUu9kYxzcVoZugUn9SL
twO1RN8+sMMHpD3rqFpSGxoaucx4taHlJ/x/lafOQ0WRu10n+2i4Q/odX52IjhSFwQ9vqDPt3iny
luZ7RpjAajCFSqxDGDq7LKNFxZ5bgCbphAOtHRW0mmHgzTYgaalvd7Bxuv/dtE9vXbDS+N3o8YEf
F3XJz7XPDDHKJdjwvfcs5PUUves7cEX5R8HG/mqoaJny+YNy3cBFeeMcHidmPvPbO8fydbj9XZ2/
SOOXI+ObQEXarX+q1nBr1hPBFaoeZ66wHZl+dfZ9YZk53ZNaK8MS7iLn5mmSO4B3nzq5yy/DogDR
ONdYDOfevXcToFPwMLMaynsIl/NSomXvOYPEvCgDt2rynq6aKyDrMA2M8LRS4MePjkNxCnOMqGR6
n6O9HogCkFWVBoPoEiOP7vRgYIS92tKihZiRHcGg63nOhdPdBcofZ2XhBbXOInu/gFZtQrXZOX3J
a6O4UB2MyiBdVUwTjPeEvWdf/q35tCK1t11OG+cCcWjY79jjLzip2IDrVPomzD7AyIkHqXLcfMw9
bFkhII1adWQ7VgeJnacmmr+ck427Dz4bAMM2QYmr0sBdjXknLk1mwAQLo9t6/PAd6QLmhVsFxbfC
JwuOpokGFpwxPYr78eoHTx9M+MMdFK+ao/0XLnPia37O4Yb4MxvN74/F8544wQArK54rmnR6Nu2n
HmsdZaHjgb5/ZBB14n51NaVu0r/5NaurfjGpbt2MfetzfRZgD3uLOakvORa4mUSPFii3eMdFPXqL
lXtNkou1tBWdWIRC25Sy30hJ9g5k3rCAWg4ZKVcO+XR3R+5UDmKUobRWwZUugy7QyrCsclRelrda
EC18N6TE4hGdGhuDf9T6Hjv605FlRAELlIwU52iiWtq2rzh+Keiq9AFbvMM/7T2vtP2zDo6JAY4k
eustKif/wglZpmORi30QX14IpKTvC8XytI8QeeYXghMnFLANyUMGBetM2bA4v3bcfoWNbbltc5q3
vo7aVjpeon4JpkSdJ3c8Rm/7zJWR8C+nW+3p0iSX01jZheajEpf/dcPFW9LdlNBO/mciuUR3JubF
eqnDN0M1ep4epUB+OY9rqckL/NJG7L1yBZw0oxEZLIIajhDI4jznzfCapYdE3uzbaSobKtot7Fci
gmVdoYQSxIPw6dQCi5jRKJlz89QlAfA4IJR5kV9QkONELvbFAjWhg27nqFAiDHtON/crlHgZtyev
ndKdCdHuWbOU5706udIuHRjWYcpfuu6sXEPeebXcTicMwzFfJNc+AeodyKDjttYF05LLOg2sa0dv
FqSy4i/ApvpUAJllIzCItWEUNCv5As9RalDq2a/QkFqyNEUaBwMS0RoVBa69oC3+ilPtpunU+TXq
JMy+jM06RCZbBkASc9rHEXQh3M6x823H1sCgOrgHpURrY29QRleltYII7DADsNU9M6Hbk159ADnA
5ufvFnX55C+G5Qjhk8d75ipmg2YqHFXYZP/IkzWM+ZoaTstYkmTnaRp9NDG+S1BZqOCqJ2PUETN/
cLz0nwVdJa5CiUzjjiWdZ0kfGA9LkiLs6+l0B2OBiAiO39sqKIn3jPOjzbqQIBnTO4tAFg1Leich
68G6CNOkRFemjR8IdcaaVlJGyIuVtRdx5/YlhJ2ULEz8ay0wjVwdYthgMcz40KrfvI98nj92jD6w
KxUcphKQGu0UQbjoL8Y34rVbzfI947j31JdIWxl2aKAyytheDH0qv7QV8JcM5HnhPKaCGKgNbiW+
ksRMMVhJmZFes9KReuRpJyJdSV9H8xo9fT8/bnX6bI6Oihd5S9f8m3aIKknvanIpWl98Mbk79Uib
GRnO55SnHoac/n3KuzzhZMdTa2iJHAWm2wr7paTDjYI384pqMuBZFLqspyXsx9gxBUW/QfvWEtPQ
OLjtlsrfb8PrAabYvdQh5Sxw/s1AxjGbtKsAQqngpddj1DhAXqWpKWhsLdbhoCpzTtxIuOppKzr4
17LPUinBaIZh0oyWD+ALTWnKxlpGicM+wZNumTanRQdx55C2BVKu5aAvdYHiJKbzzstIH1TLueFQ
uQCJ6CpnVXU8+fqd7zvgpkecTf8C663eyFGqA0CLaNrx8ynu3+nwyeRUDlzIiG6IeQkD05baG0++
UTjD+QRYc1FW9IvGW2yJTcglg504qx6J3s5HF3McrZRwNBet1UmFe27IHa4pmkrHXJ/h9fH8OO0j
f3lM5zvrftgRVdRX1eOtLxKsRHl8RpLBxsIGJcUiUxPdrKIeJyqkAGMZUhh9vgUWrJQnDwYKFPKe
DzRiHm7PT6z9ZAe0Xzn2MeRX4MkoPrMDLa9Msi8PnickAi2UNrfn7EnFswF2Zn6Z/aziUCd+vqN5
GHo224lgOw74gp2XGsdATLTQ2lr8IIP1IiJDT6ZhCB5Q6u+DpLO2Os60McLMiZ9P+XgePorAFPt5
lP7eWT1MilVnqXs8cItnjUAdmGcYFlEKOGgYahjSPo1yfzSazwJ218lmnG6syb07K+LNhZ6N4m/B
mIZK0jaS6az/Lr1ebykTlQxbj/xtKnv3v9Kc6x3OmJpCPNxO7zI30FZzpxdts0+Q411rrPdXOff2
wkFCWC+Ev2ushzJk5S0Vrr058sDMYbKXVhnJQ8xZcARN2VIc8pj5kNLBNdTlCG2XLwdwihNY5TLY
+Qk1rRbK28WZq9aU5/Tn4HVi/f5W2SiOvtWQ01Im/d9jr4Szcj2NNOR44C2kGJfX2TsU1SNK9WmC
Nhm6VgHdITyx+UOitKEHFtyeUym3DjYHRVJvN0uUa7bU+gxk05/4PhU03fzJQ++D+bWTVcbjNC8Y
pB8mnb2LlfhUW9YBGI/DupJ0fsxmuPTKGFQcL8v/7N+cPfg2Mlk5IjHvb+fI19SUfn0klurPAZ2/
BX9ANd2BVF+I69N1IbpQtdDOjysomxSo4E2urwbiQqufBQfv8xhQatd/sIfsMO/bjTABRia7chfn
gPC0bI4+xxkhG4vXxFdJpri+JInLKqw9IfgoP+SjvU3voy/EGAW4sHVILS3XikhtchUhh2JD1gvr
zxdVqbPpeeOqKN4n9JpDSctt4R6aqFAfszvqJEFmD4z7WgbrUOA3onBw+unugLtFmW92tmWqMlog
fUBz+yEgYFiZhiO1lbwvn8M6i/8xkHtewN6ZqBLtjEDm9xlEzOB9MqD3l4zOy4H+yXh6EmPR2DBu
Fyz2KpZYjhE+i7Ez+MCxHZAFCtLxfyt+Ld8pRJpP+1gew//ajzKII2W5gWv0JmkYkh6MwWhcOLSB
N/bRIWpOgffIs35srbRx5npLWpwvwwEUI6R2NbN62plhWGvJ3h5z9gWS1x9r5xoWRol3E/S9sQEz
LJWmUOJ+WPV/FnKkQhwh9QXspP8/b4LH8E7FaMYr3g+q2f51h0noCY/0P2E473Va+X6/GLIA41Cy
wkqGMrq3PAdlsTKG3/RRF0UgiyKoGVbmWfC4jFqjBdK1P5BtdRi6V0QAef1g+PndMfKpxM6t6ROS
2X5XXDDTxlfqJ2JyPrCSrpsnQY97ETumUDdcF4BIMRYdKvsStjiYOgX2E/uqXmhrNANTWlbupGfE
t4kMmt8z1MlCsx6xoHnHPSPdiWX4rRAmcPhffCcr6YBkMaSBXI2ezOgIg+sMFptu/qTKK7BBh7Ef
sNJ9UzLSVr3XY2Z7Ct+mIRPvC+DXqAl3SRnoD4ctqyVlwPvkzaqVFliibSNi1cSfVzRUsst4n795
4roiRp3wzaZvHAvcNMDv9gER4c+q/OVp8idolN5rkKqt2A4hp1V3adE7BLE6Q2KDB/eG+Pxg8Pbn
jmRu/j95DQAcABepeMMltfZ+7E0AcRSk1hkKJhqf0cS83hj2fFMLN20OBJdypm5CJAqXQ8ttxzig
sJ3Coqygqh/krmjVK0388eesRzSMEQV8h91PC3z8+FPO5zV69tPMQNSeFaVPqecwi0iJ3ZpymWP2
95r0HCPw47ET7JOLECjiljj8VGSGvcPl7KL1SiQkJIDlhBoOoSjdA0f1Ki0Q8XUuBatTMEmhGUsc
BBc6oH0asV53KnFHdJNE/BckanYMIRfoixqMRj4bZUXv8Rg3HnkCh3uOWgTxFPGJOCxqB0KuvT2S
KirYoFRYXJ4XziuLmG3KwLNXUl7Jvi72dInlWVh0woLjLd0uYgIYfKYJgVRhPQD/Rt22DFui/YHc
n76JwuKZ1wPtQ7gbsudjGtIdUMzQVJf9Zbk38MpWbqoB1i7IbFQo3a5RkyY1mxonlT2eC7RJBaTQ
dStmeRDrSd59K8m7swVwTo//kWw1fNPXzoFrnHbWG1cRXgK35SlC4vmtd5fqQJK44o6nN66H/dh/
+kjeMaP5o7H0OylD+12NMpQceelLgzA0LYaYjHn3mPzi3X9yYUic5F7p5TZ4zAv576D7jTV8mMGM
rfhDsLsiiE3JvwOKGNQM+pxpS753qmWKSVKxb8dYSjj8nswDsGynNkydOeh1Lhai+ou149GRYTWB
94Q//Jl+rQzaoNAH4zm7WweNyc3iilOylvdd54/WbeSx+IsV4gIBHpZlVYrCvzZU3Cu+3q/lcjN0
VQhPhnfPBRVt5Wz3/PXMdTWe7wK7ckgMcEHwo6kCLWGYNTnbOaBzuFZTUvrHYmo/bSvhIoyvMhkV
jWb+Az0FakMo0dJB5OPfVyBEzBDXBMXBJ72dnKlGYwX9hZt3BRmUx78v6d73Txm0QddS/RHv8yrD
0CFZpNCVRwAit5Cj2big8EXfZ4KwWLhQ+x1VFKHTiF/fMViHsaKEAMrl1U4ZEE0HYBYO+bMfFRdB
Y+OfwYwtYYN0YRrbasD8bApwz6M+TIzv0P8dF1WZjukLeTUCnMG4y8UinOiRhxUZIPA9KbE5EpKo
O+Uj69MBAmgioeXW1dYYQ9OyZvjXWV0Y/MBaXkJAS8hqo99OVRO2nyNx7qPXkgosux/+3eSDu+/f
MIV2W18agbqNHkH5SAgA91CHik/CEujwdIPd+BV4o0VOhk8W/duFoTCNHtDug/PnbjatNsLR7bQ1
4A9OQp/MJGiQ6lCUM0lpqHo1Rtz/gKHEuAk/9dX2BsW9Jl2iZs8UAg20tl7qeTwQAu3fhKMui0/b
zc/bvOoNW137yURrYz1w7TjtNK8kZHkPGrkSMK3dY6+KJ+/mi3YIqIXh/XR831jHFC+WPLVx8wWV
X/TvCsw36BqI169sWOiSvfAxexRHUnhE0erdZtrr9i4oXDr6d07QmSkmrabkRO64EYA5wft64cNn
nYStZB12eqODHpXgouSa1DJIoThZl4rhEAWW8cx7GRDrIjN81eIDfoHquvakYAO9S9LYkndV4tyn
8jbkLleXs1NpsHZfLh0OEMQ76hhjPoQg7sdFfzYCOvesSj8oRg/kEDn5ehw/vRncHVYyh/6kyp46
8H6Gu0d6i5t0yrP9j46NqebB81BHPXS8irl3OIJVvfZt7ts7QvdxPdcKKK98i4sU41RvBswJJw+m
o0CbeUvcXSUwjaM4tMFKSKgp1otRCxk/5zdGkzLTNh3SkjWCR3pQYcwKCb2hBZ4nLjGXEo1OBVQ5
+sxS1b9B9vGlz9J/vbuvV5wKZ1QUqIxLU7qFyfCpWSZ8Kv11esytfGEtz1eg1rKSEaBlFKTuC1vD
KeFuogDoAuYghXRwhlEAjnfs40eyakwyTR+U+VolUjyeD8PALpV1R3LbD85FSCVXJs1RCmYgXiSU
P3zwEtaqr+INYPpK26htPk250SyS8P0m9EYpH9FEW5i+vdENQtoqgV2bZXWax/qxCTrHaga0Vzy8
fgZuAs5nJank76qkkzRC4cddAnfkER+xco2Qs7InOV0g5S22yxjQ61UTQR53bcleCbFyXYmG31l/
brwJQVRVrY0H+14UsE+opvrzQZt1LdLjVb8lOhC6JPruvu+/ZANffGsyXy+gNXMTH5CvlN013ua9
vN8apAT5DnP4VRHgo1/+huG3MfgjXqD60IFD+qIoxQnQRWlPISEXxcxyYH8guzRydUMYqcBLl7Ci
764wqZMTfuJOCEh+oBbcklv8PITmtZbglbGfBoARwDgEXJNHg9OuIQaiVz5W6vzaWHQ+9aR2vJTV
tCHVu8QU/l2QKq1Uc+sgM/E07RzD4FqUjNVU8cpmzozxumeyzn+rKoMnf/KEjG72cy56Ih2bniZm
6EbCQKbzMG188OwhyKZeefxSsRTRRZjcMBnlJrOcjvDkRUqZGo6yDH9wKF2PD0Y44hQXrmCKfSRI
ZCpyVbMSLykbaxjNzUbu6B+iRzwaWPBjx02uPaN3HeHd4CTAGwcgHlVPgFsFKu6bRgQo7K2U5c+5
9jGRBPTfLoRMScE1kdo/qXdLWRc17blpIMu8fyaUmbIVoGJX/3xgitd5CRom5Zuy3+zlFLzancwB
MNOf5QjZMmZppYloV5JZqvWrq/bt3eCcNms7rxIJG3yCv/KAWBnLUXqtqN5K6ub8uOKdsGjUcf5d
heVStpHmt/Xlz/aZ2wlsNeyGTBFAL9E0/WagHGknu9981fPtEvkICwi4qOaUkTDugIvYvfTCbh9s
sRe3AkpNirEkMTfNqI1DZzhKx+Z9OhVv23YfFuRUYfQgyLYrMsvWOZfi0yJ59QEuwwCZD22LYW3z
k2QpDGfAPmgX7r9XfpXq+BBkoSSQTCDFw9KkRr+Qn6WqhvJ0LXGMLWsX06B6vBqwIPTnqZgRzYTJ
gQI2gVJpRFNvhS/fihOU5FhGoPqhMJHEYIGf0bP0xx70fm9W+v4hsQ6BdwlZeyI/YRRF+Z2sEgN+
5Mxx28xuVUDAY5/MIg08nTG6iPDnVVrdEBYGZquFiSjnWZrHBech6u6dxg5dZe/DuukH32wlX7kE
jfOQSYq/xXs36LAhHnPK3OX+aNpOQMmVadlWyjbAodEdNn/d8M0lgEnaYzpZBWD1tBIbRPF9Fpeg
9GDQn+V0Wt3UMjBcTPyHtNtKIjp4Rk32Qj1ItPmHSV+OTkXBHN3XujWuBSD6ObOneptQwrFxnvaO
8X99dlXwmnfkld6l7QApew0Hx+SrzM6kWDRvlpM+qM3H1elN2no43HfR1On0Tf89Mjp3QpIT0psv
beXT0SkRDuNIQvs9pf19Ej8bX8d1tNSbrpW48FRUOop99HBMCZ6Ga9RAbgUCE8WBC5gXgj0TclrS
dxGNv19scQXVqDUO/0YJeAXmMHb0ruBYSXjYj04Yl9qM+QsV3CUocCSfYkUn5UYjM29TrGNnQqAK
7PegZ6+givv3cOvT0pXkU9vJ7sC2qf7R+ks7HrdlivBS4hcCFzNIwc6uZMdzVs+2Uq/vp2HzFtVg
3nFE1ocQtY3eHpMHqlnaCR1g8w/qvp0yxlxE6VxQ8HMqu9iuQPBUMrR1Ao0fVFpxcg+SyXr1RD+c
M0fcIogaem6rltzJihLXkzbNH0weWzkWcLZrXSMxXLp/X0R+lIHRdU34jTO8TjFSYNLJMAvVhdNF
mroFz0fUjMoZH/FlIUgsoRtZd3340UmWX1IOLADxJlJqDZYtwFJK3rokrlGm94xZMV9vgoIp4PN/
toD5R19Db7i1K3UsT1vHK2ofN21bPQj0/5H41tnD0fbLLvjodeUHrT6YO09ucsLW5GVHL/K3zToY
eS5T6nf8WeLZqJifZNHzkzFbeZQlqTav6pSu2941gds1j7pFXwh/rq+OvD8hwcqsaFY7W8wTR0pn
L2ns/JuTNtvdOWZXArjZEvGV/ig+TPj+TPyytYs9P3C0fWIMBFwAf1vuALhMoEG7pgxfnOoIUjaf
jOaYxXtcNmFdoFveLWsFpQiplmBslAZQB77mdMExYg+0QGjTctTwDgfbYDBur2/KvlqZ6RRc5BoS
uG7mPds8+74OMF7PkrOuxrcJhl4EOKzeMnV51uT1ycerZT0JNLagFzOhXwS2OPNWahzCbVAHyn5M
xncUcecAPANTQ4TTLFR3Wd6hlsPjaK6MiqPb38oodKW/VsePpZTBj1S4senZxa7sc5zquC4yCaWr
MXOZswdAyYGFgl8DqVf0RMPNehC4LwjrML7x0RXLvLpf5SiSXrXE2pA662kHY3nwQYnNa28qFbZK
IFscWOrfff2I/mZU8UAqUK3PM5cQ0lEmm7xDiUGJ3G6p8Vk1TESnAAuxy/xx/dJx59T4Q0ZyhZNB
BzHU1wZ/Hp5HWoVdnmU5EvnWrkEmN36Nj7EWa/4ntIO542rdYffNsa42AsmrT13PQK2M7U7MiBqG
HP5eyc2zIT2TQFXd7btGCGRGUhhXdBFQ48/dNRFzqtqhzvZatLmn2qD5ZI2c7wRKcuxR5AYxNmvN
3T5CzBfJfHXZzBCvE0yuIl3F871sU/VmvApW58mu9pguMnNeJ/szIB8tYTMRmI8FnjrE+9VrK+qe
ndLaZ05CBXSRRKuFhzKeNadgrRiC6a0VKVLuQLLX3z+jq1Yz9kjtuOE1Z7q5tk9VJ3C6akvgGEtg
sxXUqQb4pE4HBywjJ7Oaf2rzXz4DNJ5E0NNCuR8iWMCei2Jgv6utDYXW9b/xqcNED3Fo0scn2HPf
fJA6DFfNcU8TmkU6RfYHDzQxNYNnJADh+LJrF3WOTZvakMJVmserBTYuve1gHcf20IfsrMgu1lry
2OuaO6tSb6v5We8UFfCCcCmmNy9MWzcLHkJ4BX6sHHCM9gvC2tGm/Ya/A1UXT0elacR+ul5fbkgz
9zISu65t2BOQqoKo7+1Kvk1VHPZKuv5pS9OdER9eM/jGc1ITVjaCMMHdP1RsvpDZDAzPuiubIreg
fK1SGpO+bfPVUn70AE2sXIg9CDELC0fb4Erh0Nhmp4l3yh8o7JPYbUtoq4SIzjTNJXJ+MQvfEEOG
3IjGJb2YIcvXPSiArIz4zoVdfgu2jUJlU49j5TjAAlwi03WpKv4HMS3QSMwj8VX1xSuIlhBUEaD8
kEuFd1c/M4Fy9cObc5Brzh7cDln/pQkVS88d9HziQjkd73eqV3yorJ31DyOZOSHjlDaWxxz7CmG9
G1E2nFv96yyPrySxOMdbB33jhQd7+dMLaRQe/RVGmzm4bcBdBkV4d29bfUzSYRCf1ahLZV7BY8Pr
2AXCEmBdzou3bF0f4TuPrlJLNUCM4idMMTD6Tk6vHObyi6XwY2ITKJoG2K6y60GhYssVjVXd8+GB
m5ld0Ygt00Na5rMkF/rc5tQ3rpH1vaHbIgnz1plPLVIZAaShVuhO+oZrG/tL/7hURlxZiyeaYAqQ
BZafTzgGfLQG188TUaOysxIi4VJM29XXR8OdVLAotFCYlY60+z+pSYQ57nWbrl/OhCHyca7gRsop
MImOYQBRNLYHZVCdPWnTQjKiTYGlRklt6DwfP8xx9jlif0Q+FEQ4aR1KXBI+6RD0PRQZ4QvozmTA
WdczrkB3vnexgVzfgWqAG4HYkcI8ctyw4FDLkagqSBd1mHOvmG9Ad9GgVJj70HahrpjvBlpFJY3R
aWE9BCa12PgxIxHC2rGlFjFRWd3yqj6kZjZfQBXhNGrspmfjYbWjZxj8tJJ+wubzEcMQBe0pqTLI
nwE24t19wq0vJ+qo1usCFYpDRicEz1irR4qcUV42w7Ilk8sJ1O5dhNFA+z4j6W7MeO7TV/2jCy7H
3AKqzHUJd0i7pFUt+CdAcoE/gnzNo5geUR1MZKOJ0gavKhJLj/TatHKnRnWs7zlGvFdR6rsdvBiJ
ACOE21Q8AeuiWLusX0DfjO/j9XSnjEjEfeV3mnXvw0QoP/QlTMmpVT4f9PwOWjnIQBHSJaIld+Kh
7iAL8wZslN8CrpQ9zlZoUtbPzn5puB5OxPdyT6JGJGGWT2tz0+28p4OOaNPNi9iSHgiTUlVAQSHb
9893iuwVyIQL1YFCKF5ZV3CBe7uqcZhv5Dr1L+r4EvNQSc5q7VeUu31yT8rjcBZGx+0UaPLmr6n2
AE0xGbr6Q8qJeu8FGDus75GEkQA3RuZsj5qCmRn9xwyeASWGG58pIla2O8fY9a4CPznv3aQwty+S
P6aSsvxDn0DivT9jTcTT3IOtMDsVcJvvNupReVn24nUSX4Hqm+hvTGg4I1pIoS/cSuTHx+o/Fgeq
Vt79Sct5sInpxPumN8FoQIDy5S+o4hXKDXGY/wqWt+aL9Agp3GvnvNy6LkS0j8ZNCWYlPZE48uJm
Lo1bDgr6hefj9gZFmGwK5skfSdy8IcWoj/1I8UdkprvrqYqWvmqIuXHn1p8zgR0pHX4dLlLNWYkq
vt1GZL1J10Mu66F7UH9E8IsLFENYBAwJEoNzXS6R2cPu/BzwhUgcFEwqozUciFe7ETOOcXhNc55p
RevRIjRDrk5FVA/t7GG+50dDlUOc5/uIvWJsb/AUrZ9mNvoVBAwHLX7Dq1XOLQgnb6mLdOWhnHgs
Y0TbZl+/tfYkAeI67fiUQBYbK/ZEQ2uBppdkYcidz23sAgUWOrtAxevKAw2yPJ/fCpRYOpg5ODk7
uk/8zn/aRXWVI/LfB/AWOgjRytYm/rltV9ws29sdAu11MmAXK5DRoN3RrcNqngJfpwZEBhN3zDq9
HJtVqAeCoTDhILzk9mZ7mk5aMa0CkfL8l5u12hS7VEIkfcKNdOVxlb2Q5v3HtwGFh0f3BvA9Yo1t
CuorfDkrke2MLMHFCljLwqxcmsJdtnfh1KPy20WEpodNPiVLnuDDQs4TiePcEktGoXfbhacGhwOd
1bWm6Tx+TLLkzmYQL7ru6IhsDanEu4Bzy6iAfxnS1zDPa4Ov80f/gyYwbDvY3FUmmuqDewj7ETTN
u2OyQ8C/TzVy339LcgGGEn3W3eCkNZ95aFDCz6ASaoWtYlkC+dM53eiQr/Iard4LUYfx4Qii5gfu
6r0QzAgmoIGMyM9pKigh0FcpHEGR0wMDegbCiM0OnTPpGb7HItkLAJOGPMAp042f7Wq5NQ1vhDsf
/DR2UXXjOl3PhzhFClhTjanD0Z5KmMch6dISUTvCOvzpGV3iXufnkUpksxNhCsM3sa51MFnQgyiA
aJBo4/PsWVQ/XQWK6OHOBgQo5MPj5MEWZBZUapY91DHJlDqJskI8OfwCgHNAAGhtwNeKfF9VJ6Id
dw/GQ/Y7tOwdbks/inuzA3f1qDS8N8+RkPx9EsFhRHGiSWr0pq1wAfcLllabI5URaiyCEHXdUS5b
Ecelvt3cGMWUudzT86ePNrk7oYZi1zw3FuOfdu2iDOOBQWQyT0wIftgnd9EIw9Y5M75FAc/wVWPt
leXm+qYHzwsISgyPhsbiv4d5dv1P2yLgEi/uKrHYggHvXLYqQ8EEqSFWhncBKpV//CtbfT+O31nM
aqEzhc3vDQDfb1Bjud5e81IVFfYB7bIu/uWcog2uocArVkDHr9tb7WSfwuDKoNHAE7RnXDNJih/4
iTZ41xKo7/pSRNT2dYnYwzhANuIJBP1dx/IYJhRTPVVzCzs0h3Co36K9FeViU7aOwMXZsNQamYiR
Jt8uxHc/wu9TAIaaJppDZKdoT+yWd3E385it1ozJXTr9FiYkRBZf+67emEWz6LHqjby7C/bIVpqO
RT9+Pazp9hBN3WIMUrZfVr0JAJ1kejmuPQjlIsejEW7BSqxk/L3g8/rOI5xbBDjQhwMJ3zJyMfhU
zANS+i7f4GxuTDUEaxkuom9gYOp8SYnYlpi78Qh7X0uQbbOBIcjpOMX8IPJe0Ja/BjO4E1S/DN/F
PajssmPlij0QzCxJBZi8WR8AmQBE0Db/GeiJOJ+hLmRar9mpiLxE6E3t2L0IuFhnKqdW/7PQG5i2
u4oY2oaHGPDf3agWObeDknMvaW8OqhYEH0gfx/jMGhJxRYY2v3ZjvhOj0rS6Kc/c3DOq8H5z4uTR
Ji7NP6dJBV0CgsUeNQh7Y9+KtzOc0KruUaTy2dJrIysa0DV0zbg915FAI78DNLE2+kutmA3T2bLV
r6sSWmIgPAyl/+y+iMDBj8SShL96cO/ANydFUDssMs2amvlqTPo8B8L3DfBOUwY1aKiJkMLw9aEp
7A2jTLiIhsOWq+hQ4jSbh267GjFyV330PBtTMZHeDaNo9d5+Mft1MMSQzRO8RuifU1l3z0fkkyNK
EIqk972jbHOSKM5oZ8a5LabSC5aPZZYNa7RksYcvoVMX29gGlP8Lrt8ZjdnYH6dlcrq5PPkMwtFy
PyYHo+frcw4wS/7fjQyM5u9cL1bM5SH9sRqhC3Gp9cwprhavyzfjYRmjq7eboUZr39Z4ZU9ywCnM
gX4fw9VdzSnEsH9anLLPROa/c4fTS0vaVGGQCIVzI9qtcutuNIdVQidUr05IgDq9hvt223oQo2pM
3Rzt6SaNI/9+SIFJYtJDdy/J52yGIfK48liH6XO25cfXxzC4XaEMTMLBD+MksVijiWd/RjlcH9UL
6Cq0CsHuHZIUPPMc45Ke9cgoHvYgStLyMV0+zAxa3oOp1PA22xH501CG0DfrUOZL5rap0AUVnHJc
wXjl+HKBiC5cTfWvTFdNiaD+HWVezXJaNMQwOTkkOKEH4myAhC5tG+EkEcZaKuLnLP6aNThl1SiK
ovVcOG/2uUXbds0GaqQce2GKChDb/YjfAvP4X+qYGI5+ihdOndJ4NbLImokRfRlz5mkFFvrSM9+L
QlYh9FqXprrY1bJZI1zHlRxqroAuC+BPau6OnjHKrNqMZ1z0dwkGuk57HYAufjugZWsDX7+IEjDQ
inAFZCWdsAIDIka1WEZLrAN46WSeBCA2f09/Jo6lBeD+2oDpXQ4ze8I7JOuoEnSIxh7cJOq0I7Rq
aC4Q3mOWVoDonqevOwLawA8aefAJEeQxwv/YsV1NNyAkOTJbEFpjAWmbIrpanI9zd6byyAFEitZL
/OWkkhCjIKmi44unk8CA9CyBfKpUdlMS9orn0NTr+yytD75jh8vamNo7LDJO3PvktnfAz1XqgV2o
uc2bHHOzM9IwuldgAUCNDFECLuDS7LDZw/+HFFJm0bv5eZ6VJTRZfIhmQUoigqnbqyKSfqJ6beB/
NB3x+W5++A/OqcSRy6f0RzuEBU8qatA/5nNzs6HqdaKk4t8F8kgCWsokeVIkypNEzX4cJuK/IA6x
Aan+Dme0PJ8a6HRLFH+XlzbvfwAgK7L4f6mRY4eO+NYkSGTz8fJTqvQQoC3d7AAhH+QCrn8FmE1m
mYW4xsdlEvfDCN4ToQX9eB4zhWZe7Alg51/l4YuaLeARlIRDCfcpbREwweUtxMInHbTOQfOl0OVE
1pWU645NYBw9NCobe+0o9XCLy10Dv0hyUYa4G6F0VLjDo75DeOG+XcOBV9nMqc69QJGSVQ9egy9z
W2BOJxPW3B6cGZzkpRrzMXuKdm8XIOR+YLrFdjPL9mqMl52STsst4HOPy4pDZxiUHLOe5oWfLuZV
VvbBDzAyXW16jzH3z3Jr6/xx2rWSoRixYOicat2MSvBtgMZ+RIvMbiUeGEhCEWHrca+xkWpMSRlH
aqPs1yB9t/ykWmn+KNasUzuenZt7MW+iP1E7IbjPDj4vPuFvT9cO6+3jp631Ok+FMOOevWkGAiBU
UB9yFAu5WdX9J9HO4vX/wWTn/56GKNzDv5sb8f/zgSg+yWe2Yi2N49ZJGyhy5q3+0+ARMcCsj1q0
Y0siEmcjTyD7RvsABppht6PeHe2aNrl/TjTY+4FcjqDEJora0RNmzmjBpSbfO5M0ohzeyavSRbwD
oJgO/pEML2fQtI3pxFlHky7hwJMFhtNkzaQKO+qgidtk9GbCUoI8KePvYmCF9CtpYhYyT3dfAMiu
3/IkgUQfvASMYfeyEhQ83PMT1MfI7hjilTvmlYep+jauzo2uc+g66v7pqM2MapG18dvYq6z0u8Ua
BKNJQqrRL/waazZaMkWxxQzO83kWRnXgtFc1csm2fkGAmat6E6iI/ha27Qqfpx6qPLtQqTprpzXl
ZfEZ3vFdlOFfmCinwWDrAn7NasTIrOUErWOOstz84FRxgIyYmO4eJRP9GSISEBgP0DuycT9KxbO1
YTiI2QaS17/nX2dKy5zTRlkOugThYty0NuiZZ3MQvJBdrj8zT5SUDtGXvx19YtOKjR2AZrws03Ly
tt6uOC0yXEUd2vay2Zd9c3tcX6/4Z1/tkRtrgcsO8AhaFyK4vZuQ/xux/DZUJ/jclDI84UukW8MI
l1o0W4hSzsdSdkSRIGSuEIf5gq9KPmiQ0JpFLzQX0j5f7MbF9+yvnR56Zm5mGqUj4xEZRonNmuG+
SlH+OyerS/Gk6H0DtoAXLdZIvc72tK1K+Cmr4Ts3AqHLt2jsmLDFpmhkhuM6hXX8H7gDZP/hvmZz
6x44VIppFfNduIpzR90srSLF802md1f9fcrnrhwrAF7kb+nVio7YvjoY9iFvZh+wefR8P1ehHkHw
vWSCXl98UXHPDoZZfd0Y1nqk71MmxMobnXQG84o5pr9tRAP/Gh+u8CC2DFe9+0cVi4TXaGpvPEMO
Y2R6qHR0xqJcGUdcJINCvVkWDLc11F65VcZ9CeUfOnfC2GgLhJdf1UbkA6alcIj+d8iERmDvYpVj
EZVTFNXpZczY09H/rk/zvsLBaxyagsK0HsasYOGmMhVdqEOfCFIXeKZlN3qBPcYdAWTqs48Mdq4Y
RHCNbyif92XdcjPc91XN1SpCxuzaZ2/SPv2/ekdF8ti88+GvBABjJjenso8ghytZhvA0PmgWAyGN
QWoipLagLATuCDTKaSzEcwRq+PfI9YZ6WVwa84/R6Eetk5RGtAF00mEBgcpaWGE4fAXn186ia4OP
+vUloLFiAt6N+tTy/ruytwT3GfLbnd1TmMJ9Fm17zhuAZ22G2mVMTpK+tKYnReLr9lAhp0TP2L75
nKOBJKLreooYfBeS7/cSIgXkJvs43yhUVxgSdhNAu77s3HCDyHYqZx6G6QKval8kdBE+ssH2ccph
iAYKMFGtlPjPkWKiquvBNMI1Hxmvgo2RJSSldiHU/+al4poHl1F3+P/yCB4vr7oG945yO0L2E0qX
4VAGmbw0oV5trrxTDITJQxYl2XKApm7EXhVCAcuDyDluTf+kqMm70aKxG0yR5u1E+Fdzz8nxx0DH
R5hJY3aukHyIroaSdpap3ruhxUxYVU2n7lSflrUwbcF1ixjT9KXzxoYobgXNR7AvFNQ0iqWfzaR1
gAeZzH6vgrQnZz8vEUeK3DipYAmMVOUjz6UB33aG8bFhvBgphhCwP7WUBJ9OMBGepL0f0nWFPvtz
8sETTDFyK7rc4L77T+8mwS3tLwb1zu/uouIYzoQNMLmj312V6EJga4UT3kaqyMBzz8N+0FH9cCiY
tMiZ0V7USwng4EQkIiLPKBRUUxQxYB6OkLuDWxzuBvpR5P/C8iPWpXkyLB2q6wxvVM7k0gajugiz
Wj/DXB+9GHa9hont65Vlq7SZCPq9G20AbfGfQAMiElEdz3FEgTZMXeUC2iIAEzc/p7KhunXamAOj
yLi4MMY/rM9LMVDSsCdstxZvYzFqeYzMLNeqVvVmuOyUc+ayo3VB2opkj9cjsIHKtUNpidzv9OMv
GSxXXmdceBGKOhl2oB5VjqamB5lCyYtUHmQ7kmiJ0DwiVKSilTetqA/NVzCqGFs0wfHc+l5G4+RA
dRmif/LIEqu4VUvjcTXHOAnT9BR8R/+zUE5z6nVYRMdoOFCze8ZX7g4WKUvZ2lzk2mBMRuj2i3Vj
LRRpJ0k/v2lsxKztr1i3ryS6OMJY8G99w3FFmVhwT69zhigqdYZLvCutDgauCUx/R5yHSaEa+5jC
DjJ8gNu0fpSytGdkQ+sKTxTAGyp9JO0w93Rnc0ahlw/X0UTgggw9SfswIOIDfw1SPRlLBZCCSrHT
5YrVQ+FHaOQcgYsxlwz/zzF4Gyb/Dbu0jv7ds+WHlIkzUo+helhqtqEMxRsp61wMHhorc+JknzQk
0jsSCB69Km0SnRngasiTqOFrVy14Kkwdf2Ly+ZqR7zRqm2oD63rQJgYdU91YZDN4Xx5+REfFyJWh
Uz3HzhMs/wU2z1FmiNGgAUWPh+Gb1IQqDSKSnszDgUBz+7T0A3olT7tAFj0n6p3xMe5c7ELTN0nA
1tFuxsFViUT10KI4xr33jiS3dglvkVe6v+U3OIFyOTfbNKM68Mcj+KfxsRCrqdZcozznSbyN6YUi
UL9Ll+MZUfxz1p98HdW52bN2lB8DCd6feMX2N19tUpgNyU7mxazMKHU1CSfo8UHTQPcyb3vmhIGi
wdFhKQruJnK44N5VNC2ES8jjDLq0+5TWdF0IY8Z49rv1H4ze58fnd/YbDEzevN8+Pq6A4wXTwzmE
DonJFO71VDX7XuZOpa0+0xjHAq47C4aBZwbf3dq30WX7JE0qBRF8hZYyZfr4/yNlNj3JvY2z7Xme
hVJ6KCH6Empt4fFm8/ULuaj0tMpzi7dhksYTZRC1XRSdeTCY5neYuZFTYA/8pmJmrcS6F7ziBOD9
smWeG3Skk10qOjuZ7zM3V0P3oqVe4bnZwY3o6XFohe5GGALDiPRPcr4eyMSnYvijEXivWmcszlDU
Vs4bwuieotPrtFiNmnBJivoDGfDSuFr60j4dJJbE7yJsxLmNUlumLFZLYcNhqrIe/jdNjrOjZ4Yx
daCXoHaERGtU/bfraQx1HfViwU0qILjiGV08j3138/m32CyhBm0i+K0LBYPslUnk0QhZyH2oVc9t
Zpg7J/YPoWURP+V++DRtAC2KHHGdm/rOMCYRfYdYP2ZHxdKgl+mZap8veA77MeibUEZIgdzmcnVT
m7ve3biO1MAZ6p6D323olBcpmg76RiTcOZRz/Qo/LtT95mbrrCVZ/9qo+YEm3EiKhx7QJDtLSOP2
onBmaVAgQ/OjkiM4VBQ3/N7ojoAvZ56AhlCgkOiDztXekYM0ekxzel+XZwIq9DBGsEl2CH/G7FK1
7QfqwU/riTIUB4Y/JzX4EiUhOE/HMxTkFkcuBO8dBK/vJHU8av78/gtxbotBr5CiqQmzOs/wqJhQ
o4wI9Kj6IzTW/Tj/72oAWFGqryF1bi6q/K+Tv33A6tpjYOdRhV+7Z1xLuFeOjeZmoFqCjONlhG5g
RcByX9H3sGtq2lEbfNGCWhs7t0zJCxxULaRJ7vgoFndsR4SG0Qqh8bbaSK+E7XIfE4MG9aIqVu3e
fQvprvsJxc2hO3vBmbqtrvC6msJa5s38cnWG2DGtUvr02nMCZ+dReF5bGn10+VE4FwCRgQNHYacm
fN0W3b3iAjb03qJ+6Q6fg3V2g3LxCLtw+qj8B1Qly1IjHR3rrwfxTfKX/n8cQQOF64d6NYdN/pC3
Yf0x9MdKe0ULvjdV7xs0+p56Q5sjV79Ei8jaCpsduqgywYtHhkIisoi6Jny3IH79+6Zfry13lCGw
Wx8zLuamF8zBug9m/z7PiYwws8LfJksHW0m1EfHkYqS4D4Oub2mxOAmgvU6dwvF+tmmIEh26gNeA
MXGxFafURybJr62Ii+AcUanm2mS0gXf4MryhS1pTCkh/QmRyGTvFynAQ09YlqWsLvg+8KrrLPY75
aiCYZxRlt0617jDneEh6071XZYn649Nege5FduzAVbKT6iVuzNN9+SYrFRz3cOuhtWaPSqjSfVdQ
sLf8TCM6DfKODpEJDTXbwqVlncfm34RdQvNkfMA4FKkY7MLGZqfs1k1uaikdySNlrnjlLFowszYK
9+4G0OjAGQd9z2tVhr1OHjE6z6mrzGMfoCwzm1xT42ehep515eVvzRKDNG2/J63kv7J6v6+sypHR
3nJfVS9HWbmPrSgVHgO8nPx2vS31H+wQ3TyVQ8cKJHT7FIDNc6+4xsRgy4eWoPh0a0IKvN53prfq
Qj5b57gXvjcmdwwrddV9exR/xV7fsgWkZAnZnIZ1C1WGq/Y+33k4gVBmH1AUHolsbIVVCMK8XX12
C/KR/ciE4oxhQ89WtVrUQ4kg3peCUTEjZJU32epiWuG2ZScTtEVFeehHHE2jfwXscbcMrxYHxpTG
gP1z/reyMRwzuq9X2D+LcV8ewMJX69aZUT9wJt0mrh9EWT0cNs3mreKxuMqIOd1mEsNW8ZYos8gS
ohpFsu1sHzLdmIZrpUDHfWPF547p1VBEb+JJGip6A5QJNPIfWXRxvEJwEFJb7xFjdIS/m2c92At+
W1pvAbJdD12RHVO9LZhbCYru4wY0wKSgmkJRFwTDHfRIzlC3H4MrxppO1/8Cxb/JdD9EBL++bdGM
QB6Rp7iJ8jdvRSJYF4Vma/70z48APqrheduX7gJz0okkTa6Eofw2QrgvpSh6oq3YnufoLO6mdeWt
FaTDL8xmZ/WPp6m2lJ6EyUROeThdOMsW6jVC2be1a27MqfHTuH/tAwB9uQB2PQKRhWdBb9MguPlL
4d49excyZFKJS5LA6lHpEVztAkY7Z6+VmRQwlH5UIo2qnwd2vVhVjjS/vglDleVkayAgUTMPyfcL
2XpynP49MP8EiG/eNO5AAkfESfqebpCjYI/GxZdQiiMzzcwKRxdcsDU5kvyGsGiCUsKhXVTKYZAP
bDELZn3aFImyaR1QVNNitbfMvqCyxBt23ewIJvswNhyT5hZD9XSUi+IvbkRqvALuPd3fSprzYLHG
d0jbIb4z1c8YnIiIXk5sCx/AWPuLanBNLS0ghaZWtKi6hAhrin/blD3NWE+sEwstbVSMogh7ekJh
DNWzHqmfkFTKkS1ixyXkGk1UMKS4PhEBXt4jN+5KhpScKGWGpPVjG0hRYnxgTeF3Vc7vQphWbJJI
UMUHOas5SuwmWtqGcqMGtvtSoyWc9W/4YLbOyAZ/wfClUXEHXR/c5xwUhFXA0nsNur4lGyed5M7p
4QxlGIx68mOAAuC6nAcKlUptBG1peWXLqEtTzhRJvIJ9SCPdpo6VlhnVx6UzFWJPnGjXIgNQC4c7
amJv21WdlbWmq7ZP/3UidcO5F1r/fr//k758GLbP4knucZL2tR5FEOEf+jbiKGW9XiVplUbwGqjN
ZyLHIMeo7vSn4IMhWyNOmwfkDADDN3/REbdsRXAKcLya28O1mlBuxShm1mM7jP00oViUW7M77Jn1
MUnfaubxsVsc6HBpT6jTFeprHkb70/fBeatTt6ljK3yW9K4vYMaShZGdExNSp5vnTcB9aPsBYk7T
w5fs46Z7I2fe4GzngF7qoHL9VQ5y7mCwMYCZue+lsUKRydscW44URxTEDr90Zh56OlbX8v5t0Eln
7VtjXXoi8pXVA/4s/u9uCmAXl/+IQRNpuOBVn6ZVCqVJbbf0sZBdH1HYcccippA3umYOgf9oEvHT
LZvDlFvxFJW6lIjqGC0gvpPahmyj2jnF/oxQknr78+sYpQ5f8EqPhaOBX8ZzqFpQVokznSWT2N66
ifzDlQQ7bCAP7P/vmuzr/uDHH/ghEoWBojDXRhMdk4wWwxalR34u2La6j3SeTkfNHnyxlAooJ/Jo
JtztvWPYZXba/uPrNEohwjvO569md0Ck1YfbF51salF4Kk24jSpKI8RepJkRDXT85rW+bLScfhIH
ZOepZH/5XCnta/VKYaLi9iPnriPbS0O/8289hlYFO/2xp1AjG5T4dlv91mfu7LQ/ZqskAAzBsP+C
L89ifCdpEqjnifKJOcBuxFRJBn7D5JR4BhSr+q/B56Zzm4IhJFoFuz8YLN0762EX8QVhkP1KEKdw
jYieta/PVYSxCTq1pApqILrxyhinDBRC1Lre8l1PwxsNWUX29CRPNLYpF/7EkvDGyL4VnAu/3NnB
ABnImVuD9orygPKWbmttm7Ei5/K1s2ep6IzA3JfLLBw0E5lXjQmi/R/22xwXi7pjSbKr1QVBn7UD
k9++RRe5/th9XAMEO+HwomHYqwRuuQXnYFeE//OEJqjp2rIJM4JFZkig3yjSVvkPCQsAHBz45SgZ
ScHLUEYAnksGP+cyaoCg1OZ9QGXTzkMsM+ixWDt587hquYs1pyM2iubml5ZMuMsiZVHwL9x0ekiZ
KpLfl3b/63xq8fGMjEhDTYMppjPHEujOX/NdlfLbl98HHlq8g+FJoY4J6WkqkIbt0qLbJ/UuNG+j
ImHymlgRWqPvwyIldiQjCz4rN1BVrMYi0m0TAynaCCVgOMv8rnA/Ee0+Qsb/gnLbaDICHIvaCsko
gU2JasE6DQOXzjkOpFP4h5NLJCvyBWwlOwAz5Mu8j5lO9PnhJIMtSL9P1Zujd8pUZ7iBGetQdhka
XanUOdHKVmF7Fo3ou388Nq/7J0j7n73rXIL3jWzjS+hnB784nbaOXCh1UhqX4MCw79danPR3lyHM
sXGVf2Ib41XufYu4ONmuo+18u70VScefOxFli7JK9A5dwns59tfGSmgkMH8diQp1qPVvEw0yijkl
Zgbwt4zUOBfZsJ8I/z6nX72bIWeJHfc/9jwP3ZrxFmnsXJJljUVTZLm1Y+5XvngaV9KAuY6liGjV
mbTpfjX1Iy9DAozeQSR8bIe6EKQ23jKTxnxfh140qaazd8E5yxI06QA2fLM72M+E4SAp7cNH7t5c
31Dc8F4Q1KVU+4OV70Fe+/u8ReBMLPoBhdE5dLfF2CqCH/yu75SkrZ8SZ/qbFomFt0pW9RBPUqEf
bAe8eH/vaKn1U8CqGLjRJvTSYVjiC/84Yr48Ugv9UaNnp1DfIcRbzHS5HY3OoWOowVmvKxdpd/su
A3QcP8UmC2MS1bUS+03hSdu5WCBbLzpIxJ0Ls2TB5F7jWp8r3qeEoygFLldJsKUiH6EkqFcOKiNM
9o7yxreBxC8C1lilRKu6cAZf5U/51IGqUbZzVYV2idlA0eBto/pVEl7qI3S7rX7A3J5yDWGOQAjv
ucjsLYgppWjOuil/tmei6+7uPkBv05PFtT8RmaOGc87AUxZEFcws/iem44fBmo0S/wX1cwfklA7j
F5hnwke7y98y0NiKUpPXUDwdRo2afAoMNKFvsukxC3m9to0QD6I05XzVtUc0PIyXpJRHfNdtIiyW
kPo1r1XjKcbGB7FtAVQcJvFHc05Dh7Hzbi1Nno3p4OaowjGFGX2jSkSFtyvBonKAyX1NodheQ3oH
NFA7SMd6Ri9oAYGExm7fNrDuCXpnPRM1O8QW05j86z/xnsHsHlUF/hxETkvf+Ne+8+MT1bbOOcOl
mx/82oUQMIK3zll0uGxFD2XDVOQw+1ZI4MPSJMUvnsllDOt6dmBnNQmaTuyRqss4mFOtuTdgtkky
6A+0B0vk979izY4/hsCoEUeZM5yJuv5PqjaoKG9ZqJcc35N7xvFK6piS/Lb5cUcaCy5uHeW9NhpV
hGL1H8xRAZ8TP3xSBLPrlbcwxhC3ykzqbAAyK3pP1Y67Rt5PkZ8265GcqTrHtIe5Xtp7s8oJAW2t
6iQtHoibN2P5sTChzeidPM/5a4/B1YbQhaEUvWE7pa1JSykaK70TEuFGYJikhzUuYoS2yjMOK5wW
ROMuNWz0VE5xr2S3M+Mqgg8md0abT4tebuYlBPLc5ipBBM3OZPY3rCcHdTnypHiV8AvWGQJfP/GG
LgjN3eH5IMUrq+DZObzBQcVnri4yOV7ArS2eybVEr46ReO3/+hzPCoqsPso6D17/M/Y/0UE39tUR
S+gpsUurvIPnd6aHz++qhgZwOy3y4poSoLG7BhxSZUF4ilYeX3rPjhCbl+dgPwqSu7YXoN4TRWBd
9GpI3DGnZmmcXAzd0oIjgXnN/+NERxl45YN1+CM82wWDoX3I2WJk7TEixQZjsCrDau14StkaNPGi
vUoIM4sT5WXQqAsVtGK8zr9t1SACfkcENdB1owyrQApvq7ePARXA9GFCeX65VsFWaGxXbHCHLFAn
8oENB1M/w34yCjtOvNnFEwnBFb5DpgD2SL6g7zU4vrbi/9dTGRRFwlEbEahbxo6mu3C5g3juMqMy
zOW+029Bz6KuDTJvnTqbfwXG9kqtA4hO+HBuIfk0fhpBeuwjykWhJ+QnnwsIwUvJpEang6KDBfux
JAMBaFz3LH1Qfqs+T46qmxrwIW0Ajh/9ASo4sAciprbLghVu6e8rLJ8kek/1HgkA4EJFPhM7bJ8R
fDscjcOmsb2B6OBvwKPd6TdIBdi6LshPLycLJCjRN8KOgvwrtx5PrYpx03Vh7MEX90IS6uVWEbvm
UvmMNb7BnC9F7MyZ095m63E8k7gDPJmu0zTNYAHDnkvxiiQdwkSjSFQXu7SDZmpClxM+zkLkHr1X
r7k9RTTbI+70+gCksU7Rd8tCOVFIev3TT2fXEfjk35gF9nFa+xjTBDkJ9mA0NPX69+w5qjNUQnO/
oTNqLLlitB/xPpfTB2mUMZmhrU0LH4bjowD24f1his8jyr+gosmAQfAng9lWP53oRuKJoR176NjY
vGn9GLXz1DLJi7XewK8YRQoDYuDrX6bGkqbGITpev4tZB6hDkHNjLEvyFZiB6Q1xfQI/ss/UDXNQ
Zwts6V0s4/JKB/Np3jO6ItIBOVeBGZqiBSOXRDVoPO7OgvEUgarOy9IwuNL1+5/CLPXv0HMFTzsc
2OPBrOx24kFZX0MVb/qs+Xn9+mt69S4xNUGUQRpMJ2VMj1ixKb+bwGSRjirLo//deVR2TCwlPPtN
oPgb3V/eN/drWNgMAfI7xpWmJewCZRN0MPI05V0QU4grW5bSzqlVqQyKnPNC34RN8i4yHx/FlKrr
/zZ3C4rvdub0buQMdBOXHui5BkostHX1/1XAC2eeUlJr1xTO6yh+yNtyTjJUCbcXwAXh1PQTxs1R
rFOKmYYGUgsclt27pRGyYx2+1uX2u0M241Lm+BRfbBhwJWYy1kE1TitjIND4GHsptxgZtjpYjuuu
ieQV4Xr54Zz+gCurcT4b9DnWWa5yb7mnqaAqsFo75O6xiUHwjmfIzvB58Mq10FfARPAi5VZ19fGe
pXBvq924dyzvPTkxTI8S8sH5b8IVHmsxEjvg4p1Y6CFFBpdHgMz/amgcTeLpBhRnGeeiH7qcjBzG
wrl1zl0g1oesotOYv2QeLE1x3tijwXaJNTHuVAnOKKhNOCm5Jzi4NCj1RkBLyFrxjfB5/Z79gUyO
cViOfIBF7eH/raDpQ62D729bsAp8Hid/8Z5l9nXBzdqDHhS1XpQ86a5wTFc4nimk9yLMGt1UXNtD
BJcS8YZ7CwkoJdXacCsRrtJVgB2xnAtCq09am8pgWP8f2kWWl8WqzvdiaP9eQtWDbuQSn4DQ5xl5
d1SU58Rjz2YADDBnJvlV+l2EReIny0SoR6UPi5Gu+9ilWYFURudBuMJmVODSKuVfE1AKYwdTXvpy
G+xFlscF2g6gnZHQfV9OTJg/AEHajMOoYxQu/Ec99AXkPklWByYQxUSYpKeOqqnPh9mDs//nmuoB
6Te3STD//UqBBOMKnbd423vhhQ1OYxNlemSn6umgmk6/enlxBqD2TjzAUX02CaezSYzTUbwNKjl0
/WLlmCBqurKKBR1iMrmE90ndlYE/DjxW0j3cTaBUX0y1+vzG0KFMUVCgowLTFyumgPD6dFko8PKZ
L13XfTUG39d5WstK+BMD5mWCGnGdT2WrDYzO+Dib7BOHfQUwxX6aM1TqlzjInUtVgH5ekvgXbhl3
ftkN5XQYYAKO0jz/UB8+JY6YjS3gcwJnWplUeMwsXagMqF8xf+vit8xtnDsgcqEEfgHZ/zz5vfFM
oEWph63ERgFh7wHYiavraw6l9SIAD7FUXnata4BgACAp0rLxBvd5qIT7NG4ZX+oBjqIiQLubF+Zs
FBHGf2pQZ89Tex3ATy4ns8FqlIocWtuMqipHvBvSSAis/4nOCL5Kbrimt4XuIMJx620U5EWi/O1q
Rx7lp7HvncO7SQB3/ofDdSG8B9WsVbhBsav53zQlYrKRCtOPbWAiCouXqMZ3kNjoaZRha1lSxMOC
lL8b5Zcv9ti+qH1ad3oR1xX2ZztHWm7ht1pSl+CoLm2qqiodwmWu/ARj7JEup4WdA2Pf9LCxhzT0
DElwuv6yPh0VisrnwSmbpz4F173rCiaIEuprBQRizoIFvAwjg3aKqeLIZBHskukKm+KzNJ8mzrLf
5AsJNy68qMrJpYhkMo8sKyPKkYZ7jz7QsuwFIOYaxxMcu5Kko2CL5Huos2ogC4vu4TwjVHqn1lsQ
kH7G3yrS1IJkjexDkLk+AREQCDk5/ZNdSA8pwJDJMGSyWqj699bBW2oiSjCvUsHil3pKHMU1aJCC
B63Y/AixLwL044ZySrC473QZDW5+Nt13ZYAF7FuYNVjIAmBHcGS0p1YBjAQpiCqhFcz7PkzkF5Rh
ruIhKMhwulloMcSmce7yL5zhWc17FsGCNqDaSyQl/K/PVdkdrJrxeC3sDgnpGx9X+lLOM9pr+0jt
iQOmONSjZiulJ4gcbpGUUP6ga70qkWXRY1OmFFdyC6OrrVPGHKmmIfb6T6qrBG06WzHFdJCWGTR8
oU0YabB1Pr8wSYcmPKK7kpaeOYC/dzN1o4pfJv9cKc/DmmMMddhKbQmt8rYUYveL7XmF+dlf2kAj
UUmJZ+WIsnZGF5cOzRTWRTdEU5aqdL11USPflGm3WhCBZS5OHfEIyQ1xNNr83L4IFnpivrnM4d8F
tUNqiyALNsJfw/h9xQrUyOQRNjOnoZV5e+neY5lzMBNaFgDA9lscwB0kfj57c/71jvxB1wL32iV4
wsR1hYqWfehQRq7J+muXVv24wa5reUzMpfW1aW3wZ+aLji6pMfKYw6tfg7HZXGmawhO42ntWBiyY
kyRQCy6m2V3mOdp9QqrsIphqCTla7FRtfGf63eIb42SyMv9euuG8mdmndRnn7Gh46fq6/MWCai0j
obThoSZLhvwHxXXBJhyyg7OUTHl6bTGYkl1T69eId2hjXPxf4M3Jm9AF9i2UvNHb2Mv0D5MYXnMf
mxfG11qyTWoI9Fif7+DohXFIp5veg4flo58yOHIhD5717LlPcfPoSSKSLZHzGH64DPljEehzmQzB
i92ln01IMbKQw2JB0LqSvDCHPG6AAENKFs7hjomRO0MudZB2fa3fiDkSzXEAb/vIuOo4tV1hesuQ
BhzbPFjsibL4uA2MFI4h2nQJRASKCML9rwdsZVdMnpAZPDH093F76gj87Pddo8ULwdlyPzwQI4zd
HIrriQEqOqAnJOecwPLeomCR0SnShIYAvkLvS8Rfvp6JrN1gD3SPXxP/dQ3vcrIBRfG0T37cL2js
afCLWjLi1YigrMBOJq3WuifNwxPkfUp1E0/Vwd2sT2DZc6JoWUgPAtaTxdbvP3HrPGDHgxR09wnF
N0HZsG8h0fBwT3zbtkRN/j6FK16ZMfHA03l6rl9KZEwZHQWA+ZlrKhE/7lirvIERHecm0Ad2dD6C
h+W3Tv0tqlCBpKu6yHcGJIK6glb4oTC0Gs0XsS5p95fYpCH/8fG/07+ePD0wD3nwelBMLrEhG6xg
jXgLvM9NiOpP+x2mx1V4wbcoMv3dfhSRCi+rpUXew075hm1GxhqQe3X/1gvDTEh+exXsdJtdRZTs
qBcGZwB9RMAODNcJtBj1g6xLsoITyClv8n9E5qYjsL1N7QfibY35dEs+qvjA+nM3RyFOXpHCYWEm
116QDHda84xR6rzcKiwIW6rJ0fK/tXBpvq6tRz8HfTpZjguWgRvnJrbLfKEvzmTOwE+uFtcJK5tH
Wqb1/kob/reRjQHzLX+VQVx90E2R1+FHENFfgJOZwXDEXZBchkleoAEGH9gY2EMBsVDP/a7GC+SL
vpW/jXmMDyuLpSBlWIIUh05PPGXDxHzsrWQ5hcuFgOPCEy3S5xnzyEN7UhuT/Csf4jc5oGkFuSpT
6NHIe+9t2UNTVfUJOnHWerihr1y56jg+pi5Z6EQ3vY7xbSKLOryXycrDG8c2Cw93fuiCP14vjuJt
mp1UZ0Z/rZxru587Cxile9mPo22zJQrHo0u1uWaOobYQBtfLULS8OpFG9qVvD/0w2WjBN7X0o2vx
qaoNcU300DwkZwmeAllG+4A28+BWbOGYF/yBoOU1eGC3dIBIRiYdUZ5bYJs3ct8BQ6gQ82Fplzj4
FLwrs2+ltp57E/KylL7ZEmuxT93n0NKkpXXMEo8MjvlE2XSwU+BLMzol4P//zjZT3LAgbqcmigqA
ZdVYehwUUWD+1sRhRmYGiYJbq8NpAJJv441gfBvcWk0rwN+q0A9jNajJDhqfU/wYlKa3BSeZeY08
ft/rNCHhGoci09wu69dAJsxDcNKvtUuBAFQ6JeqUnvz2m/9zHXkWFFdsPacGT0TaKHZYWf0YstPV
09Qy3TPM1z/X8y+j4v/3R/y3h+/n0Scm6PEgWWZFcof4+Q4LxOyAN9PhYfjYCkYjCPYp6TrA6y58
HnBmEIShFP4PJqmZi8J2IAujElHikINwKzTSB7O6lYxceyNM7K+0pRkhKc+nPx4B4ckXw2DTI6YS
eh8jTq2RCcoZZqyg5OmWDWuWQR2oobBiba2oFxBudgB9jyTOql+0rbpeN9KJJXT+n5RYhrDVT+Ny
DqQnUC6Yo7h6O/FCjghKSh79B+p98PsEPEzwHuBtCptMizcJP3MdUHK12sj1/TZ0OKP4RV2qRk6f
jQvo2razNikyThmz1F2EmONELu2UZ6oHWWd6PiQfB9+q4lWpOSJDVRmoYq/8u92805NHZpCjT7Nr
PoV6+n6RE8c97nk8tHCARlUw7L4tRD1KJNHU8FUHZdbet1Rver4NhsTvuiw/9Uk5CZ+jWIOPQxqE
chJloTShA3bi2sQdoxnAsPSiyupp0Uy4jH+9SCXxapJSOKtmwQS053OmM9IRoQCFFIhbYImpEesH
RLowPveDwrt5ZWKlQcAwBE8fnfMQv4WoLc+667aHyDlHgGI10D0HcShgngvolMo/rGMviSDo6+cK
LdN8HLsAiM6JLRVIzh0XupoTdaehXoqZSS67vzoeZfsiI9UO3ecHV1IAlCujijC6VX9R38ZiWh5r
/DIdVCzTGu3z7jwtCj0jJYaAorEhnk9jE4Eqt3EcxnzWEJ3bBk+5gkdVubuosw1Ywy7PsS0mVa7N
vfRRxgwNl8qgRpuEJbFGbBXBY8nwjylZWCAgq2CV8dHDyeiHAGAxiqb/z5sc9ZLmG3PHVkH2IzH0
oG5hOLOu6dBhm1L7Rd6iZr8JtDXY/kS2wq23fBFGL2G5zonYr49J0zCI7NCU+faMCOz4BVMA92ut
I2Sc1cSMtgYH21uZ/BnoMVxzmDQKjeplSbTze07/EpAPHK2IJTX6xDwMj2/OqmIDyIghow9ElapD
D+37Iv+IzmnAy3GQSpBUijYRohXNKWTGJgystxNq1raSZK4QVXBhYD76ZL9BApZ/5WLqAzU4i0D6
Gi1kk6n6eGILIJH/SVOgguvwxbQ5MxDzrC9UzOwLLgOhYmU/8/cZFa4Nnb3SoBxrS55ofXhXnyXl
xTflagSRIs3LDh62lZPRH3CGCkTWc/Ktr3jcZcILTFD8O8iGQTw2bILXsfe4CpLgT/+o3W+uqLI6
Q5J5VN8AQN1ILxHPOk1KRmzYMDcbYe1Xy72tNx0WD89mM5zFOuEEyoFJ3iwl+7UwzrdWg8uyr4AM
v5pq+zpbd5oEOGiBn3uW2tDcXvZ+rYTRbGB71iZkk8pxTLQfYnNoMRgU8Ob7o5JNdA0E8vlV8dxD
lSVtyiXr6hHGD0UZDW4/q0MUeZq1YK2+7Iq3+LuIWGhhc1hEKdMHa7M5kaT8oRhJj5y/dGsek+hm
bpWfQTZDrQQQa1HDoKtynWUUqn3bs/+rXOwy5VT3Gz0QUM6WvFiPlNJE5tZDsHroeHvP38HJR7eO
9grH5qOKURYmI2IJDGFvI5P9nTHvdOXRfx05cyjxeonMcGGB87ZI7pqAQ6gwIQw69GrerbPCBtiT
wcTL6W5l9Xdmrf/tv3qhavVhhRfw5/BcyjZCxXe6k0qqtSCQtVlGX0uoGVbvIFyxNWbDWtQXMW1L
Z5+I3tLjeZt/ycf/VvzbndLIiupFFeUDqODZKkvLhO0Q24eene55QhBZs86pU0xTbZAsLF1KusYA
WbVn0jkTLKDSLxvAk/ooUAiR4u7WrqbvOc/7H5cQfKW9QZELayhK0Uzz+b6hEu9qEfIUCicU+jb5
ogNEJQhoE0Nzi0UV89yzRxsI3DVFlOMXFBy0kPjj75UydE/wK7DL1XJ8gxgloruP16g45EfIZdTM
+CmY5X8wybxy1RnTFxtVqGjGIdfhQNvunDZKbup6fdgufpHoe8mNxOpPAqjtVi/YfGMj+yIHz/Ez
2cR3uaJ6ljl1XojKmNLGTSuDJE4V/CjFDisMZ5DdHhBsD68SBBZJgE2o6Y49toaIQQxL5AxIeJL6
pmN7mUC1pdolJfgCtU9bMPL+HWZj+ODeBD7jBpLmYCc/SUa6e/9X7lOjGDHHZ8jKBJSNYHemB1Pa
8V1aynjPMYO6uGwUqUNtbFhdeLRroL3B868sLkJyWS9ABvdmESamNAGpF/iMxH0pgEUwkwG9tlUt
iVQmcRWBAVVH+6EMDUkhHjXXSiH+7fUP21Iwl5LGDAE3XQju4cbhQFHKO6hzwr5nWBra3B0Eiu4n
MtKxTgf2hFptTseS/1KInYwPkNtFcfkUlnKbDeWE0dOk81NvpB4WMRuqSv4NQ2wwJm3+ljAQHBHy
a19xkv6Irohc7UFe7yos5zg8Nu3TqfzlV88aW7n1hoJVtkjWmlBEZWatIQR35JMyZzBiFEARD5hS
dmaB63W76kHWeAVrGX1VNIj1uhGjVCzNC3oht9JMW2xkAmFBPte/jDbjARYtq+nm4yxNXvb6BmwH
aUJpI3ykMMFeiKWWrS3kV3HTAESMtzrOBGjR5hgKRTV/G6kh96jXaIYEHJIEqagJ1dBaRIJmM2GW
GyuGwG29expztC8j39V3GqP7yQbmBFSATDcBTerqCdTik0xK1TkSFlXpzhYTlzL37FgMmCudN05v
QTRKsJDFpFFiIpYRiJPb0fPrwxCEZgZiRO0QmlfIf23sPVUhs2lGbPasH8B3vcz2vyEjc9b2RTxM
agdj8UfQ4zoS7Es5I387wGThqw8zc1Xns0ZeS+pWpsIMaic+uRCVYQaB1ZkbhMVDMH8XDnTjqimJ
I5oXnWgg+TeHO5iNMoAmSnOG2oOPj5+H+DPbwgyJ6fzhTn32OGknjohioD/T3Oc9RTgMeVDpycI0
MNk1wZq4hFiRUeKt/nyaBxRaUuJmXcEWVNRGMiWAp+huW6S3PIu9CDZf78elRrsQYVI6UQ2xGXsh
tuBZjzkKQwoX+W0SCq2MD/av2E4ycGjOa9opbFYBsYAHr2RTw+Tuk0DfXhEIxX+bWuf2eK9jZYQe
3ay4Glo9zvut1s+kMLDX21aqq1Da7CQVXZgFmhtkYjYfaTgrqJSZGBFtz7omtTER7KHzDysSDhPc
TRQrNO3tAu2n0GummswsCCPfi+nw5WMxEzCzofImD5rTxcHRaONFqtKaYOWCENNO+1UfjAjf76lB
rYRf1INI9xhI4KOrGy7umOIbHX/ShdGQl4N9oalNacclC9auzH5Nx3Wa8gzkddeKemdhlhgEKl//
5bJVjhRIt1qvCzSkL28qfmZxMrRsiAp2jbbJbPoTAiBjWxf8erFao7HJYgLWzGaMO+uNMoIlm1rD
F4rMGe4nOUbafirEUX5wcmtlqL2XryscVJh4jID6N7zoY56hSlVA/+YUAvw+gec3k4FE28z65VOd
/4CAjxBYgEUTHz7ELl6ehT+T8K416gHaBHzBF0nJZdujrZZXAuXATt8654eSbHo5I1SJNBO2/bq9
PlDFiG35ySxCyX4jarfUDNArOHSxRipjUxnLNo0VWb1GJtck/Szq76jA09/3p1c8yHMtIhIBJfj6
BolORWgkySpXn45VMQYzdhJdpMYwVwaniY7P2ccg3yQypCnLuhOCfdTS5eI9czl+UKAoR4bWznbV
bM4Qwufcn6ImvCSTatry12s9v0qvpyzgYpDGaOBE/BnORIzRQFqBdAt/H5DdulaVY7OwAcbmj/pd
ZqI1ZaBD9p0BfAYfDckE3Nrgus1+1GAwFk4Lqj9Q5vvJRaqH+o2quhmSuFZ5/gh9m6tRG82ttCCz
duMroW1bKCqYJINxrgTDpvNc/V5Nj1rh+lZjSuix4SVgqYCQF+2/Vf2zOFyAJ2aw/5SeogEmmOaZ
KJymFfL75aZtog2jOh0AYKYaDRtsx7SB6lnR7HvaZHqaNlmQLppgkyY8O5qxUTBnCcvd774yhaMl
y0s9xIyqRf7weBbRHi4S5atEyIVq2FvZPVOJza0cKXA72tohZmkkFJXsmSlu8LhnFA2Wbp290Bis
t48SrrttJw1l6NEkWuRu4NucUmTYPr45AgK/EIXhCYF//30WDQo5nw8TYcrvjDQb0Q8uyl/Di5RD
XxN7w65lmGtf2UxQNKmZZ/clBYbLVt1S/Lk3/EzklucQjTRMSS4q818vSGaXUnYkbQ6bEYIRHeLR
eRlbPRWXVm+hMWWA2bTc+DVqW52efICsK46h8U7/9pH/Va5a0qscM2/hbvN8rzuBTwafdPRs8lmA
0fp6lxeUBHdtBxFDXFfGghifgBQtrL2D6TkbB2Cy2y58T1e1ovkrrEVaE3hCrcpLree+tAc6V4qA
6Dkv8kCWzSvmLjCxD496Qvf/XxIxmeElLnZQAW6HT3hwFZDDJ2GVim48sjBXjiZxHi5DHT5hKfoF
75iMe4KZlVz+ulpUNwQCRjB9/n/VmKVs4Juldd2PgcQotSqU31syJgYH5k5DV2p63NbYz52TpZ1k
7ot69Vln+FsUK8Vmf4+1m5LS+R9OyD9Ml/KWOSZB4qcxPFg6U1lKQoYTPwuzpPI7iSFldhnd6MHS
SqN1MPW2ncxI89f8uZl2GksVqwJqZQysEBrLCeIiVgeqmr/qHI8P8n/cngI3fy3edt91Ttw2CY+C
/RdVVT5Jqz87UFN4BTLyONTHQ9lvrumsnncKvcb2jDSM5TlR7N/cdTswEggbz385QJdc9LblkYaG
8j717ItFoKao1lfPpH0lrasB6wYEaeH3jV9Fh97riv5p0aq74F/Ob0NDY11ejGWUGKCzyiTNiYOo
BZa6wWEJN3xYFh2Q1bpBG9+gFjHYDVAjBC1I52atE3qBw224XnKlctPPe5P+QjrFyde2faldP7TG
ua5+HQq4F0W+NQz5ThU3Er79RC7z5MrD1O0kmGFdeBomcIPToL1lRyMB3N0Mg9uvkiNAWp5Stpxe
Ok4mrXhfCYx2gk+5Zy92Tl79BSf5hebsRQDlmzscpZFpSpPjFvB+mSKuyeESLk8QcBpyHFwWYdXR
wSCnS3piPGyGsfOE0ZQ75vsaISePcrnVquVIXUnGDkd0iQzaajWDQONXOTmrFOIhCFOhn35cIkEE
pDgwl11QhC/Tj0gFoRXb60eyAeDbkom/z2DDFzeCe3+enMNN7JBcAtIzv/NQTthQb/xFGsZdLDBh
OtZouyPOZL3Yb5y1O5nYXjggMyLbfff87NoIk3ni4ig5nTu32Lc6ZGxuDbouoZR4UiKJ0hwvbb8w
DYe019WnyNoIa38TMEuKQOKWokBVp7MBsJdG/IrILlx+m5ignaRhig0g2EXl/wr07X5gmdjG6xIw
zJlpQv3ip4Yk148bMgP3mV7O3bLtk77xQa3l49fG76N8sN9s7r6PKfF5ettd9shjHWPHXKhqRc5L
bNtwDGYc4K1yPMTEL+ohC+8CsG/2N2wntmIc+E/t9egWJqdWYKQi5LvE/M+wKgQt1nV4C3Wi6DCB
ynTL6CQUneVfhaMB9X/iMUWfvwe6lKODKG2PbJHmN+U4yU53N9YJIFy5MmRe2a6BASiLuZTHHXLh
+G+2f7pKYNpeiz64uAo9UYqU0HLgs4qtz6vQf0EXMy38w0rbJhbUGh6z8VPVv7zgpWXazg7X5gSE
WTs311lCGel+iw+AVQWrEvOks8ZkIiuNzOswqlwpj06pkLkI8i3xXB8AL0Pln/pNj/OKTvSD9elU
Bk1ORPI3G7sdcceuOg67sEPK1Ianjl4M8GTIzFRPFnqgAFW93/grvSFTr148oBOZS4TX6o9hKq9G
nePSk9m3e21HqJGIPxJBDPLZY+6WZ0H9PEe05xsYjIk+fRF2cx8TNObV+cyiMjgXvYRq0cvInlTZ
0TprckbYKuqG+4L7C6krKX6229R8SraW6RD7k7xHE8xmoQIqvQoJloB5eHjqXFBaiDtHPhSibMhj
HnUZ5Wfy7XVNi0gS6iuJecxrAB0bfIv3tDTNowaSpm/bPRFNOTeYmcqpHY0tXZAjSIVc2G+I10jW
4jpZs58sNf2UowaNXjUCpxSQO1zvGNu0JyoA6H8hHwZ4w+P4bM/Zi2mbiLw+/XGfs7b6rtV0gTob
w0UWJo6br8YIKPuQYKbl8tmo7xcfffN3cUJVOJaBYdDSVDm14sBrpQxs4cQf1FE1rhAqc8TjgoEz
7qf00D/cuwR1hG046NdGfR53LrNZ1ZsAAED/viQzKVmstwBZofVhvK1xGGp/JjrMUWnIx1f+GfFl
86768Ubhcjp91UY5uTli60xhazmsoEQmZSlpjCvjborcjRzx+oUsM6ueQZg020NIIGNJjIlQhCHG
ZOjvCtS0M0jCeZ/p6LYyzTAyqLzOmLq8aoFH2tSzziM6Ggd8K9wdJ27ZcDX1RiL5VAPRZsv6/Xun
AujfZUv2ICynfTJ1Js7kP2PeaWqfCMD1YtnAixR5PI4A4Apr3kSlcMoju+akjST25yRcWpdJ6SMJ
R5XnyIf2EFkvsIxOw2ekkslsu4/+mBWLW7CXj6rMtZq4Xf3mmqYYaHlywzCyooze8SjGtod7yI8I
4KO4JABByTSxGlwInyXFPD2KnfDVON350msnwz/cUgqn1AD1UviyZ2Y4crjRipcFjV8CkRkTDfP6
WfMJMQG9xICMrGZBt32aF29TOJ+77z6w70AIjULd4JBqpPwX7rbpF4zqPMQO9T/f4NxFgZ1Ogsh8
xxHwckBliUHI989k1hPWUtcYpUUwDWnKKvIH2zk/NbMzAAeNhMnfmosefp+DzM5923QBekztBEI5
o2te31+hb8tYh6yG9wdIWMJ+GQmAbdIrELuWiPmx6hFcw0AeFs+RuSGier7Atwh2v9B+E+k02TXq
82uNmsVTTHmqBCCGWjnwD1+u5gHRR8dBMMdD0CB2OTfhf937+gulTQlqV3GVorppcf9ftAL8V/wZ
oHZxkO/piJ4x84vMI85txRZHGNx7+8bYXfbNZQsquLbamGrK4tvny6upAoGv+MMXTVdfkkGtpvvg
gpXPdc02GDulCSBYy4Urg4LVt9XGKvq+7sNE0CRGy5m4Skowk8YhiCxsekQv37nVgVU2BqgkBXq5
uAFxSY1o1GqOb50RUo1A35RkOIdCHLFTRxvXCPj2DXCO2TTXWOWbDV2OzVk/qCwMaUlxS+w2/WIA
yLC5kpAQv+KEEsATAQCB0JmRZJjQ3p2FsphVZRD/zAKrGJ8zE+ZI4TdiqYgF+/ckqu2G0oJt4pRj
r1qeQ1x1FxjJSl1LTILXKCQMd42X9/8GP3KOJDny25Z+T2c/Ug+LfIafpYII2H9TVbPAWzLSL7DG
K00Yo3O5jaiqNbpkd/7xmyLX69cddrM8PcPgtME3HGjvpVbaqOyffypkP4rWrask5jus+rfL0YuF
BSF6xgxmWfGC/8+YKcqFQZzoyNfuCQRLJ3xNVXlEQdFSJWn96EGBJN/g1KEfad6lVabHaU8bQkAq
fssbwtNbHtFIQFm8SAzMZev2x7tIdC7DTEcBI6od6m6VDzXzES2XvC5f61jTH2ZeIDSNbZf041s6
dzPbigzVx9UWFtz6iRi4VnMQ8zormxvq1gASwWuiEhUkl1wDuHTwrVKQvtfRPOLmNLM1zdkFooJw
wGaawKGUj/zB6G7WzMKYNpNtrNYTcJ29MAUTpsNRV/2LCucT0rN8P4xvxoCh3YtDpeNPdwMDO1WH
ncNfx5TmpFc00Ixf97MHpGGyUj0HWH7ay6NL476tteKQFQhGGbuSVS1CZKeqqAmA7BEylOhKbMhI
YUk8yIPQdFbbjLdmj3OjKshoYI4BpYY0hVvjE7iqX4su36leh5d9QCKfz3OYtofM6OzfJ1o2+evU
2FjDmGkCGEP74D77tUzjMK9SrmcxmH6rGw2DQHtnMhwqZXHizZLZbEp+zQ0+WDDN2o1GgewOXDZk
ewLSQwO6dqrIZvj4IhuIbBjvuZkMj0c4N8VTaIwmL4pqoeMXhb0u0vTws1yUF8ItIqv2XFlE1Qdw
OAUw9TNRRyMtYL5wiqxlVM0plMNc59lIOVdDnvayXY6nmN8qGVmJbmVGkmamUPGwC0hQq9mRH/J8
5D4wp4Y4oUWllkTX3qN2xbcEcAqSj2OT7a/Dq2cAwlkaB54Be8h7+X0tg+Z7vnnvUG3+IOsGpAKV
EQ4IOgQnSsz3W4aUKauUCFQQF4xRpP+Dk2LFbPu7+AFz5cCq6GazeF1Ing7CQa6tG33a91NExI9f
6kSwlmlqvRttTBmaq5GvlYPR9vNNZcCoA/+PuqyB0IBG9Bc4+QRkjmRXz4nbSj/fEhZwqY4MOjAk
r96mXbkD53X4Ui3ct9uII2t8op2m+vmu2unzHl25FAKlwc2DW9yTo/vvxwTF6YUKf++YHQpGkw4c
h21MwNd8CMkiexNgoRPPFaY1tdNIr77ctVaC0jwjnsO06TcTvMsqjgaEttAx8/DAUBL/6hW/hdta
2oULGLC9wFRGBwADTi44J6NN7pgUuoqEOOM9Ww2tC/iN6y8Zc5To+i21kUavFuoFiB4/oj7dc32i
N3ob/mT6bCeqTjxfRWiOxCPJBZLT2TnmBrBF/wKWD1wqYmuslqLBiycApYb6DunwAgb+nfcV1ag4
1I24Wqu4gCvk/2x2uBoKu7ia25XxuyOY1QfpO3M2ZCNKW7M3ILBHVxztNR/JqwRNi3cmJuKZH+1X
EeL6lyiATvla5wzG8bLI2KSHATwEcHfIVO0A8RMsmQWAH4sCPa+nz5Nh8Dy0jDYlLixwlAaez5cM
JeAcyKACOf/T3pC8Am+z0HN/6Eef0N9Zxw/WFbO5lvGgXnFYjz30DhjrYvxEHwYtdJTs6oi7PckH
HLj4Ec/fRXLGjxJld9OmUk6Ie1VtlLcunxA5LWtw6VCwEx2TtwjoBPwOwyfoC/bhtQwvSqJqvdsw
moKA0wp2V45ORWHCOG61uUjQDWzEk58iHCmPaJEnGV37mnhgGkUVblkGUXH43EJPgG5ypQ5xM4dG
3jXcgTb78a42u1CAEeTQscjT+W0W3zMuA4UR5Er/i0oJpPSsAw/XgftlVcAcx2+F0vc3JumldH4+
f9CqB2kX1K+zjO88d8T78js/yFJGkOIiyyuQ+ohVqg9PHg2BO8OT2PeGeJNIFr16YspTDp86/n7Z
YUwAdkUPA9lKO4ZCtLb5eFmC4YAzdk1YWD3krv69gkyX7w3y0Jl7TGspXtFP8Fu58Jdp2DplXMlW
+IMNHGkcu01CYvYv3mz70lFd5LunywSarD9A6+/LHe0nXXmVeakpEDCh7psX9HhIgHTjqHt0E5bj
V3bo8m79em5DAWGZ1kjNx3YG58YIN5UnQJbM/VwUhA2WYqF6pIRKAJiXTM0bRPRBwV8ssAyyVdrW
qSvUxUXePuZDFWeS6HXGnQUwJvxRsvpZ8NRnoxAR5zjJrWGouDHyubEKJHhvnZaKVrpDSZFb/HkJ
9pamig8xdUmRRecxXOSKBcbDR2i8MgBfoVMrvj92bFm9KNXErYHPNJkb4ia+D0GHVXCN1+oxt2+f
+V+saspeHVp7JzfjcYqoRyWz/3qychRgk5iE5eXzTTDi7e5g2ZDDJMF49BoRphNjkQiEZBgt2ANN
JNKIdNlj2X2CvbmzwpwrCAts7f9mlihDaQIcTbm0Qk8Vqx9lNAFoQRycN5y5hF6oEMC95VgStrEO
D0oJTzKAkU0RNJqZpZbrdG1LlaieUa0GfTNamEHqGJduvyCOc8bX6VN841szoDcve1N8zwLn/HhN
2t71MIGI9zujCDA/knTiSWOykXElPAgI0EPCFML2Brue4yptf0dX2lk9iMv50wiNyAsfnfcLA3MD
Z3ELfFHJgfHL88oOf4ZhcH5E90gWn1lC+3OWCQo2JinQy4gH+pipdNpj1+u9jOmOtK5ptnSl4T9k
ZZEhQABvMcwxNVPWAlhyG6DyLpnlsyaXxKn8+TDaIsoUFPhrHo/RfuxEarxTSUO0vhF9iJBOfwWx
qsoqJ9cW2J/33qadEb5E/e0PVjNW9SZOUlt+s4l6viVEDDB/a8+q0mF+jaDOQzzUgCqpQUYFOf6r
S+SpLieQB6Yz5VPdsTNfoMAmzEuu3TDhlgg1qBI/u/ZK+b/tI409knaK25jCOmXTEZ3H8vFz+M8E
GIpNoaNYoGBtDeqCOc4oWvZujHysk6DivlmHoWv6Zcb68gp/ktd1/IhricwAFS4IurtSK1pydpgQ
tMzIM7ONxXjdBsQyylr8rAWFX+Juad7iYZqqM2c6ke/WRDr7tr6UeFUIORVmSMFbOS03GDmqh98Y
5DRMTwD1MaFIHpd1qSYF1tYo8EVRnNkQKG4sgg8VttFJ3hVyRvOxE/kl1StDMSYTDBy2kBKBNFgc
JzNYprePUXBI7j5ZYATMsPoO/japn/yaWIl1LnZXvUnhnu0qQ3nsnk1ymLCzFWpmSaEj3jgV+ePn
NGXBPkNN/SN3jkGpGxv9w0OKzoNfvULres836sz4+XnMUhv2gLY0XGqfTFr9UcnAvXuRI6UN6ZM6
nTg0j4qj4eMsaAxrhDFbHjzQ+etDxCBC/2jepw+nnv5z+/CQNl5j1iscIc+NyRhfEQIiJ1osPwbb
JyghXBD5kziIY2H1uv5X8APHvzE7CPxMWlAYJ9MDT0YVqSLxfzmCB5sa+gu2OGAC9iwQZRHaoseW
Eh1ldwpN01uD4s4mG8Xjfw7gj87dnNoVCVk8lirY076JijvtMcw3WzbcHdwv885436Aw1dg3RQAr
0STe0f8z2i4yzGhXZfk6ImEdqiByjU3Q0tmu9V6cdlfyQ+ENNXc7ulq4QPFFucQKBkC2tGfOGFmA
6MnmF5d5T0Pm/bZcdh1RB4ZtNQl55klCOw7YSAXWMqjgMFSFA0mTXeZDsCExIJeuwaiaFRHTq+6y
0XTrw9wVhgttn751tYMEtyAM/AP5hg42Aqmse3Wv9/0crb8rWmwhJorjXdWlpsLGAajSI5S9gyCi
no7M5g52jI7rcCgNTSjVtwJjjB4br4nKkkH4rtDp8LCoHSNwnZ6X4ulGHhZT01eNYuY89DeTYUAK
dK45X0DAhLk3HNmiDFLguPHs0DABGy1NMKfwrjsZHLkr8bRQZbAl7cUz8CVRs6gwsH1p3jjkLgCS
OACbwf8Qe4dVR7MRg31dgiKkLiYXLdr+rq5Z4akZaFEZJuuBsMSiBhAknq5yxV/IA2WvAzYVz+Ur
RFAlfZioQ0YwY0CcBQEdajxQn94rHTzk8qZ8eIrhPZ8tGVbKLEltDEFAfnXwAcjBh8qvSByP6s61
cd7RjR0u6wM5OkCmXiTt0xATYodbXXY1Kxw96unovb3gbn+oxZVizbZvBY1aDSLP+rxLzoAWzU0Z
P5bNtU1BMg0evEAqeIUtD62vOZE8bFYt0P2GJoKn0b+1wnWhoEsVRT1tKw2iAL5JS0EozADvzITW
edzqOvmFlEjGBtAOjadZo76g53JhP7FFnV0kFgSxtgXBwQanzLL04tJK0x5qW3+UWinRkGjGfBmi
lDXwXjw4HXPLuTQhwZO/SYQ5+Au4tAADev0h5Hy8m7Q8Wu2ODtyihnVrVDTHwQ3q7AtaK2fBu68e
iHpP4EyYtGq++2kvrRgJ/C/e3ZG+IN1Oe6GI+aIdmpmBgSeTCqv6X9ZEbetOODdtOWfVrQdbCjsY
IcgyBMURfQFgVW6eX1wYtrHX3Ng3MZaOl5st4tDUu9P8NaDEcjyQgS50eCKqRXuqre5tWsATiOlv
NggUh7eTSU2MsHk7EVTha7Di+FgjkzEEl9ezEdRDw0sVRLCn18uttjNblmxjS8D8BrZ32E2z+4WS
LUnvDDLWbBqLHtzcULNRQj8WrddK818QchJhxMpOwOeZYIRv2JUEdC+OS8s2lPowlWwN81p4agTA
Vb9TFe6E7r74ryDfVAEIdXSylp85eBzSiP8p+bp7LinwblebeW1lLckBo9K+5hnpQWC1BAl9dAWb
Lthv3wwZ7LU7YosUG/vBSmmhtULlu+uaglVFgnq86SQc5uxL6T4vDh8O9zeWnfDeqSrb/bk6rU9x
uLFi8p/D1jCmOsNGYOchy7fiV495P8b2+WIqajwFVf1gEGRH9kJnwA9J8uL4fSZokScLyYGmA221
mmivsd6ddR22BSqMwqCfGre0McGjUTcN98kq0cl8Fu/fRzWf8Cl2G1pWPXxspmI6i9pL95wobcYz
dyy2w0AHMQOsrQ4UMMxQ28/JlsndbDzW0hQtHOKGUz79gajok4jyfnNj8PY4KFL+ejIdpSHG6LIg
xBSwbNaQRn3bU7K+RwfliEC8iu1VaODUx+HQnm2p3u52Ktc/fKCrF36yR+AdLBjbIiWkvOvzGyys
dzv2RK2NfPLIxoNsfGsu18Rzwxab5+cvgCQ0G6BIJf0Qm5BQR6g/1dWBPKvFv9Mc1eRmhpsMy/9p
Brvgaw6tKZkeuzM+/vuwZdlRu5J52nAHGNk68lJeM1+yPZ8LzIfx9KgEK0b8C9YbjMQzPHjie2e2
UI+cOBNGnCuEZqHbdGyWJs1iavuwDlx0KD3luQTQPu7wfiddkGdVbNl2wibBSbjVXwTPLNdT2/up
Ns3AzCcfJCv2FruLik6DxmmBPNSHKItgHA7q/k6TKlJlTnKcYQB0rsgjx+KVal+A5aqFP1Wy9ieJ
W2qf3xe+dYLMBcWPh6geXLNtLTwdJs3X58Fvc1PZLS5r+Fx4Jrgq3fuIi2XGWhwCsj0AKF2j8ZiQ
w3V8BCCEIylG/Wzst3gxJtGBqSbaAF4khn/GuO0s4KSaBedWRdkRQCT5LkL72EBmJcX6vGRelTJ6
WhfsHh9DGDsbtnXaRqDrYMDqxpT6Oumt1IxEo5xBFc1d/HqbJ/Yjd70MtaHGrV3Ob3YCVXISzX1v
q2cmab4GJ+vKi+YmLU7JJ5BXFs23PbZM5i/lXVUbUwDI84EPex+B2q45L/0AaEMMCRzp3e+lD9vY
Vt0B8XWLCz19a2dAyP6LNJKWaVTJLnZ+vN5/f+6GfEQNwGENqVI2Nru9HEI9Pf0cSQo7pUzel87X
v5bqxJABVx8H8Ug/4WIePHJZf2uKlzKN89NNMevS3IiBv3Wj20esi2Mq8/xP1jdep/xlqlQLA4uD
syEQVwb/9EZ3Mg2YYf+TbfS7r0QMTVxCRYkm7y9RB0tPRYveWUBEvnbOdPHD8jWYSxNNgbc1glul
Og8+EELJs+UzlBfZ60QO9Ze2n/8H0QXgXElkopM3g+sso7gHLj9t/XU6PFVXsSYI2OW0uaMT/dnA
c1zfroJWeCMwFEilPMh2HqFhL6YB0k+Bu35xlicCaAcZZz4Lcs86fE/6cbZIjTGG+lmKzhL7rNOn
rD9e9Jmav8VRog5B1ucCnJHByJIpHgzRAmB7ziLuoJwPtV7oSaDbJPGpfsbYId+zXqGTLQ6shUzq
pQssrYL16QIEL7iI9ARPQbVVfof+Qv/7Bwb0YVZE6hHA6mzo4jzcoQLDeHOtmNvcEP2vINLiu4+c
PlWJkEd3vq0uTDqUz9x4ATlw75RO4xgKxLPhWIdAg+qkmKEGqsew/xhKXUqddJB/t0eld4Lyl3ev
alsbdvtm/j1hdTFlfzmu2B4iLOUPDsfI2MZ/pVlyCzYEpZjy1mHqwxZaRsxtSUrsXZygPElSmDq9
KNpa1CLdE+ft2sgoEH0SSibKrY/7uUUFqNWaXU1ZFah6n38mLtZhInH2YJwdju3Yhx6OoL33NdSd
Iqdoz1oig7EZGpcyqOpZrEu1BuOAKs7E7d+EfUqn0yP/8b5rur5Nz9DNykJ5kpDbd8TtLJ57dBgo
flmyRH+iRq6cT+qoewbkGDuUTNnyJ0JAGEpEU0wibFAt10GiwyhEa/i/aTklu45zHpDsjApEmh97
oU6oz0u3tG3qxd2uwLHUlQdFEgiyigOPONH6CRZAst3T5n+I5AI0ddsyO/bpwD49eRaXt38V/yP1
bRKfYfCYgoCSM5+QWroozNq65wogeb7n8eMJm8vrXrK9gkIGPh41GOtZgC55O6JEjRbUEiS8Zult
suODKEvC/wsHCzVWbC3CrHC8BMA5sTeORYJkr4oiG5b8dlFA2MTITyrrQUXw6tyAXZ7YMw84OQFB
i5FzzlZk0qSg8nTR/dZRhEF4igifvLr/wwp0Yg4Kg4xP8lo3seBCDhNQ8BwxMTXTNhN81lnCe2hX
boJX37FSd8673eDDbe/YEchKTLerD5rl03RQ83S+g0c2e08mKtr4TSDWed8Q0fMueLqTKiRiFGyE
4LpVe1DY+Vk/Yyswxj7kJ4wfLf0C7kIeRv2V0ce1xVcDMZz2OwCNWKVZAm0Jiq+BzkM2qZ+DFmla
4zaqiyjnCiNNcfOgBthg0NuwHWW0FGMMpBokEJGYlf8+bXpFRIuzRXULxd+LgHsT2Lsh8ZT6dZB6
vyDddzyI5X3xqazp1j19oK1s3FzfDQ8SCFobMcUadVmldClQhdiE3krJhavs1Wmor7znXRTtZt+r
+qg/e23b2+/l8k25VyqrSJvUS6wADoIuoD4fFB+JiMvHs4JZ55TV7aViVdJVdIQOwpf7D2Z+ZnDj
aEfvLLVxApNGqBIdWU6xHBpLdSXT+JVGMPFhvsc8/JeJGYkBZKE0hxCeaS6Hm55V1X45ySZtyy5j
p8GPnkUll05Qyp2HdoRqY3hkIl+70/k07A+h4+/kD3HdYTaU129X0Kc4JWIokEaLRNxXDME2zvo2
hlTQyoZEtwzyhZrYMPUqJhh1mmYg+l5N9oqg9hIU2clsXN1ymJME4DeQXCLw/Kkvc2KHMPKs01bQ
k7v8cpyTo/CfgfHEr7j8w1lznLWSAt1LZCgK2WCZFU7+d3gDwKBF6KAKZnuXcG+UIvc0n1v9jPgg
yymJhF3MPt+J0w21GfOHI06INqp16c0mlKyO9M+2xN0UNWKigGeGjIErPZYX2xbPqf2D5SfLZjGc
yhdU5LA0AQpZv1BYl6CdY9sA4ZuHUlEmExSmyV3vU/LjdjwsdF0jdVjehwIqrtxHB9UhiZ4UdVB0
BFWWqghi/BYv/uxMARFIc31q0XT+aC5Y/kUt/VQ74/QrY7D4kBLlRJ8LzKVAzH+lx3Cfy+XjrkPR
6oJUu6BYOtb0IY/kWL/mUwZHVsWTSAAZdeob8Ws6MK/6YC0kW3S+vNJuLn53bQ3iR85yLeC8pKbm
AGXW+eQl98U7YB6kgl4hTNIlZX5lftFPgM/s4+vMOV2M6CpAueYhIU6pOCNf3bJJLRKkTHgjXXO6
/44Ei8Ns88RTOS3x/mCreWxup8J6xMGjcnkRFyBvPaCNn8DC8AF2w4O+Pxflu8K4HEZvDhIMcXlW
2qiHt4VolmtpSM/M4y0491DY9JPVPWFS0guuE/JYuH5mnodt/kueDNGipwERGazG5N8fLqmgfbnc
VdE8bvYO6fk2QnhR+UcMkVPNovRpy2jy4vzndhphJdwZ8JRzEN+2XS3AsWoxzjJPjuUNYgTGuGt2
1jQn6qFZN9asiM8hUoh5fLgVeJ/RjgF1wxbSuuBBQqGyWJKxFdsfbtrF8FNT/FkjU+iTOn14u6GS
4KAt9e0IRcX2sUWmtVjLtsAsmHfXfdNF8sjEQtB4EYYqxefw0Qh3+7WNfR0pe0GTPYU7Re3Ewm03
TVrl2QYqz1Jb12lHuRl8N0bEYCiBRZExF8W8BgEgkJjv5FHbafBt54sIhUG1Y9XT0b53RZLMRVkA
OJqKUdO18reOTjHx6MwN6RGvFcRIf1rPTxwiTBffSsRkyyvFAlSNCJT0JEGN7+Q3aco3NYGEEOtt
kVPN7GxF5LxdzHZbsa2NCxM+M+0vDzmazQjJI5ZgUq+UUoMi+iucClbak7ZNieryT/n0DDEUwarO
WQygmPOYjJHbQRNBvWEkHo19qY4ZUaUCkN81yNkosDnCmqmez7X5ogScc6/odQnoplo/n7UM4tXn
VTo01PjnHLqvEsGDScBVipxhQ3ptgMyS7vxDn+fYYWTAlXW1G4utkqe7f//ng4+7fFLl759JNZbQ
gh1t9P8iy8qtxFB528kiLQRr/0kDVaoOQtsdxPYXaRWqIN59IX5s5cgTwtQw+CXwASeCsiQCZGWH
mg3BSd5V/YlwIhKPVzICxUOs1DxxjM0990scn929oCtUifYd4WEwjxyr7/smY1V3EXwGATO4iv6+
Xx5tk98G6Xoc+sM7s2MHQGIX1bopZt+8e6UEAkK+2tDloqzfieutN0gevM+sPPCvwc6sDIPgb1cn
wYgn/2yBUrhmMivf4dHAIIZKtI2eqHly8Gh3h4pbprFqH4TjqLwU3bnPMz0QY2AnDhNPY0i997tV
OkrQKIXOkJDrWX/K2YXgw5CsydvZJELyW8y5g14CeP6KjQgx1ORp1riOycZco/4L3wNFfcuaTXWa
jwyI/NyaM8+1zXNF3hqRI5TJ0ezMRH4kSiYbSmp4fMfSx1lxTzizJJLJGhWsIY3+NtAH7SpOk11e
Afxsu93wPfXVU8158UaBYP+t1hM2aolZP+Yqmi8gU0KWArpi0CND2Mwdma6HbYQJQm2qdJhU11Rr
lLO4aR/euNqHJ2N+aWQDs3+ilXuRktlIraLEMDJz67WohMBGPOVjXk8fhymkH7KsfIbaRqo41sQB
W53xS5GDWbc9qc8Yp0L8aDT9T4iXlz6SF883E9ZEz76NtySwNFWk3KYhudRQXWME4wHaNUnLPWEJ
zMS7/+VdPwlInmjig8aMZoy0f0UUaABQ41T3vSVADD/4OmBdbTETJraLl4WZ5YVv6PEy5APpTbqQ
rpW5JDMV4NBt9IzcXz+2F2XfXE5HhZ0vFacDssCDFUgn9XgxJAawAQmr1/grVm22+EX38lGc5xHI
RZAXFwIukcKvABxCRMe35GRyvjtKMciUJFMXlz3wF+TecP8vKocSWnOy8THTwFgBG03m/8Lc0y4e
aAhTAVH16NFCcxYu0M00nnAVfU5EK/ZVRkYXSNhU/FrOX0Oq+MBaFR0fWObjC5X1VgK3pp+Y6vOo
yWzM7MaHNw/5IrPQ4A9LVFA//6RwC5psntfH8BXUlDPlsMj4HDPEV/HZaHQcA4MkaNVS/UGcbEO+
tgnSsHM1UO/lukD2xC61LDlcGZifib2wAQKP3K+soznqLNDYLfJn1BccZtSXGz9gWUTyH58nYqxU
8xZsA2PP4Y9ibw4eCUrljK7bKRVFMp72DelvdlyU6ZLtFR3UtHgJe2g+1sIamFzyqfuI/5h4gIvn
98UZD715vFZLXQc8Gz2ZNxwYWy4ApVN3AsDQ20+ctTY0VCjeKPMvszRWsEWS+DKlw2nEdmMo3bxy
Bw9cJgODNMQAQmMVuc70V3+p+lbUCF6AZakFBNuncVCB6nJuDChdncjwMCAETiL+Qnwn5xtXyyst
Owk4eh6qXyCILASYD461cB/8DDuDRTQkYJcPoOHs2n8GtKprwUfdnfIWxAfHk8JDxCoHyPaLB2RG
zgNl9B9wuFZq+rfKp1Yrfmfdjcxj1+ZRYXFQXo4FOn2bgXypOjIgdZ6GI0w9+ppkhjyvVPUlCxxF
wsywcGAAIq3ykbwSvIkC2Vpb6du+xfyZp4dGwHI4KL8PIKF+ixelJ9ERoKjbO7jy4yjudj+gI7EW
E8uMvXJzhOx+UrS/FZ51nx9o37guXvBYX1V8S/jPGLzQTvOiY+psk4QTPBXAVic41HaB/CSnRqWB
vPJQNAHTdVh8L0FoKHAq+7iccpWJUW1mzD5ZoOFKHRz812meKV0jxGJCrCiAsZNgzERSj7yfMMCx
po/ydYcTXyzu08P0Z6TQfOoYkwf5+Hevp/uB0D1C2awIgvDn4b0E5qamRsIPyvA7BRshLQsoUPIl
Pz4PTbpRqVVZP8w+MOsiNLY6DH4DKNkup00XL7ZGq2h8At2vdQToFNU5MqupfpSVHs9tlaJXDVTt
BIdFdxdIgBFXFyKG90RkR8pMzsE+ir6ETiFERTGBsLvbLeMRRJbllFNKQSKvq6LQ7mrJKLpQZ1jQ
0ks2SjYAXQfg7q++xOrXoo5lQLZNx+yeE1+ZZTWilXLamMOz47bmQe0Gqc+kLzpiR3FWkxYsbhXa
oIVdtFRhZhm+OWHq8Q+nw3PFsdxYaKxf3z97/+hYQlKoK9L8OEybOmOlgKrpd+HoAjvr1VDZSvbE
bcJieq7kk43No19ebhmq+D4yMIpG8pI+793aTbfNLSSz5L0RtiAsk5/24aWXLwZJrcXCjqbDmXMq
rT22h7TrpMrOr/g4EFWeCLH491c7D6WCZp337mht9GYAUbBhv0sHb27qvAbFilslWwNrF4YtP5NZ
kJKe+TD3gktV2OJS7Bobqt/Fz+JVU8DoIvkrXkpYULUxr3s0k4riOitbDLTLXarFQriGPKc77bC2
ikDSG+k7HF9X06gyfa8V3zD9yb/mAC56Gsg8G/rSGsN6D1rOjVns5kOMLLfxDeDm9oFe09pAOJ/L
dUh7LWXrrn9DvhtnfLiEopWf7axgPTQsq4K7UXC28hc8p1R9DhDSTjF0C9c5SkpO9VhCbbxdM2UT
4qkfRjmpmhhBd5kmQxs2fJhKiVWfQPLe3hQOWIFbSAvXw8bOJBw/uf4nwipzxvQhbJTdQjBawjmA
CQ5lAqI5c297YQ+OUp52MrYoUsTU7RSk1Hr5UB49BHT3W9f2gjNEN7cpktp53TQ7a784jiNm7yQA
XGTg50OGgOfX2mmKxJUlng6EQtEKNR4pPefaihM0hUxniXXOqtAMILRpdnND7IoAxgiuH85la1WX
iYmKyeTwmRiaPDp0b0CX58zy/Wx83c8r8aDEsfVXXUG5bmQq1xZ8ZMEOOz/uMkpPeOICEac0z7C+
Z1+YjY91imW2M974LZIqCTeRvEFxHkUfAirdvi0V42oJ8MZe7qSdJ1LxKE2pAqBRN8V13VzsHuWU
RKdwQEwPGc4NPwE4PpMYUAtGhpT8a9Js9Ov86oZbrYu+ZIlktkJba8OZnH93bqIAmj0xkWxvFyeA
CaTqZ1LdJi72oSm6t9DnUxacRh+sqS2PWPoUKsJnfMwQAakJFsJ/kNd5J8NJZpCgVoSV0WrHqYGM
+VDQw15KQ4K5Jyxj/pc23ahVUYCjLoBuGEJb32x13PUpFmrxoqLPOuwo8Xmwo27oAlg9KIkjuj7S
wLid4YokkBCuoraAaU+GW8iuNq19wvy5uNMh0Kuctjvq4MFmjZMLKKxxhXqqxLxJuilcRbxnaHo9
bbb50u+QWIasWtR4LJ9Ix/qMu/VMBXMRitG96YJgNlbZwx8QPUCQyIUXTuurgdJ3USdI7vZr8ACv
Ds8dvr/sPZW0pvql7aIgmzmF8RL3XDtNar5QCaflAsG/NY1Qn98EcYQtajY3ixTw0HBX3a879Z8c
a5Op22htXsW9UcQRfh6aWCQ2U8NrO+F+i5RKzNrGbWI/p8LEXg1LG9R1ZrtnRhhIn78K6OsTcv02
m6KTA+CoZSNt6xe9Y8wD2R393Don8IMVF2GQBzW3pB7T5YDV6pV29VQ4dNBoM8ZceNdTVdW6/b2T
2hMpY+Bgoq+kCoUHOOxtsizayViXVLrBSB7z0Glo1lrPMfX/SC53X8Bi+g7veOILyGLgvGPaNx83
emyhucKhHvxIXKEcYSyznKlIBTlpz7LLAgL4Yer9vEh1vl93eOEF30qs16aIyb53sU0ZVQhWxPlV
F86aallMgLlD9UzDTkomOkAJdiXkPtWUGmxZFH8ppzGLnEX3xNN175ivbRoKJ7pfhuwKGjbNu75y
TW9VzRmI2bfLPgGvqgQOw3pBqJBuyynY29L2MXEYNWa2FCWi/0WntU/MTTBSmmgNVNjDapi7ooH5
3F19pV11cj/yZmUQ0Uv9pAlPwES8y9UYN7knU2A5mJikzKd/u1omKmcyMzbMGtVrJY+X4/o9DaAK
YWlORFrKIRVaP10hG+Ifbh9hEUoOrcqLjUPdXJgIM4+WwbvKXF3AEcC1bbefKlXHp2okkE6xSRGE
+GSqijmBFrV3tY9k0JUR5tXfvzTt4kMWXpp5RFKi62yZ+mrF/mmALaw7JScbTYm3RS/hlSvC+rUf
bQYeTU4ryUvcpDYijgV8U9AUTezHbDOXar8Kk52NyCymy0yUOVu03F42KYeQK0gnv90lTnKcIuB+
voA8zPp6W0rQJ2Hgzhz5DUUHTq7T1TElAbtwGp/HXYepE1zuO68tqBxGrGTo4MPplufARKkbprsO
3SD23dBLW4jUw3U7OkSw/Qnx9i+xSUfuolyIG81TYKfuSfjYMEDpMJ5JoAF+zQvImjpK6UPoypg4
NtDsFXtLof+xlDVlV9muNqQ/i/D5FBf45lmRkb5RLuJXGvKTSRq6b/UbzV8JVQje1zQVR/3SsaPX
uSywbfPzk37u2IecilNx87vj7JzGBa6/HI1T9puQdTEzYdxIbWEG6VL/9Uj5H8hszooiHOodR/aK
t1aj8f6y+wbEC/A6JvEqz/8DoJFke8mhD2NefKPUNdvsQqZT7S/IQIyXHccG/GcDUIPW36NIIY8q
tm4EeINSClmxPpfWVcvZ0dJcH3mNgE6A106znRF0l50PBnybKdsuLTez2DqRvzxE0WwFTdgvhZrN
V4tAzAPQZfgdn+zx4/hDOG7W/oPfJul1sN7FoCCyTMDb8fG5vFxsxKXEzFpXbKghYSsnN0l4oTB9
acpAve9KSRICVGwm37JtzGt3Xgj45/i+4HWcuZbhwkgBc8whQt4bnN9Ow00B9RjvJdmAFK+1xBgX
elZhSwoaKxUDNdwJW2CgoRSt5natOJgtgKql3HeggeOgvzpi9nw5ish2F8U7viK9OmaiFmZ1Pj9E
NPZ7eRMt67FOxCRrUZA8gX1V8V9fZhcmhY/AGgL3SUS99//ByYcR9P9/EDU3xTWMBXaf7JZuFK55
93DA5DBpmXWr6es5K2zB7kdLrOc1Pb9Dt0I4k5JdKd4XO6zbYI5+Q5EZyP/53cWMedSJmSPZubXO
jQc2HZT6orkeMfmXc1ELgki7T7VDeY0YcanuMvbT9+gGV1/r7OxIGW4VLHFEmLG84nDhqecPKWa9
HI57dfaG88YuOuVPLeGHowMv3lDULYHfJyTAaHsn4k0qyP0k7eR2SrLiR46y92jobLtpVA8AoesH
vQ65Ls7xamCelubBT06tCdWyP6499bKEuGWl7e0MQux7zLJVnq7oaPMmb2fGxIcY072B9Y+zrI09
d9ZHnail/6eJVnYFBTRmqSVUgiJ+aMElLN4Waj+vSa6H6+Q/4mD+VLw0tynwT2CG85GxOPMLHDPm
MhRb3l0v5xyiQh2Wp0zkkIxaaFW7aqy6LxxQU5fVIjH5ICrrz9r73+xatX8YQ42CQqx0T5YcWiMC
juQlZ1UVZZlZ2kZ27QWe698QGUpB2NgRI420qHdm78qo9i+QznUhpKL8MyaHnwlpDSGCIjxegvwy
VTV4nPXoH+36c2n8HmWWjBmJI8XgaeChMoEq02LPHUUa2fKDMt4tvRxo8840xcD4RNZdGHLIhPNi
WSItJPzyPa9W9lVApWmr70JC2NT+2WPubl7tUyygkeffaQ6UAlzv5LOMdPbZpDEiJ8Gah/4xCita
DKShhqKCESLExhxlMlInsD9HpRKs17P2NTSSxM4uB1U5g0aFKwpioG+bTroI2q0HRnpO3G1zo8lI
RFryS8ANgTl8whG7MIvZ2AuUaGeYqDoji4LAOwlmdKMBaeG0l7LtWpSYbBRKbCywZl1GvWM0H6/d
v9OWTRGFFvjtWarxlAeZU3XvwSGW2mDvJbe5o+ksNEFNRcHsB3rwr9VNSgul2KsfCzwA4cLKBDtM
h0x9+u/bkigvVUXskU4vyS9Bm2tlmkq0sy7fl5jKY37v3j/6vKFOEX2LECvvfmCBVl/rl82hecUe
exhXVzMMywCgubbTlPYkNsw0wp/St4oWr+GR1XsUXGhyHaj/Tr/kosXpLOatdtkCXMrS1lE4+PR8
Yv2ZwbUrSZGp+cIljRBSWowh2rSc1zi1lHXe1lEPie9zOqItlzmLj7cLt7XkeUXX0DoHD4mboWHl
PC0ywYkp6XKgCpt5E2+I89tEYCdjyfTaEKPnahgKQ8eHTbUs7BLFaInNRHp4J2b6drzpa0wtw0Y9
jbJyPo8k9c3xRwgewDzsyThuj7w+Ch8sll9tg+NYSm+yMhvJQU0TBmesXchRf7MhgLqxtD6UJiu9
xKbI0UT4yMlcE4BAJBFSDjItcGv01m0ha+mKfxuMD3CjAxeF1Ljy+ZHBGxuUYCnMBruEBzQB7Ix9
v1VK5f7fN8c8IWC1+UztLD97ektQdpzRsj+dBqZCBdkaFwtLgS2STq6MaHNTlVmahTTk1nEbqPki
W2HyT6P4FYRJ3ouNlWKvtvO4fEE1Kpu50648FmwujnkeFK1zBBG/Rcs9TQDnSBTQuye5qWnfwjAT
0Zu7Jz6obxyYp+lTSwrxdnmb4zeVjiYSZtUHdpAII+i10Qu9tlUscx0FdKCrhgxYSu4ytQdL+kNi
+m5DJCaDDCwyK9I/hYVdH7p0TpRwmI4ERxo8DlPV6hSH+rmhB12MBTak3Ya2Zi4yajkdUTtZP6MJ
B7cIRxozH1JjCK7qayf4inXworEQZYqRqCrDp7k55M3RCGc0Un0U6gez+AigkbcPMdCIZ2jEtu2l
vo+2ykCWwJjIYwdtnkBuauKE8LB7pQTYOtvvUXK4HcghrFG1EKcVtQFVg5I0BO3OdlqECKMA9lTD
RfWN/uX5X/A4F3NxEWJN/8CFPhgroTSOAJvQpiyIpm4ekIztDjLZDAGixOCYHbvgWTEvs7xEeimL
2abQpfflj4SUFRsYUl/0bwIM7d2+ZjnL7AagfAaLkcLz55tBtYEwR+H+bPJRoH94eP1LXDU0xUjW
Mos+ME55wFzpGNRazH3+bHcbLLkT3Am8QVz91Ur5hqSXc7FZY07XSB8yETbUH3rD28ojMLrP7SRd
DpKhBG1lhBrFl/j3jmscKPXpuuKnASAFQdO1opB8DvaQquEfDaLj/rQh+eTmYB8Nu77v683yiCPF
pt1BCv+s9YWlRVjFnwuighOt+TpLaq3Z6iA8Q0U6COlPVMJ/5W2TZBM0M04CVNmfq+YGRcobalhv
YVDQ96UoUE00oPykzFD/F5L/gEjhhtpvohzlNv7Vr7plD0bUHY5djrXJuKnoDKZTWf/y2PAfumUh
Kw3hTAfeQJyd3mf0bc7x5AAyVLu2wWA81slJPNbXu1i+WpBYoqeFbol6nJlzt82occCgjH+QjOJ7
Z1few62clIsEV2x1/rFGF+cyMjMM2Gx/EEcSvIZUO0zR5MKCcChccy5mF+esxG12FgWeRXRDTQVy
/hMDoHIc0hUa4jAslHs3pKxWlHKurnkcF7Iship29/DAO3FtvW65ogrqTH5tzqDuWvWbsqZA5lqe
RZATTfnozk/xBWf1WVSLuCHePBlFucPU5xpq5CSaKFGiOW9v4YEaZJFifCARrErjzKdwuy6v2YYL
lgXyGPHcznD3iHHFGPI4V1sYsqYgte22sWbtgQ4s9qg2SPJY03W1ugYbvQklw8dashUC6Sli31Zm
kUrf5eMj/1EJjFPnvo1SSNW1EdDj6fBeDmdswQdvA7/8tHgAyJtbz8Jgctyaxswdq7hQLeZc1JsN
c0L04MrTvq3NzEMEnRAHJe8ygJpDaZTqdrgfREq4hHYLL7LFItvaNT1+vvTHE+as4+g9BCh6rNVF
XsPd74/bIMRKp2NMeGzre5tsXMFo3S7dhmq1x9lAYzvOoicjOkKgBxOdPq0254KLmEpFoGLnaA1t
sIvlAd8KzSN0k8xNXHZRKeKwvPBZYQLcMZGjUA0JfkKXIZJv54xAxy81favsEjdcBwASdVLWcY1O
OZTymdcVI5LBzOY9N1u0fWGWbiBFzjKGPnOpZoWz+tCVV1wLbPUbG5N2PxKZXibMLsqqB3gSCr1A
RBDOYDnvOCg6k7HJ1QBL04BZ+kkkCtAOkc282Zmiv/UfVmz63P3e1n9kBArfd0uAZw+6DsD+2GJp
UAP85b1y9QouX7HGCUa6ju7/5T7/e9n/WHy3hnNJqEqZs80ew+z94FBkLyVgm+0pxukhI1crd2mL
bKgRJp/U9Gmj/G3V4rwIJVPjaAj5ErtMbsv8FB2VKWami77eCUmolzcGwacAKQcoEu+CvFr2cXxr
rA8MAEAbhB5nGxUtmKi/mX8my20YBrjGU/wdsjHEjYct0jWWCvF19JID2Tb3DG5vdbO2/upXSaC/
2U81oxSJEa9KHKXC2RNnbeEwHCb8Z3/tQsL89U/LS6FpP9DtfUEiWfubSnywVmMLHOc+e/oayiDs
oT5rTnfiR6tfsGTXQZo8EkqR0W3J5tqFY117Zq0DHi3CwggVJ/iTqNDzBA3Xq/Q4od+nZrj7c9br
PI1sAOToZt86pbAorxwU2WB9Gmkdn8ipjkT1GrP4juryxJ1NwUnDWnH+2RYdb+0qWFKRFBtNQm8b
SRY/gdS2+RpMY5yPljhYssHz8flSpRWAxhDkDWMtM0PEpGlbJiGlLm80Hj3iv3AIR3vdKQhb5psh
6ibYfaYeCoJcnelmLUWJe5VedqgUYgHGc9xTkgPcPFhWEgMAtLNrBqbKcRFAvCyq+Ffk85PmIgKh
Z+QTYakNFkKimF5br2iEl2oL2ZjN5yFsKUJ/3dzKMpdg4uDSo1UF4wHTLGRibtDElSsDhY8/0Gx2
0M8/F93CHMnLFDZ3daw4Md4v2ulN0mEqES3F9k6ejqkOuCNI8iOGKvKIayJrdmpBcZ4qlG5NZqyG
dXMJphVXka15by1roSsEidM/x47/v6rZMHrVudPZ/Jl7PKX8gEIJnnPRWfTntmbY9SIMDXyQLETi
OqZYKKNVjtnE0PnRUNFOp4r02lypPciVp/jtv1FQAtRzQiTFhaCN6IRl75tFFu9DqrJGOc77WqhA
zkJONGltIZoNVe8H+QMDymX3GtlDBRDIBoUvqAog1qHWDlPN968q6da3bVqbq8258IgMufpI1Lta
cmXBxd1b/+eFw28EwAdHVF0vqxA+Pi6DrSGfEwg5hgYnpu9Kt6Rk+Qk29xbick6MK/EsPPUwGgqS
raS2tGecZy5bAHdyAdoS3g1W84mfehlnf05g+uFdMx7w8NvS5bz7/ouEjKucYUdHTdmERJbG+ZEM
ITqaWbYlCexcTB3SRc21Cb5mxKtYfGm24by1Z8vF9JLkS9cztcMKE9oVVkakcvpXT4is3VX4KtkE
e5St/7hdRmFnIiFZ36iulCVWozQJL36E6mZgrrIG9pzp5ngUP4N6RRTGNNZbkEx0TvZaZr5OvrPb
8ujYX9vVccTyPBqmIiBimx/lIzJZ7ZYveng5f98FMNs6S8W7oP2dCAWVg4HKCiOrVnLGx43NinO/
9fGumqwhDBn7tnqCoSg4tNFLbIpJL10IZ2yKGfUyICh7jH6iVeDft4wUU6x89igY9eeNKeKHljMB
GxUFR83KV19hNtzJco4BtiyuWXWXynwM6LdlZDPLpj6svrDFvXW4zyBe/z05/fhUhy316Wk4N4sT
HpjdTZ5GS8bBpuTUvLNZOjVIaWFXCKZbRi3S5Hsr1N86YUTaeLyqdD/AD6Z8bvh3WatrXVRP3dBd
PTlHPJ50s43MMTjFYLfFMRadcrvEkf3avmIcKdJ1GegMkE/IzJoXSPrBlnkq1L7WL8r1yeptbRiV
TgQRHSBLr8pP4fGK/5rON0mtb4BW+HcZl3otIQcMkaiR6+DHCRBTl/cr9oVPehsqNDyGU/MOdTFL
GBwjMF5oVZqmmRxHZBMvaIbiao2ixQPKg77SA9OUdF5zqpck57MO+AI8zXObHpGPw8Z8YSh4c8/Y
l+jOofctQuLwX8IdzQlAuheCrhgdF3yg+NF1IL/XO/K1TTLhVgCjE84acUhV6b+Hg6rZ4B8Bpf8H
LNQ5Nql35xLYZ8UE6Pitj5Rk9eAILzjV3cF77mMVrxu9EE+PnF32oSkPzS9leDJUSsgOIu8diOxe
Jsp1zzHqIzCfOEDaq9dJ/8lvCyB0qkFaEBRcH+ls6VmPmpzExb+CO/oZF9gNxhalbzPP29RylWqK
aBg/kLcKg3KmlxkKeg+hVNefTHrNszFrpLv+FF8vjuqbxAOzqrnilN7RlLBBzIb68XFFn8szUbsq
jZSTd8+8nviH7eKPOMIP3YuknczbbItiZbMFiUxCJRZytDzVI8C8b/7dNprDvpjhxQfsMGPJwjlB
FlITRc7ofE1AHRv/+LPJkRWhjQl8P0iENwMFO35sossWO3y4AJv0NTn/jtsDNnnbnRsqIAsevfDY
jaVYaSB92BcjRidvcrdTVFCTFep5+UqFIVK6f3rrmhD7bqK4Xpq1WbAZI0YDasxiwWHDvYDw3VDn
DYLvrPIv6IjSJNk6tVg5hkal7d/JN39ko5XAN2yTnYMF610MQvyKrq56WsuI0T2n9FNfzAjaU7FP
9j7DeO4ZH3NWqi5v++TJ91kOJwvYFZkmWzBLrkuuAU2tLHG6n41w9zRV5IOKjeKTVd1P1PJwDBeu
K51SCtNgJtAzsJ1sgs/5YogOWUYIALFdlYWzSDh1rDr5I8gumXxazi7Gh0VddkUUL2mBX+knjgLD
Beuj8VztgQ84XzX+bO+MK0WpxkSUcN2FOyGtCbjGGWLzKq25/uAxw3DRCHI28pI9+wC7ZFXCOi8r
LPhckPJT95MAjdssHfbJV3ctImu4aEnIJsLYlMg0RwCmr1Zyp1gA7QyPslJjQtyYvRe0RCd/Dd4G
iA57YIAK4TBf9j+y+baZZrH3/7Ivg0p2zsVsFMHO7gOqr/HF4XFgKMKHOJhnYCPMSvoT0pHytgsU
V5AVrO9AfdDyn3t11o6ambZk1QX6zL/S0hacldSnzS/8pKyAcgGOHMwEZzV7w6CF1S1UFsF3LBDL
K9rvogRT2vS0AjHjvq4Rghsw3WewLv6onmh7RGCOv6hfbJ87MYw7Mtp7ta4JGPQfgufIAQuS1ho7
2MHi3LRLNi4ZOYlxNlxyHrti1dZXGWPTmxLKQTM11XX2BnWuHoU6V0clJZGJ8M+dxU25fSKAbha3
0i5st8pnrc2Xl8cEC/qvjL4maqY0rZdaWjMS82NRvEZvRDQtS1MGq7OjWRHCdiLYfppJyKNeqKbJ
xtMSy/ZSjvP0H2cDI3IYxtA5IbfbF0ZmLWhTL0MRnbgCoFUSKf7Nce7J3ph2KgtthFbXP9zzk5TB
squqPdRT8/qOTclOtpONKoxWrKwti3xVwOFohwKAQIqPZGWjstFJY5Jt4fSet2IbNz0NgI8WDfK0
3UU06dpHZC3d6qMnELzqhhDZf+vBmSSrscR24rvUxhtvteO3cmnfhTOXTEB0LAhgxBy2lLeCZNen
NaHMG3T69jKZgbElLjJytFQhvfT67wTn58s4j0VrTWNUbpLUCab6YIUz1hOYMzwGtgWHP7XbQ23v
VEWHcUtsVbUVsNROTr7CfkTqUIgxxP+bl9hdxqnq4FOdhfBCbjnxL1hpLioRJSbjLJFDbeOc8XKh
dY3vqruHJPt78Vgwdiut8Y6fTg44YxntiADDpurUMoX1wE1P/Nhr5VVChgnpEPN2OjQJSxV1a33p
385+LrX2MM+DX20iGYD/9Zr3T0PuediZ5p5y7XBAHJviIZY2vuAhIOKPiHDNJOMhRMovviQqApcl
FTr+pDj96hk4GHzZEhERuEnm1Nj1dvJdRL6ggMrccVmmnLDo45C8hTVNkPgWQSbToRVA/7dS7dGJ
LU/oHbJOVOayRkO5sND5yOYkKomdl5pip5LKUv8zFijL9zS8igOFaeVEiAxa7Vg+NzkyckxvBwFK
3a2AdbBhourHqlTzJ/JOY/hrtN7KYeAKVxk5akFLxNJXZrwO7WMqgyNeE3g20A6aUGx5mCmKeAv8
TnpUmTkxzIxgFtFajJnWCE3M67LmvWh5acgxZuU7gL05WUD/2R10g5yDlgWfHA8VejKs1fiL7otE
SNYwRu23rWPvn4yMIgpbXEHlBQDk8HzomWspYgPfiO9vDNQA1B0rx+BwC55Yx3ddXqVha5EYwj3U
tl3ecUYQ3IzDrEpjnW0xOZhH3oqkQCHTZT21L05fx8/tpW33QAPA7y0ciHUacbqV1fv5d9bvzD6F
t+PvdxH/2XtqHp+jN6vhaKIOTnpHQqOuWJjqr1+/TBd3s/I2+wdXHkWE8VwNt3dUuSUGIG/fCyJ+
x0olS6mfY4OW8GhKnKfOqfwvsvF+8i05GPth1WI/+OEDGAvYXyo3csOO7mu3L21E6h9Amubxp/+s
pgt2fLz90qjxFPbBMep2YtLXY/BeHRw/8AtWueh/khJaUq++nFJlZI2l1dp75oIHJiV0B1JKyeUt
dgAwMoHCbP/yRSWQf76aQD+Bw8KSQDX04fcyBcltQQ5AVcoogvJqxq+v/BfXgoIRgEooZXdN2akX
MmgFZ7frV8xAtuT/KIyA/l00kvoX3ujK4+suFuJsQGZTr8iC/omPNU+VxIgDfiFE+sYzV+Bq54Es
5ozj1W3Ou4S+bdPObEy23cGqX1yKiGT7Qq8w5ws+FHW5do6g9Jz//sJCOfXsStaagI2j3JBisLwI
4OpfipGjIoiDuyKZcZkeScBVQ/WynRHlcKs6CxX7CTpsPjW89jy85aKSNXBzOwFLIfQiVKCiqUqG
KBkXipjIQFZSK64FkfF516Wcnkt3BZDsMAmn1w22TTLmZScheCyv1N7i7kVeOJuGFvKl8blZG3GX
Pa9+RlTuQ6benZqSJSQVo3JMqGfn3WyW3cW/lvCnHvSboRHRU0FL8G0Yw7DfbSERHFYK3vTdEyjF
gtX1Vcp3NXortd4Uw1Zh+E8slOisauecBeDPFrRhkKj8qaUOuQeCu33/tJNnKHHuK6W064pQSIig
hZ13ZDesUBpe+JPTyYquxsOzToNB6+VlSLtNDBgzLpHMFrwekMGahlUQdHbDqTCk9F+BXxYumuuT
V1SgUAYjF0v93it6hC0PsQBzEsWHntlXhEvkhYarovZDIlfFIONbg9ZR2WRdD6SFA/dvBr86He/1
bQ272NkK8QwPY+Su4qr7UISXfSf96ZRnmc4cKDPJM2RX3EbXHhHw9zyjZrOE8d+om8AAN+E2AM7Q
/cgLE9np0v90Uv2PKv+TvAMlNKik4y9N1gYOMeAHOsgqpr33mqYOLmHUVj0Laekbjuvwa973qFBr
NQSq8IJF4SZIv2rPDgEHw6VwxqG4qRnwC4/GbXU4s02kK3IoTAGdrUEM6/k4v0Ze+HFVRUWqhVEA
AV0jQdEp2OiQv8JzCVZ0Xn/6F58Ojg2YMzAcW50Sj+IGJJz6wQxGlfj8yDARTYf0y5780k44aqtw
Nr1aCo2MvkRSX13uXSy6YiiyoacfxyUA83xjS3SW1R8Q06iinvVB1vdcOrEsgNOMyXaPuvtDjp0T
KDOF0nHpk6Y+SLIdE+7OyG4/rIUBhwJJHZM+cE+SFteE2JlI7N2oD/r9sYvt6/+JDG3WMrSMTIvK
lbNsmsnxhuslImTYLVT81dVJNlb2gvJ72gfvXkafiTNEhIrMaozCLCmZES9rqFnduI3myb0xTtsQ
lulbjjZw0Yc7z4fKHkp74SodCtuMGr+J3V8542TpethYKkhZ6kPf5q5mNCnUawcSMR1aQpv34uIH
73KHBXajFv7TTYo7MGtT5G9kR5cRWJJ/pOB4S3uhP0ZDcW4Khlal82MwkzLdFUbmasBwJwHqxczx
Pm4aFPNoITV7FcSpUoGv85BN6WJTC3Bc3P8Dy0ikLSYL6PG+nCwq+DFrTNcXK3LPV25ymRIFlwfI
MbKTaqHXsjMQc0NfWne8X58IkKFhGuOdldNVO0+VEKwDJQAORhFv4hGlsmJz7I7eK21euoTJQ6Xy
+Orf/PAn3rhZ2D8hk0zpmOAP6S9eyunnKmZDV51dLJm9iHy/LiEKp+6nc8Zd/Dn53z+Zdd9xhpe2
mV2YCs0xlTDnwkL1DTjr9nwbpLcYIEMiymPkIacforgQ6Y6kPrJl19iHCOzg1MTQUbx12Vt0deQQ
B48m0z42lr3ln0/qGwdM9GihoGJ8OJpsmvLzdkpkfsvRRvY6Rez5Z64GnaERBTzk3Rvqs6D5JFvd
rs5QOPB7UdNICRjKUSFZxO5V28IcU3gkx/tBmhs6cYr0N31BLhOJyMR3hSad+niFvPdjQUXXK+oa
Zk+4khPq6YKYRgVpqK92Q/BjgmQOdvC5DOqm6iQepvav7clrHjFr643mf0I4rb9/eQymlDcf0pl7
f4VXzMbz0md1oJgKHNsvGmQkb6n5B/7mLh9HGiFXKDbLADiTWQic31QSZEqzAIl10h4mVpqc8NTx
f+20uYog8Q3LN7S3y/8XzQM1yLa1vhSHVbf51H8osJBTM9h+Ln1rUTi82NpvvCS1j9b/UZe8cmsn
1gvk6EYby5Xtsqb+NB6AoJgzt92+ut3eBxuXQoLWinpWHpOwA4TewdTXhAF/d6PERlWu+2pLq4lF
TAeIeRMSwbPbnphU+tF+vNnOKQStXq274xFJPcjTPzL9Eerj6ZaOfokd+RtGuaU+YOnSnOthlXlO
YAHSzT52/nfy9tTzfjfUMLF65VGEZyLNXrV5dj6gEtddxvR8Bq1U9QhcykbRZ7HJKP8WaRLFOuob
WIUNtAGp2mMbQZIhY4mrLkdziCCsDCnJ6oIMlPqO6FoauT1UcvDRp2R1j5P2WgG2D82RxJLsO/uk
2CKyRQx8btwom2Gi9qqtkU/YrlbFdu87eocNv1yNN/zF0G6lT+kVEKkL5ZwSGTskU/N2J/0u8kPm
TRHxkxWqABu8wa/8rN+R7DWaHgqmAuVw1HUbX61xk6wbYuSCF5cc/8l0bSWRxg2PyDAxFcerdisZ
YkuInQ/vxctDjYo5IK2xi9fE/YiFC1TCiFAHeBSBmUiovxf+OINhzCbQYbo+wGS6FDzXXsavvVS3
LQV4NT5FNIw5kDzybIE+N9RsBXhUYZgKJyCgyX7BjJ1d0+HTZvLfH7R3ArcpOP2QJGQy7u3UEIgP
TYw9DaAd/0obkfOhYO67seHdbIvNbibNdHmxzs/uPDeSVkbJlKSYuuVCfFAoiLCvNUh8O/SHsE17
vGOIh99dxHyn9AgSulDMDr1bPFQEU/uXKSzFgH87X1IafIKm5de0HinYNikcjr7Kk1bnUswkilIE
RkVis75+laZ1WCOHAi+ajVVGIRI+k+8zjejDv5xkTVcPPdRl+PqKsKsvD5oBk5RExdWsYAnTOQlH
+XkaamG56IqOjnJKie+aKfD3Zo0xwbWMKxKsRxE0Dum7q1ginTbUN8iy6Xjty+BZMknv5IRgOoKC
jOHTfnW1CHgIm+YkCSLp05kVFD3DOxymPaHzTV6nNtAUqYjhIBwxf2c7giaSBml7xbl9kj9lz1WU
MZ0C7r+IH0H4scNENdBtlOjPqIrKZsYEpkcZEsuEJYmPYKUF4zqinfkg2Fw1U1CTRayPgOS3GTtm
vpXnlhh9vUSU3HznDFj/3+1U7Eivkf9ZOJEt3MnVMGyo0uAqLKHFrjoK4J7fv/5B6suSFOiyefQQ
y1Lpa0ErmX/bJ1jOmsi8MYxqt0InBmpseaNEMVC5Fy9psIKUx3tD2aOncrmk1JpGv8NfW101pRGU
fyssAsfxWXInuvhJirq0KtIGUnNwgMxc0piF+gOJFjY9JWoSOigHGO1X3mTd6a3/VcHF4hyiqGvd
IAvQNXT2K0Sz7YL3ce6AaY2nUgG/DZU2NMVM78pmjhKElX3qtWGFtPGa3gbYQtppxOtCEFktp2ci
Bu3TbBMcUWffpakhxfR5vB+kNMxOFqMxmKRZqYyaCW1h1slP7Oyj6sm/CM1n0fC7m87a8Rq2pTB4
Uw6Bg6gyhI9N+XseXo/86adzVkYpZXtvgzJtSNwvqROJnAKjURWYWwlD7GlzB5/TVlmd9ombh9ue
xf77E+qlkgC8THhbkaZRetH5i8hj78JCIm9mDYTpT96tmat4X/vTIV07Hx5TsNQpc3xDeLclR8Gq
yd3ZIb7kZEOwSG9rs3je6EIb0Dxltk4PtZRyXcKxWryGfe4ua9vLw8tWmg8GmXseB/55H7sPwt0F
QXUJlfTQ+B6261+0vUaC1h4OtkNhQtq73fUyhTXZgxDi5c4LBnGgYckB1u3NeB6Mpsrb8oANedjO
88PFucOBHeV2oSJj3x6OH/tAUk6XgWW0oXnqIoUcxp3VcbuC0dUQuhTrJNAFocFDlvVn4FyZLDmH
nzJpAI0Szz8c3ZtBFSbM1Btd2mg0Ny0gPX0jVWcScr1HtJ7eIrzMn2KjsuxNSLUJ8KGV0M1S3NBa
lJha9PJZBVpV/3Ik1elmTwy97SaZpmaokZIVhTUOfF+Rm8ZFrPQlan+Smf1whvRAIgymWYs/m0ZO
NFJVNatu20OG7cPuGMBpcor4qrvnT4EnmfrGy0ybM30zGZA1HCyDdRdd9qGPZrkDBUnO/YCHaC47
scEG8SoLDQ+M7/pZeaFzEMAJSpvQplNPrK8VnFEPMy/CAWG72TpRPx2qbe9yjgm1JWCxljqfHDf7
mvJD0+RQL4oEQoaUKYRRuW5XNfVXYXAe8ULgsWely8chXlVX4iqGxlF7fdvuVWQfssvNUsFWftDN
hXpIAQzs0qFvReF4cZdko9iomToNKuCsmb5lJXIoVQ3XxRrvCHlvl+Ylv6qZdRq6GL5QSHnU7yaD
7C1WieQVExjmUbzGFDHZqiwVBHpbjH0Xpf+TMRZLHSmVSttCBdVLt69e4Id8atwd1ivNNmcFqzZU
27WvjdBt77pymq7AsdidCjcHNJS4nk2PhJOq4AyZ+bMwP0CPKjovFM2Eiu+gbmt+g8NuW5ccn7f3
qG9MmshA8BZo9ByjMF7cxVlX8/SKVbewI1JVpNJu3q2O8ZEJvw92QcgmmlQxFgsR/7fF3dewka+u
g8/21+PfG1m5/u9dcWxyfQFW0QNzMusQjhF7DZNky/5AAVgSizDTBvYNMiorZJu3VApgyECWhHZ7
NIhwPL1tEVFKQaOUDx3D5IIDc50qjYcnYEBHb2piFFXzOPvxzTbkRD2qnbBRBDrPyMeJcbElOr5X
GKIln0BNF9nx9N5OJkxi8dxuAvmsPi9TcKzKmw8qt06xw6r4yCGrkwSN2D7LvlJk6al/ae6KFg+z
dgwCwW/G/dw2KYuSKwIucQO0bpFW9HbKlHz6iDv4AlICNe/OwVKTUETKvsetIS7LvztxBXOonOuj
iNSVRYeCPU4SrfTrI37VVu/RZ4+0N9FP28ut6mMYcD/kRU/g2P3HqGjT3DCLu8b74dvibHjslnKi
W6c9t4XRDEcT/Wn8I6YH6XVQ4KblPCSBTEcZoShQmY87EcA2zAiCnVrzKNKdHai8m8FU9DVOjdV9
RoyLsE5EDHEBOBCmslqlPRpDt2hH+dEyoo7XAWBVfthK2WFihbfQMurE7ur1wsviNwULhoLHxhrb
A1HENmzQIrxSaW8F5qnIOm2Dvz82V6lwYDwCWorme38JFuU/i9pYzGRcs7HKAf+l/EDM7yPDw98G
ccZd1jWJUqAxTdmh06X0k4v7XocVb0FUYGlQupIXphnWGAXXRzfE6Ck7gZv900HlPUCqKADDHX8T
S2W9vqtxFsTGZMN+9Sz8mfW1C3Is7orHytLzo5av7Lq9N9zQlSxGxIwqVszfh/ZRQLA17dtyWkQM
OHfiqMF8IxSXB6vrdHceNZBJdJOAh7lM3aJH1DvKjtgapSoR+197Qv9yT9xBNMXVBGKcrA8Kj2SM
pHW1b1XB9qje6fRV7neQvN5EhJwnjZ36IOP5DMd+GVBhJBBa0IiaecJK6xAPGKsZPGJG1ZgyITh6
qpQx9IBAmrFn/2GOEXFCbrZeiqFVnmYKTnXC8md632qV8iAerTgbxpOeGr+9E4rwJCcIf0xWQozW
Yvf4u/bEr/s6yteF18Yq1DRYQXne/6uy1LrdZbSCcwo4osaGvzCU8z8vR6lYdv6a+hLZc5H2CibC
XEeNLDiZaPPnbiIwilYnRMu7oMq8U4o6+AkE/BcrGrkUcKOBSGFe9/Q4NK6EbktZM9qB1EQZQq3T
qcod8boEZ+DEABmmiU+HXJYXzkgvFbDTD8/fs8SNzvyywnTlwR/52stQcQ5pfoh3JT5ajzzInrJD
axykpN2hLsldhbiKoKmI0SQC8dTPD0ftZIHVsHRT/6pMjsEzb9zGtZ29fNBwg5I8PcaWP02mpB3n
xX0Fwcw65WfbzaahSGlWdVcZK9aDM55WyjoctLx1KryIUsMOdhLxy7qSnBrRWNN9b28LaQIFn9BL
Ns+c6vToVNeUo5bKas4Wi1HwM0HEPR+dGhcyz1KGxEDKZfRoEFwyxQVNHM1EX2C8Vgdrp2NXxB/q
DTEZXkIHPA5lQsO1YieWKc44S5omouRr0KnjaO2g1UtCX9NLOmpgX7GlczOVOfH+WQyFojzkVy6z
ZAkgyWSfLu7zmM2CQ/uGBE8IGt58aMHFhSIHZ+dKuZKOXmwMSF5KghHnggAbLH4FI8/msj+QjEiE
wDZO1XWe75DJk9HqkuEkP3mORnOOCIi8LRFelsLi1cLeGTF4/UT7F7DkbjDq9kGIJgeRgFuBEfeS
6HPQxO5n+107w1QlY8LoiFFkzLg5tblxo2oqs2xVo2HJ9VCJMfLTG36QAJLR2x/wnPwxxVeL/jrr
X2I78gaY+6+jiBGMi+RWxkYsQ5C1EELYK5gUfvsld9EpvFAg+XcOSa0Y9qzubnJtBdg6xoDHD9N7
CwnNdaS/0unkFbz60GFJknN8qzSCZXFHwjvv+XG6RD+z14EjCqHsHihV6goFLSUSQlrMA8yo94SE
pj8BLhuFgp9qnyt9mX6WztlHGnCdEWnPW4JqujnuZdI2WEuOpONBBLBuRn7UHPnh1C4DLCBarNvP
vjsuZ17NYTKR5p30+RVAvfFoT9lGaMWnLj3t3gR3sXur/l21xVM3Gu8yvbh6W/oPvEyHk44RMrOz
HPBH03YZyw+FXZ78d3WsROyLTpeFMDOw5vrQR3GOsOVyLY8GXRGNOWZBZaVIQMqK9AL58xwd7YxP
/2GB418+BbSeWJ+N0v50slXGp+JMamX7h9k1/cYzS6nqwdU/sK0Piqy5cfp7ckCZpU+dm3Zh/si2
bw308OYkjv4bMDZ2xshxdVLIIYgn0IQzsYC4ynM6R5n/Et3Kj8GXyCRqs9aMUgV57/gGJiKNbUZM
UnGti3dv+a6i4B6uCz3RojiQy6aMKWPtqaq3GX45B2YVyY25Ia7rC+Nm+XSfsSULIUVoxYWM2nKL
37RKNtBh5eFVhLMZLswfopH2+gNnOE/4rGKxw+3BU0hoeBvA2tP8ovGW3n1/gHzQMtYwj/clkv2i
+jNu3w80apbbDtcJcOygCriTeLf/VDMjW64WWqHPYN5B0qBL1smPHqCzwYEs5G4y1O+9/1UCHwXC
bxPXBEwkLBJCEPxgjK6N+bA8GHJhYeqGDwE4f5N7JrwBCRPi9i8Y2QK74jiW3hwYo+zxZUmvVmGq
DVLQexikpP7gu+IrpMsvpqCrMcDK6oUFBJCL3fq0DB1jtBH6n0xCkZtOmNEqqkyLQdXkFeLydfdU
pCkqGGWamrbDLcPJwDBkNNqzwDBB5yIV/j9HnbYYXgCXdPaqjC4r1U3HptiUVyANclB+bLknRArC
k3+2Rki7kVgYaTybY/cAUWciI2Mod0Qtg5BugUm4k+FTWA1Br+ih4/Hu9rz17qtIMFXAMOtZYpt4
/xP/CcXARj9ETAPMgsrmpEiSOxQ6KwwxBWZB+KMDz5/MgLwPER1OrLfIIQ6rtG54T6fmUwvB5cIG
eYPQm7Bph2VmixJj0pVSUyFfFwHdjKl+jO8/DmCqZhNYB2n4hce/0mg+NIw6EziQXIJ5DHT8DM4g
sL9ZyrGvgoev56uu0g9PEYm5toTy6Oxey4dJtx2fToi8X11UyhFekWpxjnza/2aLyjxVYc5URuhM
RlN0hdsHvnDKTIl6yfB5zfKVQ5ktFfUVXfUc+FqG+JHnd3eBvBWuUkG1M3zAH0OjDnk03zqbgcyz
plpxqTQDmgs5+2u3t13PKjEqLeHYIUh8tq26pJHbcQ6aL9a+ESacnB5btqpFMt8NRSz86sl05GvS
tU58oRtkaGNVpe8bTcbu33yNEnd0myEVuVt7Kwdv0jyq46TzGgHx59U55PCCp2q1CLsBe9i+G/yz
14uQ6kvi1dJo5voNgBfE9lqe7kQhXwQ4v3q+PPlUvrPZBZc1yMwzVm+WfUfFFSAQCCSK4CgSY1Hq
7TpzkzcdjZRxxJ79T+99lcxb5tgq0AiSPVz9P2M07H/nVV3cNR6ZBr9PmB+QBalAeGK+ot+91wLL
aGI4CI/eqMJsmRkz/8s0ZqsHIFNZ8NOhN5ihJxZVsxuixO0Ww6q9pLpjYCd8mDm7PKjSOL3XqTRD
2FwbWmGl7Yu2CG0Nj1UU4VJ+3ecYD19xm/eRU93Va4yKWE2yfxc90mCJHbCIrJG2nzmRUOGMQcSz
gkE2vrlSAzlBqf30AeRT5TrcguC65xycWqc997gns544ljI/DKRQQctl0nb8XVtr0E10JvU+qYaQ
4Kj9XCozCS85SDjYtRnWpJ3bSuHLTbjVAl+k+gXakAaXr0iO2W+mrG9rA4uXsbyeE8hwE1GlcMta
hSmx1pzU+scPLWqtOSPtd5iuMawjtWpVkX+L1hQPhXuzVRZ/2FNN6Awoy/0+NY7clgg+dUpqgkja
mhPp1aNLnn77joyOvCLJAaQ6IkiVgQfzaumyOmJD5TI9AqIxbRpMhgQ0t3/4WwVajdYTMQbYxrez
En+zq4hdjT28WzhL53h9udWqpPhYTg9gCw/dXqKQm0rqG2ORb5MbGcK0hlytPOLbQNW1So3gE+B8
MPiiCKLFRm8gAqLJfuLp5H9V8kn3CaCr+zYmqWZjCPknIbgVuj5UE9I8JYuPBziMmWztT3VH4KAs
CQ/9JRT8OaUfByNxj38WQmrfHwMyElySrcwm/YkDESce6lbV48hplMbFBYf5j0SHDaICAYGoeunu
t5Bf82oKj8RP5HhERtatIJeY6tR4vbdNlmqPI6kXcvjeFYq3xgdX/Rj5hxaYPmdGsQGzhggECUCm
PxfsykC2JhSNJ1LXSL7dCXi09eAay25G9dlsv8mlE3WSH5YP6+HXNDQu2WfxqFFwouPy1FrKqW18
LxFnESjmhcV0P3il3A2XP6pEQUkmgHCKJ7VRfG0rUMBtgYITliLH7sUvdgnt5p09he8vCjJI+CQ+
hzjegK18EjVfvIiCjseQJCDC/DBxYSNi1jibrv7WNJgZ0yqvS48NzWsflfRQer2ORtoBesNRJj4G
2SQYkazpH/EHCyjq9rQonZ01bupJdZGOtdiW9sr50lvHighVM8tnY9r8CM6XVc5hXpzQpNOv3BJ2
7oxqwBDkljFyIAkS5HfvNThqnuuwCm1Qzh9PRSbAMP2B7hhIh1Q3UfNbQBlEOPcTnCW/s+/O9wW1
5GMu1i4JBOsRlGYmxMu7bzwUpWWml0TFWb/tzSsnJyRxI+q3iQTzbigi5npdMCHhvL473cpuFBy3
wv5mSRQb4anwR1yMBFBjnPJ6BjSTuFbKJZzICXL8+AxsmpLb/iw/HsdQWn5CpNWJbmL1Lohs6yuL
7TOiI9IBCqaXXrjuVdc1tkhoKgCBD42jDEq4YzMPD0K+UC+p3tAeP/amOAro3OwtoPcZBI5aiqlb
fBeZwHbm4ja7WN6dFNOYqZLBxft16iTvnsG8n2QnlxIV5SLd1Xnp1KWFgdb3pNdEW88Ylgtnb+9w
37w8uK6DXjiygDJNlW4nz6AJv6cV1SUrNXYcLDc1D4GiaVY5GykvmoNmPaNfbeA1eVNi4JaR1QC4
/CiuIEO0XSm832gRdrAkFNhQ5+8sr3fZ3Qxn4zxqCb5w+mH3ajNsjRE5p4UXYJS9idJ4ZhrQMrUt
Q7Fs3tDIMvzflFbQjyXb6TM9rKOsevkoxCpCkf4chGDqRrhJnjrZzQXCHyd0P2Bc3WHV2Poy7VgR
6hV6cwZUTDsOybRhdb0WCa5yoiJoqYSubOcoYPteHZLFgzm+mDlqv+ej5qp3w1YlNsDKJojBuHH2
MO57Z9X97rVQSyXc+JccCeeQKX0hsEgn/L6VoF1VgxtnnoHSa7vfTieUlpr6kBn+qNYui0JJ3QM2
k7XPBi4MWoFFomzCJYDv5mkvs+VQ8TKaGTF1KlnJ8RAcNHbkHeG9q88AZLFqgRQL+YVZc3l3G7Lr
oWJHSmnds4Lr6C5HEaEO+1lXCxmv8pkoWdM+X7opfmXCl3FZ8vpRyESEJGRZGB/5bp+PhKS9gQ5O
EL/yH2uApQLvU5hI4BUlcn45UsT1+Sw+FHSlMINP+lMV4xHb88I/pO6ZZQCJdzboenPs5Y9v7Jx6
37QsdmL8gKCAtiiABQOLUgFr0C+i3pDz5Lqikx9/YN1Eune/IRBCNvkW0JIUcGQXNaOLzHEth/kY
VGoPePfr1lJtcNnLayMprJ4epA+aPeRer9FPA3utGvyg+sKukSjPMWbUkZZ3TXL7ZX88ZL8IR+9a
xM/6ABHWefIPV1SarV/1mD/XEfKZITFhMhGg1ngrVYrGpzj7nF91WjTCzQ+WgiHFgde2LY2FfLsR
5AqCtO+YhlMprCx/F6qMbg30K7TOFGWELEs1XrPTQdrG7x4R0JIOt8+ozv97blGMnQNR8KUH2PiS
oYeIDvgqTYWUGC3Jv0unvkVivTr58HjpraNTlm8ZhBeLx799QUONjtezDLVX9PxPpF4bYuhMtNC5
OgHzWAxsl3L9mCxDPC5Et4Yw2jvyyI2gbqnVb4i+dqFkSZQzBbpbci/ItFCGaz7jN+AW8tHe7dcM
9WWqgNtTnsuwY+p0ksbKJLRgozUS7CNqFkzZwqLXdyjTICy6EI19k/OrYFTFXPQAzd1Yp5f7DraT
AcMCNSDkkzUvPehoIKDm5mFA7t22q/qj12Avytq6SIinOCxasseqlb9N6rRUx1QnvnbdhIDW7YjB
zTVnNRkUDqajlYCXDdu9n08eG45c14mNjmvR3hPfdK59ZGexbSKhDEJpeLDHo+ebcvWIpCbu07jv
EvMVrRnu61NIrvzlVxAR4F7+01Ad7FUILWs+7rxXSbf+F/Phb3MgHLBKmOj9KufbbvAfLWGlsLtv
W6nBr2cyDIgNaJPBQ2yH63EiCWxXP2CEbevv7nW+hfW8CNv/Hj/4Aut6oNuZjpP3VUaWSZoibDtj
Pc/HjHEP/Cu3avzlZ6/7xkJ2qMd80MikIRua2bHVwv6BQvxlzdzROG738SWcNqcOYHL4fGgXgU8u
OV6Ddl+2gP0dcTJmgqqRal5+waBv3OIgP/46Wh7tslMECkD36oHmj2VIwyEzWqUUaeLPM1ljc6+S
77qGxRvLaaixUjzn76g3yQH664j9P1NyryV6n8dVSClS+wQOploUnTljgWbMyZ16dbW1of2Wmqk7
KzKIqTBF5MltiyXpoLmRkohZujbIRUqHUdk8fJBgWJnx+nJ6dgZkVxfi/1hoqeiBzf1XXO70QvvE
nwshZL6lMy0RiFRKKuOLgWyjMdH6DQD09TlMAF3cPCrmdvnE3TQogUlfzKkStu9KF2dXxMIGB4p5
50lR48ZwugYWOJ1WReVXq/68gepDpZQGE/j5Rm1CRkAs5fqFpUhPcBnyKZnGxiQc9lpN3QsLAoXt
A/Ih37ycvvoBjC2xBJqO7Bh5r7Cq4u6Y6qTSj/lYbr+KWLL9GcshvmKwBzDnYoVdLr260v/c8R6E
E3gk/Ou1Cu/jvYwEid0hXZ2GOAOHiPx67bFt8YuDEfSNvTXXTy7PoZfVhYwFaNZc8XKxlQ2VXqoK
5fgellTJSGbCp9dgWX8Y7+kkiPR3kfEgobLazIFJvcSdsr8V6sUnj4DXs3/AOqkceUhABGXWdeqv
BQlR6rwetceY2oWhh6qOheU6cLVreTfE0QrI2o2HddZDgKThmtFtNmlMGQ3ZcOni37ZKdjnVtjPD
qvONnUgc8qFmznn/OqqqCm0LmPQiSJRE8ZRYFz8/hhViv8/EIQdwRcBKUFRyfr01b+uaBYdapds9
5OT5jM9jkI6E9MFg6pZ0IBusMOmcEGa2AQ6m7ZeRzD96Y7xxvso6Sth9MgXtUsb8uninREZmMCcx
RZLAWy4CUM6YJXOHNKrbtYNkcxIzD1nJnLAbKLmdkIxNimZeC05WTcE+/X26RL374hLQ/UNwD9uP
DtBms5CTGyI4CkNurmM8WT7LjMhAhcEJ6uocRjU+D93s+VKJVrJXNwKoMUJ3T7/PMUoQ6dldmbI8
rO2v/LkaNniO2TZt2GbyCnB1zPRUMiBSBFdsIuae7D241HUOzOFiLZdifxxnAbsBTUA65fxufRyz
2ufH5XZUrvHOi/644UZ0N32sHmExoK4hNaDa6yKtWTvQ4ZcbB5g3bSywFCoArOanAnoD6QRB6XHt
3ON5bRW6aNc/0gTI+gt8CqZFrJC6e/KFOCDylnC805q7rlm2NF3QBYsAtlHxVB2t/wYBCWFPSRFj
akkWYJRh84ApzC8cCHueEDW9TdkFRHuT1BUm7NhWh7HdxdQhPUDx1NkF7AjzGLNCivaYflOYtSbS
Aitd+PChw7itOVUiM9zi8lss6iFO9ijiEtGqT9kiHcwOPQwWIkVq07UyQRnLSRusadzMxQXifKJv
GkGw+jYWgG/c9Te+Dg05Kz/JeMUh9bDoygFnKWfu/pWdloyHUQ5uv8mvjVzX1y74NY8HAiSZ9Hbj
FVrfpLDz5YCDC3NoRBv9/GFoy29KWm01SC7a7ImWzJHa4Qbv+Rl7clEYwBtKRSjDrLRX2o090vtA
S4Q0KTPY9a/nW+V69+6ycwmQJPTa14wAaMUn+hAd58hcVqmvfSCeXqOFZF10kFPUUXwS5DsTnRwF
6CyzJQ2o9isBNcz7s8TGwlJ6ZyeRBXiF9S1fVF7n/NT96dhuYjeeb2WRFfjUgSeyfdJdKsBM24BX
o4oF9z3PUd17XbyO1XaOqZ8xyw/wBpck6GbuuAI/KNQ9dPXM7mszke12BfNokiK98vn19ETuy90n
d89G2cozMf0TPvXOzobYAhZfWqUONX3BTUTPhaWAExkSo5RY7dv2T4tzwFbZP8QudwDapcIyBD1M
YvXgkr6YHOXdD//FrquhLs1bkGG1Xh6eW1g1AL+tnWxYsUFXReIpRHzM0A6tiyp+UfGL++dg3wP+
8wjOMIXh7PxWwzJtv7GLktF2afs90imza8MR+7/k2L9f/f+2bZY1kWLDbxWERCMZPZqGkYx24Xgf
J2ZRks5+SQGa76fBCnfeV1pG+tb1KhHya4RuQ3ufgteXHKD3LlBxSyurkSsLWb3/6mZuxT81Xxy8
cYcGhifn8sP9TSdCJGXaJoxopr/yuUB7jTxKrwZT4I6bH3auoAn/tL/wC/icYsAIPZ/lifSVYeda
j8Uetq9IhssqesPLyrfux3jpEYt4NADznVCdRnkjqxeC+fy08EorkvDBn6WOu8+6INp/RsVXXag3
bPwB/+lvBL0RXcIrkjZTXBIzGkOEr4qB4Y4tgX7BRBgWT2yZXtkpZMLUh7QJYZoswwHod09ffxTu
iA6dm8PlI8ETXzJOR839Qz9v4hKhpyRjHo2wpeK7669LGGNUfVR8PH4hBTWCUBHevM9H8c0U8CVb
GGgnWB2vl0WphX28ML4aLZNUltYPolPrfAzFWAR1vwEO7zX8zMW1ljLFUue73SSOPmJf6MuleHln
am9GcydACdvXF8Cs04jPtUDnGfBrOeGSzyL6fUvYwodtlU1iKuUuMcqpQZhaKMkgVd97rCpoO7y7
FsPMT5Va7Iou0mxw/+VHZDw2GN/TcDianMI9dH+C5Dh8IsvRB2JOEeM7OErIUmPiOMJx5rXucFh9
IFz3z8Yd3JizsyQpfIXQBHgy5n7HKqOJN/43pykeD2W7/WRldWAJCpa6qK7OwPWzeuwsmG0ruU02
uOr7tWytMOdB0bhUb+uwmsSKx0GtgSBcbn6+Xgef9okl2KZ3W6BbYE16Bz1wZ1fDMJuotLEUZ0c+
xXOx6sWH9bESBc1zwgoqM8LaD1x5DfeJkhlhZhN3qrr9qK9a/lmCNoWLzLH5gb4ho6EuIHGULy9y
5aTUy9DLxGLFDd90Xzhd5r0zBkwdmdu9lS27Xtd3S9ixiTjhdUnYGM10R9/UAEgq6BYc+oWWjEw5
LQo2IFCoAPcAgz9vlUtDsQFpFWXEE9cV+TX16SzxG7lcgAxM2VrHFBTgj64OBTZE2IGSEGmZMYSA
H6aEKUL+UdYFCviKQtcOY8Rxxk3jIhel/vCBnQkQQEJqa2NrjpN2GnpdU6vPcctY1rx6t9BY5pgy
9egpHXCIo2MyYZwrIExm2QQ8z48QLlESbbcNsD1WFsvX5esIX2K4uZ1bZYDUYouy0mSIxYZ3iVTS
TioUR9tG0R5kvP4pBHPMUK/+RXk4gUCAfC5iGwHug4cgIkGJfk7ffr/TMKkuSwhJtg3f50T/S/0N
0A2ncGtdPFOuNRzyNaToHpYRVA9yRJ3JJamyNEwUesNKbHR82jFuh7yl5eRvnoXRzhtIRdnz1CYq
La1H0dACztF7HEPhvwrqbGFEzsshCIBIr6qpTAmPIRoPZCjVowfAMqm+MKOIC6XQ/dzzoTVmVY2F
1q5ZeTfSXNb7xR53yVNFqsTo7JDpbVmAWkyKkR+wP/lb2Wx5vBMFd3Q9a4PKLFVrThv6786fLbks
njoZ/w1lx6i3MdeVhjZ2Ti2gMxWNvrlWyiALNkmu7GgMr9LoSvVFr2MJf+/ZjgfHNZjZOURKmVeY
8rPH8GXfoIClVZhzSpezfvBsTsqcWVt6jiyLCVXgMMPQ6aWlk8WTLbbx+mryp3zvpzGKcgU28U1/
TMz1WhsdoDGxZiA9JlFV4DaAUSsOvaUrecgcckjSi8PYRwNz/rwSoBGmeCtKvj06NBW9LBVXchk9
IS3L9vTHnGKSBz+l1akDqFB9P4owdbcan5kddcBu8uqUuK7fE2tDwDrosN74+W1bRs6yo1AzUUBz
rwAc+LpOFHoxGLbSsEwmdnC0BPAX41ZRwGeL54ei2yOMZDeQ2I+vkvXRz0Bbh9wAERE0MElNvOpz
rEvl5ZSzugaHVSdvJ+bTALcgTvhCESn/u4GriDeTfK5bIssifa3y+W0pkntnaNb2hZ4sLpqxcHJj
ylRlI+k8vk7rm503ak2o5FZCAx1ylIBaHM+gglMYMOCMYRktvB7Cx9L2iEWQhQREHbvh9TkSHdm3
kV4PKZkk/uK4V9rXN+fcxt2pmBZtRpE96mV5SfkvD9a4QLM9wQpRB4XD2VdWr9/UHlVzP785Ftne
F1ywS3+55AEnXcqli/bs8zLyPgDZEDe0iZQgrrgvS/QrBVnN+ehS+ZJJyq9+Ci9Oo1JlPwYai4zG
Na72GbWw/Z265jWfc7HnPvmjqfK73Ff1I7ZWhp+2r1EQUYeO54W/D0H6jbBQxg75vBa/z+vZKUby
npnOdGvZ9IhZKYIRvB6jS/VzZgARuInXa7CjoAFiVCeB338o+BsqFpLTjPYB4u6Kcx7wnfrOt8NL
K+HKP/k4ylTNTG3tyW2dXWqlAKHDz68Sad9Gdjui4qtdK6Cpsn8o/LX790mdEhQKs3hq81FK7xHj
fylLfRGUwp0qOAmxCiA8fX/T8JEwQz8q0cG9ilHhKXJH9jUg1ryVWhi9PDQG7xwwyXQrZGmZDKkw
jueJOpEcMA5ZJwQtAouy8oPlYVWqoGjp2xV/H+hJ29KJ91pjUjOExyFRrn+uXMY6HaqO/hzN9AeU
6mH8xvpDCO7P+aSIP1fzbZvs4G8RsXDIzkPsP7NaI9Kqg6c75kiu3XLMcQ74gHkWSFwaOL6MATtA
cSwN7IDLizB+lt61+IixtP1tXct0VLu95GsVl+cAkcxaAS5dfuyWBbgNM9NXPXvmngZ38FMOA1ut
vhctjfdJyGjUAP4uWRLptH697erSbhnFJRPNNuZwUk4MPOuwmfAgeSodkM646abchACcK1oGRN1j
J7GQchRfmLO4jOKXDo2RJRgBRCyKr6zY0xt5Ch7P1G3E/vQLgJicVMEZj7yZPxxCT5rRS1eSn9ea
50Ixz2h3uGC7xnhWyie8bwCVqkJDOGYDt7+gSjWlrPEyweCeQMDG6gqtSxS5j9wY2FpE/yu0/fWM
snNfWQaalpTUIGwfbfuf0wmyYxlN9YDroqsT/aR440A2+i89ySPuAmxVKebQ+mPcyc0KJbSW0Nvp
/g2YwpFiulrLwUg35qU9lWpFZBBxPfc/naSW5fvCKsdV04HOkVpkm8qRIMNnCbcu//2S7+1WoU+M
a1UFA60AO/HcMWbYnZvs1LvxarkDr8Yz0chh/jmI8Ko9CPXRd3U81PuoCvFcS4f56AD7seZ1WGB8
an/TBO2gOZjAvpngvfX33AhFr2nN9En5OU7TUi2h1Gkt3wXlrBh/u0jLOm6QTngG+p+GmpX0aQCj
8Sm6nUd2EJkLQxALdItMqlntC4Qht9FPoP6Y708LNeLUCKLmKdbbZovb0P8OhWZKxK/iU6gO/9bF
un+Q0Q1M4KD1hxpTOBgWBYCFqjuRbg7PcXRZUTlTI3ydL8I9NwtaWgxJj7aiVaqhCbEjdJFQXEwU
lv+X0/HPkZOp4HOqeux9jVl8dx/Rbmtjyf8XTR2NX7olHb+IvdQWrvnuzl/cXQyymHYiFk3IowYO
E2upCfPhs4B8MjxivNtbmYs7PShsheFsNW+I48il+R1JZXMiCDPPHiOaB2D7rueHrMhqTV5yCDLN
Vm87HuwY6Z8cW+p2NhcYEJINuF+2gOJ1wJarp8wrI2AxLDFuvCwPkKA/cZ/HtzpGGPVyQXTIB7Jl
030gjyV5As5eRotJlrFETqVzxboNJZuMaEY7ftUGwop3OnIN+WxTcjPEuVBWI/NyomZpJ0oR+a+Y
/b3YOdTE8pMACm47QSofNYYeyHj7tVrE8/anS4IxCoQwaCO/GFnY3v3aS0L+kff1bDp8KOgkajG7
5KLeTkgth1KQKmnxFeD46srBW90jsbeYXBs+o6HlmN++pdWdZ63dRRF6rsGhj6woz7gDOrDrwVGt
VVjo4wuYO9EwtoIuHrB4e+sqUZLIULdOC1D/CWJuiJSbaY2TaHMJwCsUj8fCUuseNot67UfPys36
UER1L2d3kMtrxglLkcVHYLXIfUE+4JF0ksJA4TlRbpAcvJrUUZ+sYmKoY3OHrp8xhc8FACEgVfu1
duaPgSCAs8Ap6Ja2DOuFqy+qdaODgBvZhFzHrEOKmxlp2WM46dyVQHCow7RumayZevlFRg5459Pd
WtoinyLr272fIIEFDET2XPjnEoeBXcwkgaJfNyOiXMT/y+S9m7UYRkvZP6wvCc9DInOeJ4GZiYOw
QfkaNwA5zhQ7JkeM6+GSykenjadzydEE1liXdEq1iG1/nNqV/62NV/TV8+URFhtsZuvDgLpAkZTc
8xeYApSBiU1tCQMxU2HfEsDA5FLK9nbpz6kZyi/NbafSUhN+B+giCEtK1/0ZoIMa5E4E1DKfyk09
iZXsAmyw586scjSaWjPGVAncoWMvbPZ5iBSLctwGQON/J6/Lem5DjUgZqjsBBIVWYi4RjT/tofPe
f4/pZwGnmOCt+JMxrrxrrhUtDDPcMBK1DF95mWA00UftyOM3aAarGVMsgYu3h4BWgqZquj79ZG6q
G/VLVUkdZjYS33lOFkif+J5ctRk6AszxXsCD+jtNqVD8quKI9d9WKbir9JATOfkcPJOMf+wmG47t
+eqlpgrv24HBLPeS7nUdFkQKpfiGlVSq9FikF8Ik4FueNbnEO4qEiG1vAkENw046KFJcEE0IKWsC
ozlM7DMeHVFvNvytn7Ur3tQEv+ghoS/pAYqu37y2NaESEivEjnNknj6AYcAEvXh3r1hG4Jk4H9ce
7coj6REWyQSkhIzOauXhI+cyDIMdMVwhfHfjrtGOa6uwgtdfKyAKLHAqw/aSpixfOrRzYYgwfNhQ
XvpwSuq6orC5/smazbnCK9zXL6VHqKJPfPTXKyAZ9qaTkvfDpBJ5X49pJaxnPiy1leVynwutT//m
eZOCRPWXgaLmmISXNGrM0/7HOLkC6zJ7t26spCc4BVUi42KMwWosfJ7zArHadvIxH3ffzZfxdMWx
mwvZFw678BL/C5onaja5iEfY1WjvW9edDjGTgYIWNCk4uJ+ojYp5/wRzORputZfUEjxhhOHSbJJ+
0UscxRHFfkAOqqmZ2gy/708ZO+fWMSXdxnZ7c6xUIp/s1Zica/3teAVrb7b5qcN2n8TywoXM2BY8
+ak97foaBD+MDsenEeGsMAVdIcMNGpwmDl475Qe4jDT8gUH4EDPnR6894WlMGx3MlkAoH+vBoMiK
6kXKz4SL7s/I9gmX8Hi/0+XgZR6+MB7n9hSasmVcplNKKCpu0kyd1v+9CVG9JHP9TDo3owTIXjNi
zAv+gNyd7DwEkqu7gbq59T7Op9MHbq6jgqa3Jd8+LMSSyhhNbpHtsjnyPC9752q43of8F5s9dMT0
/18bZQH6cOwbvUEtecM4ZUFw/sqicOvTQbonljUUbvQeciw8Vr2CPM4I0mfDlY1CGCpWuHMHYUSJ
0KI0HDtthBuZRF3Hsc45sf7GIgSNLyhDpN47L2wFR7GmM7R+0Yar3XFulWa10lM4Wkhp1FDmHAJj
VBsJ5FHDYTVyTgVVCsogaFSNEuaVr1TRHP9+2TklUHMBnCOgnUZFhQ5e+lz0lwl6cIIpbbEe5uzA
rCcjf+Zlq+QY56Kx7iEzIAKpW1w+y18FJo1jVZ3HOF9sZ2298m+7xruEC5IHUYFMDiUHGDjjyxHC
hGSP/GCUq0eMSFcDR1TKgt1Ecj1faqOka8wqcb5h9/nsx1Ah9N4x71zMq/Wp/JehOxyCsJ8RxkTI
Znw0UShE+kr6Q8do0aWMxrYAdrkScIsXF6gHm7xuWGLzdNnioL6+KVxsGxGgJ7XFf4DoXORU1nFP
bxprM3I85B5SGhMOv+Mnw9iMdgBJyzg5T98evmSHmgd46dTGbdIwcAFfGAsV05FY/4181e6Uffej
vWvSg1qdEtJb4FXD+gm+42co0jkkD+pCocD6LfTmlYV+Hy6ympEcNNPOH+Y6uwkxTOzBsbVcsN01
jT3ShMqgN2hr/BRwFvXlOClv+z3uyTKXRTDTJEmG3fBqf5buDxaq/3O2Bz07XHMFfEr4V6W161Lj
yhvm8XIxuvwTarkQtr2kK+8HNvIVSSSu+DDH+BB3GNVmI75BOYo0dyphgFWGE8TqZ+FNR3GDmvgR
8yipcFbpaH96EEBTbXp81HUOBiaU6AryYeVcip80oySF9ZOsnmw3xGSGcVSVIFsqOhv16sGwZ/LQ
X0GXXoNWp1cb9FPr7ZhOxjPnntp93z8L8XFlk8RFpt9N1Ux6AMsz2fkABwV+y6Hi6MoQuzVx5E3E
SECtZ1ylLKDtJchPaoe+mz+ED+3msHCgQrbtWiAZuhmGNES07j67L72ZFRFEfnX3Wa00yCIlqkOD
hxy84XUK5uc+Y9utktmpxN36zmaOMOy6+G0Xpbnbt3viXm/Ts2HoIwLBmuaFtqsJ2JZ4i9IjeoZj
JXKEqtkQEyf3kuzPIcU+A4qWf+a371+D0RA9mkqI0yXCduoYYJp7YepmsPHC9GOeQMXvYZUId2up
/5PxmCbJTiFVkznqJ412UWENzsAZWPOBUAQMXE+mVmiwQUIlbhsTNbW6MipuEZSaWJpGuIafEdX4
8Hm+2izhtAFfK0ZDgwurL+dRtO7wDevLvWJOaPKw10uHxMbsFskflzj2TYEgmnNYV5KPcCPQ0cSU
INYA7RODTY/4MTY97O6W3WOkKJz20Nvylt5mfs3GVtSuDJ+eOvTruxJEwqmrMBB1UzFuuewXBxoP
MM2kZZpa3t3KWDN81ei4t8gwfXkQzgL2Y+r6AfPtrQR1cICEe19SEnoAVIxyE9N/jykQd91VtbI8
3hv+aEieXAvd9djpuxC57JcpySqD6X6KM1pWqmH54aCYW5Mxd9kAttGnxy8oLDoenrmfTiAkhEKB
H951m8ZWscr/hfwmypyjXwBTxakRbFZ1phAsJ5UpTWnyU1n+NxUfHxy6+M5mfD/DYWge42eqT72b
nN0sDOgX5Iw5SLvqjjAiGxxgKpS2GiKwYJ1z9aSRLM2byC1+ZXqOcmjy12rnkBP5x9bCqe/ilOJR
2HEvdLEcmyVOV105V7UwOqZGEmDvGigY5Z3Jbig3ZRG2CdaRsuOypUp8kSXkdRSHImMxLiqBq/U0
+kmWGjQeCyoxqkWDUFvsoHt6YmiTZBWldG7v5tHoBmyzrjqm25zdECdzR/NrQhjOag5JHi47+nLP
sia8xr/9QDwgsk2QN/RiYMkbpQwu140IvNwS1bN9VbZLfI/CEDdJcQDuSx7jYEcHIILIY6qcM5wr
1q6v1Gdrx1dCaHKoTBzXT7MN9OtY/MLfpIu1W4qae3S78ZVvPMFomzxHvueVd7KWOhAphvMY7aTp
ub9TFW308RQxkmyBp0E/MMnd+zlyhZzPUG4mHjIjsrz7Y9Wi/5Sza2zl3BzTM5zuc466p9J4Fj7G
0lMBOgfTDNDDrRngwNorzvmuX9mmo8qlMgcA9vbje+eRjofx0O8cu/rhUHqVh9GV9S6fgM2qJ7SL
HRuaxdf9PjXXy62d3UVX42+tNaKF1AQBR2JcaarJg0r7u9XzMj6GZIg8h6U00PnipxD5bEtmg9dX
gQSRqMap5DO1kf1yCiAXou+Wm7J1bcYkJdVN0uB1HAQGEuCmXgbVWqXub867WMsdRrbrYw6++Csx
VIrFyhOeGIGu2RAdrJjzPTDUa5DTSH2dEMJfpYMNul2cfXJw33cSW7MG0Eics4pELLdrG5TnLl5c
uRFBYQ5PWFmR11SPIRAcmjav3k+TQjsMKbBcFHb1wGp0bszsHLy9eZfLpHvsjgVuB9i/Pz3yDHML
W6MdjdcG24Mi/Vu1fLtQp0wFiJhYBGBDzZr/z0PgNjG8zd9JHuD/ft8qmqpdtsdL2nECP1AIAHN4
hu8sPT8ykyTuryJbWAmXJLaibXqEFYyx4hP11T8aJjtn9dsX7x2Y4U2HfLplmqjzL8HBBcP04NpV
lBQU3Aqc7ANuNk7P+dY5HQCVvl8IZY37ujUzEZ+nzEjNDJaDlMYgYbEvqViSb9yD2ew0H8A0PODQ
9o+2QLFNX54YxqwiQ+lHClhwSpSYofdkch1GkIvWBFPWBtJFLJqh6X6hrVuKUtOLvAQ0o6pFGXQh
bcbMkydtP29zGanYsEGbOsLPMS5X2ICCrSgGsEKLiARlPItlxThVxgKWUUnMzAC+jPpaZhmd6pWw
xaaE/GCtigumX/tHsGrra9szaAM5j6d/0qVCxrjwxzStwemTeRAb+PVkaa4qghSlhuSqeCCCH9th
tM6RxqjAaorE+XrQ++LEEYPpQS4TPGBA+q5ITPhrZjCOOtxYZFgtHNQlalJy/6I2CvuBzHyBB9FB
MGboE0j52YazFWtY9BPvZm1zbEiqOi5mHqFsd+8kUTojRlH0GYWOS8jrNBV5CSXEznZYi7H6f/Sv
5jltsqt5ZYkAQLhUQ/hMgGyeArq+e2n9pVRRYZHYAWoRHVAXUdBR3EcKqSqQi7r/s+X/hZpx8rOA
i93v3LMZGHaP7BmNPZJCCaVeA3q6K0hsaBrnW7/Q3FekHiNHWWudnBZvJyog8P6IK1ycQaI8CIHF
IqLQBMRrETY26Yv6IQpmNIlV/mzkJyZxTpAawAPKtOqTIZuZiQHxa4blC9ZNYuPVVMbJibwWZqo7
DWAWzb2l3oEx2TnQ7Y7fukuEVY8GdWGeyuihSkxZuA2oeTwbV95ccdiaG2gcXPZItHfQxMrY/dYZ
Xi95wEaOelnzKUiCudi/wckrWAKqlEUB3MUa8f7uzpncghFbP6WQ9wNBMq1oPxeaiAm3+NPB8CsX
XPTtMWDD3EiwC+oPhKHyOGqrqg8vAXEkAxqMCutJU6d+tAdWkNsjNTI4baTPFHgsRxOEYGtdZNr7
b30GS0piMPTahV7U8hHslN1Q8lvGKMlzJDGJ0geDtT2iqblkWbSzbjUp5pnsOr3Nb0a8u92oj0WL
nryiRTCBfMldREWEZUWGRcViT0ccLhkQG2A7lu7tR/Xa5XRsIp/v9im7oSkvdYsmaulBP/PYMWzw
Cr7TYH1g8WMX9bhn1PEEPSrKL7mSfc0Jgw47U9JTQvslD+dFiIOJrQe+vGI330vApAcdsdTPE65K
4rR2cpI+ZJOXLna/Rq5LKFdp4Uq+/j6DAk1Z8eK4iclBPqcjjuAvoE5LWchbOVnFasinAz/jbX7n
3DSEkqY0rfbMuyXz4XXPv8UpkKgpunRwMWLcIaYjEIDg5cphMvZISjklJHjLsxpUVMhHyxPO4B77
w1qemUj9704lt8Yi4a+qqWKSwh4Di9qN6sSYFvctlqgpDD9Re4q0u0Y9VitHLzb2qNg2wlsXbns8
TiN05j68Z5dZF42NVj3/d1u3Uj5qg2s+ZoZtGjwC9/6P/0vtK7MLrbPei1WEfQH8Ptp2+TO4emxv
kwbgfOk84EcscNQh/WKhFruljzPyfS1RCN8f8BInQhoiujFkMqzOvFuItsNEMc6X+FymAlU6+iil
XCnIG5kuSrKV9RzCyT5B2r9xPu/XTL9o6NvyefkJehXDn+mrGM0o0bxjkTmn+aB4Gy48eNoxNMAa
F12FzYrHwzLGnoBQXwugCZLyrdcwlO1Y0+Itg5zFvyBJ0hfj6rq/5qsqZb2Q4fDlkk1Ik67hBTXA
i0EhToEBYqxNXQ43211zojRSiyobBnnvRndAd1OxzHxl+J9tPQuAAd3EM6GSibYOkimg8fs1EpIb
ST0QtQ0tVm+88HmM5DoG2i3VNoUWsyLVjGw7P1A6/ZGIXx8H4wifwUnCfpmsUYcWwiFv8hCo2GIk
feqcDoui+0sDIFUUw1Ds9UzD6axBHhx7BCuufzNhdPUc7PzET0xa8rF20MLX27baglnbTgc7YxJo
FwuTYA0KH9dNjkEbWIkGykXxgx14X9eI2tMNiRGeKy0cJTiz8FG1QE14Pfl/8uMGSzsYm7QG9SaR
1Yy+yvVoNx+lx7IwkA/Usaz6gu5vyQA3irX0pmxlMAY+HSaGndbAVJSuVQr2Cxaht1VU+oaM6Ony
IuIG4UcsVf9emzy/ZdrctW0Nb/owqTbpLAQoqpBFRzs5rLszgrDV5oju1QAvbBtMdMjkw8wJjRzF
gXSqRMBRiGISrBYL25i4D4ucqgBQOROj6nUvtKOgXkkAuhi9QZt3nQ8WrypSiXAk8TGH72tqXleE
G3TqPBHl+pyXJb8MlJ9AeSKkFwVXZX84EevErb7/5B+XJ+fZzPgMdj5VudJhQ3zR8Fn9457VgWXQ
DnMrDlo0+fQZTLYrgH3orHHMDbPfm8xIS8b1KNTtGHK3RpiWcz54oaYQnNSPvHlXXx/aN9KE9bIC
GaruTiUXA8TjBlzBLt86CGEfwi5yirkFqZfUDMmSLqH7aB0bXDP7cZOiy0phCcuQIqo98OrPTn9o
/bpy/cd2R5brF96BMqkaIGzH1MQZ6SaOK4pI6lUfLfrj5rpO7MCfQ9HLBjeFjuJKKQfPid8B/zZI
9gl81M3ZO6ZrW0zBwC1vW6zVc+yf1/nOLW7641kmfR0R9WwOd3EOa1rkCxFa1/19PZ7Xh+KJuvFj
uBbFH9uIA9R2t9dBpW2npwxXFK7+JZEvMCdLcSV+ogi/Rk3xilqSdyr6uFF8GQjU+E5/rLzRp1Rf
hRERaMvxR6l5cWQI1mAeo6yZsJ/rKvYY9dYw3gQ5riTeuMEOEm9s3RtmTeK/52p9YCeRKRkkWq/G
ClEW8MbrGvG5sKRf+gdTRASHbqt3FwNu0wDE4d2MIQM9dXspUd0P7PVgsuFzeBc+cyXq0DLffRYt
ZUcdspgtff3MyPKoGEdD06yCMLGxJA3z7Qd5Uvj0Z9MqIidWCVtmVXu/+rJee80VC7U26COARDVd
VfxYfvsCQkYywNnsOErmk+kUFu+B9ex+zDOmv4r83bApW4zjcd5jL2zVkB9y/K6r6obOpYA8lj0D
1kBLl1QicucqzTTukL3bbsyu1u0HNuhWRPKBH5qwZn1dVb6A1h4in9XEqsouXc47feo+6T4+U0+8
95BK9nk/lCbDBWVSWR1PhRRBqXh0Myp32YgFoWDCipDz1a2Rrxomf6szCdAVM6N/X/sGGlzFMia3
gNdGrKsQIoHXNByEgicCuZ0Ia+LG3+rqIFdq7c5yGBDNQlq8/Bq1uOg8gjzimffXpyOzPIRrjNkK
QAvTL1NDoVcIZ9sQlA+Cr0wPHlGAAF0Ni3BgA8U7+s4b2k/WAyiubh0VagAAAVBNTrW1horEJZP5
O42lmYCKJWIfqbets+XdlUv0g4tXkq/7mzbi8Cb4sXvfKUIenEGThZ91mJwXbFDo4E2tVSpugAYe
ec+ZtRKJjPAFOlGLM2zzN4UHvBAvLlu24l2GhH3XwFjJWkWbLCwwEzW/OAMZlR1UwbFIzmrx/L8c
+LJjsszlEnSGWCh4VlEGdhM3WYCp2ng7e5SNgJvAPvx4SFqm0HrpD7/pGJG8t3APPPTlx6o9LNbC
2Px/2qFs3ZWAmSwytcL3o5Zj1rTyINfFlaLGadgdblTfV0nV/c7/FXTivwAGTjJQ74FXmfdwruPz
AjMfA1WwgkrdTbcdrRboDIAuaMdYjLwM8AsOnz87c5eRjdU6KVdYqjmd5WEZD+O7HvGOND/H8Rvn
kZWwNGGhzLUWStDtlypKfQhS6f7uw6p+2XzNzsoOCSsnsYvXlb9q0vDV/q/2BPvanuH8BGiwVVeX
FOgJbLMbDyJQ3PX1x5UZDxcGRtL/lbUSM8qMTlSjmaPZh5uAj77wyn0+rSlzKl4Qavdfx5HXDAh3
trWTkWOLqnvdvD8eQvrX0QObyZ6nJvfTl1EuDBnBNJuRs1ybQKfqOgMCYcIbvtkl4/KZrpnQJp47
0tWGfsBUWtmIRjWl2rZDAl4K+qic/xD9OBsKiFJklC4OqATrMDO7In+D+MNKe4ZGMl96mIKJK7RW
fRwuB8fqlE91SaxGfQ4kqMKzrHJkaeq6sITdgWGjJaf2Axb/Sy+aqQtQc0/KWIooE5wy7eCqzbZC
YUYzTdjoNEB6TgWWENWctVdxPXjgq5cAPpF+bt+amDXPuJ3grofIQuRyY9V/CtS/syWPFNVNMMEv
p9jANp44F/1zEyboyMdw37iKawrmwf5KxIS2AsVTaDSCRdweH7tR18EXeZ4UTtazsG99dqlj5qiF
HWsWJnghF8Ct68cziVB9/AmMrVP9NALZPkbjSwbmzo3gi5aRYR9NqNCaPQGf4ZUIuOcioRB6CKdZ
sisUOPgRRO58X10w77l8LM5RwJXQwkgRZHrMd3S3DoG2gKvr1WqYq3cWvRxbretnClNLH/GZOETx
y2/nlIVp76YucwqOjSWngUk8gW4WI16VKAgrOP4EDCsh2usWIQrOJsAiyKuA88ge+nrMkS4VcQUo
TygpBk/tyGTQGPbhUwVZyLxfboFshaw++cO2/bVSqweKJ1iHxgF2dOXTKMFxjUR+FlPo9Cgpj09D
zJVyb00eUK1IE0ea7Yj6iXw8JxAgiBdoT/vIYzCLCrRntl93Rqydblxe29FdSz6vIjxle6x6ld7H
yi6JBOO1EYwLM4XgTF0S0QHmovINxB3fEK5XwYglhidp2bhe5IkPtccGuhapUJv3gFK6TCNYUPkp
tLJF+CNo16p91LvUd6rZ9wScV7+DL7xdVQtLlDYAwS/V8MOpRKdLGIWp00KD6fMpSzXOhg/sIBgZ
5JTA2eaDzbehI/mNMoTDsPoCtph2RL/KCS8kNlX/RoFJzSy3F+LUC3lUFTDM2GxqWeE8+6t6sIhN
A1pEOngY28bT1yTBtWMLDxbUKyE8PJPQqidpcMWLWJ7F5Y08NFML48U9e2kWShoZKnh6SQratdzM
pXaBGUrWL8+5r2f9MTrtUjqr7SXkI8Y4O9esmFf5ZB2FBQet7UP740HSEMm+16LW0yjST+I7+w1z
+zgI9WNPcZMzgPsLj6yAJfzjLriMlEuNTv8+lXEk8TyO771CjGtNQESoESfo5D+ulnEASlaiFyIu
AIszjV87BuFGcb9vuLetlTcC+smohoK6OJOCu4cx/StJVwkVrMIAcVVIa253xFpkbCCEfT06Z7uK
9RcewNiyMx+SfgtHo7vfjspa48toAhWtv9ct5gZ3xB7hIbBqeSMdXW2gmUimdSgNXY0T50ACugBf
ovzSJ/pjZ81yvv/q8tnbBQ7fnP+lG3F9xK9bLYg55qmiGVb7RfQfrGgD7Rhzjm5hK766tZ8rDFcr
fX9kOGMR6p+APpPunwzMFy0MwI7YvP4SW5Qivpm6ft7m6+bHeTxitG9b0mY5brrHD9MXbMTE3VTm
+jpAoJoVducinF217keRutEZTbrKQnpfc9o3xKsWzAGU2BjiL+KntZtec6JGfay7LKNioEXdVG/l
6nyRTfcSG1NMKi36wR+DjM6skYXIfGCV5Sm+q/2Wtm6mXxqiI+BrigV8Jv7Xy3Xw4nLKSvsH2uHh
bsbZYAxBbaFpgiYoCvrQclvLuiQX3RKmKglqn7A0wLySepOoLBMeWxjNYFmrz0gVnou1RsXfEejU
flM8boFSFM0mqjfP0yQDoEHbxikb9MWDEM17J5nXv7fmwEsPDfsqCA01oO8KpNXZyIwbMEMrPTL3
PJbHjiQgJHM2VAQV7snXGqBHxCCpKGKLy2o9ouc2T4BkKfmLjRQaaAvAXyDQUMw6foO2HVa5BH8I
Tmh+hdJJCtutxaMlGwCZbG1A8bQ0k0fh6i0M4U8lsQ+QN1LTcGCEvyCOkTn0F3fvHmvSPvozxO8d
tgx01lBixtGQmJGp81ZQqcVvSsT/QCrH/inRUFKiOEV4TDNcit85WK+hS3Y1ZXB+E/uE+y8ia21x
pkoi7tb0gPf69zapNSiqjxIMLdBDRwQMeQh1uV328y71caEegq0bB9jrKRMRrT8HYrnPBZ5AT9w7
0tbCibesZ/32pb2c+ZXlre+1OBKZeNDLxcTdJFzWrWq3XH9dbwQSAu/4/OIVFsE+odDsst5sIcEC
0qq0phCEsq+wTqplLbDSyW7K6lvEfp+I5oTtmpm6klJbyZU8XU6jSO3VGjU1sHIszzyGVndefohC
Vo+92Ez8GD8oee/UPYYwn7Go1UyoFnJWW9+U32fbkOuIyQUie4LeTzivuYj0V9sWCSl4P1ZTDvjr
9rPUn7NU0tfoBsrPIpZL3Lq1KqDlKTwegw/+3wIudww6saas2Juc6khM6Jw2SvLJqTAZWwFCYvpg
6J2R2uvy39cP296c+szYrOetB0p0Fu8EQAmx9aotqc+kPG1XWmd9Y9ingxcMnaDtuJa7q2v8dlmc
YCHK+r2O7f7txREpvrV5EPHokoMJLvPDZZvCBQiILiLAZEZw2I7gIX1lEh/hfLGm4dKT+AY4BMew
HtCSe0hVWoBcPV/BpbmiSPye8pTDqDFMrJx/C3S4C2SVkNesldM7a1/l+jEG8b/8cMwOU2Iar2yp
z1tkbQmdI2HeUKtIdWrJOMU+Xh7HosPKQTYH/6SldpQuP9tAOgLWVY9c24ilbN2pSxskfujIdcOK
R/v4GyitgSRGtOZNgSZyp3GZ1Q97upI/rgdm2yoGoxchSK0vpPskU2kdhRn70kc/j9rqhu4KHyhP
Rjx9wpZUFDrf/fydqgNYN5RxdU5IxNFuWB3U6UJGtJRy0FmqliWH9MADsnNyn4dgzEskVwFXPIHu
P28d9549Qj/646L1LsRekdgGGpFQdKU0AgeC4Z5F/vdIMMOALI9wx8s6EYXbQhS0LEkjY/S50WMG
WiiSroZZzymWaT3sblPLl9agBzzjJ55l9us88WX6G6bS8ZeF71YEu4KFD2TzFhgN4PKZETr8979k
jXqzJoDH4xJstbUU4jj3GebghbVJGp35r1bxQ3As+9Qeh4G3sF+w78PRdB3Gh1xNsa1PZtPeN2MQ
OI0qm3zhcXK9khBqzyAJRITonX5/PHK7BlnhtTaqQ+If9uVPzmFA2t0/12mxMWWA4a5lZroR4QJ1
8RP/XlWGtmR7p68Jv19joHarFs6oi+wHo10hY5Tr8g6lCYOSzUAWD7GhGHFwgIK6nw3YcV1asmno
v2ZZp/1OaWAEeT8mtKXAYcEMsJF25Ml5S3V3yfm+zNSgq4eHDvxmcTbMDi3fHmIRD3e+9wlHjSK/
pdWdJ4ndK93WC/zbM7QLzOS4kdW84/z7nc3Pvo810UtiWJOKbaiWAqKWvIr45sDU5XEYKrAzlcRC
nqpU3pC19zyR69DJFuDr0lfAdUfXQ8WpXGG62saq/vu0cvNJgYi4jDBaBW7bD+QBsFU3oTCkhjLI
C0P5CYT+99LY2jB7zcIf9K1mhjKI3p/EWi9YAhHHVFq15AoHsUZuHkPqOZ96wiGT4/VJn8HQdO3c
s5Lt/rV7H/tPbXzOSaq9rALdaN9OPysl3/V4LoeRsX20+xWoB5XW5Qs3mvvxOaEkDXJshO5JxQq7
TheALDSYMkI/ozocqp6VLHOW+3yaXLmut4YqB6oO8lMhUWURh2Fa3CO/dJIyjulze1UHOTAa1TS7
xFH4RIWZ6jqMY6arI/s89jliQn8b1F/9eqWBUgdZu16dZ3OToa3j3awmYhdDPamHqeFvCUwkLIvo
Uw8OI0+nckBuBI/2WZculWs6cUZBf2JSMF/hxWTLQnwN9yGhEo9ZAuUywuXS/XQkzOSKzdcnyBd9
qev+Jtjvfu2Bf0IgI+0K8dSDDusm3lAEpI0iGlYEqPMoEB5McIMbjEgUmoxghyTh95y3UplFwOf4
WjS/UqY5C+rurbBchegWcKX848uOZH6FowaNRZUonhI5n2v03Zgy6rtNg5ptXsyxS2tqLLw4/HVP
xfXmgp/ezeFDnc6hKUYQUu6FXwJ7Ty9kp7SfxCGQl1OjiQY41Blv+p8cjTSPtvTnhXRQOFDby3zv
bFPE1kx8s4F9PRH4FIfkHJm05i5yx80oxZTnyZumsiVVda5K5DxY8c3Fz7/Hi4fayqLa5hyPdmDr
h3PdEPnl832T1pPjzld79/5vLuKvGl+uH1LycAw+mOuQl+lLkTzD/z7T+7rMHg/VTCekmm8ypXdZ
H9NBfPT1mIwARcJ9gomfwfoBlfh+GtDck3VLn+qVT7p3I3sK2YDbTitGL9fWXKzBWJn8sSPq3lfb
NlWN16FEc4bFz4OfeDAopyjGepPFuHoH0mfPwlIu/9Qf+JB89FfB+gglSq6EIAIEtjEk08Px+aEv
5Vc47YO0IHUnU5p7rCq1M1CSKvjUEJJLqEsvuzbWClmxLOOkaePqloPg+8KDeapXxzzr9ujLMAgC
WaU3RK59VsaT/uyWvFAhqcziwzliFNYXBrDE9zLTIqJMS+LMoEzgeRsUKHgqx5ZKTXjHq3bEnu0t
mSR3aNIolzp9aH7r2bHKxwPcyW8NsF3ydLko2tkwEIUc9evNwSTcL4Xc7edy3OJZnIBTEP71C+C5
mQmewvLbtazhfzFqOccQzmVIDF352AtlfrfZmoG5ZntuuZEfUeIlRZ5GTpIGAAu/OREIXRBw3X/+
KorS2nyX4NutvsZ84U9A/X9rgynsAX/LFnBOSg2pkREsIsSRnyxtqrnIAADvHL6eNF773E908qAm
4O1EUC7NUW7jJ1FGV7NyWwxs2cSAmvuCllGkfK9aJ9+A6XUod6m4hixMdiHwUwuRYwVTiat+BLxo
xWuSYwqA0pNpZrxeY/7c0RcW8QZ0C4h3Hsm/jlauT+CrzVLtQS4zpBNXaaQ8Cxe0KMXDIxrp3Vhg
uIeg+2iTZ225VHnu/KrPoI4Atl1ISCwzayIOBSMeoT6eu1FfuB4swwoGc2c4My9cC0NleKUMa5r/
QMFjMz1dW1nPHGYWWNItjDRuwYWobsskMSkWKnN82aG8LH8dK5ri7d84ABlapvaqmbKrVdR7INYb
rI45OMIpTMvUeEhR39boJACrpzm/WggTGev5kggwf0vBUO2/WP9c93Mqms/oTQbEX35tjOj6q31B
1MUZmSSam7r82Xt71cfZKapMrATy6jLwxbpPNtHrqt08LuDJwxTPi1Mg/b0SLZFNkd6eTGuqnKp5
i2oIVGI+9HH5ACiEgxIASVjIi0pue9utuaKZX3K4YAockv5Gn1NuTNAFiSlEeciuf+8Lbz1FcYer
v2KegCwpy5/OrYpvOeg2yyChKpc+/chssBnQTjOc/BaKJkNTM5JlarOTYlL15GjWa2Vy7uxa77Qr
GJ5Osguqo4ul2/Y0gBjomqa+Jna17rctT+gsrmc7m3eYmBuQN6XZrtsdR9ZXfUTXeyaidkyKx5nM
hBE2+Zh4o3YnWJjVuwA/Vco8c+zaIN1Ts7iYtrDixAa0WdQBBYEyGWma6BEDXbeTKXlLiqXlNgPg
ZsUOysLd2LRmoi9S/uLRsKIME6jEedV8Ht3+/83EwaMFZLEp1STo8zKsaiK+lTIuKl8putuDgqp1
EguUmhvI0UsZCp0F6jH8VtpgYuFKc/Mk06vuIREVPRXFHdYV+TYwp516Vmd/L2sJGt4NTAJujAqc
gfr3JVNn7ROIxosa1sERZvdZezSefj5SWQ2dzrjMeULfiKqv1uTL05WH9p8y6MmuspcPagqmUuaD
GbL3exnET2GURIFRobE4CylJ2ch/UZ/pnkVOeRacDBl4Gf1s7yvVoMAImXN7Kxo/F8ix6qehUxDY
+lbTonAMkABce7u96w6Nui4un5oNx7Z0OIUn4QNPZYIrRXu+Jf0mGIG5r17KTa2otjx5SOW6iIbT
2OC94yZzqIWtqBRDHIsf60kM6iQfP1ADm8iweoUFml9hyXwI9rsov2/WDpyM9eOjJJlasNsVjlw9
qzqVdZygIBf9hD/lrvGxoXPsr/hQZVb2JPuXdMmBq2X6JVKVge+Te3vBJjnzVR/UZ81tYp2q3Xv6
slKreI5gJEMhyXZHOnteuIRHqYWKR/DJxr/V3zC+WWCnWgakfaLtrmJ2XvQaFGpWSx8iMiJ2sX9p
DLfMlWHtlRQfv9vomjbyl2+AQcbPy/xkdBceNGtbQxIps8MxaXArpn1tkkEByVg9T8clyIflDhEa
XIL+8yRxypeYlcPQKFOK52no2jDW3qTHDkvyBAVdfwh0wGP0LeUdsXXH53M40BuOo7baXoBjxugX
3gYB2xvQnbYLh6lwF3ZnQ7Lsu2nt/V7snVW6WiX0Clq/EJuKSxIG8qxPa4z6tffS9XcBBw2wfR5H
iHg6zNoFsgBTWDpHlc4KkybqXMmsweYgF2l47/XVLQ6uVIMZ8ZzvZ49FIi8CwOzdWyyOyj5SdRRP
QMGWJk7t6d7bFjkUW3qRcqaS1MjHej1Q42kBKf7GIQjd4at7K7BLx+J9NC11OE0A21Dngtn9K2XM
zq/RaT9537TaUcN287hY9Y+1mZKhIjVk6GvzLVP2uyRFqQo9Bsr+tpfSVYUpoFyElWqt5k2aAu0R
MJJCDpufD0le8dU4mLJ4nYWrameZRxNJA2QRmTkjB3AsPHgU/69PPlHnCcfaDZqyO9zhPBRXwy+v
r5Efn2eAR62Qk8RJphMeIkNw9kuD4ACv0ukbzehCQcoiIqorfvEztKJt4W8OPd5VaWvd3MCWGaXe
QUbc2kmpPCLL43IVPBAlQHUtIQPhco0gCOKgrPTATz9VGJ4+XoDga29MiEQTL4kk2Y3QZvFqtt6v
txk4MCjxt3VlLVfDcTMYJQXFPXB4iCuNrNjQHi70aCvHC77s07vKkDbWEblyi5zxndgqrtAmhHZ9
KdTAtc6X6R0V6fVDEfI/iWjBLR6Wtc8y3bk3nLviBQ5tLDrJAM1rg5k6gkEiEWYDJyn5Fv8BU4xR
DlQLQAekl7AExVBAxNmriyK/3rS7e3LR8Nkages1+YM3QeMA4u9qyGnKs9hd9RU5JESKCY9SQ8pl
F6Ou6AE1859yQ9FURGi5AAIkHtqNq5DR1eD+3p7q/GuLH2HImalJcBHmUFrTRQcXQfTZlHwxVvAc
iADEg0xhCEqtqr982iAdVB+4mdkDESk6D2J2RzN9fRcxWVj+JtFGEnMcYdbPpHzx7AKG1PCBztRY
sXuYYytHcdoaGREoqgftA3Tb07SAjpMv6FjSKZw7yLbk9tEjMUMe96+ZfsrDwxnxcAuPT2o3bZYW
ndRtU5aGjFXt10FepOq8IX13OkGCHqxrXXRNt0SflauyeVKqzqhuvOtw7mDSQCuN4SVGgU9qwkJT
msT1tOLLcrIpvW3CimWMfoZ+6tOXdZt8tkDgukvQ1OtHGqBhV87RrHQbTrDtvutZhb2sS3HrJgt/
hvtpJ9WCQBwrTMeUb50svdkGiXwgOkebvvGqBbHZbxqShT6F523lzEx7oEQNXEyS03+m5UNuH2wu
DLIuVg11WyrIJZI4uj8A0ASBv3wcDfHPOY6+BHq0M76fOAT16yYAXrDfLwQYxuuCYn8MLMUZ4xrY
LFDvFfxYC+by2HoE6VPc1S/NwRHzItHsqU0Gz2LVKOL4gZzOcz18DGnFMBKIIdXgNMftCYnnl7Xi
nzkOuwrVLcfG3YGLNvl7PRxTfQUBdmgyyWktU+ZOVM68xhaANzonOwdhQFp50aM7pDyzar9OLmXR
4AZ2CGO6xWBa4dn83U93xXPtffEvuiFuaEfvWJuY5FGC87um2FzmCDTVfruCQ3rITU5Zi+int5Mq
xVyiKDG8uqZ8P+scAk6Z7OeDnZHiVwSDYh/B2dwTjLQy4EX1yHTmzJxQzZCWyVUc8Ef2aWDpHkNa
nSqEnCeVd8TjLro8dUCzdl92BvAzLpKYSHUTG/rijnhbe0CkN2unaJQCBqZBlNxOTuUmW9rls0bU
Q1ZcHOJhsKbTl6tAu74VVSL91PrKyLRoFkmQBFlMxKdm4URBdFsvHv5rKys5e9zgOf04lNrda8IF
kjXZ5BqeWDWEQSSDcQadDODy7+PK4x1LzLa1hfhpoBTxelHL0uIEtdS/9RIwEFTEZ3iXRxlR/co1
xmerYGyZ/DeMWUZbY5YZT2nvR/PAMk/iR4IsCORNqAIjuWMwtgTc2GZaR46JXZHaAWBErwTqpOpl
c3gEIj8WwVL8hYZ+IR+fW+5XjGMnxMOa85eRyNmtCx+1dnifWzCIw1+n/EfC7rZ4EblngqTK2Cp5
pNCUolZ0sfkLDIfqPHj/KHc2vwrijSxMNoGTnw7RP7Lo7OJG4yAOsic5ZTnD1mYO+c9g8elxouw0
iwK8Z+Sd3CmBB7xBWO3/F/Dj3KOtNV71iwxumzdW/gZ+BXsaWezHr4gOnYiqLyhFxl7a9vTq/1ws
OcZt2IJiEUUDVfoFXA42o/fiq3Q++3b3+eAY7bsT/lZsiv1UTVa71LenmlMwnPwdkLfM5qRSfoIO
f9UesemZ5WGfVsyD9lWVrDOBZV5CIxUiNrCdsOyPXfpRzQZajz0mrtX+nUpykHN+csjn09Pq44rF
Ug0EZVegIQBPASm/ptsmytdUuzUyOeIDRac4lWwtSW8d961A3FG7KtKrdd/1thV7JVxywcjdp0bB
MUyHrQqBK3JF0udgwaD3FzCVeYoYTlDHorMI7W7by+q1GDYjTBmiTnE0N0tTqBNEONYOAJjVm3jK
FqnPThe6k5sAboqV3wFEGJLd+1qJ2atTOYJbsX9B2wHaIf2mMzp5xpGY7CaXmSAuTNV01jflRoNO
5VE2SgZ31cbHKdQBRVTvlcyP4sfgIMp/dWpFdmQdnEELntAlxhCoI36zE2T8jTD5/v9nSOnA/SEm
y+m1wUiTrGDeOyYNIWK93nTYftccoQnVruorgiQIBjg0rznfifF1X+N1lvXtNC8zVVtN11VHpQAH
vACyXp4KzSmH0Tu4CoRXLL2pFfLpjrrZRRSzOZ9+z42a8eEDGxO7si84ypvmgHy7aiD7yomKQHQk
OqVcAMZgI+iCpS6e3A6O3wGp43B+luSAY8mRqAilBNq9TH8p+FSgEnYT2NhdqYQ2Y+b3NVcNmLs3
TyECJFtllii0BSXECAUaxxFjP1ugD9ILPq/3mBFeWmyAc8uAFIH4YL5oUT6YJKbRoyuxoTWcF9e9
x+gL927oM28QB2+y/MYadm91zvUVAwUS1atmYL+nN+i6w28v8824c5GVHeEifA41UyujOJbIY1K1
kAFYED7/j3+9Iw5zdGDdSO1DLydrx+rtLKLlXApZWNqH+BHZuybhvHAFZKc1eFlg2hToWHSooPkF
OghAvAtExqfBsBrulGtM2AYBtAvCv1PdGDRqDdbEl6/LZXOx5lv/bk//G953yNkwiwUu5KFVPntT
4PGBrCQtg7I83FSjLS4p2KnnTSA2+NdngsZXZ80FN5Fx9LlpTuYORqz2TKOTjpR5dXvQt0mc2yUW
uVxxZgYJdGrAwJp/YFe0NUXr1QARuHQe6hiUeQEWx6N3mKCbRj7lXJPQb64G7z0cWn2CIbM89bEI
/iNIWz4SjZgiHG/M+de9pzGNQS6eaGtIRcA/2pIIuAu4tZrJZxOWFLobFVHUZBxrY5hhZXAtQSQZ
KCM8xKT0AeLzTrABcFSddht43qfAQj9cRxATisrYhddmrIR9u7fCmBpAP+q/ePxPgU/u/4IMLb3C
RzFS8fvBFRHKS/v/DhPwcIyLPt8PtrgkvyYSM4BeISCUVhU4TAsqg/LhFUJwDkxJeXW6YDPprN+X
8a2bUbQA04PzPHdb8ZZvpMzX1U3LO3qlevsZO723uKgujIfNVmDQ7OAumfYkQY2g2gUqBwgAAn51
M1FTFhKJPBUeCLX0b3lK6YQzprD4QuQJUUrozRXcu1dNnZacGI8NNyPPh6rHbnVPDAr8rEghWS+G
eP4ZsG/CIQdGoJd2W1atXlMdVYDEMj34Rlmd53RmOXlm4ZBWAvxYPnevdXA7o+Gi5FVNCrpS8wUa
0Rdv2wQ75fFpzS/0NGGBXwPU30XtsoNc9GeMijn9e+qLTrG2NRh5G8Hq4BdIjDQ8XOEZAONmFzoP
4cuuQcPZka1qQofVkTrU+yg/PIfPjKVAnwSkVkfMQiE+TkQfvqRVlJb5yGvBK5tiuQU0iWZdnQUT
JYScgbFxRVZw4x2+3klNNRUzHpsFhYKiQDjgZqGboc9ubXKiLH47iGTEA/H41JNx4HSdRmwXbWDp
852mRptb5ufbsE+1M7Br2pN0j9r9Pld2Bk45OOdQ04sL6vkOPlBcD1SMnG3SLfd4oeOnVwimGpEu
o90DviQYuLyIfh3ZqiBof2QY7iul4g+4wg4Snc/CU1AirjmN7jbB3RtKTonOZEtG5+EDvV5wmiuS
9onNDI2DtJvCKHaKzs9BZCQiXLkwqzBl/gdJaggUoLWo6vWJ/MNIYwALqR8Svf0mn1Y2w4kehJG8
LFJTAVHv/nTvj38/MuGFujpP/I4RGmwI2BVyyiH8Kzu9BsS3lmVu45Pgz2ttHdcTevW7xw0FMgkK
BPEHq+8KMdvk4J3RCjECTd3VfQpQoXc4I2ReRn7Ei/y0wMV5nv8TKXNCOSp8YQq7OsUmFge0xwNm
blSmBjLjWMsT0Eldg9XaNr95xGXKFUDWJ4ZF1NeEZrXIPmMjyi1KXlwnYXK3ZkbvZGHddJj/GgP9
yhDVFwj7YT5wAp2CH2TzWcrorXHDfFin1KJWBus7s6bntQhiDE46YTKv3unzfl7L9UzvFbOfmF5a
dW+YtZZdQDe1ntGS9MkfL1XGlAl1xTQzRKW3XQFityU4+ZT1KLeh8fnO/f34goANTsiL7lk69Cry
kJMeZjo12wx7PNe7S3l8bgHb6iMVgCqnZ5/zjJE2n5XelDbY0W74QZfDHOBao8mY1RSdtF02DG4C
yJzc+G/uzu9ZRG8XqLIsg56td32DFCuwSfRSxiSwdxmSkPDs9kG6CwrrengyQGhcM+dvApsLAMMf
sd1o0gFuNcu+lP36T9XPLOd4fhMFiqi+9PyYqGb5JMuHneTlePB1Ag+nfG97M/+1JPaT9ujqoggA
GUXzCKfdyWWuZXiT0MkOAX4ZN0xVhYF/r1I/oC4Rv70SjLVoaAMTlmIFInMXjgUsxJhvlZjgagNa
XvSOdK7IvNbPurAhwCT/6p11P6UuOSymgKRJlhPqWvlo+g1DqeZUCR0WLodPzuOCU5u5l6vexO0W
f9iMThMGI8OowtaVZ7RtP7ohEY7Qo46VD3EnYRKdDixqaZd+FjxsrHI3T3P1SZi1Rg4e5EYZ2j6s
5NtFa86agWZQlQm9EiuEirzV+/WFe6+TFcqxBef0RuupsXDyjYzdRudQqA+9oYp0Qo0ZzuFMBkB4
3v9pWSNehAZ5SVRgAaMpdeQvSXb1VOPxuUdcAX44b69FrwD4lKv7tpWHPn9fWS81FUwsJzNFa8f2
VrPt9qcX2T2btRASkxbQ1k6QQ/3bKHxkcEX5vxrsdNuPFugr+MtsfIktBpsu1AoAMZx5ki2hrdcR
NPeTsMvgCpOx/6Pd7ggm621cOP7aQGzz4jtxVLLKL/tjc8PEOx+GFNyOmkbu84CGo50w+KA3Y2B2
4TOfMuaq4wySQogE+bp6RIYtaENURVaQyBM0o8fVqMpd8mYCz3dq5weDAxVwiaNuMoh8at9Gjueu
PpYAZnQD5EhZR8ICVrFEznibV4BlM6IZZ85eR4z3sSijk7Lq7knZZnx8BKaVlHP4YACEqCDAWzVw
SZsMCyAnT2YpAamDjerymdeRy5QJYJUSFWId72f12R91z//Ek935HYF8QHUip5MvYBTI646V4sq+
QtFEQDkP4WPA5J9Q9mgP9n6no+4gHxBlmgmaJ1tbVVJ6lTiuSBGPXH64s+xYP+qxmgHGjOQdNEDr
hDb+oPIy63hB5qq7zK7Vyr1ab4izvJAO8OlEU/kKc2vmd9NZU2Y8id84SdYTeqppXY/IwYi74Vyj
43+L8k2YvsNwVgzxMPu9bMlKpeRpYzxlQvQzNIvmkxNuxv/Kn/YH75kjGM1k0Y5/i42vOjPuzwxJ
m+t5O0wcIMnGt/uCeCIVnFmZH/8OkTzB/HDAIIu5nURWHLKYgYwAsdAbJgbdION4tQ4N37oJ5q/P
a8w9OxpUj9pGlI9N/UiilOGtIuQRGnIPEZV+dB4PAJGamHONaUDCDRmR0e/TknSyw+MebvSn99sa
nZ2Xt0bAdqEMv/J4PiV6YtDdTLRGcJ26+6tKFcJPVRloaIIH7gNhfWZeYiz+b7XKzWaHAqnDzEgT
zyKTdTMfISoXquTnZ36ATNKwRixqFahL+c3321FDFiVYhZDmAek5ABco9EMZAaj0OzoZi4qP6mKi
aqyNTWW+2dBMS+k1Fdl64G4SUIXRlRxnyVk7p9XaQ1unsaerw9ftWMlTHQlWjEsSXzh9gT+LdZuj
K1yO2lKeZSv49vNsUwzm0Ue4P5lQOSwNuH7dKiRwqHoN8Fm89AU5OV8ZFffUHY3i2OWnFpbDft3i
YtyJTodw0H+YzvI/DsgiluDQ7ERXQgk9S36i2wl+yZtyqOUlgCgxGeLBRdFUxCl1sznaAoCMPu4f
RxI6PPNLJuJEf7P4b9LRCWNag+fks3jVJ9w2CmY9XqYptpLgY5iuEhgFRNvVZyqpQOpi7fYmJx8O
u6cHK+aqduUxa1axso41G6hIJDL4KEWaCOQx/V+JC0RhAJUiXugK/RxIrsqfzwPZlw4eNLJbz0GF
ru7bzE+KPNrBlNmqTWXrES3AvN5e/BEjNqfEQSsg+APD+RraaiX0MdoYEkrg4DL64f1C+HsydlNp
YXgt9bDfyRg7OC+z3DW77y2KhaibPjilcyoBV7JjRFSNEK+knVlyaMQ6IlZG9kUCnzAaVxPVRG3p
nt+8YSKFaPKLrHetNUY3+OxKSJvprpEF0VTftdlPVCzrqDT2XkeH4vgKLPnndiHkrYNMLyFUFFO/
S+7NVeoTAXHY7NjYFALTmwePlXJxOGI6sUnVpVqPi8vgm+C0Xi0GloeZl5Q1L5kkootfvu43s1xi
Y23mmo7/vUxw7quzpI/+ifEE/nn/k0upArvUVUIzYGC8d67IU8/27zEedBeRx7nKnTWrLn//WSVk
D8shtO9Kauxkd8g570iRLT7fKwLTPMM1lSY2sY+bRmKXIixxOSU1ove6DOVO9aTHj9qrKqxyplLv
GGnK32z+YdyR1fIxChkzGbcFQFjZWRi8JoaMRDU5bz+dHrzQ61ekMsjYrpZwkOdysxfG9Pfqzs7M
Wfv3TPq7wcFNF+KbG9COMupZsNjAl6peX0h7tZ5yA+iR7LVW/jwx2lUrp1qLgU+9nY+0EqJsTNQh
LyywKmiIJgIN0t51doPmH6dOTw6b/aSMDpXe07MqEjvNyV4CI1VZ8rfuYlLrhSGad8mLP8HpdGT4
42qRnXys683Sp3238q4M32syEuEpMqf7nDhJOMpC2Qgt18hHfJnftE5J7bgAyFe6+ri1uBPZwUMM
vPtdKSSl++qGBnN/WZKN325/Ao7pDj610DDiki1p8UMjT8APj11feWWxjYxDfhUXhJpvcazE2XWd
dMAnn4jhaPRQhytYBM43Z2IYvQGKYV3g3S/LQJLZ8iK1MYSfH18OIH6WpHlyoe1R31DQiKe6C141
QzXUs5/DGekQ4FToMkfllLp9O12DgfYG5rZIvldNOXmfAs0Vw02VwHQiRNPKuQrgnmSJ0n29htJc
AAj+GQM+C3txrI47q7NLayDD2RTjIgk2IIBz6n5rw45wwiCjYHTiTq/+32DHT4ostZ1grIvyFm4L
+pUgudO+h5pav9ksx4D6vNl/8lYcRqY5qXGnYc2k6jgeWIKHTL4cW8AAyHw3Biv5iIdwSmdyk1qa
je4T8ZijZqzz4ZVA9CdFT24CGwN5XE91RKXVwNOw7OxRzd1UK2mwr9vIiYdO4cYX1pZqBc9G8Nbo
Yj0dyOV+ng/l2K9ursiN7g1P+waaEQaNbziM5ezpsfE3EAShjwJcKtUpabEB4zBAeQ0ypXjmxTUU
FSbVl9cT6FXLVUzRI6taF+0dctNubAQ5eZgFMRHWjFy4Q/glp5AT5twApeW2IhadijP8370pOG2H
ROXWz7HMJOmkt1B39pIMCeBabL7X85tyeunJr6V5qooLrPhqyNvEMv3MF5zYq8B1JbrbZBCtI9SF
Mkt1V3KOWLu+EtHaM0VVZYyio6wjpHY8e6e1xjFJIweU3f8HZxLFRYUhaL5w42sQVp1K/SGReggR
aKnNUyct4Grf0J9HQ7n6HZ00zueIV9ikZ5XG1NsjdPNbLE9J+yszRQ1ezx8TN/2d6PsdVDNA4pVx
vXwlixqTEmIsYGavfl6RNFkjYj3xb2S/h64oiKzl9A9Gu2FTrsoqC+ssB6YjPVVmZde+kcquNPPm
+qbLQO4QYY2FtYcNTmB2lev6JDPH3H+KFD/w8qOx8raGT/FTpUEv4JIZCIHH0uPFkZGxF1kpiqYi
u5FSCHf41o0DwNdoKGKSQc6BMRKEeZUnTF08R7znG/ZnAjJgHSj27YLSoQ5f2IZ7b76xsN1ntK7r
I2QJEphEaFr+H9HXSVhrRZRycLTkNpGrHlLoRmDVxMukdohRJNyijW6mldDayn81QJ6tWRJTKsRF
CIjpUqy73hVmBRaJnUP6l/LHhoxSZfirUQx4fp+3SkXVqc0i2pJVkj87AYIYnkB2QdTN+WWQE4Ph
oMZk3ZUbbisGIofMR8BvpLdSPExRzBwgwunx2Z+2A6Tk5Ubow48NpXj1Oaxy+RSd23sFxYylx/WC
qWNjDWVWT51az0KWqBMuhgmFnrrUAlxm31vFb8dGK6+KvZjaCc56x2e6WW/JY/AkZaoqhYoPIyNZ
GFSv5KmMmXwNvSn/2Mlkbx06SKtUqcZ3SAEjn8wlcZc0Gacm3yvngKZ/xFNkZN7GJOABVtmtLSpz
zsmvuuC/2cMUIJhrjaYmOuVAHOJal3y4EwhpfaquVVbkcA307ghKoOsN9QHy3s5JOiKOyf762C5K
CxC6fRrLAKDwF1Oy7c7tpLXXB0ZfvPdZqhepmoTcuzQ/p+Ju+ACo6UBUFrXFKCsqDhBwBzWtG5Ny
NsvaYoFMOvrlntrjhr4I30q5nYOBEflIvsW2k+rmtofBegzsICczBMF4XKL+sR1wrt+bVa3VTjy4
tzDVYNIt0OCb6vJGQT2dIUQKQT/IbauYswLa41J4awYNHMqH27Ce9WKkFfMFu5s+u/7XWaHEd9fv
4WKz3+GjiO1A/wYX1AnBx48Ii/DuINa6Nw5QmGDN2jk3YLEPyHeHR5nwuuQCFURGx7jzRnRCq25F
PZtZU7aMlbYTf7waTpcq7QKXZ8er0JWiol/Tu+Ds6AOikZiTfEEfDfWSNwcU5qYsKfnMmCwImN9r
8gvgddk68xpVry9uV7K/UUBHjVEpLHZF+EwuNwP+aH7ozBiW5XOCnZElZUINInllMThYvzt2r78O
9fZoJ0Q0O8a33RMWoFhmSEtwDusKj2g9iVFwTIIIinMg1QSQ1JOQvAI9sgm6nh1JESP3nIVu6fKT
Oqy4c34pgLL5xvaC3jcFGwDLSfF2AQlbBXzLYz8daU9QMvLGbo7BxBQazGm+10RIS5TkL3YiyhO8
Qs+mtu61Ezqj54317IhRP+xxxJI9sIelfdGc6hWIWUgq1TfNpjMbCH/Y9Duh/Ww6wqphi2toLOYY
6Sj6HVmR2MmgahZTxcYHC0sI5C7HnycfBGeTxpoj6S5cHf/NdqOf6++Q4Lh2UEhbAZCN/Vuqdo+e
dmEUWUIebOS5qhcd7zvReWvPSP0SwsMrpjH53YwSprGJS8M1WzK4/dWGL57wQ2/lKuCD8mwak/1Q
uFRggHdfemrfoNW/Ful8ZeZvbDp7G6DCFStlAXLvgAnFOble0myo8nEeJR/LZr7otSQsPpFt6rdz
lYpetB3CY0wfdjg8sooCPPcWczKwhws0dO46KVwfzKGSukCEYG+S1dk/IofBWDUO2utxwbduh3Kl
LlgN29RQ3SweFFBpcjPEbqVdKMb13aQq4rNRHTed7u9B+ZYWN7q2XOlRLEy5e4aiaSYwQ3g6Ng/C
aMnn6SJve6e0DEQg+TjvRk8z2Ys6aQW3oWeNQxbTpoSzQFRwOieSpdq6humUeEFKw2e4Sx1mL5hp
LBfDwdfFZ23GN/vDE9jpKCdclmwBJvwq+/ZcT0pl2M579YYGo0P3GPraogtEBH/1jNxT9Y8eD8PQ
V1p2pt5Ptp7tu0TElo3uMBVexow1bCMx7gQBDPhIuYW8xiz/at54B5VxnDGW3DaauTj1TUMWjIvV
UVyRHHjURtx2R1hI3eaIGLcDa0c7tqq/3QEpcAPJFVHPcthkKOKp14ZcXtUgR8B6ImO6jM0Axhpi
pWgm9jndMFuPxXopMKGEQ3Xs8/maRT0bL2OZQhmvVDCmA/phc3+zbjddm3J+c66/JXJ+0UTm+OG9
bc+i96idlw8AjvtT4htKgw7CJLS1sgNfgNbHF3uRYUU7BXEfL05ICWp3ridbjJvuSizv91ZPFa7k
SOT2wAJB8081Rt0NVr+fJ5x8/OUpolJLMUg3kacWI70IeGXI4zYTUFtPlLKFQCzNZ/hVxRMRT/LK
nuZYm2H8Nye5FMv1tasuzN6+Ce38sf1iD05/nDrWUeWp4AvwsVoJjVWgOegmz/oHL0Gj0QlNDq0j
7eAszFSbz0h9FZRJ+94s/dLXtGNJg0QpmrBSvpldZjk+wWkTC4Jr6QRrfRZHoOoYf6MTnyufyh0j
b4RzQXTelDs67hhB5KsPi4RgwLVotTMCF65jVa6KJkh+RG4u7KcBltdJl4iHNqJqYZPz5b2ZXj+X
MOsJk1YD56SBPbvyNyhfDAyjnkNdQVFNz6JpbZ91T1SjIwouScHeZEbPz0QSeOdre/MO7+lKEqJy
htPxyIT3rFCTwUBzr8ulBB5/wGq8UjCVErpklvMx7Kskcn+/iTj6Kq3r1jPlvJaFbQ6ry1Rx2IeA
14mbrgH04w6gJxwNe9RtTihOhhRcDiCyTA4mSiY2/xFEA5DuAvtMJ525RUXMFW2rzWvdfD+X0ZYV
aaRLN3tZjvqhJ+7xmeIwiFHIz8h1lPHzwkrjtxvVA3SLaIbhAhFAzl7QTAbLCjb7+X9Clnz0uada
IU9sfyNJd6RcZaQAanGfWUMxRHhNPwtc4jPm+MJOjFdtO4D+NK1ogZbe66S+3m4N/CNp7RMedXrB
4IOLcGRwpO5FtwN7ey633y2JNN+JDOm1FFZWS4EVnOga2tsi0iKz3uR9sCtZ82GBj9GKnPeNdzp3
Riu+2DGCa8FbraFS67Po6yjUTR1FQDFknu69DiHnQPZ6dRz0pdgA0DLy0Rr2+H0+RL3Y4O3/MyPE
bum5QE5pth3g3Cx/mYQS0XzuSZ/DPpXL7tBeI3mSRc0RhsE9UUQBfuKju5v8TKNXV4u1/7jY1OB/
T9inLiP35Zri1vUJdTHhC4HLkEZ0qa//Jr8cgYKpgPPCuHgatob6sDpGhkcL4K2SZSxU1qvqGn72
OlmCgb+R8ru7ibPeT08WlVJwT7OdcxFBkSqDJXTOkhBIl0YyUNBqel2cnCe8UHu9zUfjMPCdTeJr
W1O3WDSFS+dqLEHvVhs9R9xV8l1MwqhLJ7O/EF01rfs9+uoyUarLcqwz/l8fyTQ1YLYbd6t6G/jB
96Sknn6UBiuG+kCWvePcWV71/a1/ZGfKJUs3wQBZtlLq5hilbTqQDgQiP5olB7+uN7nvy3PzPHqp
nYEQhFAjqEAdg79UUSfE6j7EBW4OYXEtCC1m6HjGnF8CnMMjAxCBFIzdGN/E+SWyKAr/unr0N6E+
Cm7WNaAZY1GqjuSiKBKpy8ZLZi1aHtynPWA44DWVPqXG/VVYpT2so7pJF0mA8gzO6BU/Mmf33BUa
F2pUhmW57IoDYCNshTp2jFONQo5Q484ooOxwdJzgFEEznmeMOoNsZkq7ZvtfklCtRxdwtqNcz+U/
7a4LYW0LujcCov0nWxZnNNPxRu7PTZookBEs3wNhdf3ueIVwM4xRcs8yMrHTwvW/jAXFxjsKcvyU
90Z9d4NoDdbTWz/iSP6xrCgBfYl165sfnzDRWf9XguoTm6myJ79byEBzrxLWzSyD8gXlFfWCr8fa
42hYceJ7DyixTLuW0VfowcEAgYfHTBcysEvWXKznOU1pG4jxN5fuboN76X58lc3pCGF6rYo9MMFq
qJkuoRZsjQ6BhHKo8A1cMY735aJxqXkA5cZpgSO9qRrmfmiln8z8EAGsk3PvJjwBiZ5mJOgmK/Iy
CABSbv3EmQJ14bAoXf/i8s1wY7bFqWCfXq9OgAphhCjntmwQgGO1y+hraJsATkAYzPoCLlfZBizE
fcfB6HqpyKlVRz69+YAaPNSs+0c3Q3SWmlh3q1unbLCaH+VksADXZIa20e8Q1oHAxjkFYRzQxQZ7
WAHtfyH+Mi4RXFwy6L+c9hJY5OQUzE2mRfDGRjuahI48s8pSivjtZ0TFlyPBxDkdbBa3I2NGOsij
2evGrOyqS1Ua6C5kYe0vT8Hc2gjrC5ZXNmWlYnF6XTLpDZ70+VIx7nR8i1HzhYu4EsVVuGL2g0Gk
EoUidn1tiUyDjs7zTDC0AdlUcVHcS4QFSVcP28QEAQkGIiseufgykBLkAa2Z9O+wTQcKwYfTZmaC
ECyJp3k87rGvWX3P7PFI2jl+WIwNQwIpIo6zoi5x8YPA2ILHWtbXyslkNJoObXS+zLvbvslQHIpp
LTBoZyzU1OCwbzJ3MfF/tmKh5Bnk65JI//K3UUf8WB+HSldr2f2+yGVTGasdfAllbIviE3n/BQtR
9IhDH7EqFe+kl7pfgQW94Ixg5xAG/QJrrZbc+EjsurUSm2BYMImgJFNutbwdDVY2LZSA1F62mVdw
jbWyuMS2/VakkR5BxK28eu8E4BDyceElFMCNcmT0GKlqbdV2ex5QmmwLY+Z+BZDVmVIPQZWaUIy9
GqoGDPaZOLvA/Vpw41wYiAkGaRBWpilD+6UG3jw0kWocPeI8Z8WRMDegorwL/K+QG/E6FUDKFuuK
ddu3WmFwnKn58t9eeoGA1M4Us1lNYjKK0M8fL/4rnKgJbu7e1+2yto60uRHwESiCWGD7Ic9Vz0mU
Km4vwarD+rRX6Wcf99yEmBI+LUzrJvGXPssmqTrYKad7ep/ZlULPyzcofgx/BnCU1E2z0zwoUMbp
bVbjZkNv6Z16i38L5lx3lC30XQV+PI2aasoKlE6INhQzGExFohrwUfg3SJsgHEBNFtHlpodY23Vx
udhyfFJVZUH/9fHcZEW3n6j8UaV6LODnP4VVNpWeE5xUjlNCIxaV6msqURDqUZqKyCej1PqbDRWW
n8vbrCYhHnlZzjLyMUV2AIRlbEebGM4DuLQwa7is9cks5V/Ky4NVa6Hm0LyCuKU4ul3iJRa0/BIM
5iz/4E9TDC+Br5Nh8L+edlx8KX0TLIZrr/REsvmPrtUrjccBN/S6r/CUI05iZsRGFtf1ieeU0w0Q
PJRRHIW+j+XDBuIiGkI6v0pM9Xa8dZj/ElwRNgZjAjna0FX+wMOxci/eLckiJ/DsSUtP1iQkSYck
bN92qpSU9S9vdwabUnV3RU1t2mgnpCbWSM48hkpSt4wPPCqL8YZG9eBWHtA4RYT9bPjQAY97WN82
RoZ6Y6GIFH7MxfOXfhc/7ycyMyApKgg31XaoLDAYdzmukjP1CDNRJXN1nLG57eE1CrwoL42FXgjd
/4024KXtCD6jogtoiYxMt6mEq7oetZ0/36GzdqwGWtmyIoZVWsieibgNws0xUa/wo9rI9Z/RChcF
wy7WQfKpbar0HPDxMQd11WgaUMrj94lzBxH7T6oBSHU1rA8oL/26KgLZ/UijsHRvsjsfGmNcvTnr
LbAF2I/mAGrBPQaX2mqii771KdR4GUKjPiyxr9c1eQ248uIIKBY3tmYJj/X99hXZgrDEeTzlHil8
xmoXtAg6rQ7kUYXWcItEp6sXLGd53uMtcNWZjz97qVmYii/hKvpm2GjLz0L2wMsyJH98g/nrTTNk
ae2CwJxvLc9mgoXQEXQPvQOyyjimHa1fOnLoihz9Tq/C6YMSJGh9gJGzYTByIg4cZYlMr9l1xuLQ
DRRlg6Hzzh2X97uzFVJr5X7+5LIsCs+s1LCxMifr8C89HHaV2wqraYIyfD/6BvFUexHwQncR6fwr
LB9eO9CtrZbuf28KJRM5msvN3Y3HS22Ww+ENccRtovcHad7LQZSz4am5O1KtO/VscFPDdbqF6JMT
k1G28wLVObUmdFJ6gY4/GkvK00J8LS9nBk/BTcR4//Ui6zy72kzwzN83h9vN0fxHkkqlz5rYL024
bNTNzA/8YUIOx4rM7gBtJwCHqDKC4GSHW1l6o7Q+C5S1qDZg/O7crPAxMzTQ+PGhisQoKppGdBJS
aew0L7zKojuHfqq5+cG9BGGUz62KnGPtcz357OawdsW3xWO1lGakzO/MCg+X1fcsFSuhANqlkmrh
nnvY0S60eMuJ0Q506M24TBqvJ3WQya5X4Ci3G4V5oGkLgOPf5X/4kxkCMirytABjEev/fEyyEY25
7rsujOJWybUfx7wHWJyrnARxThLdhtrTaSX5cwbpGMNNwYoTNWn16CZluJgxGtdkpgRlbliWMwp0
ljZ6wbTa6Of2SkHtHaJBFmQBhP2Kd47uptSBsYPrvv8A+WhSN3PrfYb3yZ3Nd6pj3UoU7/h7nzq3
qQEJB6N5TTzWDkZjc7v88t5CdnlbXIrgxQnT9UkQZ5+CBrAwSB6u8bbMLTRML7bFs2C2XX8fdMhs
w0IXveGNUNFndEEnezjH4V3AcbQT90CtL9BFmAy1Xjjr4YMi3aGktsiDx/NZsrljLTw0AjPKMEaP
TiYRDQOXVCbsXJ7yK4YNRA+k+SS20R4BaVqK4mvXipV+tmtWfnyiZ13IgT3PlLKiQRUs5xfQ+p0g
tvwWKmrRx++DaXgIdmBDswmJh+IcIBeWlTSRyvpnsaTbDdnTIWTARdwB2KCWDY16T1FCGHd5Ns1t
i4qVgwSJPHa3q+uA8do1Jn22oGL2oqAGBlBLy7RldK5DG0lcMVSwMHjN9+vHE6ZOxdnbR9S7CjRQ
CR/vcPAFLw+DoTlGfP3XzthfObT//2b7lS1SFIpVTxePsBdw5H/C9oL8bHjUKZ/MZ8HuFr/R8jZp
cZ4tslpvgU87pJAQkGhImuNH9AgDPSfn7YM5Xo26YmvNFydRn0tnE7CMpFGvz6R8JE0xyUKF0LV7
nyybSBgC/AvxXxaP9NHo8MwMZMAzSPYp19WbKc5FptU1kKgDNHBtb6OMwkSrKLDTPz4HerlEg31J
CZWvdUgae4rdciqDNBzCW8qfM5W4KESe03tklO5CIb0RH5Q9OPq9C7c3cvwKfF3LUyle6l76tR8c
nd3yMpAbVsv/JzV4EXrbOr3bOILK+6JvhJZfDAQCX1Ykm9nNRaTjteiVs3fYMmwkm6BDcT0u9Mg1
Pyi3eHuGC9wQ25ozEK1I5BOtfHd9vLO4mz4S5+8aMdib2DBaABHE/tTzKFalA6woGHeihLJ5mwpF
rAfQFlI6hxi1ZIngisxhBfObm+z4OX7OiRgUlIvvnbIyV3jKAIrX1OS1bm3PR78pUIiIfjpMvV/3
cFODpYrtYClVV7A0USFUoiPSCwkQA6tA3dmvSIpzEMn8rLfVXguqjBhLxMZOS3pqhLyYjTZZJSNn
L8Mdzppq/9yqXfziLrNCUSV9AlrjobvMgAWxUgfJGKl04G5GRViPUEQbcaZwsA0EMKOjL80+xHOK
t4LS9174mphNP41cEkPVfw8iDmBnFh+yH4rGFq5+N7/5AE7emelkfPxWX28SoU3FWS7/VVZFkEFr
VetA4+9GQ+FvN3/uXbVuDZEqzyeSIYMgQfxap3tfAc1fcE+a37zhAcbvpbapEYl2DxbzNkPQRAKo
57RALqt+q7pGS94qRvk1L9rMCLYJYCSpYwevcGfUvqCwfpYbPZm4p7IGcPnu/RAxyYZJy2Scw7rW
pPdylYGjemKHUEzWhC7i0orh7m1JBt8wXMlm1n8ems0P3X8wISCTa735EIO+cluEXE+O3P1X8wVO
68nMEE0FCymi8PgAWNVX3+Eqq0cndpjn1Awwpvai4e2T5i3yH78/iswDpmFm0vlsuzPtylnmitCJ
rHOHe3uvrBMiwa087wLD+iNdHiEUS9W70RCqZ4gdN/KfIpxUtq3ZJ4Y9VMMj2k5y5dORvUdYCGqH
pcYSm7mcpuq/MDvd3TbAP5oQBLCuoNNm58IUrLnRpXRbAnQKgvSIaR7M2P1I0/5OUhh0pmc6J4eF
wqvm9AZqk3FD4Sj4UWtjKQ1dcQLGPUN97l+PHwL6ogPFlfjHg3y/JbfjPDgZAmJA7VSimlSqNy3g
MAd8ST0ukAnw1Lxqw5lCbbykiN96VECkSNgb+rYgFax0YBUs6a1woq3Ou3J9zsDkhG2xKa8liHQ9
dZVD4AVSqIBYihe5j1j6Is3Orcbl7qmyx8YneVP+nc1WNlykbeRAFyideZVnbtpE8K8M1anO09Rn
FEC0n2QeQ2YQ57NElXFhifO8d4fmeXzhoQg4UkyAsLnLvmq0zFvwFjDuMfMk87VfFHlFUGkHy0OO
ypazQScpRz9EHM7QXXJInTaokFqhcunIDQEzeOQUcRMbD3SSXocDTgPdL8xEum9B9bTziTAxrnMz
/uTAjPyXtQh0N/Wwow1IOpNOqjxaleic69dnDK7ORh63pvQTLC+sbJPqCP1DWe5Oj18P/YAOS1fN
ys/7LhbHZsHUNODBe40Qabzu+Qo49d1buKzbX6My8cBzKIEyyHr26UaCH5uvlwC3ZvwyXCJwAL+d
e+Zr2zwpLvQEI5f0NSYYfuO3Mue6IfVYyQjiXFgEhgkaISEuG1wjfAGJIAoLZsOL6KQ4+OV3uoyN
xFNGakZSO2FgUysrvtOF58TGSn6c+6fp+xYnb4MxH+NW48fVJlbXs8VQJgcU0i3mT8SxTgZhPxc0
EUUzCTBZ1HyoX7XxryaYNttTOxE+eRIfjLUg2J2ayf6M0L+2pWrZwEcdxdugymmiPDTKRICj2hx/
FiEajcd2D/pc5+sh95dBcj6gDwsCgl/V5vjLauGra58hnXU6iMrHL4Q3CsosInUI2vEC5VR4OAkE
JoOvYlNfN2nryHyyFf899Pz629wCn/ScFTclYLNdOyj2rDiugOdoxlPBKW+JMbQQuCRn6crzhycf
Jqhm5gQCk8ikN7qpFdPYNBtq4zaluuyXKK9au9fxvCG1i8KmtLRIEYEogHn9T+W49yZv4yn7swKa
GUIpO5kUFfLtXDivXtD3BXl1yhTWjffZNL19SIUxbRlRBCme5cM2ZpYQKGF6t8dZLjMrqVMkqNMV
j14TUFHpFYP+vGj3bFzsNRJZw4Cvu/2KrcejSIxalT6Ay94droUDK8qX0xTHAHv9LtRn1rKJsIp1
5eaRdt7Tn4TwR8QMC8hq4EeWl0rZ5YT8ovoTOxRFqA9h950BTKxbN0X/fZ2DBa7lElZ/UmWRKK8F
d3IXZYr+OY9WJVt4Ma/WgO9AvJ4G/yUOdpRFIRc02XHqLj/RaM03Haj0drYlMwy8nUcPFDW9T8kA
UT3CqiSw5z1gf3mrz3fIjK6KxPNlPNZHCpllJ9PKPnvv7KZwGuAZuSvFjDGtizrTmtL15saIbUlu
VZSeJprrElZgz46Z/8z2MAmKur95b3TSDrXDaK/8cuXJtfxobR0KjqaSuJIF70FEAWV+S/ZM7e08
0TKa1Y1cAAcb6L972or9HixuSU45J3cqQ1jy7iFMhLsZ+9Ef9OaXsPFj+KdAT1soCOqGeRACm6l0
vbrvt7Q8rwxPAfQQArKavToN9Abzd3kJapk0K60T+IdRefaWjDE/zzsp1EJ9pRYDmfJlnm1oE/lb
/azEBau1xogailTmHez3RM1GklUqJ/DJUWqWM3/kc7jfcmkzVZwDCJZi+OJpmM8mOhQ+c2kZ4j/a
hXVZozyJmX3OmNQHDlqeWc3F7Wjws5TDq+nYNos53Ulp1LYkEWSs2KtH+P2TmbPkSfgaaOhyixb5
SNCO5Io0VMMRdZsjiLHaFSvlWX9FAZMCokHCRU/UtTLvqvsKrPQIQQiNrGYls4sIsnqGNJICvN+n
wIunZd+9gh1XTriSCySFIRgRZfyIubH/pR9sa/5RfGVbdGe4DskQNK6YoiQxCVDp+v4mstlr4DdG
9XM/ufIRS0Ihb6F/ULt8ZZgFqAVaJIjgNpOXAtsYEaNNwYf5aaaMuD9LUBJBKRajlctcBb9MlJAS
/iu/tJqCcWk90VZhGGEtGmx0G21feG803AMDAu6PVhdMnGQPneCrsooKv6IGT4u7D7KrZ3AynMnF
d3nxMl6wRPUy35VETF8u1qGvQ9ytOaYOXtG49hHKov9VraA+geyTRVypUX9KGKoKu3OoWtqUQLq4
pDWHCXOxS3YNEk9nd+z36kOTlZeDobJl4cg9rGTP6OqSNOH2d8IXKOdVg2mx+JKKu6k3UUqq9FZe
lcQlpl3zO0/4htvUs2GYTi8F+7yPRS04K0iCdpo9+t4W2PaPVZ2gpoWn8+43c2dC+LmkkoUVChs5
TDILS0O7TsC4x7dUq7akozGhduGHX7249CG3wh083c+y9IaPtlg4VwyNojzNETBPp/dcYcmG1MlR
9u2PvwRukSI4fheV3ZLuuT8Tp3Ic6GBUcO+Q9BFirPDjsNv7X3jpUkYfk00z881VXtqmx8o4McRL
06vTJTAoxR6mS3hA677rsui+i5PjcDLUO36LMNNOuIP0e5LOSEtK3lt/nA3dOh7LHbksJgYiCIW4
sNJ1ZyTweVZeANMqrqmehsqjd/XAgz44R41DPn0Bvgn4JPLZ8aOEUWCcx+5FfmB/fZy1f7onGZRZ
ev89tEfIT+QJ3WxlgcQ7WNGeNBANOMWsceEIiI2tzWy9qQ+YNBUWVfMpcMwJXfAWTZTqIhH4Iht+
IpIpd8k/U5eP6JbhqBrZveMwLsOARbBVoP1U1GWjOQOw2KS+kUKHmwz01BU3amgI3T8PgJTF2afY
mx9O4SU/YazZTvvwuVQwEA7B3JXbXwGrGj8LNMD+U36mxputhiCD26fV2ZGLNZ4YcPojOtbS16h5
siVOMahuivBYxc1Chygj8ElcPEAvVP7nsV6+2MiLaBu49YRM2P4uGO+fDC2ri0so3vfo9rc95c5v
3oxE8Z1tUEIal7WeCs1w5bRk2VnIjqJ+4enRJCzpfK7YBWPDY7XfsSbRFVCHpDBtynVa+dgSJWXJ
M3hFDk4yApT4wf4S+pzQayj7hxXQ01wrm/z2Vbs0d1oXmOjCExfDclhSYggC9dewixxhS87uqYCg
GCHnu0U0/PI90Zpb7icm5JKl7UW7KQVhv/dcIuobDhFwCDFr+9tcaXY3vJE0oqURGLqa7W2PzGva
RyPbN+IB8jOgVMK9idnr11Cd/R9LJq6NtAmrsQdj+I9VO1YQ1QGKhj4tvtkJz6iDqS/iqpBibiRN
F2UskVdbhMYIe16q3//pkT4hP/4Ppbiffx5rt2jCK2FYpw0LqDz3erGyGYo9yvYwSQrwRbOzSQYo
HxHTQ1onzRtRhT/EMdzI/YmfTxp1mGHI9trTxe38y8ixEjpIu9G0m47XYduuVxOXQJC4kWVlNNqS
2NSs5juPTIsLQLe9fDiqG3C6deddmYchJ+WcgPltOrLeCPC+cjhrcjqdGhJ8bcS3guOjaJHJxXS/
Vq0htPIBFT2bL2ctUyF1omly4Y/WJUU4Jje8ocb2A9A0xqt/+RtRqiyfTpvD95hPpq189zZDrnuK
RdJVqjndnQsa4cwGQoQBItGUXTsIvkyJAvGjCmSCO7/kFuUerScCdI0wQatB3vo4PE7dEEDU/z3n
Tml7lIPUO+u2pOdRZ0Xz39UPuuBD6J0VZUxtLfYHlRXyCW5Kxey13YoVK01f08dupLSvSEq0ZFM/
HwEUwlmop8WnnP1zWmvHs38VRDF1eHa0Gce0j8rm+09bfi/3EwcFo7e6FIXGxd48uLcZjjPXtYQZ
igGd6/3T0sgynNomiNheVcR+smnNhZxe8exa4rmdQqqx/4NdHcXV+JPhfx5Zum/hIhjKbOhfmhoe
2mknSELBF85p2sD82z4dcGpu7jY08m83dbaXuz30QIgqwFTqoZ+rIHqHAqz15xgDwErHo5CJNgEq
O02EU/LCdb8W3CISw9L0iLy3+7X/qPbH+BMex8EyZwkiGbDUFjpdWZKTP21rMKnlP66tMn66/MQ2
CnvsfzRlY2ytIgcwDTDl+HnllEm0k4DXjalN28GJJrOcsnvXFCirzPQgs+FzUrNe30WoxxLRnzXu
VOJ4DNm46e7Oc9DCTT9EFdDKP/n/wMWf41sIrlD7r6D9owPbOJgFaNGjV9UM+jL5tCYUk4lGQ7EI
srFk2tOrlZbfwngvfSp9ft0aZ2biKtnXyYd7A/JWhIvWNfcWxiHdHCE1NYzeTFAp84nKYjDNuwoW
mtYQ0KEyWmvGdzLwwYfRe7p3Kw883pHXF4C4AydnwPwN1ySa+iOBY+c+FKBDhUtnPKqbZddZbLUe
35gXSkDV1370jEcQSyXI67FM5ekx0g0Usl5c9UXh3nK/7aGnzqxjPn0A+5WGlKGPd6iF8deQU+5c
0X5C+qb5e0HeEefPFqWRRIKsglQ0a060zIAoc0PzOCAaRpXgXGRtBbeDNQgwsP+UyncOlQHzDiPa
apU+km3MVKx4bEEkoF+dMz8Zo4IM95PnhYeZufXOUyIHehha4iFNOVTB98+gC3kH1873cPN1UKMo
npILF+ATTm9OKwInhg+Yrga5nGpYjepvKWVw/iqkqk57TgIAGhnqUH0EbAvD/0XoYDk4zQBrJp/z
fjA1Yms/GDWduK+xbYy/hrep4DnNYQ6ejAw9CqNpFZEZgj73baOkS+jj4F9xqso0qvG7g06nFGTP
2IPgdPAAnF4LoHe75KOBh5os7zhYoESDi4ilDWVEtAz3fJmPn/0DTP/cQ/wWvHrxHXJB3eZnqSmf
S7VvXvhJAMcj7bwB5ZnImafFliFrnXs59//MvM1N9Yrp98b4kkWF0eqtHDeBiiq7L0G6qyPXEpLG
nj7WAdlIVsAUXs+3SAbl42aU2FTHQwnEcfH1g/aPoUQMulWLqjOeAf9HI+jasSZX45k0ExrSHjQe
scDhowlj4706IwlMhsMqCMHgT2iWuUg5JGgcXEcKrAsgPFWWX8HZWGOPe8NuI45cWUd0rH5vhPzg
/IOkS3GPwIuXU9IxSVTEFJ2BaB8W8Bcj3MjnLyudg4JtpBE5UMZqPB+/+PZFjoZHaYez9w9/fy4p
6U5v0gEjTBUEhAwEGWAyxL2254fD7n4W4WQqhk0bkx98ZzCVox1WlMFPKsBoTerF05I8jCL1pawz
9cMBJhLLNvgEXoBbhfDLuRw7Tvh1psBZ1Ijr6K3+y8ptLbnIrpKuElCwxBVw/Uzi8twRk+Z4yt6+
t8a56Z2s5YkwTwJRvGDuy6NPg7vx6fGIRyY0x67Th+2E9dcR+9FIaqMy5C1uj2kZQkO31S5vhR4W
Yi0+R84BTHxGQsnr17jFg6Grkb1TY4LusIxIX+YhxSZh37VB6Td3srNfW0t27Qh0DG/3srhZfTJ+
DoKmGfs6MThBwBzqY6fje6VEuqLf8yazx6ac+PRcMpMdqx3OxF2C9DoSDjrtxOERmMShJ/Ww75Yh
PGMh8zUaDjMzGE0pwi38i270ijgacdZbZrhG7LS2exzQXLQvLnsDl+1XoEqo7CzQ8tOgmmLbjr9U
oMsbxKDa+WVcv39FDHgDFhsRJOgaswtgudtM//ULFx9lZcypGF66QAXj47dozFjvBT/irvPuJn0M
20YztTlmsvUGuFRXpD0OXXCOyBsL08qkqImPr+6zEk9y7Xv0S55j25bWdHvQwcnq7GpEwQNPx/Hr
y7qCdH0CjsLzs4F5bw3y9vi3QEEt3UKru+ghXWPxSSk0lQeAw5P+1ohwgUuffMG3HOn703dAwncm
oxCOSmjvf16B77HbVfpexkJA8KKTtaMSsyRhg4hICSsWtLK0qZkexvJH3X3WeeZokhcVuCPXKWGX
LhW8Y5fkTVE2D5f9tcToHNjGUuXGfA2XrXpHn8x7KzFqcfboyqyMr4qig04VG0nncffjtmbz9KEN
Zu3j6Z0tq1XzygP9Ns8WfUHUv8oEJ0TpRkDERMb0X9D9o4+CwbS0V4XYBNZOLA30I2iVuOuI9RUj
FxXYLeZb1mEb1I5EFQD8NJvYVWOiIQidv6242EZYonSmq1RQilAn+ew9tf9rJLv2jUK02PzF5WOJ
HdnbapEiV3riIj+GBYoI40o2Zw3hMnjAbbt6XcZ8U7v3KTRmAyq+dwS07AerdXD7oBeXSrSaWBG3
ZhXkURI9CDlzz6pKneMXtgtc6/MVra2svOMoeSn6/867M2tRTWu3+ujWF2qqzwL9Pb5HS/vhrnPa
7tdxJt4VdLSz96h4dRXFerL7raf6Ub0wLKssKqyFjMcDn0yv1J8vJ1PS9ozoH/390nI+vin+M76n
o9jAZDodRYxfpWDyKkUIqN1ZWpSbBVfSgT1ZnIpGyWQ2h3hzQ7LcABqENAlIDQgQvmCy8Iz+cpTP
DmJ94Qosk5gEDM/j1hVPtCU4HYsSIQqTSRfZZcxtG7dpc+XkuqgSkUd2/TsBMOOfNSAnvSE7lhmF
DwuZ4tKWKu1ngXxargn9XMfrknQ3ZZz1CxF6c72+WmQ0r/N3ozE4An5Cb7kn0UmxHT3r+5LifB74
5JwbT5T+2/KOJc3V/fBE4WZF2X1ROPsLoqE6+0MLsHarZR3VDZ/FisMRY1GyuZfFG5GkO0eMKOB5
+gTbhjtLyRLkwMYFHzBj1Rz9Dcv7ZjqwynnJlIIh5TrtxEQsA8SZc3SC+e6Ze+Qxv1qtamjyIM9k
TJPyFdVW8uVT5ShZv+7nmuNIRhp/0xtxsoPgE1nOMOs0fpTlh3kWaChxV6VkoB4N5kWPTRLTee/n
paXatwH+7f4FYRWU2yoCEBgzAky0dkUgse5Pa9Z6samRbSQRDTtKrc9sJBBWQkNXZregArHQ6F05
tUaxl+D9Mvqo9FJg5YkVqSqStdc/hliO0YHVI/XZ3kvmb1EiEPSmDL4quxzPfK7oet9xSlXMHGlO
9j3tYKB3ZC9j2JhwP2daYUJ11vYoUZu55EHHNT6dZDHq3XF7GRSWwE6yCPtEOZe+NBU1VhWafgaQ
kzUI+xrRM7TRqooYwvRS1fbitBHXkENc18Z6bUoud/W0JcPDxqQApc8jjiPpunFlkzNbyyPf0yCq
5gMhOdw2831setE+W1hq5SSqoRFCGVo0epkWRcUrjBRbaQTYLmaNOOvlQX1o2C/2+WZpEQyDd2nU
GdlJX1WkncExLSIrPV51Fy6z2g9o185YiKVBgibORKetwBo2HL7nraG29otyY6FOqCi4RINSbNFX
VYDBihC/0LB0pXIUth07pGDf4SLTErqFH/BmN0wmbGeJ9koLO8nDU/sFrrhphVQRnieFw29qAoNh
ADgw6E1z0HRDDJQMtQeoq3O3nyMUcYGucei/+UKK7z6sgRagXiUvaN/+5w74EpRMVGm4tIf0/qAK
8C+R7e9nt61LFWfBo6fWG89iwjrTVVQdvt+x6+Xr4fiECdGaFlOr1GF9gxHBD1BWHv9eo0pv5uBj
dht666U7j8De3KOntApn9VEZlaJN7cbLEB+BKYCEw7XZbmAvNmU/+lLpOMnT+W+c6/RASgHCMGtg
WCupRNLmzM1hL0EkqIX16XD2NFIYWlXstPWJylO28vIg+56YcmE6UfZRGvmeUqyHzWmWW7QkD2Io
94qpQ+xX1B083buHsZQytYvOtxyJEGuQ/yjSMKTv4V0c5e6vTz3dOvqjSgHSh1OdrdB7JfAHUaT6
Sxft2yYXpfBt3UBJhQBhTu6M+hj7N764/ZtmNXl0w+tFN524CFNfvuOESc+HwWO9kpppUvG/dizD
GjMQvxPamFznNzUCWdJ5m4vfEmHXODcJooSCI98g2oxGuuOLRx+a+J0fQZO+BQ4KGTtmat7fqAp8
vKUWX5uNpwOq3GxQS3ZuRYCT1Aq0EPiO4OEhm1WpiceglrcwjlnTpNYirrYSv5zZNBaYKjlmhE1O
SfyOV7RTsahJ/ZiD7Vb8Jcpd2UuDV4ruJI8vnnB1d01o1C11QiItrsMyW+pxaF7uOvr6wE2347oO
QiIMBn0lSXNZHLCrRNE+MF0YtS/WDjCNVbiBe3mFn9aVex6zNbbcUO7Vcm7ExAOJMTqmlrKK32zO
0lLCRXZnBZ2k8GKzi18Omi7KGX0AlJBAtNnBD3iV3fO/cAEfkBlgpVlhQbAVdmlktvQMBYrvhJ01
AgQ9ClsAFWXJ0jFyXnaDB0eSXorgG8Rww3zujt6o5HsBo1+DGbzEdNgJBar590lFtDGPmLUMudr0
Nv/oRZMmtafYzcYjbr3jexjCiOvbjvyI5xzFQE8PinyrW7n27etFl1oeL9QxJX8RcRdtFhrP5d4j
NQPnJB1hz7zOxzhcQ9SU1oqzDd05QyocYL17QfIVEwPfS1FScld6Sln8sQnyYApdGnnVsA9AhR1g
RX5O/n2nOiYXwQcJCQX/xFHB7rJ+5jceBb+cBpbVi7aXZ+2CiSFQRDYdY/TvlV+yT0k7/ril2W1p
1orWXRqoYPMl0jP+WRLyA8Z0HG5OtgC0vU+slyNmLirNr7upt1WwfXE3UDJKzbojZTfndbINHYWD
cg9BkWmT+fEBGqZpnMun1q++H3aWvn5yiqkhsPA4KNOPLJ1x8t37NnASykq6YCkpUxB6+PzpovRv
F/1UjCl9UdLMfaZ4K4AAG2EebF4WJsu3iVD+wZ/VrJMBHvrfgNsYXCwVADUA9vDieIbIg5TpXYU3
tpPDDImNt6VoX+c1dHSaK2Rzw1cu3tAN1T5HixSUCpo5gTXeOdnQTnvYOQYYcLl5e25er37fIaZD
muckXQlzJ99aGMGmroRsh3C1RHuGY+ek3rnoJu5F74JFmEu8EUANoZxAmDacYQxCSHshVdCA+IAX
qCWwK7w2eUO+qei0OjzIlTc3gR+P8K5Ns9haL7p4843hMz+ZJDRgNBghBRxxV02Do5ui8u63tIwh
4gYLTotcXngyyuh5HD1/jx35Lluxs3Ojybep96j1oYKH4IVJJBkb/+6Mua4izrjzcWWDBH/hCZac
zYmewudN2w6O/Op47/YGlB/jhgtkbdlxbGm3c5NzweDdzOK7y5hEkDnPNp/hmNXI2epDNCvNIMOX
Zvfmdis+7tsSzHnIK8pFnFxMFIZDa4SX9Dlsi2TbfzKua410e6qM5PwOktEt3gR9QbjrUYpBjkF8
JsFqzqp/M82t7L1YMqLyBcHokobVo1pXUil+XNx+AJh50DZqC0rgPBwbDXJW8nhXxMpawt6g7W8M
Q/n+SQrdMj4ePSfQ/FzqXUnVEry48lf3lpIZXl6AGYlbelX0IdnLKP0c0geX9a+monpCR5usC9Ul
rZ/KN1HNNYqkANa0zd75E7JaSmax+qoAHk0x4yuFipfkU6iLsIQmhTABwoT9/6UKx9xJSkel1eBr
THe4hOBinTtvwVaE17IJaQSPcAoeM0tF5AlKbQrDESStC/ocPvUKoJgHjg3BS65nuYn8mJzprV/K
YeCOzH8vP9eND/s+wYP7rMnRTwKCB+Q5jLNSghXEMWuyRW51gquzV+AKRjj2O3LkGzgzH4BKsr0i
TgBc+Y0L3pHSM5Z/Kt8cHMqznmaBbnDdE2860Rgp9Jd+WIcZb8t9JW/jgWf9xeNWUBSZ3QfekJOU
qRieQRotkRPVBy5iWdeDyY4pUUFnkiqyQeogCuMV0jb2GFjc73I/BfmOwBslrNBIjMt0HE94nltO
Wn1gx1vtFfGlXcOzBzzy93UC2HYTuPUadwtNKQ/rhJDQ+LAz+oXlrWBAGiLhsGRuIcoV9Ifr/Y8X
iJk0tJXenD5PN/AkKAqlpRylfFnrGepnbJkJl0C96eiv37DXeqvjhZWHjaXztKKQT5ButQqNnzNW
AGQq1KxAUIO//ILMgikw3a4Z4xO4o9H+xfJHpdMRHvD3oGfwWfY12II9CjX0RNiah2eofg4tXsVW
lsv5775dkokXpcIzlPwOR23LUti8myk7ZakCUwm43+3X35AVLNyuLxAmxQu/KDT/Shux2ZdH/b84
lOF/DilNyeE4jnkXzowlswI6MHj3XkB3a4QrNrw2jTUJQKNnJNUDT5YytWjsu6G5H2vSxhHeSqaD
tEGueDWAYTX0ilxK0u2eaPQm7vUUvkNv9nHlS2eysnfQlQlAahAfj3GXD9Lf1S+q05vFNQba1Jk1
bptDyU8KPEgytdcCC+1yCpgsl039ITPIqI9iBTPPJBqYMaYQknts2vaIoVcrSzK4pa938p7S0tMU
2gNer2o9o+KBerXycJJntr/TnK/xXdo7oQoZkwyWe7ExqFW3Tjs85jAHvjt8w5Jlqgn8PDNEmOSy
ITGefSWoU+4Pho8PJ8z6jfqMtidowI1dJPErng4tZ4EgaAqdC4ik3x7s77WQr98IkIDwSJajD7dz
uktOM722m5tDZ9bI5B4O94Qu0wROkmLg4PKGIl7kTx/Pi+NE6r/b63D7ZuHvaziHuhAAuXeLGKJi
H50jnGDF/wB0nfXDbuIrGC0HYLK3fiizRyj16Akef2gTtzNs2T0qUvA5QUWPn4ApzFxtCD9IEnEu
nruyqnK+RcK/4RC5C/1AwhNa/qZM8riBKYNyaL2RJuv7xAoJQ/d3U3T5kuTG1VLVheeayzQHG8+f
X1rSKBQyCGuuRRD1Sh02gEwEr9I/UaDJM9NjbCObWOJK13Pp7lz82zy9Q8hT8cZwZQihYZf9ZWPb
y/53oJJt7L6xccPKbl6OkRGBg9AkBJ+qjE+qq/H5T6FxPE9/Rj5Dlqg10WrMjjKA/BRtDQxRamVg
oUD8W+AASazJPRq+YFhAdZu5jIMcQ8b7vznqgQlhygDTY7Lw4rRXCOKOh4+yoZoQ2xmQH6l7He8H
z2FjnZrsnuJif2Y4Pe1XazTRdh28+latykUUi4hWGgIAli318OsMRKLim56Cv612gNGJRT1sZo8G
cQB2JolFZqZkFq8zXyaaOtS57YdXyJrWcNAXnoEcMDetsrpV3ApsFIKoUwLZ9zntDOL8f0SXP3+D
8zFkP/3rjLgutddxkFcLk36lCTAxG+8oxUxef8FvJzl7Bo31zf3PpPL0iKrFmghoFZ/ad14/V4tr
Mgh/9sNSDbNd0UKixbOrllZJqMSLAklZNekIrmT2s3PurA8CYvHb9zW17ItqKZJIOgq1MgFG3BnD
X9EfjVCeM5/cXU8aHoGE25/3fKvjiEt/KszP0MDw5AZAoJ5kQ+BpdLF8wFSjV1VvrEQTXkGAAVRu
dgahfzAWRv8QjoUPDe9ApXtJVxra1Vb+S//EVFIpi90oWxJjIgV0iYkAoIAMHhZ9Y1gMK5MMtjat
RIq3mzIZS09ToN7+UxzY+8GY6iBhh7w1sAj/brROXWwojZZkbVMDqu3AYfsUarr1l6mtIS6WOO0m
TcEw+x5HvyFh5MuZSC/v4ldzh0LTYVluEh/XzKwfPd3Zt+tVtHJDyTz0Zu2maDMJyAHSrydlOPU+
1A5IBPJIGvGGnGhbH3GI4mlFmpH22RlUSon642bem0nlzJaQp7nMfohrqk1PI3tEUYS+eAVQ0O7/
uE/egQ0H/2NeJYwoAHRPhU91Vsn8czZ3SrvGaV4L5pJjbicjVWGlCfmvdaZ/NhmlSv7M+YYOgz34
FLhBwtqYBeaMzEohrSPIPv1hPgNtNiXiTbs6XyA7LHcoBHjxwm7278R+JB/jjkn+/rkb/j4xcq8E
9ZB/DjKP730iA3muYPgw4DPGfl8V3Y9JN7FxjFLGhfEK/2vJqxSWgcAgNf1tXW3AXdgBxyQO+lDO
Xy87WXDyJNSacc2bvOvro+HKBLv7/fHjWT+tt9VeBj+E4zivYeJTs5tCSeBNa4dwq4jfTqyLYJ3i
eC+K95Z9FrwVDI8JJyx/wXwmi0FY1AkFZFL5XvuGRxyCt09F3vCG0dUc/s3XLADknHVf5e9RAV8D
3Gy6zvf7oEOLq2hPtJjykDTS1XanVTQKpjFSYS+fC+OZA2F9NYQJEWC7RY9u+5b0t4Ay2ujLEkzx
3F44IMf9wMVTzlNTPYhHvqxswFaSODdGRkTnC5ETCM3QkrxhXrFJIdrCKahyvEUNeCpS2PESfnpz
UNJx2bSSS4jTp812UMdBsRruIpW9petdRnj158sp7eqeNbiYsdFHZiIydL6VXvc7oILwTxakJLQP
ijCdew5uAszSkAxjPIbGKc8bzZIGFYDufSpbguuOjYsKTBKOntLC5eW6j4RWCjCgoMZONFtg6LD9
FlLSHgl/uq3lfC87FVly/PbFdD/odgoS5Eashv4JeBBuwpHSdfbtfCelB/tYa+V7+2QlolvA8XPO
cyAnbaEum+40nwK37vwvQKBXCeFHO3jyHzCsEwIu6gvrQZmj74V+t6iy7V7+z5HRrsXzVFhZeYxg
7TnZlBeebdirbXHVTRdGnwYYzV2fqvMjo1oKyaC1XOsfAboUCQyE0aL3gItv84+C5OzDI/GlCmbP
Mpm0Lrjp0fyfAHQW9PTJQ7mxgtn/gDfVZI0fUP+uNAM1VG8yt/Wh/QCuwrxqhVAEIckXztWc9Tww
Kiqc+DUTBG54Qj3m/5TXSnsh6zoj8/s039mHqnmA43o64XIPG1Eq31OTT6fTpLg3T+hlf9M1AytP
4LmfCJ4Nq3T3ojG2v6MDH2E6ImPt62VMm8cZ5LkqVD/9wj8Bkqj0Y1LxOLS+JEh+NhQmInbjBfax
rLtNM42IYY3tzyb7yZXYnC1jbsWQRLGd5Z6vFj1lw63ZTMyIAqvn7Ta3DmKPPq6I9/7cEiLVOdxO
9teJacRxU5o2EPC9dky2D5F2+OVcBcYi5Cewjg0EyxecSnDNruZ8xfyLwQG1jX9J7NGGTbvnuvcg
3Q/8aBQJNNzOyhrMAcU7NbFM65GHZU7L+O6OXWWdxZm0NIaHRsh0luZiNI/WJYjfNsQTPHEsBH4j
KOel4NE7wd9sY9v5GAE8pEDEUdPkDgWI7Y1S4wV2VR0iLrjSNeGrgaeg7EVgMHV/bN+DXWlBJHQk
X4AliDLdsNit88/hxUembtQH4d7njCzgeO4umz98kmaj7N45BjI2MXPQlrWAeUxqXuxueEdF1wNP
oUdHGuqpJdpP+cK+T0FRlQXU9s8uhQW+n424kfFqtWi+ACvJKDmnF5WtPcdjRUQHFd/dlbVh+7B0
5hgN6V+kzmDkhHdELyjlkyvy60OhuanbMi/cahVXHH0WRDLasI/zJt4qDDMpz4yLwMoDCTs/GX5y
IYSL4JZA/Zb2eL2tB9XwHW+XMMhpI4uyQfXl+Je4akXm76SDf2DVfS2sx5WJ1AwpiH3nMalWqWOx
m0dnuSzwbym3KLmCAUQZmulnZL2KVsBDmtzHMfrJkEZfTLofErPk/5RWKTKw42RRFkyF60eq/xH8
vRpZ9dFV0z6FGGoVhMUO7WKz7T5WyHNVRfhfCpV/xnCKbdiP6FOSDNYCP+U4vnqybV3Eh7uDW9qX
rnhbkYsL8BSgew9ShYBxKuHhQgcfIrA46CUJRiCFG999+0FNbTQYrEAe4/Mv+PFr2GkPmsGFHqh/
CWD7C4usCk9jgieItWc650oPxUnddDUqkIascsn8DdK3CAJn3lNU+sqqivrmZ0//O6C6Dv9TeU+h
7JvSPQhwXQ2tMkAkMYs5ku8DHf0oknp/g+wLDG8+dQVI0V459+uOyFdEap29ZKX+3cwK3CL3Chr5
ZgzPzm288SRoseVAbAJEFh3Eexy269cBTR00J68cUjI6lLdMVRWZV1j0YYH+ufCPG6QunLwjQJiH
i6dlw6MDcDC8eHTni8Qs3vB4j6fPMVsr0dxKz5OS5Li6/J6kayfRSN4LRH4BPE07EoEuiVad58AS
j6wf4Q84ktaKD18cqiDbXDvmlRWcxx/Lz5ek1V21p5JdpZz+DtzTp/75g7ThBfth1mSBbki5mOm2
SgV1THi9J+tdUnis903ZoHYwktEZeRS5Ix/GkbsLbEkUS7gR+V71anOsGx0uk5omwgF9aRShStlL
iojSLkdEuk/tN9V3Dv5XAPhY2upCS2AZZlcpFZVNKwcLNnFjyWdJdITuuCGyR7vaJPC4wIB9fLOu
M0dSAGHe7UZ3eKyeFmecRh0qZlUkmCWv/fWrYUpMNQqAexaHdcg8sff0fOyF/Yuv8iKI+fvVtVFD
q4HBqZEaUIrD1KpZQFmSPULfT7Yi+ySg6M8MJujyLfih1+rNl3uc6jGxqUTciGeOszwqb6wLTWy9
AtkMdKg4ZWG6mW2A/uyJv3pccJXEa+g6NiSnuN5E2JTPEROlzB51rNSQdz41WyovchWVf4AlB0iB
XKCGiodv15aXDSCrzpbYW+6SOmagAnYRDgkD2RHgjc51ru/DZlHhAMPZ6fuDHla1sAQh0dOqVHlo
J45Lo7wZQisIH7x7IPEfA93u2ebeZripKYTXWVdiukkohkh40Aqw7fs2qqXs8o2Wku6le10rJOjc
O4mXXMvRmCJe8FgSWS1+OwyFUYK1l1QNyttXIsu+k3PX2mq+4bt0RXOmgNXj23IR2UkJAcepeh01
2f4Pdd2/9dJpAu4NZCTVodeVc9hcwiUnvW9tfaRnv65ezRtycvYENKde4tfTOyjRt8SLKk0JQXg2
4G7OUX6JFB2RF1jU9WNwfK+aSAIFw1ecArfRMRKsMq+SampITR0T/4rGt8HMd/iS3VNoHW4B65aF
UjE89bUnchepXjjgKM0bnALriv7xe/fy/6VAfmia5B1duHI/FxyezC6HFoNSDpKpTBekl9AjssjA
A5vMIWaIU3zc4QdB8Lviqd7GFPwS0tdKuoM1Q0XDxnOS3Bz9e0aeu87DT5x6alVsrFmTAkhKfk/F
nI6SjrWK6ESZkyeYb41CTdDBBLDoJ/IIf8PvBCZSp6M9esEszaQcTeozXJQUeUR/uMUHy6e37Vzy
+89zCsS/ETNHzspbPGFNbueQC4FkwBrl0LTOd1csAazEgGaINNMKQjeIlaHMMA5NVHZ42BjWo5HS
TsiZdFn5eNnlrHIPvpAh4auj8xK85O/5b3Me1KXsYtR6DFxeaxcjNoJ6TzuXiMF0ELjFjCEpMiG1
TZThS2KJhGhmkPVDtRUVanHsNhIDykTA0AzGbZrjM02WNWLqGtit6kIv+CKHMScksS1sgcK04TsW
T8Bn6pMQQVkaut8wr5H9R598lyuvmVJpq2p5NYIZa4ycDSgdROiygu6GCDm89PU4GmHtCAqrrxOp
GTXwa2HcHEIK7SOo9WasaBvOpTgZFZjC1K0x2PhDDPvef72+H9gsqJ1YTIQCvJUkCIvnWQ4pk8CS
1brY54lAhU9s6AO9YVYb5W8TIuhpz/f7lRshlQ6MIIwRDB67SWJE3i8I19OQ2riVFKh8+HHBJAE7
0ip0EgTIng/0+KN0xQCpF6tAv9EesJw+700QC5NSzYc8a4vlQuMAq/Ih6MdX1eLK0mYYctRQzuxb
0UXBZQGpc6nQT2dcuQu1UhYYfxPqVzegpRnT7zUwqPrNFBbX5EWMALRAFLExuIXFjvVfl09/X2vH
Tn+FlwkiDUkZ6JXFMtiXef5Mnc64eWmzC4fdMJ5tTRTHpXwi9TCr0HQHAlMoIi7FtE6Q0jSB4jYy
EX0UfzQZcxiZEpLA+bc5FoEzMAr6a4OBLq4CdmC3Oi2YULR11AHYHl9XpjIbVkkd1ivAmNXUFRt0
BNbgPQrtMqt9lbknlP1RJHSxtsgSnCsoiZgmjRsJYdoVj/JwEfmMmYMB8i3DPEcxDSljObxCWLdF
IiNMmWEUGIV+g8L9ca4m6rqiDnvXIDixzMeUEoIaKIORWX+979RAiEiTRDFwNRwF0f8+R7n2OL+B
N/eiZChMlXaIu8UMW0AtEPgSkfA58GRP63eef3fmjyH6LMXK+2AT3OQqfMvUTKqwhXaVMVQDnd78
eQObrh1MQnNHlXYiYwM5Jkp8muRbEn5yvq/sfEE3uw6LdeZjK+mpnHvc8RLgIMekb/3azt0loJLp
Wz087QeM/ASLcVnj4zPxTjXt5fKGeAjNFLAQQWIj3y4e305U8e2Ag3+aOisc518PeWS+vb01PdEA
KB1iiva24rHkQK8bJ5XryFEI9+pzKpvkgDzRdmPBQ/rxOg+ub2VpPQ2lpc5N3RW1LMXkq+VRFbfT
pLnjS3PbmIPxKKB/ENXZFGBPrSP5z0PPl1tHZEAgMLRFmYJPDwLiKWmZi1GvPOQDc+cT24V4eH2P
IxjIpVBC7yB9/4fFhUlJmqOluf6whsImcBp6naaUSBX/TRSHeG/5TUHlvOONn40+nFGaEmls4seU
wRF+C0XnuNVZ+vSWdWtHhq5lzad8sqVeumGBfLFK3IEWXe5jAT90+pzQhHOH+95+EK/Ajv632/QC
IlyzCZ/2B5O6ZbS00kTnEcauPBYeBSmlwyk+Q8gyUePUnca0qdPPFesSW//xZTWAzPW9NLfHd/cA
xl347fWL9b//S1nzcWamCcA9ckt8K18NFKudc7nbdx9ob4FbtuQtK1GqHgWiUPUADAUKErp6KkAb
T7qJv5lTLSfj0rka9QMgKc6ojWzRiPjLFoTHJ97tHNI+2Cbv5uCY8h1P5TDxYx1n338hsUcSGDJY
nejng77M6b558EsrJzX1LSZBU6t2WwvJXYJg/nYQxPxdFHPVgWunlQ+B95s/fIpz53txeupjmv1U
1pqSL4prSz0X0L6Dg4ixnlH985KdbqEPxEvQdm7rT0Jw2G3Y9jNDLZDi2uv83DFGAQetkNMC8tWQ
lUgqfd0GCBd/h4Y+47I0M0PqmHFnjf0RHrkiu6Yzq0Oc0d4OHB777L4vkmnrkpZjG6sJzMv+H253
3k0rIGNiRoQCjG9DjpjEsLnV9lHxuxZQrx57MO2g5SYIIZMS657Kp4Zy3cD7GVXMUOTEFgQO0fF9
AEoXy9dj42wFJhMGV7wv30XwaE8OKZuIVL9K7zqbrjpbYpqnZL5buWp8WsIHQjgFf0jnw6v/ICnu
xLTkhuI1Kw51uzRiHzeWS1vumVKXXlCZWs6ERVmNrnig6UScW1hofaatWmyrPf//j1MglbI0HUOM
H59oj/8BBTXxPg2ukNK5aFKNA6d2dzg7YHbZKVokKu9zgVpGP0aGeKjgB9Nqz4KUr3jpec4twgV9
1peuV//u9FTvGfKs0eahZegtkuIY9GFvORdoOzGu3rpNnVanSZILbKLhLXtJFm42ksgkaQTFsIr8
PpmSwwvREJAy7etaS+wWEViN4u3UyfYP1So4f7K4P7LyVn8j1LghFbVZf07pSF9/kd2/nigRt5jL
3/bvi96jpHboL32NX0Chz5qsHqy0zVKyvXmFAmvJC7voyUpJdIQ6OktuazpXzH8SVPo6ni6npa2k
MjUzqToryeTobsU+BzWR3obtrMLRMqwGCPsAHVH9rG4DS5wrC+2VPgtszLIJNncQ9vCnCTHGoBAX
Lx6kWCDRw4xfPh9g6lK6WLfO5xBpN8OAhhwKlMwk40IzdwQkBYp8T+M4svtud+oc9X9zZZamb6qV
J+2ZhKLUZF1snw4pGnZbMJqyg3YWF6SB0InOeoOQSB+DcWigoCzSpWSy4GgmWuIMR0iOFqTa7UYQ
1i5i9CvKz34gxS57byItPftiMnG+1nFxtPMyW+HnVnzh/IWQjeDO3lC8s+kC3sHo5yuuK+t3zlVs
VqQoVfvgia8f7T3QXKmG2Z/FWrP475zTBoyGB6GjqE2oSMBM7UkBWcfuARFCPvRKLFNTSJYQHE8C
PzpU0qKLB29AgwB5ET+DqBc+dWboOedTOurmon1OQ8nuk+wBcoZcgJJuGrpx3ppyAuBz+56pzRC7
coauHNfXBbGFH9tEmXZh4y+j9AZ9iMmyy3yQ6VJMpuiiopANLyrZXsLA8cH5d+gq1K3qeuni73El
DCCAnRt5HyosgkOcZXaoj01GcNSOcoNUCPBQSIrXCw1DnUzzIPnrfCNQAH+NCN3QwEWdj9WP1nI7
7NWFMNYuW2vf699U7pfTwa5JCZXgY6EJ2jNrzWZjiLTXUHs5qkv6CTwo5/4+Cx+GBt4YZLffL1QA
RvZLKEI1XB4F+vMuGua/OpkavhWnfXrhJMXSTzcAsO9PV9IsIGtlwmS1c5dWmrzStaQCnmC3hSBp
tih5hkXmfIEabWAL/T2faXvfGxCuuC5rSbfCV346H3M/QJ/AaZm6A+8LHhCRUsl7z1Cwla73dLwn
iHg+zIRP+9d/2+tpBrTm0OT8JW5lF+OD1+QIbOHRJO9kKgG/P2ka68ivKarcNMHACRRMlYARU08b
1/RHhghj8GuMOEGEDGu3r1N/0RqawGIzY15fA6iUwtxaY1B1N1LfbKGO1KE+nFAI3BRlh+QlKBxT
GsyQgGCCTNc7qMowBPyeWATPOrHgd35DPzNf+198aZIiUD1gszVqgZ8kfb9SL/pMGA1sBo+wjhX5
gNcy04nc+Lv6dXXbiaRQhwSx9zJJSbEVFeiPPxl/Sf4JZu44en3KNPljSXl7sHy3xrvg46acnh2X
1OSfhesPHiZnoMkpdiABmSOg5uDdawoAeXdsGPX8naBWoCJJDi2yWsDXWH0Fp+sPj5qLE8fcJpml
OMY8Dcj2p2j1CtCQBpVaBgcBqpPElKvmSTDh3yNzM1lZ2ZXAhi4IMBzSpxur6doqV0i+gCD/ZA6V
cuQlPm2WXT5ZIy1GrbFCVHT+LX0bvWn7gKWex/UJJ5rOSucwvSwoucle7WeDuNyPIkzRU52VCXR9
e2Cj9u+9mTN9xWJx5zSrwJxKS28Rg8LItMFgjgbQf64ApH6nqc/635pQlaWShogmkxGd759cUZPo
Pq5zS4nMYFe0FQRo4j4Ks+6aGVHlhPjEezA2z9gvQsBnjFEZzXKMEzE1qTLXJuQ2hX8dfIXU5Knj
0ucr/fwLCjzmtP2IGvtROTUOOLELStDEvHVjjYhNCIgPXh1mwHafDByL4KhalBzoedUgMaU6aQ+o
b6CNxGetp+D0CRUyXYOPGXfII/g4zpoOQPiA7MhPNY2UJAKqUUtQozneDBUAGKc9RE0JT1id+hxF
EbvuVl+FSQZQLsWTMsEhhrtzWw8Shdalf4RGLH5MzZPm60fCcrmOimIScsaNh+FG+F9jmMWnJ32v
QwYHYsCC672+rzj5ToJCB6OpxuIewgWJ2F0HnnBrfMB/KHZ7r0i+/XQ8X2es5HujQK5zL22pfkPj
7mZen3lPvgz56G5D+3i99HWY8sqkPkQghm/zGa7YUgaxangHHH7DVll1j+bKgCVCreB10BgJzOj4
ESWqXPnwuiB6OmJtWTirCmbooniLcNZomGPQaSWxnP0XEJvBeStAg9UjZOp0ZNrTRkZ3GWmVKfYC
20neiI82tDZ1+JL6WMp5WX0I4PmK1QBFVgV442FW02Qv6bMOTnVM3jwQrc6Y5q1fOfPW95zQOgzQ
Tyn98Tofp3jhrwnnGVcI4biHYU6BiwJRVucxusB1km0BZq8GW/8bepkIldwGQ0iyZLcpbg74sLoC
Cuqy3KVbh+j//tq+TniVUBmhPSzuvYnNaztJvGmHyymO1Rxoi3GxllWcmzO9POlBGRDYXlmTOjBU
2B80PR8SnrsLT67W9EL8NvqQ2M3hGbOF1k7marjABJjMW4Loq/boyQtuFhgGShcIeBJnL6vW5fHm
cMLo/GdnPLW5NC35bMSJuF6lq5PlDr5K19TNy9o9lLbCQm9LFhw8cTZ3oVFREAZXzHaN5AedSJL5
6rAzzbkvPrFqkWsRe0Jfp7n4gTNR9bCCROAlPaFSK/75nkrHz/By5c1h2k6rxn7Z1gTV34CxwTPK
xqaC5mcZ6qUsifaS6bbPd5zIKAzC57dFZSXH2LnO+bwR0ugs8ik6VQ9VChUr+kzWuNKGm/hsM2bz
hR57Y1v8btnXU6WnovA6SHb8wgCA75oYEcB3KWR+lxT+1YuI5Wc4Lv7Brz65S6dZX4FtJqvZKDRc
517ie9KvlKeyT5fx9KN7drY0MhPg0lbBihnRSOVbXwayGIz1XerRuH3oOsE9/WOLKqT0BEtwmewm
FO7h7vckOVq3WtmZAw1zvbVPb7sPHQzbpp0tO14c2tYjkYlX9WiijBwBgqIAwa9zZzoICMryiRlM
97BIn6+NSPnXYugh9/y9m8RRwJonSOWwABuT8ybZzqNdTSZSwfMv304cXBZ7Lw6GFxthRxyiztYe
NNjWGhiwOLY0UKShtCxm/BU5tMU6ujxdk0NsaxgCQEjB9rjrtEgxulvCSMrHz/SzOimX6ZwaZrmb
BmwPZnUL9ATM9SlPreV5wPaYK0ZJ+qDziOj+wZvNTvjuPnyaZJXMd8qOQjJ71+3ephqMmsV73ien
yA9za/42qxWZ2Rp5c6FdLWFwOKhr/h71z+aXnt6rbtroJBCxbc6guZ9nmXuEqtniRAXsF5X2NLj8
ulpBOkKGtW/Webkr8nkDQcgf4RWT+Wml2BM0+Tgp72chIeWtkYYLRJ/03vmUmoIJpa+eAWXh21F8
+Zj+7++9uHmUzxy2T44d7ub7kOu2DLtvKJpNPWo9Y87nIMfqPh47Rn9tE/s9q1oaEOj9KdXIZRpC
14k/7sR7cUxAkaxQW0KDAqz1wLo6yERhVXjsns7C6rjqbI8cRXMsWH1t1WWiJOnQnibfKiRoecNq
82TZq2uTQX1AwDw5oDD1MtRPmCODSEbfSyjC8KvX+oAXgYC88JrUXB+nQtdlDayJNF/XedLVfPWT
7a6YBcqI7whMM2SNzzUjORjYfmrJWmadsNc+7EHpSsEtyplz1EfeWBJ2iJEBMcmNy3D7yZE80xUr
VrS0Ym9uSHeC2GJ717CLA5DtN7PcJn1+7QdEQXN+4EIrLxXHYTyhJ5OQvYb77ZIbIoj1sfsanXVf
QFKB3UXRWkbo+qgf7/oiabAnHWZPnazr15kPL6wH08BnBMaFPmiSSwJ+X2OMIDxnOYvsT0luP6kP
UQH8qzH5041qb50j55GPM8Xkb/ToCazjYw74def34bxdHnlJTqNItyEA4DIN4+ICFNA5SJOD7dwl
67AE3/9ROtvXNyS6ORj6WFr39lRNb0/wJNIEaVMhW7V/hNXzS1U06DaI5jSvDWCNFqJ0fQOlQyl3
DPtn8R0I06JkBjrlYDBEc6nR6/TrIsLoxQOvq/K1o6HrBMJsrB7Gj2gOhrimYN/GmeivOxk6x/DR
JnKuKW/ATBZJC5tmQqdGOQQ+m1rhbHWS7fZyAlaSUla4XWss2mftG8uq8mF6Ohh8W8mIsNy7X5OG
Nz47oNgiJGGSdFLcssT8aZnSfntcg5FZHYqhT2pPmyBCjGHqGFu/DppGe9RKjS8Njg9iDFEB5723
kB9J9d1Lx0rn7vr2fUVvpbO7k8KKMTzTj+Y5I9NqO9AvKADL1HYdv95ZgTI1gyaIsqjWCOrrVaWD
pxj2ubbjApau9vCkeCbPnEbAJHEqeGfbjAsYAfk2tM6XAO6Wm2/i2kyCqXQ6mNDx9zd1dDFng1J5
nWw/j+Us8JKaTqALF251uEfY1tJy2X3eEHia2OZNyljxGNfdjGDCUougQ1kPs7e+ie4P7AA6/Byu
CAxIg62ssAjxCkXCj0YRu3yuEcyh4QpIZphjwT9z9IdSwyz88B6x8beQJcqzZF6DJTeOyWC6dlGN
xytu9hJxaRMyqslgPXmsr9cM2sfLmD3NHQT/3sQ2ppaDn4lP5y9kXBG81qSbPQHgnXjfkkuEvgYD
PAFZH77ne2VMY1lgSRk2dSBsqqHiYyErsOMfame2GVOC5mfyHn1o1vN9nZ005PQFSNrukw2L8n70
v0raezqFGQkm375cfDZBL+Y/2f0raFZFYUNPkn7Xc+DTEtp8cD1QP/g9SgyUgOsqUv1uJLlwJocF
c/uGOZ58xAZEIquYkEg004OEsxLKCNmI2TyVJKN/yIPYmRjIbrsSk8rfdJgclzzJ8IllqEEAvHcO
9emtoeUAGvcglryR8VIklgX+/a5ujB6HnQ9qFVbJFaloPSrOXZfNr419AYdv06Vu54msn/ySGV7G
w+1/MQV+OfNMj3CjaKMJPBNpvl8+ovDj0AfzVaMOam2vAwsaUxe6Gt2cqyNwuen6yJk+c7Srwhaw
4glmJZshnffVZuuR0m07F13ef1L0VQsO7MGFnVM38HZkXNBnzTuSfXVJmUro/tDSQnEmDufclBd7
KKy1K4FEqzIj+gjJEBevInTxV3S5kc4BNokDbUjDvXpB1ZLO7QmDJ7HgsvLXgcJlWcyj4fdM3t/N
04dHbGOQvgEOHlw4yDQjRKwW1z3oSahOuh/MM98FLdyjxGi3pn1jW5SOe0T7NXmb9S/HTyBfdQ0v
JPyFtl46hCqxZWmYQPVpQ91l0Pv6n+0laQl+AZDoRoXjKBzF22OGPi3ZmYY3O6PUpnE16UiAkEux
TnwZlS0NqL7/luc1UHaH2mkp9E9aReyduWgF0jTcbmjkuJTASsECcDGkiAFhvFiXUhG50/YeXrNP
WPKxuiXGyN1EM7e20xKOUq6hfE8rP+Y5bO1XXfNR4ViGC3a7QJ9rmXml+IhLTEsPX0zBdKuL52ED
E+9K4Dmui7XC/VfUJ8/swSmKUbhwdO3m9kAosce1PPw2wrEZMhagZo0CUiMZl75pCyBjMnKVWqF2
cBx0mLM4aDLF5hqYYPXCPYj4VmsrG7IF/ydQSgmpwPpUSd3hRG2dSXwp91vvkCRsxON0ntBCV7bj
w06LAw==
`protect end_protected
