`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 483952)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbB/zJnlY9bLi0AUFrGn2gHL2x2kzl
0IsX27FVgcMWfMl9OdFIqozeSXmU2Cn4rzjESnXs6sgVgzjnzbkmon8bqAppdChymlUeUXyp5tOS
roiZbQGvOJcdEVGxX0I7tr4Ukx8lhyVsDL7KMAxNSstXvy0BRYMUPR0c9bfbO574MrlTltvniZ/6
HLGdXgC6XWlW4W5V2qIoLO+J3uOACngXdPKgdUklQLVTKz1188/cj+CB51Ok91ICh3CV3cnsWgPQ
0kz4dykKTv3Wc7BjsaRCwMhNFXQmoBvvXz5qBPQqYfwiQjTFsVoIFHSEUZA7sjh6/30/J7A7n00Q
Q8UbxL/+xjTt+enLda63nEm/ZhT757ypDpo9Citm3tBTcZpZ8rEGZ2mLMneJddgnndwOl9zZt2Go
vofjf6NJW4zTPAeFpbb7a+etRhJuqeIZdYtK/1QhE8jcaIi0BaSB4L73IEC4cypCrbiG0kjW0C1U
xQ2aWQMJFq7FyJvPt2owmMS5aa+gniZ5Ow/s1DY9Ep6c+k8DrRIDJmd+c612T4ReX4GSgjmgGcQT
lWJ1Hs8n5/lv9RvgPKsdAiEWe1uGRdeVJ8peCIBdv5ZHH6SAKzaeRnZGxMqaK4dXQTmySaLMynLC
kCap1nXcbl7P9uPzCu0Shc/mgsnWtpBzVL8xqzc6kWZkXsahjXtqFTlb8sTMXC02cBdD37nup8u1
+mHN3h8bLwrFBLmZMp9eFkiEps1HHyeBXLN0noBOT0s7geguNpw1tF2I8YssQ2B/F/C8Tw07Rfrz
Kou/cza5XDPFjWSkZ+dzdc/5zWrFpZU/EntJ4JXXoD+PtBFzCgBf2S6aNIYL4Hsu3tdMvSx83Csa
cl7/D/DEaaFw3mddDsmb5hqroTGJw1B4YCl1sEaOZDNlypn3Gz9nhQqXkD0WXVbz4ARWRTg5cGgo
yTPb1TyPk7gRC7ighh7s5hGsKkRkCNlz/760z0RzdXx52IydJAN24hW3zTfjyVXOzZk4BKO/f90N
6SPNeT3i/6XKc6/TN1WCT1I4ul0A0vvDscg8in6ZT1EZTUQIS6Cyoi1B0VLQFVw65NjTq03VaiJw
+JtZtEpncLbZG8jJXDkufLGtgvwLRPUNaUMpUlbDL38wZJSr0g8ZJjWJ6RElo6kb+cDcOMZdKfRy
RTU2l86z368XKlJ48yRj8s+ycQ0UO4KadqVufMMDxM+20O9osMpLTIXKzgMTBH+IiEb5gi+zwGNd
cT+RambsF3lyIZeCutMp+YJ+PMA3OYzCr0Btme2CZq/35Xw/4NXLV6Iwm4dnZ7cFbo7JUhiGZ9vs
SJo0848DFlVyrnIYo7X5SRRuUljVK+7w0TCcVoB/FEt0GsL3IcEMYFZTfr2baSNd8gkLX+vQoFGM
8lNv1yX0+CfKLR9/TltjTj6vt9ndUj2Hn83e3WdDxyuwTup1Nzu527J84mR+RHUjEkrF75D9oD8W
OkkdqHlmwwB8nX1qh948LgoKCoqjkLwinT1VxKWbA+jaj3TYWVsiO/AbOlqj20UGSTgt8BfGhkur
urGeH0h3jUkI/N3tKfw12I9dStxXdrQPdLU4UgTQwnUm/BTfRHBiRiTnIaantsOeRJFfAY0aA5Az
SfgvXU7f8hIa2tqKqDrYvd0oNCiIZbCOA0Gl1f2FlJfyk1CE+JKiA/5DSNFr+V44MEEbH5YxkvYb
yZxq684d5P7EYz1/RkZR/2B7dMGToBJ4nD9ZssyCVZ3nzgYH8YWxGPUTvshzhCWnW7sAkhMXs/M8
C2Habamugao1ChVHrwtK3gQGtzAzqYbXymzelUMGXIaocilPyyfEkxf2ExBzxKx4Ul9HiT/oKEe+
s9NLBl4V/hiLn5c9PGk2OD8dm1u9MuClS89u09bAPIVMRxLZ16bHlgk5YPQVAP9Oq5loJwuv6dsD
0rSBvrynFdh7h1q7WHFXZtRjDM4yIzTjflxbealqEh/AMFCTP4PsRdCx0fy8rP+s7oCTsv2jj03f
7deh+xvirPkJVhX+V+whjiPlxBA8YyO7rNKVv1SQRYpvzGE9qhH6aXyffTaiq6IF6DxR/fmReWv6
Goyw1CDvfAUtZx71FWqbtlC6+2Os3wuzpmsYSseUyL4JUDFK+O1hl/dTL9wbKuY9poxwsOfh8E5R
LciwkJu4LTzAe3hT35jXYnlJRZPxaPyyW1q0eCZQ31c7dcbupofu9MiEBYkChtpvjDKn7rthHm7/
H7dwhdLLugBP2uTi7HNRKiBcf+SV8Xod9x9TicxTUgpmyA7KI5eLwjfe9Msr99WthAwpn3GZSefi
HKRxJiuYNX77ToyG80bxkswjZliPRO7fJ/xCAkrAlB7McbHSTpJiXBJC67kFc7eYvz+n9jMZjhT0
/LRhInb+ONfrxYlLWPi4YxroWV7THAHYJJaeE71sHqlRu564Rz+yC8UJfA0ANwkfJxmkLJ4bupMd
P5rbZZDWyfMLzL447jnGmTUfaILBKS+LC8Dy2pFW0D7JQX2X98d7pCJQMARQ5ht21rs8ChH4UxAS
f7LuOIp0ATDpIg1f6UuMcH6I20h5p2ckzlIgJ5GZFT0z6b3rwyf1lhIDcYc9IQps/1O/WojSLx/7
00BbhZWitbBYYL3P0n4JSkelPVlgNaNER2FKJ20dRHM06u0ur5p+8G4Vduh4gcdCCZ3IEQnAcwId
+n9PYhc1U5SpXdXp4mko2rFM+3+twKO9AzMirOZ+ICGNlnooLprvDxY+O5KK6WJnu0t4zbzw5n5v
IVPgdtK1WVE2ZugF40zkUcekSccmxm40ziScDYtLCuXz+T0EAWXvT1oSc6kQkHx57mLA91VE1wjt
HBAzU5JNb161vz98uEqVl4SYbST4Ykw5KEWwDyQ22n92KapoDxj5oDHGN7Y04UApsXhzfQr8BffV
fi0bZDq2G+HlnRp2urL4z9+25aNtMQq7hOuWm4ArLNuac8rHDWbcaB6g2Z9CKkDimEjOGol6oVpT
lyDLwpIu06CnnSzYy3aHmA2PTobEE/Qg1YPrUR64U2/GF6NDeSlxbj0uTA8AfAhWrr5JvCTRGpnh
/VVkppKCB3K0q5MeG2ewRIIFNE/Wx3bUzE49TnMGQJTExJrzeOl4EhWkOdYxh/f/Pg/siTh594aR
3AUL2ttIPgFxXz5cl4WznOPgAob5QAxJH7ozPaVrNnp4HDDLI5oXjAvc4bq3KCfqtIv2fHex9JlU
RzDnjeIlad8Iw0atFXXWGOZM7P4EKul1/iGoUFwrHEjgEYFb9XGy7S1JpnsfhUxXRUVH3rZq1VTo
nGz+1h65sZrAP9DZjfLp8ilQOevteG44OyQyg3Y/vgTNdy+N+0yF1r5v1y2TW1EN+Y/Qk48U6NTS
EH6sJ3ZhE3Wwn38DPPX+ETY1pdewfyFmtwHKYF9vi6uhPZlRNkKP9lvFNneer8FJqtzvrcPeqrIE
vzXheZ/e904FBB/keokTc2b73rPWDQD9+tTskJ9IIsMgb7wMW5MJEUZ3zhCRDWcGRkZLEBgb5xo6
gssSBXNuyB0tr7Gakf9NTBf3IirvWoJR4yJjU/w8f74HKjWS+nuPXn9tz15tc6n+DvvVONCDj1uz
SLj1JyYdEGAr6MJyZMZbwhI3ArLgQtlrl23VtJ1PoYO7d66aqBhwqzqrI5E937Q+zSIzJszUM1bH
FwxBjgqUyFxCDEN6Qmz5oomgk3J8AfaubfuVMp+GlJr5DJpgOL4IchFjrvwdF+uxbL3gH/n6AwAX
6bI61EzF4QbUXqNKaFvLwOA1QrfoyB192RDGg8DiJ/HY8NXlLjyC2WMiR4CIT4xK22QmjrelfHQl
CmquYWj5tSX+5FxXGbIK0z/vTol1h7SGUor8g86ipRt78IaZKRzABNKX2AiVuYJkBgE23vZ0Xfft
40HFcpmktljtLGQzSKMdGflt7ATUe/TswOQcBk/E8UupuorM+BgEE0i7ZvX3YBrt8fDOMH9M1jfS
rxEYlQQFq7HD1oVk/oFlgunuYzmVjf4z/cqX9nlSYcGZjonaaLToM7FBJAfeDGbmo9ZrjWsljHf2
/4YQgWNxXCs/aKFFBiPkZMX/Pe0traHO0LFfJyxMSmll7pj1RjmhNaJ4L+yLM80EL7pZSTK4XkRM
5TE+6zzX2XS/8s3EbSf+MVg2AEQzfmBq0zcBs5/XdDOQW20UiwLpog1yn1kMtLeBLkz3eRP9+qK2
7uZsMmW/uSzAE8e7R11ws7IUXIYDXAVRFyXfHhqUBvJYzbJsxWnjaUrRW99we5aDSbqa69lP/0rE
3LomLRkfYlG22Bzu21OfSEa79JL85wvp6ZuGimM46IHd2vDvGuV4bSG9uWlkN4MOn931n4CRoBTM
geaFeICpbKD4OWn73YLP0+65DYKHZo2bgXwlaheVTnffkHypO//dal37XI0xr19butHl92BDqysp
C/ewmjhuOG4HUZ2rL6guYG6nwHbcWRZr/lUsdyXk/J+LEV/iMfUgWLKxWUEypxu3UTxEZJBFsDW5
vOUsaYtVTphhTMU1mD2sLPR3qrqXa2X3xugyFHXkw2JeN+47vxzKz05aSHxB+zhTctAn0pXk2+Pt
EyVNkMdKBBKYYenU1zB0okj7dnuZiW4OiCcYRjvE89bLibhBNHFZPrYkjjH4r5mAp8FgzNh8WGmx
30Zpypfd3GGVqiNtEa42Hu3TMoJ5QmDX0kpD6Few/3RMkQ6ZszLE9NS39BGYYZ2h/POoYralDW2v
5gI1Kal7Oc9puLHbKB8G+M96ZVX+A7Ha31b9+E8V18D+nSgyp1rY6IEUv6oZRnrW81DuTEL4gg2s
psx0HwVmpfczX2NXueri1uadC5yH+cDjqtQytzV/Ub1TzRe03bwtHy3IjisvVvbuiV531BVRHdRT
YjNV4EQThGkQxWGCxT2BPxDdKHXN3ldHjYLaRvkSfddkobj3Z2fEw+FnO3BLb2EBubMJETNDzPLc
HwL3bgy5B7Ks3/Ca0whwTF8Re4/DbevEJqjNx+tcoFBMhbvIWDpAQN8Q+2L/luPZese/MPQHB0q0
NSytbxMGjsMDPR2WOFFGOiWDYaLkLeLM48p+WOMr0J8BR6BihGA/QqV0SbFlymNQ2Y8St6bLU2Vb
6zJ/mIA1bIKsk1fP+Qvvhw6HmxeiZnobCMoDOHrP43dTnua/N+aJUs4J5WaYjDrTikJAtkP9QY0t
NxEBLwAAO35uO+0oGqzRg9H0u86FjuZbDDFR5YcukByg/aSTQwrhpZd50MtozwqbIXh/0GbYlYaB
hcLIknIpmDT8ZHx9gvwsHFfKBaXyrSYlLYNZSyy8vP6YmKGdSmy0v9BaQCCQdpsfUnDv1QKe54w6
qmx9YFRD8J8H4hYwu5lIHgtpCoUR4eSVxbNdM9rN6SH/p9vwVTdE7H6b/AkDiGv6LMq2hfr1kjZE
y5HnjnFhffdDBA2ECXsEbo2/T3BD0bkNjDQL86qzGcIzKh7NH6JTlTmY5Ns9Py6NhzQCsele+/pB
eVyLlEeyHwaPepe0ehK5w8PZv+wc76aPia92sHU/OLVcjvVcAf789E5HJDxP55AKhpRcB3gS/wbn
oLLXwyMPCKfMsF0JIYIaXIhO2/xVR/BwW0iTullDaifpk1WQZCiOECjAZKaxKdyZFSnRTZTg6wnN
7uhpdQINoC9Mu2z2h5AOTk0nut9s6JWCF8jpRgyQZCGpko7Hplu7G3ZgWnytIlpFg3a4bZL7S6+G
zcZNj/uR5d6NCgu1UkGgYKsTXB0lckEO7aeAVo2P8fCu6cqEIINnMxJNMBPlG1KUpZzphzOSeBRJ
kf8Mn9ncCgm+A8PbXgGBQUSLni7ZLMMExKT/Nsrum81/f10+ZaBDjRvKbU7WU6+oLWKy1vYSV6Os
qynOzN6ezGXter5jRP5Hj3fc49ilXINff9xmpefquhf2FAUi/vCVkDeMrZhVbh6MXRZyuROgYZ2l
4q8LHBn8EUyvFqicJ2cm0MwmhP7YJ0wbOEeVhQyR9Idc4hCjhe7Ft54M6o5Buvxai4N+D83RKo6T
TmuH3gR2GVPCnKOLEi+n7X8cCi2SHV/IIyoC3gogoTND3hNkcsxD7Hvpz0LyZb0dXDFc9zRvyVWX
J8sn5o7wNCV0eYXTX3dH8p4nUIWxz76/O1QgpW0eT0IVtTp23PKjpJpZ1IsJYhCJJAwbG+4fBhX1
p9NGR/KzjkxXIZW9sJJ/JXFVshw1yX5mfAR0eedoXvMw008Q9CoB7R2pRlPz57qDJCBk4KUe/+OE
j2x5EB4V390ZdRrw5KpXCLW6NqyhrVa5SSa58oxckuSpSdZUnJIhiXxDi8nPVqfZ6NzT00EzvuSa
gg0R9YYaQVGCc/k1k1nZe9ld1jy0ahCe3HsJO6Bzi2munWFt7L7hOOzDfwfea/AEStBLPlMX4A/u
8tgZfJRYog6wFDzxKvQiQrIc98nGjl21qLE0Z56/CeKIhIIBHnKzQdaiuhhRNPI7gZG1ISgwJDCV
ruDmRTrm687kgPP7sezAv1pze6eqFa5554XlUR/Pab80c9zAHZpJ8Nj9AOYbU4ILEW6z8olGFu5O
z/strBAkYAnYKBgO8/U6AqtOck2fBvdfUCS6xhG38/B/V8EpZ01knCbddsP/mKsAzwsgW7IgATU/
epr3AG/4PKj+mKlDZa7zPp7R4MVaBBHYGC46XcAtfs0lJRXhsZl4oGlvyfcKuKGStFP//GwLsK7G
uzM+Zu/9uQ/hDGOcf0ECZJM/aKRgHm3eaAttA4o5J7x/DkgmcOKdhGqu48G4lbJEpmfmg09wcO21
JiZRrdDoLqJF6QhTeFZu7XtwF68B84Vi5IOy/Mi6GpdSFpfnioBtb3sOMlCtkmadDzYj1zOWWNfW
uOYOepWrfofNi9bgIVLDk1s2XfHS5Z/huMBnxIymvdBo1Atk+XEqSmZYLcfA1s0wDJpv4xG2Wwp8
oNaWxdSC5C6s6zuTEYCF0HaUmOTGIXuLcjSzqTWU3m1j5+ncRBQIO/LtHVaY6kvBi6nSfBsWcOJ6
XYouE2oEdumdOTS0trXOMaGVDU0FcQbQ8M3sPj2G4LtOcfJ4nO23fjJygTuXZBTEVAa63SVlDEz1
gUNpC9aufbZQEUwKQbv77bgRN/xOodBU7E6OQPqVqrpxRfT+vzJYWJQe1twY+41mHAj2vTis3tQR
LLusWDu48ga9LPAqsNkh9s+CD4+RwClNAfcMNOakNdHBqvuu7lzB3NIpQHF+aKctxhgFwRxaI+Pz
91I3RIsx+usjzFhGJwKI2acBZIwAtCvSChfzCBnnxPep8Le6gFgwD579q9SaCzExlbmQzI/aGVKI
aAEo4VBduWERoQWnFeR8W9n0i3sgzanbfpjxiH8zcKDiuvIMvKplh5k9V7dbSBwueekx4Xi6NF2f
iww9GX5dkZqFUVpeAUTptCdwI7SiBuIRa0e85MNUYK/2KR9NC+5n1wbflK25tLSwCi7mWRy6fdic
jlv8MbzJD+ui6LOf328bmshTKAxeZVlOj4bc5AliObX4c0zNXdgYHa/FzxJZ5sQS826y/vWc66pC
JNf3LeOajLaDIItpRo1Bb4d2tS4Ak7jc7MrbKnwe2Z4nlNPO2aDz4thtzgdyjYWniyDr9+9Ybm6F
M3OyV8N/GBiHOXWJZD7C9KupSY/PKx97MwAc3l3Hztp1h3OVHAh8HK4pBGL9YrMyEKqYlz7Q2mk2
BLeEBc/xtQcojsmXyur6fCDzMD9jgUAl+4StscjU0OYh1UeREcaeh2QGdhVuI5k8hjDpiX+JM8VM
gZ/8u2lP+977p/5aSXB6lL8fFJOmq1Dhu7BUh2Qvtk5k393+JPa9tHRG+IS3QsJMmlFD1/NmWl1i
eK0rMfcOg5jAUhMBKFbHfN5zLAagycwuXfR/xEqjLEHuJy1hQg0/0oY2aEGHO3w4GIXnk7Ze/zI2
zhwBv4URBVx7fVna6aGJAfN+KvAD0iwGqfzlM0nMX0rhHD4GrHdXmI3HpevxM2DI30cc75dq/vAm
o9aIaN3FkZRlb+RPCsEEvuwmBmgBnWkxuIBD/Np14sH9IAFkg8PgVJZT6IzWjt+5Is2E2k0DhuVP
h3EdHnBt/UC7QezgMryadTJsk7m7utEX7qyWSfWWBPA54ELqhTy65d3FIfuAk6qjo5GEsF47W69r
H1riTDL4QjoMuuEgCIRq+w2Hqc1QaDJvSG8yz0F4X3hLI/YXFvkYa0xt3FXY034/KXCtPcmDQ4uV
3iKK9j4mm0EGFhbwvKeLWRmLDbtOwIbXGs7ncQ4ciUI4tXe+4Z9rtWWYNmGDDTTjtuhB3p4MCK3g
eXLX6HdDm9X2SBwvRV3hk5wOxdgOvpjhfJcVfgF7odXebfoLJmkR7vKnFLI8WbxZ0n+eZuo6Uh6/
JA4P4ao5brg7zVxqSEqHTcSFDo6tZwHJLfDgzhyAPq+awHwKewVVDDMV4HkJdcSZZeV0fhcnBdyT
HqTfiGBxjrEkC3WnrXyXx5Vqnsz5ygpJHcmogXbEp6AL4IFZq+6VVxumDQoWdcF+3STaA9DkR/zN
OyPQZ2R8WWU19YdudxfA2zUmBYGM5DmCxMxMCH6hFb4PywAdYlzqR4XK3ZoctXgR2RlS6S8Yh/So
YbVzI5kfqOTvygfI+wKPgGdFZr4l//Mfj68Z+x25IJfDrJL3nTr00G+WDws7MUgISYmq3zKiklp4
XmxyAPzF9m8IIk613ijOBqp1HCeIomwwSpXLep88UCJOAAjSY3BmZzA21tWYqS6nHDRpMCRShUjG
SIc91t0BnlViTA/vV5vc8i3igpmppN/c7sN3NsQ3mLdcXp1xZHvpH2cvkl5HfbMgZsG4VWrw2//j
AQpjrWoiLaKC89OygdYYyDjtd2rE/qS9BEN9ljPrBJGNNrgqp8+eqx0xwMu55OC4bAQ9kD3pnue7
xlPLnd9uYDnNiRbJkqpNNCwXpSZkK7Eiu3OURDUagEpCJP3gf/9nXqneIHIpTyvqMP4ULanoTVHk
KxSHpSVdwpzQc3t7euasNOdNlOxHbrEd5kkH2tyREVap1mND0WaNHx685vOMJXuUvJheVpAajzGQ
WTQQPRuuLY6bfKnSnA2pzTu3DneIdAaQSDm1EVXx5Tw4CX3FY4qoxkApVuY134snajzVO8f7Zzo2
gm+Cfy8CxLT5FSKH9+CdP6tAgfL3PTcOyjjCCpgbDJufpYIRMW1d9PqXb8JrdCMELswo6fOO7ipz
7ZQJy/i9GO38ZnewQI2EQPUsffWaRGWVZb0ehc0VM0zzk90prplzhy38p9DppQ6XTarRBOEOJ4St
5EvGxyxgMpMsJ70V31WxUUbKGNVEaB/l1SnFO+rzvQcDfJXw8o95l85oeisDO+zjgynZlvust5lD
v16z6ML4cxSQeUVbtOaaXAHXboqtNbsAiNtf6aXvv1qxWMO/v7hGEnMYd4uK6at523FJMOGn2Vn9
iha3RuH1n8OE1PSYnEMMhJsF47A3dge/F9XaY+5lwT1VUTXmFR1Sxya5AOC/tso/BvSht/WoCLbi
fFkPA8cxkkaDMfvwN0PkF4SpN3UO0n//8/+Kv2NwtaW+S4GlEDxU41pXxyYmVhZl829qYwULWneH
0cwmSP5oQQI1So0xRSPpm/CpcKk0ULKirxIgBB4yaDdEjDkTwXarw1VvRyd5B3Q7eBA16nErRBz1
jvjSpJwThjAMQ0oMPCr/yniSbpRicsACU7xjkUMZcWwwsw35VyTNy7QEZHtSg6EXBusmPw/02fb1
uaB5ZntWaD1yThgjACndfXPUHY79xcII7Xs0BaxLgbXk3IaJ857/Up08ENLIN+DOppoRmNm2cCY3
FwLoHamEb+lZwbPUkb8thwm3qxOXA+OKXifeQeezPUsRtYvWInsUAro6L+yPjS0JAU/mRvPbNJik
sKE9pxxWxagSWwGlweAiOGhuaMqcdlyHtlf6RtoPDSTvuVuyhAXvTLocaeT38NGh/DZaKK2A87fL
GCust+BBzI2VJsQnuWj8Ki08jfYAXKD08Qy9F4twiPIf1h7JSFKdNgCo/GwfCOAbl5iImFGdvG2X
5yTL2bmAMsAwztDUgI1pS81dD4eefclVWlQHgt4GjlF6bkR9Cz5SQWrWO/DPzJgX/bxxcICyAcwe
4EEN6A/UuU/deCgWy2f9+Km2W2px7ZL+UAPcsNK3RCvb/Tvnjj9q9jZSYp1Y5wecf3RtM0rpL/8L
nboyf8mhcLuPno/XoCBa/9U0FlhtlF5daLLuy35670mUKORibMS0fFd/2J+IKCYZAjaxr/6SztLQ
vfjUM2eXN4ngzfXYvIqtVhZHCbNcPrW5p88knA9Ni0bRD4n3/C8qeL16yMXx+yvp7JrHfTlzYM4p
JdydcCypEkdtcxF9XvKdjRyjdOYGygltFgc6Au2d2Xhzi/yrJk31Vu5O/mtIjcm58Dc6XePAKGQB
davzoGZSRGEpD8nswuTB+jdcEAVUd7VtqnH9IDUaCf7b00g1liNe1B4+eQNzm25HtIgPnQex9qNZ
Ev1crkG0UgpdKfQRmMiHiflffbnqEwHDuCFXjb/v9IqK5LvDrertaxPetOxdc9avnDrEQUkeonf7
KXW+0NKy9R2l4zWBc45MYAt2Utm4OpW9VyTb0DKW8nfximN3cD39+UjKTY7xSOSZ5UHcHjvujEFo
E4OH+G4ExGV+aofOSPA91PB9nsfxU2Pd0CI3/9YIwQ3fr0J00v8TDfmYuPYAloOs+z5rC4gycsXr
fPU5sbiNHaiVMx75vzT/clGuUrxrhKKyOZ89UZsx3myDgPw4++rYTM4j1HZ49QSy5UanbyJURAkn
MH143eF64qZz+aRNi0m+yI1okkqp8WTcYxKqMEDqWb+2ui2E4/CoYK7f8+MZ1YV6hJfFgF4zvOYc
kdZ0T98SrSlLhFOXp6U4N/nJO+ays5LCbbT12A3ZGGgl30ubHlCLYOKEKn9TlrsNei+Xug2IhoMQ
jRMDqWKhaLhgwwsrFODIbpmI0IAJ0ZHBnSKujWTw90b6d5Ko+eIPouQxIqM38URTmRFKd9TbzWNC
78nOZQefDnvDaliIqqFd5in5c+SwhUoO2yuOZU3mlfpmvkGKOUBykg3Nf4gGBU4DwIwtYH4z6zM/
ebzslxaZyC8bbFktajF8Dd7nUXBizkP0gY5hX0sI4xyka2oaOB0gxduhnHc3DneUVf6+ySpZe32B
2PKHTbv6lGUhTz+6/uu9oxYay5DTCi8BdqW5irga0yTEwVD1BpTCfdl8GQQwt3+Ceol2un/8uvSF
UVozzVVtJWaK0YwQjGVLoRoxQrfZNhy8CA8WUG/7BEn7PTWuQVBdkzuwy92jx2nWMHyGEDIW3xip
e6DtFXl0xtp3byVjfOGHqMLDVSWwdjNKhGBrgBvdWECLWQa53Lq8DnhL3ntlYPcqawmMQbSv1u+u
IhzBGuy+iV900qzSzHqkTfZ/sCHvVDVjJGRidwhAgM1WYr4wjr41hY725otx3GQcj8cLcgGtauOR
m6Nq6RMrBeuOakbQeUHaJdkz7bKWP85AOTYflTkGJtOuacdQp06phLVmGpGh9T5GCWmdAsP45a1/
pBiRnJu7tbSlNthCdVvwaLuy47OxLtI/1NEScL4gQWk/G2eaab9bnwZrqXS8mwlhyDZBLfDAtpMv
PqS6Ri1/ctCwtzb6hYjlbkWZmVjaypgeZmjXga5vDIhphCD6ArlzZ5v5k2ItOWK/lNH1gnD0qmbt
sAJezipGKY+R9HKd3A1NfltwmxZ11mZNljlWeWNNr7TcWqlbXHeK+lSUNrOtLViW84d+/r3mS6Wk
MVj+GxduiDWyEexCFy4f9MUBURbSOT/9bUkDwqNca5inT0cOPaGliu5g64o9+LzziYAwS8uQ9ISz
RNlD6C0ZTmCtXskOaw2M6a7X6hh/ly7h48xV2w3RkyGntkwZTALBNDZZwyMqRcsMfHRhjf+ILGzA
zRHEv0cI26Rh6XJIArz8mH2HNIej0jjxiCmQKRLL1g4M8Mq1rKSNGrnoUb5LDuDmJUtYRe9pdFdK
YJTydYq/TVudScVNqqvDpCyi6p8c2EWnPnVH6+tYHvgDszPfMUVBMErWcCGDV1DR/MFGlNet0Y2g
DtJnNrGqvf6hGe0Enk7wXGsuBkLoVpfTacBSknFJXROPJdfo1lnljETlvkj25NBTE6H4PFZbL5Si
8NbSUzRGuqGDn8Ve4QFlbKY4j0EnWBG15jx5+cBxKRcvBMRlBqY/xntg1C+SPzXJmmN2dnkxdzUs
Udy3VSdZjSHh4rptd0KvHQaUEPpyQHnQoUlv+nokScaMFWfwP8I26LcpaLhNr3MH4VuT3TDSIt0I
UGEi5Tlokhf3NiutLo3w0QdRbkzAnjIxDoSIZzuxit3kht/Spt9/iGaC2iAj3g0IWv3X+fs8QY4a
w4ZIaT76QQcUiRG0+anUnnq1agg+QfhNMZvRpA6xRPD268mXW5AADZXeRWYdi83vfZyxqKnh5P5b
jsIvUBxEFOBeGh5ihWKJjyseDSBp+SMwAARhN0t/uwKHjaduLt8+ftnGkkVH8IxE+Wgu8xHqktoO
EnBKVpUbSyiI3TZ5uOf0p6xoadcuaWJLPCRwO/Bknssl4sFrAkSbCvGbap1dI3OmYYtTxtgMA1XB
Xwqga1q72kao/tUUg7KLYDW7vpNMyb2QZ2FpmcvIDDsqrQXg3hz/ugwh4xP8787hbyvsKgY4J2Ix
y9QTBQKjJJ8HEtcAjU3L3b9/Jjv6d8Kfo6LL47/sCuscOCwCc0vkYz7rJpzrzpxg8azdxBcVuery
5Bk3DCdHZw6N+Aj7CL3Vz61ipKzC/0YyD5kYePR0N0jaTEaV6XbHyZO/eYqHGunemp97n3fWeCzl
P7qVz7XaKbn6CD8iq+WFQIynRRkBxFgRHHRw9OJfr7MBASG1L6NUaGxaXvmTNRs1F4lvAFgmQdZR
BCpWyiic1n1ylJj+9g6Ul5moUl/epyGQKauw5rUMMsOCLZiie2YGNwe7KskZmWqy5yII8/I3KdlI
p7Lwr08zqFJD2MySbVQV2xddq0bYCxsEEvEs+MLJpgS3DxSbQbhG/EeEyDCXV57SaUQ7y0HoFR8o
gP0dKrZEo88iSvKV+RmD4rRmRgCOrBNSFCWMIe8Ig6SE07s8aiRqh/yEfvKs7+W7JJsMX+YpfY0n
Bazk+u9+Jndcl+MS4eO6yvgqBVcTbKCkb/f92z374IWJAY/TbBFNhI+IeHNWmDpcYcmusGgLEdKL
/nitZ/GYeUDW/kuXaw1Znrq25hTAhgue7X619aURDgPujoxrRqDXrtAvlZcdSCu2FTVmygFdvoZM
LtkTcK32+P8se8BykJCdeOvkwiP75Y+awcI2cjJblm8eed9HYywBLfB7cH6JYKXdQf/SWMx3Z0OX
w5qJijiDpvM6OI7f6EJXlmTdaJ9OZDLazJlDjh7QYEPD4iQXDyFeVcFpTvF3wy04GKlW1XfF+bSL
sSlVZbQpRlAhWmcz/BMXeDnRjRoCHNB34/W/IcTE5tcyIpaknffLT9oSO2fikaAfCewP9LMgTppw
ai+fxuPSowlcKMz8rlGj5o35UAPA1qPDWmD1S7XLnvKx95dXEvKuDYEX0cdQsZscAGNPgWvAPKH+
fQc11JOEktmFd8EuN6YYnMpNMF5n13H91FmoRq3wo+z+19E/iDmdqcjMUqTOJlXS1Gcpq5r8+D9n
cx79ON0+jUPyf0ZEHXjBnG9rd+9VzCHLbQjqV9JwXG4n0mpr0ROl1oPpRK+t/fN5QGNarezzui+B
66E0nX+RyBpSNhU3po7UMarfJMJpIDDFB1UGfsLiylk0J+4jsgPeW8JT2nmEOVzBZUHI94krMC8h
zbGvyQ/Tfwp47zqeIlx+eidRiOtv6tEAdW+o2QTyWEvDo6oS9t8bEAJHrJjPmsD3atC5N5Rfg/eB
zA5ppQCptlEygLCKLPsN9JK4LIPwBscsqn/hLzbYII969en2qPNF1EaOIg+hRu5tSZuc+EqrmSNc
mmb97tGZVHZIQTdrCgU6sCdB7glTyMeHGN4xNHj41GGUmQlq+5g8m2KC4Bxc+sGMSXNDes7AQj5P
kclGAqO3wt26e0071Mj4Cb0M4CpqpR5xUWcdkDDAFB5PpgDbos5jA6vrHwLHsQ01sc7/bkiALXfe
yRp2uZV2B+CVeOyb4B223wumJ5b9Ekb0JfCsJTk5IQ50ZvUboqZ8PzR2qsBuH7qRJycO4zEHC22J
3/4tzPJIaSLaou/tszSenoA6aCjVdHjPZ+ZDfJ65gBf6jocDwrr6AS7aFd3rhFV6pnk5fzkB5Aqx
G3z2N4o6UKjPF20gRQtF6FEvHSdWEx8uXFRAGcDCN8/qOnFTWJR+dyg3MMDMmuQHvFjmPn4rB9fC
g/d6fC/2JymdTI52Klzj5oJopjznZCilF+ZYuYGQ/+jnpOFRYmJq+C0nARrQi9ciWt+wAoEVj+7S
hoPVMK+awosBC7vdqL4Qmx3m78rMvdUzCia3jUZIEBYw0CYtj9HW4ibI1kNt2X1qG1t2Lq+lleSd
x9OawkEcmmFu7Q9ovYrpVjZ6hiXaStIQ2OfOu9ELjQtJaeEBhGq47DNOeTfhWRPIjgPumXSP+4+x
u4u//c4trHf2M59L/Wa862A0jIscIdET/mrV2YYYqR9dAQJSXjmIm4DXA22DTasY8DomEKiWaaEm
pGMtnr/xEc5qIxbcjq9ndw5YQ1AYAlXfbZqXuO8DxMt7gqxUjfKmFqQet7H/baWzU2Z5cBe6+bFM
MjTDxXjNgrnkpxa1DPPKLX3V2Yrx6BftGPUHL2izoW0yWyh0LZWXVVxUzFqKaSYzJlGTcaGIMWrs
aCKaOpcNqh6X73CbJXM4ftrYdhNfmSwClwvvMYyr+qxSImmByj8U325ZtDQktcBU64th//9oIajD
Nfld8j0rdFlJ6dXx0uky4hCC7T3IcFSKV5rRD+RdrROsuEzki9IDyKknEBc/5fkkKZ6YSG4YfA7G
KpXx0LtMBKw1ViJrqSP5fHkMjOyPIQdZFaQzsM/9U9A+ZXY5xiLCR6Uusr+m0ZYx/Sc905IDXrcX
9cwJG0aaUJCdfMpXh4y5WMEvRuLupdqWSHbNXsgyO/nscvtoBOTgy4t5bSYpxZ3XM1geDIGavbxK
ntyVpSfr8ZLSkduRhPyCa7C1yxup0yP9AAXTdEuHoNzB3v8bojeogXs8iz+Wz193H5j4S25hVMTs
6xGwNgbj3VbP695ZFu6v/s1hDJC8nM4DUH0cLatXcUP0UIOgcyJcltMyeBR7bAHGqNyuzsmDWYvC
ljD+ZY32Jz0pD8njC9SiiNhEiJUw7V92XjAcExfsIZ6hlY33KhLfioYfRAZF5ZwDsuIEMDdcE3ts
wnbg+SNNmuQgcJPlUuhfFf7jfFu1SW9tTrBtLMqnizmN2Xudm32rBRxcp5uyfAhuryjXkqIRMxHy
c0M7Xl5vU5B1LZGVJHMXBekSzqjyONgXHtueXP9BzaN1Mc2BL/AblIJayMiNtlEPvbgY1V0DejiM
i3yAZLKF2e1Gzne0h/zWCuXOdvWT3qrb7b1ZZAP0lmu3XPWJUSLwRQPW0jEhoJTDqEEcUaGL+2FG
NLP3iRhTVrb1I8tBG+w65e9Fxj0UiZHpK6bT8I+OeoERgWob1UeCnrgJk+0ZpJ7FjNJbTDwSpVX0
dM4Wa7kWw/Qub5QEmYxEu/IhzUww39eHJ4vfpJK1hlpS5Qiledwt2JIdR2uk3rciv2N6JLlk4DxA
V0FW6BQhZOuqowQTUnRsJ7uD7St7OYBbV5aEEsZepeZ3zxSbZTcBn/6SsDiP4fwTeS5nQ1Tqp0wA
pAahxvNGmxT7TBTmvli0iurqo6uRKDMUvhd0Q5pCZLfzlW1yna8DowXtzVqaH2M0pQyStjRRFHV8
nqxrq0RNjI1Sbp5zUnmtq18vyjJU1+7uEXXdc2m/aUw+eDl+rWu2K3dwzgu75twRwRJDdlHFdrjN
wI/mmbh/YI6TFu+L2ZZlQ6SUZAQTx7aXNrLHFl2gpMNg4zLaEPABn6u3dgQTPZNKtMx+JdIyWHEp
rTJugCF4QFLLnfISc9DrlLnv8sUW9hdgUJqQqM08xb3/Qvtkj2+GR8jZp+p6bLiSrzc2KKUXAi+0
rd0Nsi+Ne0W92IBvF7dV3MKO0GEcnpHKyDe8YhOPXzmJEWTAEJR7lRkBcGdUP7mC0LV4ttrsvIpU
OqFSLkYIZAU2RA9aDiAYMY5M3Hg4bp6H1bTDMnGfPZlKm+c4c4Yl24cqiyy9RTBy/tto7OnYeYdE
eKK5yYFXTSk+gsDS0I2masnKUGHFxAG5YxJ8pYVEUdBZbyFx49o9KtjPNGEqTt+oMyfkY91cxpEL
f8WGvmCKcmKlzGGf+BeWzikcWWmpMCiozQrtfT+H09fW84AKi+34ubRyqy1y8hP0mu9IUY0iKzAF
upclyY7Cp5UkcH7SaKjee9lPlreOni5q1pTpA8qln6QngnLkrQmnTA/LSXRBcmnqr1Lk/aP/s8oK
nudf5csbRciFUCSh/WnYd7B3D+bZmxXP/cBNw8R6MBl0O/ZYVD6Htpv7DTMuNE8ZlUCeE9UJwa7X
bPm4WmbUgKxXgNyuLipsZaq9KzMhhAvlmmvZedeA6KodFDoEtlJUfONhflL4R22o/H1KWE99Rrb5
vh6o7KM82AqH7NJB4UTr6C2ZbwqBPjbxuquhYyEQdr7tPtoEzRT5dpsw8C/yGql07dshi3xHWHtx
uNFXoXSAQQz8XX/UQcRpm+iTO7IYq81qPyXXkwLgsGuVYW/Y+tnhoVMlqj7Zu0RpLUUwiGz8rHy6
utSP3h2uXRgWe9u0NCqF2QPZ6KoUBU1jbhzmvRchmqzKZUOyRWllZZyaQxF6/FrxLQA+q9u23iqo
0IeFCAl25rgHPN5tBA2FeWEr+UGheMrk8nG32Yid9UcOJOkzvhn9esMyNz3Wcd6RJ3NJM97Rztks
ktLxy+kEuOFYrHhEhgdG1h4FQGNVnL1eyQoDs8tfVn7jYLx0mQMpdimXzMVgdLXarfsrmCkwuo4/
nMJdMmwuTCvlap70GU2nxyikKJRXpAyCH6uEEfTNC6bJvV4oa/LyPhSd1VReOuJ4MDmKUwBthqIH
xt7/ep3XbmMl745VNw0P7xaDrPdx91SK/lJm57hXON6dLtVg3doby6xgQ/7NKku5UAOIv34G+FFR
Xctn0CzmMjJ1HNt0cl58qdgssewdk+wP9FJ+AABPvH0Jdmdhw3enHL8uposTMErtUaKPyiFn138E
hs+7rev+CxB9BmzM1ne43HyDvxS7YOyoBTLLy/xpRxvS86zaRlL1tuOP2y0LJ3q4OYliKuGI8I+0
HT7kd+HOQO8AlgKW+oD3xXE1EwFptPuUOwtJ/3aOfs/kW4wq486lx1x1BmpXlGAHcm1PKBNTH7yp
nXUxtSYbXoApVjXyxtrO4SNTxl2aLZrvnsEA7dblCsBgA08cjC6ygefmh2WQRIp0ZMAVb6WEEPt3
L/ltti20VAiGrpJub6o/kYib1tH7I5bbOBMXavfX7DDqJg3+PKO8LWijNObFgkcf2ehO+Mo9meqm
v6Qn2ZenfSixOwBjW1G1+jstoATy5uYHlfkHvkB/CeEhec3tmKmXSvS2xrKdnLwKLOS4Fj7kyUr0
WjG5hxEbQXhnAoltILnfE3wLNut+TF+fkCfqgDIML08j2TfsLlBgkLR586sA65FLQyV+qsg8lBQE
nWfLlDKx65T7mbL7kYANnbD3jaRp4VqBC3ggsWlg6Joow1yY6GFtMXl+QjJ2Y/KnCNKIuxPrK5k5
n4yLk4/y2N5YwVYsHdVXgRdkWHZktrooCoP65rm8dsbGLAs/hk1qFh1HJ01giOIAISnm8lYug5NN
krMmten139eoVsN09dVNtxITdf7hzxH3Iw60IkWcku+RkwhCEztQ/ODx/Jp2YPqylHSx+6xUnHPe
EKZiqU6su1HCaG0fhWfrlXIw+WV4QdpqN4evjcXIvqgKDjVZcq0Okfd/IMdF/hj8dLNcmXwGGfOc
1l97ny35K27UwoMSBAieP7sQ+T0mRn1oDS2eRTef89Q8I14OxndEPV1UjdqZ1g/k5mib5S9Yxzh7
VANAQKBRGPBSajUHp/EjDpyaybKnkIk/QHB10oXRrChqT7TMe7oEtcM3/HVo8+ypNpaJSKajrPfo
XDE4278APKdb5N0U/x3HeNFZeXwhTzAYiPk5YlnrwYWxgDTd4GrCXSeETxgrg7qxCFpCzmPy0ZeL
aY9xG4GFWOC+9qvTnovFfYXJOgFOTu+qPOfraGaMDYBwxPeX1JFs6w7ZB6bHRzRZr6ftX1adaQJ/
FWO1XxE2ZzgLz4NV4PlfxK+nHFnLbY7LxayESvL4lziTLTR67tMaBYjtntHj2aQUWM5X4AJJ65Xl
SrPhf3vRi7+mnZwV0fkllgWmV+4d5kyn778kgp2HJE0WlLKGZnx52LNoqBSB8RUpegB8XSUE2ycY
jujPqGBsp2LcEj/RpODSBSMT+zST9dIL4PnH51RcGDQlZrCPOuIuoPYukS6QI4S4sOBIl9oszk6J
KC59U/6uN3hg9fy7tojtPNaYeY8kc5FZzCxNjfBSK2nB3o80FW4ARHpyrAG1PEB+y64vhM42smoP
WQ7r85UshLlXHBe6TGfeGtSnnx38+mpEIfCY0bF2U4K/eM3KND7AveaxxE55sfH4VEOcaOnF/ClP
hmTpZBf05ju2IzLbEOV/Eao780H3nIKvVujn8QHimunyCP5jrQDhmgYi4vPUPPeHpNHcIlM5rtvw
tRYgbvfAsMC+ZIYzn30F3LUO8zs7zJ7g2zxWiMk3nmTaMLcLYX56+0YJ9+kTGCe0TKDtzvvuam3Z
uOdKjj+PkXf2RK/O3tXSWpZJiEmF/ikwKTY1Nt1dAwmAr33s3V/j9JaxVd2h1VbUobz/MqItqyOs
EvBGatxvILAupauku1ZhiPN6twcTroxbzg4k8P/FxwZ6mtkWvu4lsr5Dh7DO+AG/g/ygXz1QId+h
XAQXruKdUojrwSlREhmYYRJt5BvQVjVShbcfP/6WI4qk+jUTbFBa/akcem9sPIRE3II7bcwEBCsM
paphWx+dLD7liCqghzkvDY4o2TFYCsNXf4npVvT0QehYXQIqXE3quKUV9FuiEoJxFwF65id7lLSc
6KZVrCqdj3DVxso23kxrIQAZNFAck4PW3enmHVYuN1V3hAEZcxznmMRhgR+czBEOYEIcMHYHasJL
yfkW3+Maed/YZ6pkZLPV5gy5hjv6z66MXPh+YvV61c0SaqMgv+dv1jt7Wpogs16RLVq7hKTwY7TN
ev5eJQC/FSG3AHtXCtlwJMqyjmGgLhCdcQWR4gqcmePMkpCZNmeljNwP5Hgdx73RF5GlaQpJzZLL
wxta+BculgVLDZbWieRWeVRmblD67NA77xYd72fGLpe0TDcLkFUAbr5OkxlLdn9s1bsizy0Umi7u
Td1xcIkzcNFNxmFew4zgjsUEeo09fPSTAHmgrGCF/rCkzogXvBOpTObyX+xyzot14C4p+popB/Ku
XUwSAYJGZQDcc78ftp+m2/+Cq/poUTLAsPjRBdGqHq/GEKgUlliF/Nb0VaAEyITz+IAqJbYlyMJo
/HmXKRSZou82Hhb0OTPigBJ21VU0HkEpDG6NRkFuJrJzbTlrzRGMXPtZBEnbKf7uaFslqjmvFgq6
GcRDxEovsTjcOut6L9yI00e4ayXlER72JwkSizPyRtEIeY4HW7xbAZvWawdUag2XxzrZiRkDMNlf
8Boe/G+Y5FsGIsL6p3LxF53xBoL0mg/Fiikb+n/hDTQyOrpbtS5gI+I1B0wAC6XMjklFzOBYMgU3
91ravxergF7zk+XNyd7I/cC6luduiFfoYXkQnhej0mEHE9CD+jUB7vNXu5CAatF0+C8cdhUXc+12
/EIR41qvoR9Dpiw+RB2y0KeYjy8G9e54Kg8RbYRiw2T5vuVh5WHynJBEAv6C87JntPnMCdDwaY9b
cvYBKc7fsvwdSG/o1eTIK6mGUUpLK/peILtD6MX6FltL9FlDEYmPXycUmKGpmPXO3+ULieft5oFd
h2xPbqtzlijQeL1wTV69QxxzVFAqLTqM3JOBeIacSC7hWUK2rOPT8GJN2uR9cRAymJ51iuKAfudN
ouktYeSaWWVv5kz/ijKrlMkuwyPJotFoRP2ZH7YqkyJd1ffINP97TXl5y2lIDw6jBzN6OL5upWWr
2OkzFts9Vajt7f+2UhJF/L5GWYaR1TQz1LlgqQNz+DrdmTyizeJpx3l92MBglxxbhfUmRoG2mcIT
C6chexIAbKAWyM/+iMUxQxCgGTnn62/ildCmfiuTkM7yQHYlFZA4qRfV6qPOl+zDljHjN+zbbI6C
o+XucDxp8MoZPNN94FGpUZnRH5YluzH/3mNpBPIWyXMxk9NvBQZjAkfTIXaSQzUZQSeYqUiRlnXJ
9/kTzGbNcSuYO3CRNe3EftqRe0FH5eA1tTYWv7tPKwZLk1/4eEMQkhfk2XCbSkBfm2zx/MS6JUpp
Tua7fdOPPfEIbJs+Pydgy1snmGHqHsLED0ZtlfQsBjjxi5xewgeEu3AjDrTKCp2Z6UrnT8846KKh
SdbdC13d7c/aMubvo2F3WL9goeebFNyT3QDFf0wQgka1wsVaiV7ooCj2XL5E8+gUMh0oJGlpHzH0
quA0L497iGGbdLzxpRYPyiD8/yFhPilyMjKZr7HFh95IvP5X7M8IiY4sR6wt3oTx7l9wWtqGGQ4p
7OSmQtOCgJhea6ELucJy7iCM1fZimTf72JB11AjdidLQcwmFh7vgLMtYO2pItuy3gREe/Yid1Et4
WWCRFi2EWINMxpGOri0IAnjfxD7a8saWXYqZR7czGc9IKCj2uvDw7DjDR0mTHfwdPl+gRt5P0S5k
LHyjPZ5nAjwDyx4GYht1q3vspG7fvLeyYglNzpytLrN+KhNB1ukajGOKzHibaIu3kLOV+8Bj9OQ/
yfmwODSau5S6LFKZMCnWbBTs3TU+fsNjDUmkbgMtyAFdKgdnuUF8SKcX4J2UMKO6EEe8hT4sHXIQ
aK5yMm1555NFW/wY00SM61a3sfVXgSrz6LElGjfPdPS+PUo4v+OSRnLf/7gjd1m5TCam4RxZRKQ+
DyUFyOq02I+Lynhj6iKD4jqTO35fCY1a57trFPzHl80tO1cXunzzs97f2f4xXdjKbDWmW9VzyW4U
/j3MSDBorn9wFdXchtH1Y13dVZOiMkkalMmSxXs/oJI1xputNv5KMXL0mtug6ORtFNqoL4Fxb/vo
3N+SUzZPG9GhPQ2WImOXuVOzlKJmViLM8v9YHxRHHvGX5X22Nfp41ynQ1ZskQF5WHhsbj9g1nK47
MQhXM0Br38oyGixCtCab8vVUngl8Ufukg9Tc2lrYSr2zkP2ZhAh9QrtLH+QZxQWy2mKyXps+q8xM
jpX/Y0L0SCuKpLwDKYbEKXU7wvtt5RZ2gZRZpVKM08chh4dqqStu/IAAawcvVpljWIFcD6kSYSyr
SH/9dPpygw3+0RRCIR6sC12ZfGgHpx/wJ3C06c3RdiAKyYyT+szlhVDaf5JOISZ2Jdzg08GHROYE
zJc+dOjayq2bfrVInfE954CTP3PX4bWoAq3Kby4bedPKPEtbsp1KwW9zPZo0fYFU9ZNHZQLJpnig
XnJ0xWdjs6rd8STcq3sgHjylEChb/QNWmiP9DtikMAQL/a9IYuzmXEgXhVXkYvtCtGmSD/3s+ZBj
N4GwukcyVGiL+tmrEpaxdpX3PdsnJ0sVuXXCylslKobeM6GlEPfY7ujnDPSqtBTxJxmnSANgm+FG
ywfTyg8Miqlbf2MPe7yNBak5lZN/XQXx3LYzpEIE1wbVnA0OourXtR+2mT3km8UkJpGw4hVwthFI
mxlkpUkuikoTp/GOg/dGsPBGbOXTDHkm0+006V0n3rVMkmDSvSTZBqBEJ00KhspU+RVujwh7mI0R
lBm7af4ymXo/9+CBIxvubP7XezLYjZxSkgsq1UZtNsuoHWFnIU9O30CErpXrenSJiuhp8Fwjibzd
Yay9W4JUuLf9yJ77+xFtakpBVJNPlpEXFNKFcqaQsrza0AKJ8bVXM83yJYrvgQT70z6VBvir+uIU
AoFZkCnrUK2TZs+tElTl7Vmzosp/GKufBXyOLremJz16I3XoHDB2Fj2T1XCyczUSO+u4OF5M7GCS
0ppinHYuKLdhlHktrg0VwaAMftNEIhJr/BBKelnL1LthTg/pBhXJYbxYSdVktxASAdLnVYD30H7b
FW459Co7chHMBIcznb3JGieUVvrzzaF1swaKHG/UNf9c5Zu/hPBvndqHtv+RdpNaG2py4Y64rmaQ
xAY2e6WCuvEuT4xAaBXGb96cU2KpVKcISi6G5LgEZgJsbc8/tyHkPZXa/rvUMDxTXIsp7wLq+PBy
e7GwfXbDr1NYMR3kFlEGhBlnuXkFaNFSPw8U1Em0ItnyX9zq7DWam4pOz6hg5hx9CdsbkBxqsdZQ
AgnIrCaHoXsp1KsC5lTaTayv5R+sO3tx0MWxat8RTz6xaTPYXg6aqugGzmFUjdN4CMLfVcz2/ff8
Le2F5sWlxKGPOYasVpw6hzaJCBIY3nt0/+HRtN2faP98xU7hf5twJJIPw1auPWYbyHz997qVb1u6
aQohEdQQgQ5Any42n5SZuB3MejzcdYrwy6OgG3ZD9vg1BqOo97hgCH9OxCB+GFqTkkhqxjhHC9DV
fQFLxSiHxxGR86eWNG5gALcYSa0HhOgHXNn2e1+WbJFAZQh86u2Spcw2qSgMyBo9taB5PabAYH6h
ktldI86MgseFR6WDnYqIkIAz0KdzsKxnhmdIhoSvKvc27CvPN1Efx7t2u2Gz5TgWL2nmSyyNFf72
fGatl6rMPJ3bF95t7woEzPz4M1bvkJSPP5Ez2fvHmbAqVSbqzh4hEFE0GNihx8SDDRoXilr3MILb
aYCdF4VbZaID1zbpsgfg8JJA//Mih7tDBq8Wfcggc3hMlD2xroOzCNZ3wrWxKx/U3giqtYncF+Kr
BfNJLfBv/RS93AczWrzTB44QgetV6BcbcOqTbgpLHTCPJUaUdUxuHhKbpIVlYi0p4W3wTFnfUYOc
JzDSxik8WTwZeVkoBZIfiunE7280CaTq+EQkptvkTYyHVNw3H/AD4jZum4uVbVdqkzaAwQSQ2Ba8
PHIfqvnNvoFAUNTkl+wbfiibHCOaKahyRQs0i89PJygm4SNS+zNDyyaFlLQdGFYa2+kOy3UPyxaz
19QodRRGy7zRvYkgT6HvfRCnnA/rfqMvR3WGxwygy/D9ZPyrKcCAu2eY5/pgEj5s32YVP9tGJjQo
ME9t8IhxhkC2yF85zr+oim7Bk0pMU9+j/M/VGi6uo031QqbcwlyUl6nw6G6+ATpYvgBq/gyXJ1kl
UxAuVFh1fGdHMRvVvuHk7Ut/UBYvGGopATAE2hE59vS8nmBiF0ECU2bvBzM4QWFuPpeDkH0eDbrw
mHQenExRACutfDDUk3YaYI0AJ/Xrt866typ5IlmFDyX0xgI2psIXuqNn51nSQwplw8DS8F/ozcbh
F+HajV/pO73cDYEgHgb0p5PkQGGbPSQhOZf0AsfzmUlHiBn3K83QgqvwWs2afLj4NcGGBZjZgfzA
+pFK1SshpLHz47X3p9p3aiMxO58qpVUkPOY5BmXCDjKENri3h+gLH/rDqWzIG3vCtkz7/6sbl4zk
GmtlWwqkdtSrcGmUidiKl2yy5NDnN4CMSQ4SCYsDdP+ChzavrH/+fs2q3AqGRdQh9HKQAKrC3Txd
icyjBRtxy7aQXajL9ni2l5O8HmgJ6w42RrSs97XSCjGRF+nG41NRyYU8ZV9ZHDb7znBa/4BDyTn5
fY67vVnUnl2lMPSti6mjDHBU8s1gGBc0CuBSznyvwEp+BoInMpp1i5su8cHUezHLyktlkQ5wvP0t
D61houxjfWG/0sHqnKxYQ8sfoiMoVy4N13jSSoRq9/lnPDeG3KnlGhdzY4+UeiwTnIzAI51ug62v
EQFoxtRTl/6jtPk88Yiz8Ut84xPp9nuJQfjUr0OnkiPQH3iMjYHH/il52qBeLD3Zlg2bswZjlyfw
LnmQquaNBvRX9gtOHo82SDOqpiSxJYtDS4ZdusLyZe+WQzNH6mjPEvkGd/HZ6EKd4I+L5NIiLO/k
P+r1WhYt3l6ghcGhALcnYL8rJ50gkxT2z9nib1lItdVupuRLq1DcCNXXjllo98gLhuNSgq88PdPl
g8XtnB0w3x1hzdvgol+9h0sT/0r6LICC9DEQuulPq7FSm8R+7MpZ9bUUtyrAogViN/ZmfYqn7tE/
EZV9oRpYcFvf2EAoortX8Eu23HW+vGNQmwithfBEO3GwC+ouK0IFOH/N6jF8xK24iiP/INowb208
ur+g+ycBHBjcsdCLaNWo2aX+HqbQaGvioMQguFAbmRYnk/vbwiPMfkAv5kOfOG7C7plZIHmuhDxi
42cXQv2AH31C5W048X9GQfBM9c3rIogV4ArFhJN7A3iF7EF1W07RW8RRkMfdph/CszkXlRpzL/AL
0KZlUPPv4UIJUhbSwSrPE7chgFd1Jdq2qTPD2LK7Q1RgFeBQTGBYAj4mqmVJ6MOzqhxwx3/wc5Zd
Ju2FbYspqhHMdJiPphwAAwlKDKH0QEmU6GROO14qETD6PrywcjCg59YDueAzm7jcBGCPQHHXqON7
wxHceoDESs7eHmDQ7iCQ+MI8spk/k/3VQqw54M2EZBcAloPikM6FH70j0gQUHj5rA48pk5CRZk5m
HafQi4516J1LXm9piH2iVsFSz8ucG3KvDwLoQd7i31qcnGZaFHE8SpcON+mTfJS3kghxkEeu58Bx
5rllRwi55r1e8ucuW6+ka6nMq8GrSegkqQOofOqrWpXXdqsVEroE/AEhZe89wpfwrZdioJYpzeqY
NAcI2oG/k1J/Dt4xE7EaqzLIM34oBVQEd2VtOBQ1MrJw0Jhi+wjqIzzN+V+ykknl8Ni84JFIxFl5
B2i1AknBh7IGwDr91heZAwucUr25EC9PB9a3yY3bPQmQoeRv0rpe764RD+UZ2sWI1JddQ4lK0yiz
nGK20M7FVPEzzSzGQNVXA3zFWFnjpiQch9rGIpF2fcaEq3ntlWzmaZ0O3nbzKPclzbMk2KcbexpK
0+72g4kFqRzdjc0oeXzmDQm4ou6bXuYR9nUl1hDbtU1enLZ+zMGifDBDx4v/k2R/uEm7Azp6ti2g
73WfqK1+sdJHZvG4ZEOjHObZzPg29ymGW5jSmP3ns7mEkP9TstS+jlC74qJD+ga9yvHcSpVCWwLy
K/4dEM3apBoO/AnzhDNqnxT8DHC38AED26ZR/yyuJakEyFQkorFPUWO38jNe1Kfp6UNmrjuKIsvA
YsJJnedqFum4d63mv64jNUWppeA0tRn/ywtX9LaZT5rYhcQCQ3yLXwxX/KLmLAfcPVhoN//Tw7Vl
GsXN2yyMJLHwVr0DS14qIAhB1Mduzk7kDprUS/yXp7xNSIUTyApcwQPZdy4uqq7l44i/pfBW9T5c
+rV4Gda4UJfHbO4ZhotIqZTWvQyQeip4lHEulxxesCS2O0aya/YdJ0cpzQxZtw/Ae9aBY27oRp8d
11Wl6UR9RDaoRLcO5uqXivMCE7hfRwBPsOaW3JAX8mtoC67yn1ZD6N5MpyJkMr1hr1vy4KN5nesd
1SJNjwSumP7sLTksXSDzTJ6+e2qFASUj2KsmkPOSXnphuGnWOphTBRMdIva3v3VuwhkQfG0he/dN
VIXVtm+F0mujamh3Ac7d388Dm64kN9/mBfNfoALkkc6kdoAX6nm/C965lL8l3j0T5y4IpllEU5kQ
IqJHFUfjNHeCFN2NhrEik/CPnLbXG91f4DJgIbV5rWORlwVbhCcnw4AqXWidBtos9U4cxF26BKb1
7O0JItPxixpi+PMtyPtWtExUJYSDlnekMsskl4z04J1A6TEVBTxRhJnzqEKCf+ZT/RfiCymvatb2
rsVpiUUpb5BXeC7u0JRjtASw6i9NjDb9oIJZczjFtDJCS7An2aEbsK5dQoCuix/F9vM2hILY+FP0
SUaPnrQLjR6Sw/c088bp7x/cFjcQQDqc6GyIucF0CnmwfgFUNIPYrtmIyWjQ8HMemRBt0hdLqIgE
vvqbBncvj+9gEX6gL9HIZtfNhlIxCcFtCr+4XrP7HBjkX48XJKEnED0b3pgXtqfizU7TiREN2JUv
BC9dyhXgEMfPEENzF/Jp53qJDLofRRmfPFZFOYEGwvdb28XH4AEmYskq/RLfMih4OUzYirCjEWg+
Xwz1o2Im0zr70T0kr7WkQUl0PIImlvAqOjTJ/6+J/UwGbUEsQNARzpN9U2sUKDEx/Qncp/vFVkZZ
YwMqFoBc5+OXOfaVgh1suWiYE/oiI4+jJnwGppMSW+EzBWEVMh1tHd3LTCqZY0N1x8g+hbFhyGA/
AUUMP5K9UqFThxOn2oXtRH+mtPY9GOeyTHa6VxlhvR4IYjTF8p66Lhl0fBRbJ3xvD3FLVklzuI0g
wk2JKiKR+k3/HtTxhQ0QnVrg8qlmf47qCIomlwisyX5rRSvT26iRnvUECjwWK5UZhoMdMG9UQO3+
2KTsGwbjnwgoObxTWldCLmuF9H6xQCjF3qQzgWJMYqLto+UTqTyropx9fwBC7bPQOv9n1O3L86w3
wEvP1M26bmIF17RymTOnqWnvta94bU8F3C5Gf/HxxgoFJR/ccvJiyMIiwltVx6o/dKo7comz8tKo
DnoIBHhZuwjHB7ZE185GwpcAjYmKp5/6RDcOZyFJGvOn8MaDzT+kGnA8hspMTIoYvXRkUyLyCbzG
E3vYnyFdcWj0ANN5dwS7iWC5BOV4yK2mS0h7ux24DG8T+OJAAWY09yxZIew6Sn2ShoszRCvxhXj7
pGvTs5PuD+sUUlPMOLaNAx3nsuzX58g6sI/L5/65vu41Rmu/RGghmFAkGoJJtM643sz6EgiAFjMw
z66volFilzmzQlpWjUl6LAEkN+hDm/fEhLKaD76lUUZAJQFrM3lnEs+Dw8SoSUHrsGS/AwU99jH+
BQq6ZziOJNroa2NIBmsTErdOSb16RjjyrhYeN+xBIvX0es+YYNHrokGKNF6Yq53dNrBlHT17zPUt
0Ui8mCeG84ROg8s4GKxE2p8YeV0iaPmtbGtD4UA4xX+OFLYHjY6or2Du/g2yyETrPw7a5sSW5APX
wYPidQq/XUbm8utSqiqdlcUhyRbdRCghzQ4elFWoNX5xhtj/e4BBZtW99agd9Amh3sltXDMnmV/u
Jw6tjba21/fzRv/0V3/HTut9qBDIhhOcuoL1/XiSvGok02+2MCPvrUOikpJj38mWBPHjz4Hjo8BG
0QrLNxM+RLLmsfaIKKc7MKvffWYqTEZWSFVbkN03TIq1kK9NFXHBUkk6YU2lQ0CuXyBktjsa6R4U
92g+3QIx3P0S7HBlhSRzd/DhlGcNsQYWHfvuzD6Slput/gKmL5v12LwLHlrrpHzoIsuTj0UhsabE
5dFWekoRrPBaoimfbtrCVT1dsXEYW6ffUiaGtS/BJCCUsFAaBNKj2vRDiqBQMaMfibMh9d511JLr
UaWxda1ZDiRBrnE5qJFV53Q3xXbYDzVYeGpzgmNUTLPPv9pr75XKSai5T5txiFHA/KhC/aOtt1oV
nXL/SETkFbWieaAq7G9rX6BRPjz3NtRSQFik2ZazkOGbLP24nLLgSuf0xTLbSy3ubIJHk85yHyfP
wLNL3980EbUx2OM/XXESg/MDrE6dGoYMivucHhDp1xxT+5L/pHBz/t1bKNNKagdlPAR9do7CxUq+
KUT6OQ4B8uCqbo2JZZWkSh0PQIOc6A28DIJ1FDWnWdNS0qClH481H+zaPD3yNJwRtLXeuCpJ80RZ
CR+dFNVIZiKJftjVUrHBaFfLo5lpswjB4JhQ4YmvCwd/Zi3zAy/KkxD+KHfF8NK64mANrJcaaoWY
L1k6BsxSCn/JnTl6QU/PRZY2MSRC0Kzsctq0MoQCwe5IN9ANSkL9+NqgbOSiIHKcR69xFo7MAh7F
wezRZPbVm34mzj+Cpfgit+Fx5tnwlWZVdz5Lf9wmbNCzbo+hdu0M5HOQna1OOuIn+LYd606PvxxG
nys6jhQ3XW1ygHU27/xme+OHIRhKVpxokDbI6hl0qgrkNGYg2NntLRgp2AkFj2kymMTVQlJb4Hc5
/PAXHSGAnf0T4oM17qUnYMJAuwi+uVHn0UprEuA63ToMLBdktZt/L/o3eIOGMoesMvvzIb3g3jC1
oPoAcrUHaIoBabWKsrCjg36d5JKMUjQtgCVMUFSGkE8DYmZa8QI6O+c1WteITTygJ0v1tAWJhlrS
MiUlHyyT5/e7LzUr0RabtmrGuwjdOjXjWtOdXT/XU3T1S/vD/h7ZQY8iXfnsnKk0wbo+wL04uiBQ
OJlwN8rEmeFe2PsEGCton72sJ259vLKQt5lFVVeFd4pG6eSjF83Hv1avYTncEG67o2hKrB5Cmc86
Kaw/M8Qy7nl4n/KpG82TME1obfWyIYX81dV0m5s9k0CmsPSvFtiiQmdVoqZDrjXuSw0E0lV0roVD
wPB0w8YxsSpftS/+akALN/23RKCmof4O5uIqRdF+atZlCkpTQ19NuUvRlbCaWXzeBwiWqZ439KFY
QC+WZwitvRM693N6NwQfWQpEhF1MhEaSEtnxk4iEsvyFcgMh5evBl2N01vDrBRUvaSMbajWlmGjG
LqN4IfQDuzi/akkzmsZ6H7bb3zaQGc92Ky2mGDnzaKb2plznpdt6X6EJh4wIadB/M1hWxUtkggs9
HrFiJu5x/0UrKtzPVsNn+yHd8XewGMAlfqKZnN3hx/lQdNbw6LOa9C94Oqfln0rXgUX0BbYPhKCv
XPB+A/hh7gOvGCAB6yniln6sOqRkNebI5ey5VbNWemigA/YGNjXZcAmsbWjPwYl91YfiQgFq0yZP
mESrusJFI9GHNjyZtmrJBGa4w8hA1r2t102jNK4cCLBdn4y36t1QMXYqcYtpULJwEUzGoyE2iANd
h4AiSfyUx2yjb/xb751nojVUzC5qI9n7iSy2W9Navn8J2cqLzXRaCmHF6t0Kyhc3wgHCJiPUE86E
fgJCBrMhgYHlW91EHjU+PpHWYtPzkGCmjESglM/bcNQUmNHObT5qvpavWRAtOjYJBe5ObBQrRejv
8t7q9PNcmzND4ZbF9rL8hyMx6CPVK/fuP9U6h6oMrR6GLMS99ArmdX25tMrdTdLj7Z/+OFJCI0kN
F5fFEfbMZvgaIZVVzePVlCuDZ0fDx9/74ZS7I/qp9XFm/oq7ZlvQtzJTaWbaCeSx4ffvS+vz1SO/
fJyI/FcSAnqJRMOVV6QZJRTyzRl24zdcwu3JvQsG0TflAfeHfr8eo+PKd5T9yBxtpRQYFLKPToA8
K1XpVVbqnsVEhc3ErwQHLgiVGiv+CA/ikq9Go8Mhx8Y4DaHQj01OeBoh+V4pht1GBlCx1yfe0q/d
QEFMnFLozd1gw5CvJdHna1amBWpSopVOcFSwVEbAyhV18t5W88gTwjh6okAPBX15Op3LqXnn59hp
1hofsisDi2MOYWkajSyajgvLignPmJm0+VdDafHgWYT/hB/7Luyq2JAzz5c9ZcNI863FKq5VHlv4
+QtZLxCZxHG7SeUoDOdDQ9Eu0iodKEfs68TkNVp/wL78yhPS0677QCfGaivxCXYTH1xswp3HqKKe
uSiuQRgyJXni1DQ4vYPFTwOvpz20YkxfpQgsI79t5/FqPCOdXTJ1TeTi+oLNcAAKjj58DhjDIgUw
4n2+qD4tk51fwoYbYMW/u21cJiSHc/RIA70BKGy7hu5vvmP5oB5zj4PAuyNps3sX9N5/9kek+gkU
eLt1Iqd4PNKbqY4ft4x/ylmh2iHhbBkAdWd0Nh0zWb4JXjVt9SVrWgQHDz6tulhtRnpDLHanpEnU
mXG8fbdjvTKXesXA8+aFSporlFkCHyDVPNY+4yUIv16Vg725txW8P61ixma/O7NCcb3dBQhzt8ME
d1IGoFXGG8xFU3Wa+XLf+GaDbv6QAMWH2Cu8ADSNTHX2k7oBcJu6qUr3zEjJMma+3l5+6G0BfK+c
IzNWT8mD9VatuejXwQv6d/VARlKZ1AU9YcOXCqSke+G0ycf1Pd1VTDpo/+Xxz7IUtmWXMMRyZjXC
agaUBiideUD8owZWsLwXKWlpIm4AcU5XpmEAZq9fK1scYH57ggu/CAsR9UPafILJTIPOE7t8m86W
KsPUiPr9O8c+GJcgjsPCQEi982lcVO2Y3JX+abSRq2Nx9v6w9WkGPfGeRYKJsMLlgpmgl5qeGadd
V8wbRJ1JD/C+cDXK4m5Q4/p6BeA3oaES07VkrPUrHJZgP6ybemrxvFNJGI/VqoBEO23tEJ2cXDSf
znJ+swYULk2EvQOqUOpS8lgEC+OIHnDRyortdhDlm9DueV7GflYyVkM/SLo20RzYYQ7e9w13PE2+
bWYNmwtA2w3qKUdWT7FQ+VvDTgzT+m6jpoq7B617JtFjg7PHnW8C8OqUDhcN49ag5KJ3K3iLTeVi
1kq9336vOmmGL7dX88JuzcdTGPOUM/uDdlfvj3U8byztkP8jx5IhlzYRO2XOoruASmsgnQDagp31
jMW45K7ieR/zsLuxyv1+lBkQ+a8uNbarhM2GhazzCC4oJjbgaA5tojEM61iZZky08XshcAbxg/Dv
5bShm83VPsB8z0acvXi9ypZdAEsfK+YUwXlZojZ65wzCZcPwWdneH4Va6qXIfLedgfp/NvdjTYqx
wGdDuuNc5oMIFmnFHP2ZvfUk2fVuqMDutZdIaw3ZG6Ljf1zDx+O0uuTzKg90SRIE62QkA1uvP4y5
h91VE1ZBycbriI2l2CvcIEZKASkcgL8eyVj6I6hq5/mNcB2Jaa61t5bcDE+O5lVmdCnJxSD1HMdh
Y54qGnsVkYvv3GQ+eFomRHkG+7N+yu+HbvkK6QGihNFsAG5GzPc4K2YRLyrFG4VcXz+FZJsvktV6
50yY/vv4jhoiOzZ08tCDEk6+7Pc1v95N16y3oN7H13J8uduEtYq6iWVBsDNAPPRXvMyGCh97vYPf
Fed4tf2tMz2x204sdIY3AaA2ZmEpggoAuMKLq3ZudC929GcEsNL4njPtuU7IkuZy3gsj8C8TmMHg
zhbcfxXKuZZgpObHoPoRaAsLJRBCUarpMBqXvonOiPDqrM9qvXnik0bNjr3cCojTA8N2J5vgkTSp
Af6gfBM/W/vqQFH8IIKHWfk6oZEQuGigrZqPPPKPuHrhAIQwCvfMF0DCfYgAainKmQbUe2CEtBUX
AbFjS2lL/HAjCpiOiT82+NQjdaWXmdLUMtZ0X5UrfC7IP+rTLgCQiKuKphxoW3eVbKsv4GRYsBi/
UGmxsCcsPm50zZ/Ht7kDDQGhC+Qv6k7s5c5bT32astHot0tPUWTBvx6BeyHUKzMZi2q0NSC5bIDF
1AO/BL9RbuqVeStWPkxzEGim3p+t9ukVyouZK/i57JIkUbi0QDL0LNmCuVINFLrRYOwQpUHCN8NV
mqm8KInd5yld6U50rfkwbMO1mJJy+5kU9eGhQ+RKd4/HTwJrTrS4YCgxX22N09ufdYk/mK4/VBtA
z34fHd92UOhy8iK/mIuVl+hu90YN4r7yiI+XIWEsuPpWm6zI4KNICmWRua2qQisKsRbDei3hcQ2e
VC8kMqChAFiLSHMdtcMHQgzCtdqiRUsrVOuY896BapGRbQNwE8QBILN2s28Sict51MWzQXUEW1zF
2ecFMDl5H1bt9jBJ6tyAOZWGVQpEm/duDSGsT/f/NxwwK1n1/Hh+C6pqzNFmmpeQzaTUnezXIFXW
/WIhPG1AgAUPO+pkcJoxN0skFpfulvmHIMHbSuWQ0Y9IxNspQsvDMwQbFVtxjFmpahDooMD2qegg
g6L7kugeZFv+HdEMy5kFfr8b+2413IAu7lDEXZtL7Ngk4pnKo/7/DxWWRx3Mf9mlAhdmQfUougCP
M45wOp0KDealA2iwyeZcGP08IfjHHC98FcuMY2mw5t1qiDgdUXv6Ork2se/Bc7blTAy4SjO3t+Q2
/XOGJ/QPry+KmYNv/8CjDHQXeQ1E0r/MudD/UoolVUi5fx8jcqCAAtk+JoiXoK70UGpG9jlrfwX5
O+wU4clM8PP6pO5iCDHlq2BVwLL2+bTtkeGhJbBP9d0ZUaIrKshB+1zMqLQK7BgeSEXBffy52sUp
AZ8W1CPzrkzxclAaVfJhLDHzKhhxMRbXtJK+kd/e/7lebjsypCKkLKSX1Qtagy8gufJaJ+LIMj2v
WyfcvyIohQ/kO2CqbtG1PlGCnARDZmvECQqR6i9Ga4lIttbZ2uzRw1DPrSWTpXUZ8WTRQjMpES9v
amUUzK06zdTEZnMgCiK+jhY6AQWeFo8FkRyFHK8LxTVRuUwa7gMZuon4UeAv/p6I868BM9omzTgy
CsOR0GsdGxFF3rc+35K7MYh3utcI23OFeLuOK6ICBpI3imBb6jYElxkt9SCsBU5qKbxfRvrUACqu
OREttbE4eg/LnXVoeIg3hH5rC1ZxV6aAPYT1+EWhkHPFrXgNWCjzV2g0zx9L3WQL1i8fiSKwnO0F
CJneSgYSZGefx8BpXlacNrcV9w72n44lwjudgp7/KVgH8+nY+/s3T5hKiXlJHUfvFHKEqifWVpF/
Sfjs4HZrPsTmKcF2s/JdyoGe2/LX4dUiv5PHvhiYTpmkhFBXq3ydLR1V+hQtaA73ickofi3lQONM
wqbzMGtqDxEBKk1o+q0Ax+lHvU/PxRpnjqubrp2HVDsFE4BMzQQPQOHf3pz9DZ1gQdrVMREfuECL
dN0OJY41zZ9PucGY7z4eOUA5VAZQvJH0QJ3XIDUYNSIBy5QHKhdqvj41SNLuzvS2rfNDoPecDjoh
900BsWIdWahOGrp6izFuiaSEly81wd0P9m3RAcYS5208XrHhNQaDE4MEQ8bgtplHi/r04HNUf+7+
4ki6mp6djs6G1Sih0dkLI/FJOnrkGtMnj2Ix2onN5hQ2/l9UsD2q+7zvEs/RUnXP/v7N26EhWEPQ
EWO33q05grj0mkoyucGdFBEhDXeLMG4UIcdAM/RGvevN55NLFX3Xu1a3FY2tEJ2GcGcGXDQMEAE/
sBrN98Jyr/gI2SX0VA99BCeQKk2HKFY8aPTqcG5ZmxfLcrk5k/ysXgCKVcGJ5gYlBlHLRjle0QvO
AJ//jF0gE0O7eP/dY/CaHnd9URu44qOVa1xng4oqIAdbjpIe1SQYAxTvRphlwY9WmVDqggjXDVN1
X9+Q1qiQZbFdMB2lX/TfLS1j5J7qD8nCwC6HzDdhK+AMYIarLIoCuBmGI/GC1UUg30OqXp3UbWnz
bwj3YliT0fHac3XS1MYzgULmKoVHn6/Jm8i9MG+4PafRGYCnCpW2tjj8isg2BHdkpLkuCXl/RKU4
+KnnyIdnGMK49+RIb5FU5uYAMPIZxFKE6bXHa3N3ZpiHNCQIYkt32mauVsdf0Cyi+A6d/mv0eTp7
bqXGKl52VXrn3LQ286oKiODvBC4dMUQbeJJKOz51omi0L1cQEzOfXeGi9nIcFeQxcX1fqq0SsB8C
Oh39oC9tNIHiQbhhu/VWDMFpw/FQQu4o6+V9N8FDvbstk7l6Q4lIEAoxTnUq5SjfRWElTdSzob9I
KpqsBrVeY44aPbM+WcozaTQwj9LPmsuVocF+UMS1d4l1FbzOYV459VodXbrP+njWaKP0cQNO6xlo
IxdOYznOsTz9UIxn22tbL5MxtsVQnBTB0o+3s2u/OxyjY/KkH3VMdwnf1/yZxTIlXX6dzRSbRE6k
M51GMO+eZZWZr3UNPxsO6urKi+r6qBA3W0O7baeHddUKquVvxVhIKe1rojfxEEhnlQhnTBV09yvn
kydLCp8I3oJGwehXoTgBjzK5DfCHWV//uL3cfc4nmFlvsiPcUdJWEsG2vpUWVIbCFZpyOpvZVxUO
px8xCjGDn+IyeOXYxE65tCv73YxYtJRW0ifbxbVLgZU9N7wHQz5cORngRMqHjqa54xjkkPyHEIvr
tbtT/QcgsDZL+1FCcVNWxcNSP461df/AM7mcYXoZE5+EeXjtc4jfbT8JXVdq+tqc1EMNHHcXC7Da
Qk18f2v3QcXIgwsLknB6+4pT1eDOqaqtK+KZhyzxFw2yWFXUXwIsJV/iM8e0XZTMTcKzpMrtRLrM
ALS/R6Pz8BTCKLH8zkQ0J7gys+N77Pimw6W+YO8DviqUqQXzb1HRqOWv3MY6dU3fz1JWwlA3AbOW
LiLWPhQW/oJfE3CFR06SpPK/POtWck1m3FdSx2YCz1ecNTGlR72FuFBzHlhHb6IfQ4D7LZW+vYlf
KPUSZ9gBQdCbiCockdL5MU/MYjvBtvwWzMgjXHo5mKPiq01VhZ/ZyU1ySWIc3DdZHhoF4c+w6TVW
wYLPo/TgE1Vp2Yqq5C9BUGOEmecrj5WoZRTWjXNf+Ir7FLumeg+08dlNdApPpbugYV2x5LeBHZWj
5gx0eLb3Je2issnTdjg57u6xdHyIzBDfAUlYJn0goWoF/EDtXG1aYsbCX1t6osgVxA57X0TFpgGU
uIBNeqq+9VMy3FXVMHiAyxZeXzjfmJ+SboWeyALSCyJbkLELF5unSZz8tF6DbMnYe3N2QRfM/In4
Y2V9YDbYt2dGQmg1iuz23dzOudyC6wd63yeGDficOnyen4RIWPpVYmn4dyOLg/SpjSuh51M64Z7u
LFCOoPdMZye8FV/CqJGEKP9z3woiUKds+XBxzu8iCrp2kiJltJ++05b77RMoM+/KtrNTYfjDPD9x
8GNRbC7OQvbbQCPx6uikBmfEJCkYzVBhZ0L6wp3Dfg1o1/6B2cmGxxuoEVdQ+UiTZj0MJnKVQ2dv
YoWhcgMzBE5rDbXBXB4W1/Om4SGFq2dRJTxRC4X4XVJxsWqtK9ZGnDp7IVbmvqCvuEkAOxRn9PZZ
er7e2ydjGhYUt3ZipSaXRaMj3TQkN/FYWPvRWYU88BRN4itPtNt19vAuiyydoi3IfnT4+w1TaZz+
y7yylp0X/5EzZud+FCzrUZFPrbysTitWYNrJxG/xG2ggV9yEnuqCFZltz2DtmlHbYFYsh9KhEUCk
OuVwafvuRNEEQl+S3DsLnYoj03F/G2PqUWPmC3xo8EOELB8kzhG5cEYwTcVyMTigeLKJUFgxXEfx
bgOIBbrFf9JWbwdUGCgR7XkkqbiJVuklC5HhGU8e6fndSZL3xq/U7Kd+EOlGzkFWPIHRjc4AdqOo
mX03nzwq4VH10KY5tAJEc3WpHqEqGAS/PRQeWoYzHehCowth8siip2DRgu0kZDkiRt9RTt6UkcjJ
PqudzJ67Cc0TD2AKRztPb3J5cxAQYWp+9yaat+8aSeaWGAjLzO6GTttL4qXXDa8zwV+4e1MHVmBp
OZqQEGPliCKd48XT61R8rN/WidHVAcjb0mV7wNmpWG4YUdLU0xnePEuMSo8NcYXJMvPFTA7Ak1Eq
7wDxw5ziXQ/dCgS/JP8L2R/x65Wpdadj0NpLDwFtvIqTE8ax5H7bLPhDkFYS317QNYZ0Ail7EuBJ
4BINQC/C9HdDIxHIJLvileYAC5B4TzCUdRnLo8vQIwzyH/6yzG+NJNNfuze/gBcxCV/G+US/9vqA
GxhPWxdVU1d7NdAvp/zgyLWYWd2cwgTfYrF3fcGPfiTPV+FufaJshWDsgK8Dqba1ID9skubiHxOO
f6BOKwGW2eb6jTcSoluYq351SlSj19HR8zqEAGpufEvzVPY9FA8q+d/oh8XC8HhKIjZt7eF+bLSS
mUXASDVBhqlp9lSziJqZEHsjz/1FM3HBhtg8jAdTt6JhUDb9U9yhsJybfVZ9crnE+RxIE8WKVixI
qcRd3MyRHEJSPmQRMiMWJ2JI/zCNIBoCrCiWBPYCp3+fi/NG5vbJSsVXZBC+ma4QFCzbTZTlCz2x
+Zo4YG6FpJhjpceW07rHRKuIBAt6mGGtgUoCeMtYTZVpFCNWZN2nnMmMTzttSWwmRPDfCnqYLfxd
cQgZPc6yAqnEydT+RWqyGbJf4UhzQEvQwlyd6EXU0gFwT3ywEYwhmGNj8sk4NQzlDgUFGSb+Q/oM
QtDJuOFWl3DRfAyrRsu+jJWQgsdR6M0rPOAQmsMMcxlHcaUzHjOiCXARRgZVWhWTWHJ12ov8oBGS
39JJ2oE0IeIJ4E+QBiDPQSVCNg68EsJ37hyqocbSF26zH5S94w1sV+vzqu1DxQAZqJH9lM4m3Zdm
9KpNcHVas36XeY1Y3dR0uQWG9EGoJdNzQxpBgDaOpfUxeSdOu3kTtHYcz3RTrgfw+q5G/P7cg0qS
LZimPCNkAluYy0b9mlWoEVWx2j5ar7Btd9EzSeJez0f0dEvg60KMuppu2Io0OSRWeDfrClDepvWu
Q/ZIWhHsakoqEXUipQZZjRvngdqV+zKv3JuKJ6dKHLuOkC/OqRgA88Z1sUVeotPMy/TyKEeMTb1Y
ZtyVWsexkeo+wsp9LR+501tZwR+ZsimCTot36guZKXBj5eYuKpnEMVYyDJ/OPpRdcp1tKxHC4vr1
Hb+sc1Cvrj0VzZBBSARKhN5VVmo0+g1Z1RxCpRGWmryzfHc4DmZ/4FG2LFfsZDQKBZhIRbFkCUgg
eyQzSgqOnAsq1BawLX3SHcxkmX1+aWmuvJabGgfDW0HkxzAlaud5mj3XZU9+ehx9hnIYWE6xt1W6
wxfmwnJiB9PwST3zBOq8vTV2FaPWXRIKPENG/lNULpErjQXfcEEv2SqwdaXxHcNzGJdnWf/Bw6dc
Jmy4VdkHHyQLMkDHdrg1UfCIg8+mbabGxP/wZwiKcs+b4JUXdnVTm3uaJEMR1RTiegnzpTqn5Nqv
2aFBCeVkA6Njn9ePv6hFo8G8jb2sAIgcDkzTdp613CNp5otj6FfBkchPHcb0uyAi9oyq6hO5mO4g
Xkq744jOH+TZY1zD5trY/nxN2sxrqwtvfOorLm146oxMlTLI5dfHUc525zUV9436qi2zk6bfWAQi
VJl3OXl4o5IZPg6cm2zLl/NKIiqPXYWxQmvm6nuospA30/nPO18Kk9wEXzjmvsFrQGnpIw1dcvCt
nE3NwnG3dMNYjqPpMFzuq9FWTMAt0YMbOg0CoEtJyP7MsbZCoqVDoLBDBZjy+bkb7EVtCateuwS5
XRAwokvjn1cvt2oaRi0Aw/BcNQCi4fmnQkxS/uHRQ2Rv2q1wapjylRUXi2XiySRKpoYrrjkgFhxX
8lA9v6ttd732NKFpTa8ZrSb/wM3pZD2DVr4PluewqGsb4U2idZLriChAURVnC1f7i3NHmzkRncde
qy8N2gzeAqQS8hgKkWymNpDHn9HvrMj2juLjKCsY/S5hudDBGKy2I9Y+HGVtsZgL5rD9zIIJr43r
oFhgrd5hyoHE0C2yC6lDO9mDrSlGtsCBTuaEm6rBJguWeV/dAGSKNPiTFB/h+QTeR8yLIYhebsZw
cRRM3SVlTch+JHi3KW4XZO9B5D8vJu+oiv1PX2dRxkY2JifMMhe1Bjq1bnYdDtQFXohp7+Z/EBSk
jhcpGTTnY9+glSP10gW5kGFleuIECDqPLPOZz4Rg6CAEnpjwrraMSghjqwEJAwrLe2zUWiVF3z5e
izfikm3OrAz9OdWYSMhpMjxTN6UF2yCjmapmRJMWgPKtg5SJoAU5gWKFEpqwyytx/pmAghiaOwyO
etDPC0urRnDRgW8riNXc1LTCgl+U9MgVD4QBVRpAW9NUAhuujPzQgAreRZ5aoKDfN4/AvvTQcAqw
qWfg9MCoh3rPdx+UlkonUy8ZszXq6z/wAEvPL8w1hCuFrUsZ57NkDl6mIY9RBWPnafQ4W4wS7+KZ
lFNkcTlwRjGTedOUEpHbo7OKXTLJA1f+gc/i3IOaNsa7xXiFO9TSdW0JfV2w74ikSi7vCCTyjKXZ
nmW2U5RL47pWH1ttMz0Dqhfy8TOeNX8aoFPi5D8ZschSOnYGx06Qmssr7NCCI9l6Mgfib4/K3bpl
RgTfB/HVbg9cQi5ieg60n4uyS94ibE8Ys1aAS/BEz6Tt50xsRG/7tTvZyq+g7Sgf6ZRxkqKA0tis
8XOOTG/U7zJgD8T+dW+3tSn5wrBObD6sxVlT8YWHS+fZl0zIpZPotUJToSO0rK6imrnO2F74mknx
C3bjsgttFnbxQISh5OG89JyI6KNMbvHzR3Y3e4LTWKS0tB465K33ABamuV17GIYZMfed01g8FCsl
1b+kczEkDPezHdVeSbm/mJBj1WvqHGpCCFilf/LlzILW04RI7u1ECFIhe+vGx/Bd0IJHm5IdJO+A
+D/XW/8i8FEcZaRdaP+u8ysZQBQT19TbWknqiIc0toRhLxlMxePm2AfqBXGdfOM48gbFJhwstIo0
RB9Rl6dne8XZhmSnUCFih/eWGNgrj3SydirYbHE1BqCrnfSN8tX5PDcJlC4yLvPQT7e3gQZOFaJL
jhrki98MR8XuivvpOxfQ4+OwR2STUa3P8h3qvTYsXsItqH8AJ6n21fQtbbQ1BCJpHpeD41qIKbXd
cxDagxgOIRZLuvvAHr8T02PhzwyOsMWZeNJtq0D4szFXSjBVr4/Z0JBjXrND0ptWoZdJYenIpHvc
qxmCnD29Qa0iaJg2qr2KOEen4lEBcNxsJZXpYAxOT+oUjswE7ioPecmJ9feOIulTKENL4VvCZRPf
aSmguMeoz8bVqsAKLtIvUZu0Nrdcp6HcuzjEZYBjZDVdYrErblIi1KjkVFxL8z/wV6xNaKmcpqks
7Je4+uGoRT4YZRkt/bN5UHD8f29f2+7Bo91M1cdaaQJSBJz/d++EC26rUmBVUYxKwfZO/GqVOb5Z
ZUioDFtuUD3KAfOBbIm74njNXFD7IV404ZwhIh95iliDAvTSTLBClSfSHMpx5ih4kU/O5TRsZF+0
SXYJJwqLlCfMTyD6xt1DhZ7tHSXv2sDdEb3a5PHRQVi+YJX7pZwL7+0Au1kfbshB52jQOYnbYEco
VCi0yiSV3c/loJYOIrVfYM9G+9+l5hO+fx5URAvoG1xs7hrci0fymT5ommSqsqFm66DVGENnjLP3
IT1ohGnYzYBk5f/cYnNFRtHyohK+D8qtWIrSvnqfyx85nzTULU6ddsCUky2e9fQHfOXyR1PytTXY
9mNfIDHGsQh5cZEZjgtFwtuKCyVpfCBjfN5YBisVyvFo9Qfqs8U3vHrpWbXKa6Wvyki3pc92nVfA
cZPiM/1zhjlgiOLx+Qe4qHoS55RAGJFLdZKI7HPoHSMx7zOrOHesmaG4domY58jjMj8LOvf2Mxa5
TanpFnf9OH57cEWlN6d139f1bQ0UyKGZ6MkkBcWTAOBM4wwSCpgmGEQXL6Qe0vmaWvEBDZKDNlGS
17qDNXCHvFG0hnPq88W7goXUN5RMz4TsqR5I8jokWHIJpWdSxwbSs4sXohpjs3ox/8blPXid3fap
Fra6FIoAyQ11vfJ5IT9s1qDVLBW7qGb9XgWgPfPk9Ui32MibRLMc619dNmxKcNibwNTdovg1W5qN
gVDfn2YyLvVNM2jrWCKJnr3laTYGCxkY0kL8RfAWk70GAnHGfoUKmmgZWDDHMUXeZ8LOnSqylb+H
Pqf0ecui/G50DopzYKLsA5HHlRS8/fZAWbuCmwaOfyuvGMIv3jahnpEmTUDUgbIzpTQR8tXMvl5v
JspCIjULAmqxLQELu/syWMVvGC0wnCbgLoOT2RahXnxt2iN9Umfi6oR/uFJ7U9VX1xvaAMW/yM6E
yoI4n9kdmqIZvNL9yJ8Pmax4DFuT24Re3pWqAAfzhxwBCbP2KTSEL6BU2bMi2lo7ucZt69JR1SI7
IhnunVTD5sPDO1k0eT2T0s/M5qwqvi3IR052VSSm1kmHBWUVmCrkH4QBnKh+FuDXL88w5YBEZvOI
f9OK2UF0avqYI4nkDbhZnliCJ2UnziqJOjrqwXLnv5IYL62aXVCWawTy7QgIpprEnoWmnX4PToVk
miXlJLazgCjeFH9ZyBssrC6+3nPJzzZjLP2Hqd8okZA62Z1fxvgpKPBNRx1IDHtOIej71b/EjTrX
PmxSpB5gQbMk5EhHGmyXLiUfpg+scefXBPsh2FwQtUZWevy2mojZEbRlCU8Ub2N8K4RVbgsj9LYh
kie31iBi1BGiXkC0WgBovHhlDh2VX3J9QPW4rcjE7lZ7AQldtBsG82uM9p+ZN0XunDFtx6+nGKMB
2m1nUkO4Gtd+fRfVYg98YyRg0f8ikTB4rQVxNXohT7ACgK/3/i51LUWTvxITc6ygGSbtXahLdql3
FqXvDhLGJplOK0XM55gdMSlJdf/1CKggOugr7BBuV29sza39fZ+If6TYH+Ewb146tkyVFtSNpUV+
ZmfBldIimAyUMYDA64ZwmQJhzzM6wBSKsaAIET05X1ciSPmDyhewyoqJ6hvUoOb+dY464mxJFFg9
bKBZz66PfCv9zDZu59EJAe/FWd65O4DCmpqbNaOJFsPcMYhyRBmL690hFqaKeMTyCWNvVH8Lth61
MMhXxA6OEh2rpZvxYqLeWvMNKRsYXRmsaR/erDuBd3Ed8VFoweuFPTI1gIFtPF5Q2h3XtTTI0YEI
x8t7BxzrWO2pRzGL8t4cZKoDRCBxbF3gcFH+5uk46enhBYg4R3ZqYb4HUF9iLUI88y/f/8P0EmST
CNX5GbZvz828yLINNXMW576FVPD16N7kvPm+CvqB2PEfD09bfchLrNlYjiuYgdTCOexmhvsnCIuA
4jTx7+fEOTRM2aenLi7+x0k3SE6xuQ3e2Wd6ytBg7X1gycb1zt8pDHnE8DcEzZ1MG8EVXSveUJpD
Sxepf8ytnc9rKovVPq6dK+creRkT117Z6tkFhKfsyaZjdAlZhUe2rh3V/Usunba+lIJsrjs7Ie9z
FPqnv+iAthdMTNRS4YUaT7CMddDZIc8qSPIngBXfxTZJ2jqBK5x/pviarJ0/raf12pQrOMO/Y5S3
MYQ4rZlsR4B3NwPF4jGvFWhTXutDnCTAPUxG4Jc6wcA9v43QBMwrscyyW0i8VH+Vq90d6XMjNeSc
oxbp9t6TVzP1MyrzvEkEASAoA2pdJdqdGOuKdhdp01Nr/0ddt32nS5CCIgrE5v3zMT8rMADnd698
CR0eOen1nMYr2EJ7PrhUM3Y2WQkgagPXGIske+iJ/zKshlXIVjkUBnxj/znmKW5Xm+17ednfm704
ydAxWT3Togsa+jWMAPCCLgf/acSKred8jD080dlTB3HTcFEUqJbaW6atqklMjR5I40Z0CYkLBQYP
hgU6WMJ2Cupm3zOiyPPl4vYHGvpYC+TXVAu4+o2vD5hCjFzIHGwflzs6V2IvC7BEmzEUm9mokA91
ZiPA4sDGAqvIsW/z0VelrqAb7CIXHo2X2XtnNBgqtZqDCON2qZO7fwrnfetdQ9DrsBGkqO4WoDQG
UQ0qFXIJRyAoi+tuFyXbAbhMLE12Ovz7AvWYwWRBTgJcswqYACUhICXCOsZSCmkFfmWZwUq7g0Rl
y9eoZy2H/yHdlro/+RibSrPOqW/bZ3G1t153SpZccxpR847uC/WHjJZqHOuTP1N54Hv/kWSu2sod
aXLmNz6ahHn2BbO21gIQFgqivsoNvIW7rrrtMIbRoWUCTE9NASDNLn39ZZQ1yTxAQfumNK8VZ4oW
SV0HpV4QGUMc7LE/ZriY3dkGQrThMymfJAcBKs2dMOrchU9QAtvnYwC8FdQn7UoGGb5hStD92DRA
ur9fog97HpQDBklt8de/jNAMjfNZSP/PLCx7MvNaq2c99DdvZ+6uxRSkvtiwymc4i9KghzZHA4fI
UslatT6OHQTJxEiAo0VfgILF1h1w5F6V2elG3LrlF488RdEyaS86OAcvPdHCY4hPO/lZrz71c1d7
AyMKQUF/C1au/HKBDAbtGbxlhouM/9yTPEaOToI1CrKBvpdJdlU1siP9iiUe9DuV2qCRYj8t1Qfm
Ibv2n6dSF4q8+rvkv6SShOzyM5N6yD4twt4pC3dYLse5q8EEMS0mohxuXwh96uFLQgmTIb9JsRQg
QAYGCBfPM9NBTVqxFnal+dyLFW8VGRaPa+8XipPVvQV++YmPGz08ecIILJ9CM61kJeD4sa1MadgU
MNQKKm3BPMoTrHaOTgfd07h1mNO6l8FDwDcmk2X7yyJWwciAaQGi5XxR/xw26LwKLZco0sywJdPN
bpWXTO6xmsZxdE5LO8t5fZ1D48MCazQrPL1YyNKOCyv3JZnVyjrMenOhaiMO8BTtNwB4IyZqUfJe
Mwm7TDBfDyHaMpdFHENwNDfXWSbGinaSq+F8dtbhZXjNp38Ve77rbK4zeX0DihrH1VXYRvpVrY4e
dc3AoFLRPCLQOJZrwV3ZabVkMZzEexzjwBb/8h09r9zpbcbvN0TLYlml3Xva2j5dVUjjxq+HwhCp
ULVLjgPvzGsudrWZDw5xWhjnpFdJehUlgJSIujw1crjAZDAGUxHb7B7Q5i0qr0+/kIRvv5LyZLFp
VEzKs2epUlp+w5WFp9t+FecSye7rtw5jWc2eR2MfLEuzFWxDx0Msfm9xrr2NTx2U6mU2ERZNnLZt
7hxKei/JCpfJqr5wvfcnui+6SY7XuXGwSeydmNPiQHCRQ1RQAvoxUEERDFtRhjU411lzlwYWHWMa
WH6romqFTxaKlYciRfkwpuqnZu1JtU9t2qCaF95oRDUnZM+J63y27KsjWFOLy8HSS3len7l2B6D8
VwlGCABfBppYXgvF1pMWxGRqkjk2AvzjOsyCkcsAyLkfSV8Ju1O4VfJ4PmqhbCtbhLBp7LfnbsXb
eYcvd4hNwGVivpFN+8WxnHMieGSSu3VmGVqJnX06KrMAyjg0spDr5cuFAjHT4KtTOQ/ArjuF9/qd
fOWU8qXh74/mQmvH+WuQhdYPzVXEhMrrvrf3+j7UL+mlqcc17eeG/exUl7se3TeM3P47ZUaOACaU
zQxDtodCIFDGZzYrNZFrooFxsRechtD8cnzv2TiTaLXGamyRvXwqTykbTl9QEeODlftgnKnp1iaK
ae4gPKYfh+mKxEbcXtpqg7aII8PHvGZ8uTqtxa3j5+eBL466J577YtmoPSs5bG/rQycpRhl84HO9
2P3b53fsnJ4PPgyMIR3yD3cNrUDNnS2WYE6VILdtm5As1d6eFzNTlh/7Vbwt7gsp2EfP253ljznh
ywS2IqK+nXrHPKNcBjVsI2jNVQfmm6gnCRU3GRH3mEggfqLCOynW8gnFROOdHNr47eRj8+0LAqiC
JBAbj/NwcMV5Yky6kjXPCzi3x7wes53GerkCzscub0keZZBWiw/93mVybjKXIXL59HAsSMqekCxd
ab/6ng8fslLiCoQwMK6+Tip1c5wVs3L7k2ZVJTQ1PR8kTbd6zrtVlhsrfuulG47tkLvdca4jARW7
9Dm3lxlA9ndVVUQ9lbCP00qyvU8bxCjpYX9zxQWKd1WEp9s81Sg1xZOZrqk2V4TFTsZUT1vW+gXY
AATu/pWMYW0SI29SZ1mvIBR4r16TI1KEE+njtLN2cZJbBMnWZV949s0+BMqSpZ6R+q3nLu6cvPQW
QA7HAzAdJbqJNCov+NK0Fwq2XVBbwhD034mTcVZeP20LeNJtWgBmnDJCmU98wwnasQTAH9XM4xcU
3He9/8uJn6sJVjzMbY/BOC4d9EFitw36bXiO7LjWsIrP0pI5E8FB7kQrTHE7icSsq2MWcl1h4lIw
d3YLZ0zMUhc2pXU/jcE+QCgQ8d/SQEtzxHGWcN5jYMMeS8RI+QrE/ve4gdPagDDhSXdRUq2llBlz
2UcGrb4NWLp8sc9h2vDcX6EE/0pRXQ82hLsjIenfekGYOo+yWqj/xqv0s3GNMtyWQuW6SvunhKvU
zMygK15ZmzVnP+Ssb+/Q28EP/gAFWSuGZq0Y6R/n225TsSuKPAWxx+sBzmppBXCzrmpbnMyZqUaY
jhJWrk91yn/TGrJeRmFFsDHS/r46yGP7nkG3j0oIl7aFMFmGSTIrkkQyaCfGVncq9YzTWv99SmxW
gGg1R7VGQndKxLRy2maYuUoyPKh3Ix8nDTOEnAze6e+16FuSzM7ji6LtSmPqs0A8yRdqe/q3AW7T
N8VLJK1xQh7PJ8k+xf2NVw8oXJXbX/A/Z6tDViyFqMrC2VQ1xZ4dS9+aJl+K7pc2pnzIBdDRRlrw
RtvMlgKIVsrddR45sMo/zEIJ0P7ax5emd2eLP1h66w2dZtO0tAoO6RMOYCmCjDlBfNVOCM5UIfvB
ElpNgIBk11in0CIaGrgIxm4PRu9HVWT+ybS9Ua/NGkJldSeRK7vhPPulhSv+FUxjRrZYQ2ae7MSe
g3xGpsYoSJBWtwPh00i1/CF4JOZZtLICHKzwm0Vwr/tDyUj8Di3K0+oPwFDIIHEA8wns8ROHMExG
CT4gzbn2fjn44AaXa3um8u2Imp9hPakqT9lJS4ycCXD+zH6cAyhR8/fXIqSJh60wrG0C/lRyYlh3
XQynyA5hMqCpwo6h4tUTXIcKHQWoZB2zJZDVxRv/U8Zk/Bt3C4qDgt4wPtPNF4P54pJv4muUwury
OWXz+iOwtPWw501MSies9jsUQajNy5hTzVKjbP2OTjW1SLHiFvI7SsFdy2cFzh1rjswFLHAB0uNK
pPJ4AgVHHcslgzFdQv6zKyvrW2Ar8X1TUkaG2Z2Xz1wzIOVo6KMFzaWzeMKHpW47SVX+P3JdF4mD
ziNg5gG/hetH5F+8d2RLxA0t8/20EaIEIglhlmyq54iCw9XrACz05jsVOouorRJndynsG6v/GFcE
7bGK9aPnKjm4FJxvsJrYDRSmL38gYUTIJUSpXo1vHpEAeqABcKVtlmaIHHGdmciJXCCAdsd7I/mx
iaunsDsUGx4hDl595XmkPF43Q8XGgW6PQVXH4pWC0llvI9976BDud+Sbtssj0EXSK45SWfBgrY45
k3tVeQQ6nkyihpTr6fbGMXUyl1RpebAUS26YXhGnR+n9ysP9KApnFRCb0p3DFrhXglphVaYe4PI5
9WPf1mRehcDytJhfYwzyUtppg9Yt5fXoGteB7SLVVa4LE2lSaqEOwZpW/SjcNBew5d2HA6b36e1B
ytRR2ULDe2sUMu5CEQ/HUSqkz7yg0lJdx19zXk7prq39OIarikcOIPocyEFA5PeEOyhXc7MCe/VZ
gXdOIv1UCy9i8hmrjW0UttGWPYmD3dxSloDNHZz7WS3BZ/uX01zhCVRWq0z+220U/mDBbYl3ugWw
+U2Urx58ASOmQdc7z2dh3mXssDZ4xFBvB8jktuH/fymmMoNnRHLLoTYeudr5Rku1CIT6OKN72zXB
OyHee+TEAYJfJj8iiud7MZ15Em62o7A8yYg1/4PBp7eLhWG2T7Q/SkrBIzvPopvnzro1sHOG5QXL
Lc/Z0FlTdV3JNbnEQhman+KWEEm/Pq7dF/YQ2G7m6RZ5iEv8CA2xvgkCHMnhSAVNA2zuaBEwCGtf
lZQ7Htn8LG5wmXVyoxPrnsRAlFQdyyrvU7MtsEDsoi2YIbz/zd2BUEIVkdvreno7j5GOvYeJqyyN
Lcp1lFOwhfiWAAG/xjKR1XHFoXSdp+i1JGqoRyr5WLYBjvD8QpktgT81aoIePDxBLWyy5rN08eYY
ciCMcDeANvyT5pPHYhg5HHkxuQWlm/FvtxwRcHZ+n46osIwHYh1+JJ1Sd2wA6+v8u3ff+2k3juNI
HB+tqbcl/PHNwCN3HmiS5PwqH4nb+4bkyOd115FCrzEIsqoRhnfJzw1h0SldYMzr2rGBwW4r3L13
Mv5X/lsDpkehIT2seMlVSCPP3tP/uITRHKklmzoS5aFe+YVP/6L8R98vzmwdfTi5V2Vxfg7RjYBm
kSEhrXo0JU6+WzjK3OnY0FYZiu0ACahbcHQJchqDIt3VTajdiUsikT2HnOfZ2ykmtFOghyifO5fA
/W+CK6d75NqdEV882E2ytuJGgSGEAPtO60Q7oF+6qRfwQS+ZihUkEsQVTBg4WqPyuKa3NEdR4s+P
0n2LJyKAbcOgylEGpd2fr7sXATaa0QHtz4SsvOcbLT6t6WJCtOC2l2rl9ocnC8lFUa8a5DcQi77A
HirAe63SEbcXIRpV0M5/TA3WM1iuKeTb3M/1jewdZjMUpzCl+k8xtCghVqrUmmG2Zlj+O1clFtu0
rwTW6SSsIsZC/bumab/xpau7f9r5pS4GWg3RM49LYshVieUJds5yOpS4wkTSp54qGHEjwXU8ezjP
wB0zTQbjUmjHFb31iL01Q/sWjxMnaw5BHsZ+ZNtk1xhw84JMF2VHrtV0mF4wqYuM0vf8kX15DSwE
Qboq00qUe3EjHyZluTGzncQ1hGRXm4pxO1XA6UUjX9iPUI8nm09K4grAUcLU0Y8fFQyeGP9ZZfb0
j74dzKwoUIGSeWMgZvO0xHfOd5EtaBcuKXg1oLPVjXL++/K6g1nGhWFLEnBfFMOpBVOS1no4XGXI
usyU4vH4NR0EsNG2CpnBQt5/2j748n4LOdPxMOQmNUriywKsko29JioWfBrbRCaNV8m7qEG2BKTJ
8SsnSnDR4bFS0GrLNPvW68mK5/PNmKpmnTXh1P1dHYQpeZBwSkWSc5FMNLzEy0T+3kuxhZywzsqs
NXzcjS1aN4awuygei7GXRI/nHbzfHcKdEe0ZJjGlCnvGuVCcGA/oC2SeX8000YLS5vhws7OtOA8Q
CETSF/brJ5zFW5hBcaOZZVtwMrZciDc/K0+0wbi3kPbhBhh7E3yzlFFERmXSbTAsixcZjSU8RRj0
YppdTDOmp04ccii6ZopoN6+1yewMgcHtGyko93Bo7l2UIGOYJZjc/9yWVucBN3YQWi+gGuN0N012
fzbxTsN/1kGr70INwiSlB55yFjH88lFeRJKGixSA+rhHK+y/LARJwLGr9uo8PopY+w7rsjbfr6Cv
igV1c3OtPzbLHT+5wjc15ge/cAc3tUbawmSKwOpBLWodv830cgg5jdUxJ9mT3UkvK7bPgNHbpQ75
LdoHY9dRsUdkKpH91oEJh2o5kCryKAt3Qalij7i7vWu/946KJfKSu+D//l7sEdyP6WloCUpo7xen
jDf7iLSlHsWWgNbGD5r8uAYCZEJVL0qWW50b2/LBHrA1x7wsmm7KLhSpcDpt2RsFTW07GwhGx5Nf
q1ntbCpEg1FUChAkQ9qqvWO7w8vZA42X785gwTeSsS2J/q46sx6zDOwyMVyTOTIrViPSVuzQmHJk
9KpTOPZufluH7EEAaQLCk7l5Qgxxc9iUVc6ny1TfhBZRngRV9CBXNz5n3YfYM7ldB/hlsGX5rGTV
fo6lpx8gpQUkEgp+fYI/CA/+uiTlatOr7oDChlAWWyhiFhni7jCUANrpSxb7LRn9usLXl4MTlPEG
Htr3EfB+Pqpt4u5oJ9d+tEopsqw4FLr45LcLyHtbcOHuZwndSzIrDgw7sRlzfgZCJM32Ch4g41vC
TI37sRrk5eWLXMLQjbgtaKY3lcWcfMB922o0M4LCIEERqJO55t+Jmz2kN9nuLxngxuQdLtdO2m73
j56IH67/DG5h/7K1vBfSyzReJsixzncDVIXJ5Ut0AUxH/0jUpYu1AEwEFnYBy42TXZYa/lUgXT9l
i8fMDTCEtYl2DcceDt8lkYjOBUYFz6DKka0Eyt4jSLGKxECYhOxooBS2ejE0rpZC1NktbZFEPNTZ
jk4FEj6szAqeYykV9vAEYnEWtDMVTVKUhM14nV0q6iJTi9+kzgbfE6IPn9Ze/7G1aBEnmVOu9pqB
gDC+4L2bU2MQNqwIJ5CzpQduFWty55o/NM4Nysi+F62YAiEky2yenRYPrxWWdde0g0a/gYFq8Wsj
pSQRRmsC+rRuTbF/oWOD2sJU4Tl2Zpg+hMsrOgR8nYTGyUl1Z7ip6ALe61jLsGqk/1Tr7RzaqFaM
0ZDFTdT8YaMOmxC91I7W73xVrTDcMjrfHtSZkccG5mb/1gAA71W/uuPZgSgPwM+OpI+eqI/L++Mo
NfH8npQ2vultABg2q5uvpMKHa/5X5KlgzUkB/ToQgp5dGhhbvXp6PjlnfNe3n4UkXbrN/1vBASWu
loAH0JUrvDnMP4B/M4gySkHXVNMQDgwrGewyelcFjHcOSfKeIdKjajxdHXLeXOBKm0mAqNdMBW60
wkwo1xoHG+ir/NX5n8aaJUHKM0Xy8T5TWUh7h7bWGnCHL38kzg7Hp8OQOfQe80W11OixbbNqJFL6
FeRRlyplVHEzxooKE7iXUmDBu/JjToCGiB3HyorAexr1c2FOAqNAg6IQ2JIoDrMDGc4QZ+h7t+yi
y1oThHqsEKS6hKBUvoMmZw3H9jedMNWiwO3wGCrQ0DjoBJdYxC1xNQFm6KranhgW3k65dDnIMJCY
WuEGcyzqqkX83812YOO7A8f7nLyMb/aosq5Ue5VRh3DQsV0P6Y2sxAPfNBZfyOLmv1lp+xaZJUUa
OkzP7PUD1fgdxPo4zB2jdHKWOkEBjlejZlfXVWRR+50hdM9XQQYB8bxXFG5TXGVpBTIm25vLIU4L
3OyU1VBCJUyGd2c3tscYAs0Q4k8P7Lc7pPcHWgmBMF+RxPvIS/ukvJyul4uy1W0VBOpZMgK7ijD7
qIgXsjOUmiCZMF+bc0iejI0a7a8wNNkDD9uBQvC54DupYRNoig7V2tPzesux2tpEBrdSFPc0NN7p
etbD+j45VYqV9vEObBLNGKuXGNOAxdL+iyyr3VsW8wXr4KaDiywQo+xKSjU+kXkUlWVfi9MhPFWg
yBxAoXeiiVgKh/tmnpmIOH4dprWMSmvTrYrAV+CsVJmto2DxDLic0gQgtxzFAoVa/Y+RKRCgMfuQ
KOGG9Wcgun1coV6CZuctHXMIAyfIBmK6YqRpSw/jiCPgb8Wmwx4zjSsbObX8LaeTD20VAFHwkcHy
2g2GC4DscSCoC8Eebr675zlWKe7UegPsHTCDM6Cy8qs1tsh58OK5+OavH1xVk+clXqhwPMTl8FXA
VZLgORK9O78d4n2k/9gwrtMdhdJJmokjB1Kwnivh0hKAhB/CIxvSQ2/r39/FXt6EsU0IHUy7ZejU
n2J0ISJewhcYXY9PH+5DTyakDIDG7v9by23HOXS7wNgztZx60X0yPy7QKDXkaNibfu7i2II9/HEa
Dih9TstgPWN31K/9IfNWwNNwr6By199bVDvZHuKl1YlPqEEl9SkldyT0uzoGcIgoTCTeeYI9fzXO
m8fluCsHY86BSCksSVLNmCc+jYpvK/U9K9ORLn1HG9N7oNlJbob5ls476qb1i9lwFdAxwQdDWbtO
WjLirJS4YIX54RIHYxz5yJCVljkfOHOBxyoU98y9yiIK/xN5pAg6GfMKprjz4dRBJJ0ARa0kf3lx
UnTJXTwvs1mipksitFy0oIHMkfZUbSzaMIoC5If0AqUISS91iXN5i15RlEUQ6JOHn9GAic6W6Xhs
JjK3cYijNgPJKrULLdPR5QJWSd6WehI/m3oTME0Nqk9szK/a7YcB1dBlRbuK14sm3wp/wfA1M1L3
chMKOh/s2Ph85yBVlQFYVlbFNFluT7xEMeKRVDZxpSOmrUgktqum1j/Axqz+6QEcPKRxbhcR50VP
7aXF592dK50arMTWvB+ff3L+jIRaGsr9l1Wvi5YPTx0oM2mGyM1tbfG5YUWIdO30ydHxa98cDQm2
JPhn1wYJoVNY2XQ5GwHX0buZt578oGdnejf62vajwgHkYYV4XnkweVP40AHTx08tc7D6LOKwBLeK
QOoXrDMJKI66jNy8dmg7kl/ABKkh7zl+Y9L3liCUgo5pmyZUfw6vzMSBLFN7BPPUpnjpJWAv0ozK
uNXeB0xPD9Vat4HPdqQlE0wU+tL0/4qVwfmctQEYCS2zMQx/zw6hpGAqePlJbJl9qTtWIVPDqwtL
yEa2v4HFASkortXpNBsxH4p1SIMVHwQtdXNfK5pj2OqnqcdiWCuirkb5Os3898lEFHMSAvQ3/raU
8TsTyapldfCpC9LbU523z7QaipSE6FfGgq1slXcZlJooJXqLnb6Xe4xJ8C2tMJN4ovl9Ki7IcrVU
QjNTA2fNd8I2wKmNL8bvxzq3lL/095AYMuSmqWwNbO1JpxDhO35/B+VPokiLEIWEJi0okLzDOjRw
hFAtFRj4VdO5bNU4cZ72ynZhRMVtBzKiuZTNiOACkQT7U5LEKurnu1pmxodG0AUkjYZPztRglbc4
/ZEwcDof6EQpH12ihQPeQiQzlQ4SR1nAYT5OikHAhWPGgcz9vtphpp8b5tHCwg0DzoTQH3vEQNU1
ydwmjDiiRTDMvT6Mve2ELG0NLS1jN6mmMyEhGKd14QrvcNNMSO9uYrk0pSFWK53UloVbpQxb8Gj2
hBNA0egIsmOICAwusKq+UuNZo+HlkdCCHcjtLhBsIfOfB1a0qbHhaX2TH72/E46RJCGYMmUDLWLf
PWiX+rtXSokPrd0b0aBEPjwuFVno/EJyhK8op2is7P73+xcKwQn1ir5+tmcY+pw4vtmTchDo9cB7
wTWBbkZZuNOwERnxsIHdNru2pT49IYeJSlWlym05LfJaopDbPrD9Ilumxt3Vn4i9/dPF0lDnlQsS
cEsMjeNilSEgmYwNdjRWmQH5HOmoXB1Lzj1RDI8A6gY6T8FD2HHfck407BWteW3sH4GH/7IenZUP
keTZYodE2vM46OJomNT5mqw0221ea3xvCKC06GwQAMcgas0FymnNXAkobP5Kt6D+PXKsA0OVlRlr
MJS+rSIPevo+2RreK6BkhVS48J0wJ1E7cepTy7M88R4WkCe+IRSn+Sy6Gu8MGhMm1fiwehRzbNNS
bko/atzK1mSiRqkBeOKCBAhp9+egquOgr4CmF4pVGg8wJlqJU7a/8wioCgn0r+liAxjpqKDhYL7O
9k+ISngF6k2XbWvSpdCnSxJ9u0Qefl82rHVcIVW4OdQ1DX2uQOSC4u3z3AyMHsWB2hZFMNt5Fr7V
s6Ob7lUfuXzDE6CWapffg4Xq2nBTCI86kJ+gdmkLxIrbnniz5aKU9USUHOltvqiEdvnoXGbBd6ut
0X8Q40KHB8PBx+4ZCPSCYzFxpTJQ+Dp+eQlYyf7XHoOZUYv/uNnf7u+IfzId/ocJUEkBwU6yxunW
NVhFTOUcNZZv+DuWKgUnq19SPkpU6b14UogaLNcCSPM2wynwWiwHWAJAF7nqCdTdW26mcHE3bKIB
GSI5MXqO1Y6q85tdqzJK2f7RQ4QzwVc8F9FFYt5TghFcfzakYHMUopRWvLsn+OzXnhztea8PvAil
uD5Hzil76AL+zIz+4iRobAlSHp94n1uCOPO1SNfSTi3PTXbaQ1Dj7WpHjolHjZXw1a+qFEt9R/2l
fJYi+R7ElWGhM8T9pyYWODVqUiuYlMhfQDIn/vCKwd2eB1cuFNyJ7TiwJW3V+Q+Ua8mSBKHq0Q5R
+KLVemxFI3kle0W98LF4BTGyEe2Q+qI+NsaKnrLFlaVD/eWDDsnC/AuMvLft7dCqvwXZ5XjZA45j
mQqn4R4VnGYFgBKyIa2gKrwK3eHa2pHNOU5Gh5/nWgu16vfiLDWL9xlxogxmYVX/Qo5b9ZNwH/LH
RruWEDk8q6ZncWtyTGgElJ0otsXsetdgtP1AfhlIMOkzTLn/ur/lXxxxZkEtq5Tpgz2bgQCQmk/C
nlKQwdshV6hWtDdPfUZnLGoPyVZqk3sjIwrIVazNM8zFMiAzUq2ExtMfUpQuSIU9rR9CvAgy4shq
krGfe/g7q7RKEJQXSHsopflEL8BRVuEI9CdKMju2AB39YJEmDGYPCQi+tWijRvbTdL6UxOG5l9zx
ZhxLy3/CutjhfptqwJwFskVlplN0xFUTk1AlEp9zEBhbj8ZeMg50S+BLYTrNNR0aWWBQoj74uug/
+23QdU7B7IM8qEym1zBMJenA0Q1BWFNIqQQNCj3SxGqBtZIV3BWF0h6PtFyVR0uM7LBoqffAuprw
NyX49FjisFl0g6yNMiToinOc8Z3mbvj/n7n56eEkSBKchyyPQLhdMzGvZo+h2bDjGwf9Yem48qFW
OZvZij4SN6JKqsCTrhpB4nYGMHQm5YVkzkPCxCGp5CHMum4MtXv+DyBL2XiR0HdQZ9ccuwt71+LQ
bwrfB4MIwt2+6CjNjEGH9eWLpWyV4OIm69KWqhfyxZS/ArgneY+L3rllI+3WV0tHtHkOjr+gDJ7t
V7HzGqE1ULgDwu3NxLvG6u6qDOaxGdxnk6f78zphl1AKDi9XSSOcC/JpMSdyb/o8qHz/kC8xbS5r
Iax8CPv+rLkxiszXNpE0QmcFSSwI2VCBsoTPIwkq3rM/equFzPoP8UDaLiXvsD1vE2XrIK7tgn85
0lNucFTkhvSCeRho2cVbVpQu6bYFWsCPfI3lAu0OnoI3MmmJx9t1BrEj8MrQdt5Msftd8aDNFUeH
0GGPoee3QQqSwCP05r3xR8lordXYhMQWHFG6nXQuTMfdDI9MTESuc3sJev8S81E5YW+xnY6EpmbS
N6iumx0JLh+cZSviOVTJi/b3aer5xSo/T/yKHklBaIwtf9RUHvfDNAmnRBocnArrflEgp5SQOHss
MD0JQ1ZEyMYLvkXkcyVZroXaJNrMSMo4oTGNZpq8o+u7coIF5V0TB6HfkIlj2QAg5vy7IMbZZSs5
FIxniw9TX8CFAlUe73T6RzMmdWKc3XDEcJprhDqDGNeBnSWphqpoo68PNIyrmNHj4TTNSWQJyVgU
90r70fNnBxZTEJiSpxbzHq171BUhL3Uw/gafGf59g6HC4XZhIurPjOZwWAJmar3Fgm6AHGcDjFnV
F6NiKaLss6dGv4iIEsF8hxWuuZPD/FytOFUysn0DXMno1NThDh+q0DySMUay62oMc/9U9S+v9zRL
g/QSsNsXRQEvWAlH4IU09jA747l+7ZJ0pwamO1liU8W8vkAOLaohT9RUvZ6YjfdzTsDYJwwsfGlv
J/WpZIh9cp3JffWoSn/HhIHckVHOIAqJ7yJe2N5ziA9rgvkjeRuEefpq3yPFY6BjasG9YaHc0Sut
4kmjoZmt8KKjBRMsu2KglrPbK4AEWjiOs6TvjqKnqM7zzb/GeWMFLGZjSZJ8A1EHM+Y/1kY3FZSI
GN1uT3qgNRbNEBfODGZzMRBTPF/By5GXYNbCzrSs9VsK3b0cIsxNDd7qWNsSLHnlwhxyBDiRhxA6
oas9QIUUVPlnJ507hsk9zVUVeWE+cHgmSvLzuc9l1Pk7jKhpE5fXscheFaJ6+ls9y5oLy2x9A9dS
8cpAUP2n0qJIC5VULP/sOjrJzMf/13NwXTgBnO2Kg4enaYPK/lBuS9EKuCQUv+QOOdQEp4xIf6RE
UgMsqBVGP0YczpmS9HNBePSO+kPSaMCbL4M2HN2DHJ3E3Pl3KmviDMcvHqnIqgTOCgWcSfVjm+fU
JIG36M9a0yaNxI4yv2Y9R94Qlp5mAQgsoPq9UblpQOuh2mH3MzEJ7qdnIZwWWVWG8CSbgAp08yBW
n6flnT47upCuWqOO7PP/cMYRwb0Tb0OplskfCKppUcEDLNfQ3cfXpvbPW2YfP4Dt+4ONybpRW5ZB
YAyPeSZl2zVoz6hElgnttFe3wGuq4mhVzT9LOAmSxzImgaHJUn1cCjEe0xXSidOheCGizBMveEGa
pdrqHFybzdN/mtd76bi/mkfsmOGgsVAxgqhKKRZXo2ZjytksIGJ8UsdS2qHdIp/E2aHjkKqXsUPG
Wupfj362uEyJoxWvOjPVKe+Ot5OgunJgylD/fBoJ8XT4yWAwb6kDvvE9WUXHSL7NmzR/5r0Az33C
InK+wo6T7gGcV6eLiBJY+4TQYANh1aMQjju6VdG/Debg/9CkzXvGb3ncsVqkqNg8KyncWKa70u1/
JeYC+U3ayyCidoRGLCFHE4vaxEdKK1Nbih3GFnYvKJhBac1E5gzkoC3uSRf3E6wMqkBlC6/yYfhR
YPu/rtHeP2MRjYUhRckWnfhno5L4Xk1yvIhLaf7Sau1kW3nHlXUR9zoU0XopVnEhl7+L3/0jW/Vh
7J+gvEQC8Ur0SzcE40pUs8CWCklc/RO53LG8ci+InUdsejboz+n7Oc5eyoS1ibBzTXOMsp4NzVPd
fzdsHG2t2THOoRENbKn9ssTyPpcbrEQDZrbcRDc3y8UPBpaJjCf8BYRbx0SNk9YQo248xeLT5wrn
4L32RRyQ0vwQ0CM+/syirUOh/DFtfXGEExR2ncQzN8h/LpWHIbGRR/+bCmYgmnghgqxj3blg0rP3
JXgZZQrALAX6fLZhkLkrhxxZ6zVW3XAFGUdMR2Oposkw6x2AiVAB1m2VEXTZDOMU7vEPSxfog0Ld
HPI9jwEWQ5igI2yZmcAreXPtk6OVS8b3/NKlpQr50m9pQHjLfdCU85EmVc/ftNOkrrcQBZqrDpI+
w64d2f3QVMNW4dyVpSiCpIlPbFWaXtOkwYQkt+X2dO7L3GYXi286jU+46fHLJUzowWhrT7XITuAJ
U0lefo7xjtrIxgyq2NzgyYTQtpzoDEG+AVI7nmdloxGKhhfYWhFhSO5GKFW4nawHjx/6SChE7dpU
k7KLumGgGd7nXVEwFRLyuNey+0oHSNMUG0nCSKPEruUwRrPYaRUMWYDIJ2PxE74t0H3Y4OoelTGb
aJkvc2OMNRXkGytZvhThFZO2RwuJ+QytUzi05I1YBcmdw/kCwJL3IM0KmjydnUFAvC3w3p+5iOBI
vvLYSAEAh6LxI4yG7hucFvKHw43pX6w2OAcdY84PW6YchVLFa870EDwLF0k68zJWLQIne9hAUrK/
AbkDh8uMY+SvASab2VKVsln1Kh6jl4OJoUMe8sPidy+3hL4wKNWsOFLq8WhuxFAUjZ4TVdRM1bCa
x4hPpOGbV5WjsRz0O6PuxZV9tIh0vRGsUxpcujnOq2683WnA2tXrinuRo5HrWBdtFS8t4TlelWUi
Jj54PC6mLMHDqmsSJKGoKs2fkJP724MOU8ggPqJzk1Dn6n9AI4ZeyuLkD0AqOjNWxMaXYTFrRNnm
y+JtMXslQAc4BbbSRacOyGrmdjOMCuZMKZJECaL6zW3z2AtNC6Tkruz09ZNYS51QRaCfz1rNe/qy
TBWA+DsGqP2R3yyKVpjKN0HbyTGIC7aFaVmNQgN2H/vm7Tte8OJGNCTr9yWsk9UPK6W1uwzLoh7C
s4W0OSVv/IlqzKCvjTyqaAoSD3h7LONbh/RCmR6vwIiSM6hmkQRJW82FPUUIecXGwTPqDlrvZsrF
U5BNGkAKTn920lWqG0Ze5bQW1tfr7OdIiohRL7quBx+H3bDKgwytM7SMMuYZBVbVtuauy1NCBKeF
rqHtVc9xKBl76FcGBw5K4izgpwYb/Z3KfLArYxTh0NzVqUggUsIKpNIHG6VYjqh+W+5BTv7uXshd
bnqVQlOWyyibIBD80Bs4e09O0y1zr8PYSX6A8hArVFwUFVCFM9MtCjbt0Xr5LN3ZyVbiAYn75ekI
+ug7poyruFmRwstn5KEMSFMWmz94fUvHUiZLscZkg7HmBLE8pntG2taZwZpXled+W4yqKIfW+E8g
fD5E5d3UQRXOpJNQqSP8ShYtJunaItsUHCiOymm6pBNCsr88Hd8uy/LSNoYcAcVi+/DNvR/bzY8g
vvP8aVlYeQZXXPSRuE237mXDBNMCBO+ZN7q3N6u1Mk/DXg+t8NhJNlkPW7GIVY2zMoXmH0IWqSM5
i9i4Xhsq3wiCX0a+CLCc5K+TKlyrcbV4DiqrSfd9C+VLz0NHUCVB3MYBBPYpun5AWb1QB8g+gWXC
sDvcXMIOARaQbd1eiJWRDyEJfJSQ46Px1GI67XN1+sngKKfOR6LukLMxiZhN4+KVLDWxKttiHjx4
3f2gkijNaF+sh2I5g4Zxfk33LSEb0YdL0VxwO8qHtkwI8ZgW+WL0I/fm3fG8xOh2tpgfvh1uRRdV
eAIGRpLKAUf2GWtVORUvN/czZUOZySaU5ByIxcjIC2b4MiMrxsg28+rfaGgCkCoLTa9aIJvobm7M
jMvNh52mhGWguhZa2GDi8ZTHsIbJI3tAFhiRlsCjzHEF/DEbcSyEFfKLp4wtnAW16k+kBN7qqMPa
45XyAwy02EyqhhKem4OfKltQVG4VJG1Pl3n6byYdBy6nnUceQ6GbNWDgVcnN5qIiTRyEmXywgvhx
2nbBuuS9q/BDOPPkq77PhHL1QfdxI+Gig45H+sFYxfrM12ITxVIHvrw0pzV6GRmxV5JaMm6obMjF
Ihz7ek/zC0oxnTLNSUW9Yx93jNeLlCd4II6Sa3/3voTtDUgMblnvIaKX7ynLEAo71kLmARhVsRK9
Aua4M4jWbtxqsOghj6+484YY69PKumu16rlg5nF7znTUGxbX+Q+nBYDQ5FJWNxIKdkn7xlb4tvf4
st85+Tvn0/bd1e7KsbeuJoGDGKIME5KTIUIUO33t6dN9r0xZpcUqISbHW8nulrHSOSA6cUcYuCrK
iEipcD02mRI2bIV4jg1ifxsZ9JC5Cozh0Zn82zT6muS6RxGBuXIGrcjj/gOVjoFyzgxpH5qFnfOm
MqF8Npi516cobwYOJMSqwz5jks/JbjZP+n1GiZ2by1Av0nzbZKHsxl21tdtrHAqAKtPBqQo1clcw
VJQh6rrUTCHkXtuvckLKo0+cUi5dNDFL97cFEutyviiDbQWbGGwQ8PFQtDMu7ggSsCxgrp3KB1JT
3TxpBHr+pbRE5n/QBx0bs7uzpvqfKT3YxyLE9ZOfpVFnrLR6N/f4yx7Yt59nRre3wVybjcRBqbmk
7CJs0QHuriSonblh1E46j2fqugrVAyR5yF7DEnx6F4DFwSB3yFibFcB3mbc0Xa75qJu3IoMkeSe6
s4ziZxEVLghvc8kd73ArUPbnkrykP0BgmOPrFHwYNVzLSomD1kcOHafNNxRWTp0Dk3jAk4eK3SWA
2LdD5hlb07jFFtX6UkX8wuQ0GEWRJ6e6xtkYNIqz6TV5V8JFpFyuWYpbphv8Mz+tlYEzuW6Zn024
kPN1Kwu/iMniCee81n9d3YwBSMXhADHQ4fPMngOlEjilQlYiXl5MJJnviX5WHYOj2C5ZUK6M2POr
092RnF9UX8Bo7Tx4hdIJT0iAXWrB2s76TvFen1NYgGB9k+bESkK8pSMANOfDNcZ+xMOehZYXoQWv
4m0f1v2VUR2HFNVMSn1zvCnUp0jH8kk9xN0gWm6nfggU3qMy9FWhkE+AALaNpxZjC0t0LeJXdhO7
gm4BZLaAHKihuqWU8l0FFRJDizhbj0Y06U+0coCj2NBLpl5L5UacK0csSupJiDNK6aDYbDcDANK3
zZ+Hf62X86ZP0tRb+yyQcuO2Myip+wBQw0YgEVGNQ26pBtt/m5DRho6/IkXygXbQy77C8zm3kF3U
xvxYOgPTQVYLqy8zU+Fv1cZRbyl5/Xj99AePYmQFMovjGHqLm9q2m2ooNVo3K/HYONlKzUJkxJRg
ImPGX8EfPLpl0uTnA6dBRWZKo1gejxmyRPSro4MkB+hxEfuD7YQar9SpUc5M+WqcG+Nr2TISqSp+
Ec2si3GmQC6iIOBqFvXeEHTp2arK+jv6ZXWK1jANH28nnU+QxfozClTCmwKqHaIAHcPkJN7yVoj8
oJ7pQ4vWRzRlJMgQi2/VM+RU+CrOfPtXHFTXTd7yUmo+tyhACy0XQIOszEWlThOv4BkUnB+WCETF
+lvX8Aec/6aXGe/SQ5JD717bGArjynyC+tEtoaIzb0l9kOsbv9xhWXSyaIz8c/mAzDfaVn7Ri7gr
K4ww7UBQ70+qtsOrnaiNoPKK5Ktfk16yZDHyGzqCK+LFhnYMYsjV0XEefm6Tfxak6QoEckAH0VLl
4gpu0ZJLel7+z2QAOyge6wcr2E5Wwd8M9jmuLVq2HS7f3r5j2bkqNyAh5AO3VkS6uqx2x8v1QbUW
Z/zijL5TvK00s+7N+bR2M+zvyVXSO+fTJexxIfhvRjueX+6kO81/lXrzAqOSgxrDU33QdQvu3g/h
r7hdpkgt1984rrc94cRD1GGGGY1MYkGTyVbOawyahKTIRK2bHuGQILhr0GRrN2pGQ6tr7Iu+1Gkx
nDdkDgxP2/4Vt0FR7aJuX4Uxxh2FYRpzh+yvWyiJlye6Gtbf/ToaD6UgYRuvLGJnWkQKVO1BFKqD
Qk9uvJNvTyZuazV0vwDK5Wk5KCHD1y7xniCJKtmoAGSH46jL6cKH/ZGqb/5mgau7AcT3jJJiOQUi
pPZXAtsZjQP0E5y/mU7kltXqvWBxqQAwNCFBtQcq/JNTG0Jkmmd0LJznbeWs/QDOucU9LIICqdlb
+EMykNewgcfCPvZnsthYQonYdAHOF/QVBielz7iD0OtgvqjEdJWBtx0CVIMmgZbB/9SoH6UmcyJt
VDQdbKVbK0jEFc531z0RBurMmXfZC0yPt2QHES055IzoO7YvjZpFvJsuBHkCY6IIE1gToYqO2XV7
pBFbZfXdXRk9uWFavz5IFZwDBUNNPj8l6pda3aABJQuZTprXa4uVHJJpZVJ/EO4IbKbQqylf3/0B
fj/txS2QbjImXYfkHf+07K1gA/K/3NVkVK6DCk3YwrnBcddFXyiQIcX/BIb1mSkX/BP82QxEEg8y
mZtbzgo0Yxo6Iqqx7eMAqCvcFMv559la9Ne8pG4fPH/UcFE6mHMA1uyTWD/sUAind+F9dXafAzF/
vl6/sxyQRFKh2PBb+MSjluLNcoaYvUcHYDcdnT3VqSL5fdHnSpIaOen4DgQT0d6rft8Fh7hQDl8R
1s5oGW6B0uSX8ef6iRnN+nvwdYPuohb+7nWwWqs4vlFFkTXt3OTuCz0pLcUrtrCFvMD5NpF6v8vr
wMeJgqeBMOS2045t7j5xJR9wENQbRHBeMVdbwmy8n67mEcGH/evLiOyKNPVsuWAulFu0ANGzR0j+
wv8A2UxaYJEWXUvMR735dVj8ZIYZXRNfFXEN7hXCLItmcQwXRCK5mghut2wMMD0PwVd+kXxK900o
iJBpob9ZysdpDKuT94/2S4XqHS59x1QVgq5SsYp0oH+RoN16NPQQ2AWpfqveOOpdbxfpE2RT9nVm
S/mZMt18gP4sQvfN5b/JPB1LY+DShh+EsYpJD8/QDOB31SzcgcePZrnb61JuvUoU1wIyksRR06gr
ujleO1fPc1cg/xKNt5Q5/dea31WYxuL+miTPeU0pyXq4t7QGzcqxQeJEoRS/tePOPAokJyqXCG/8
4EeaO7QwxlT7tUMIVGn16V3BgsM7TGKYds2fawTgWFFjn/JPZ2ByKpA/4iwPMYrhen/Oeb+Lasaj
67nU8kTVFvEXj144NO9GWY8BepOnIZxQYlDWl1iTJ+LAHuqMkhAlzKHELL+fee1yncouEm7Rmnu3
cV/cD2A38B+JXVNj+qkr6GWX/xI0A4BR8ZgQpCkXDI+m2XFctEa5ZEpluBBsWPtzU6iDPpgnOFkT
w7OOmaEx1KNte2cIYmwFLtIVEWcrf/pidPfJ6yAbKxaDFxiAhre9V8dvhyeMM+RHqFsSfa7VEueD
LpFKL9uc8J1cls+qqAWAhDYjtKCvSO+p6jJs984QjpKeeFeZj6qYYF7IUgtIEsP/j0nl38qTvrpR
8F/tv8rq3evHe3J9BO36ptz8QBh3iP/8D0OyJxFjWeXZIx54BJ+gRJdkSui9gZZDseH2uKEY8uEv
6rphwWYW31nh/Dv2TZOQXiw5kWThJcLglUYIZnbirJFoK/3aFaFYCaYsBum+2u+3zbeq/vngPg9Y
sTzh1e/MXraZQgtX9fxNjNMPtDxNLpLYx5Hcv/xZwxqa3UdbGp4Z8EGE8/6b1kUxNim1NQt1KlGi
CBF37Q5sAPpiDmboOR/zzrUtuRszn5jtlc0eGrHbavPgG6fQS6ezyyKnwNQDtrtbSfcXt7l4CS1x
MB3MP5BJ8kN4WxA2YJZQ5Ht+M9IE8qPmMNyN/JozufdEYYUmF/j7NsNONzfdFq/wYyCCKXVJ3mSd
TIfPyoEF8+7uGad9FuTqVq8VmzS1FVsH2duruOK5gB2FNSEtbY2PjL4ZrErYBWJOfbzsxD5rRCxn
fpqdRDtp1wwX5EzRrqJH6DfiPiTRU+JRCgO9cC3lANxcJqUBeKc+Hv7EvmDk5fZv+c7dCojmBfnh
sMQqYe3roXn6rtY8SKbZaM7DhJZgBFPr/sm9dWDVC4VXhhB+h4fzO/GF/gHbDNEylrLQPlFZqFSJ
SMBFeZ+UdshlhNzwDx9pO+7x0utiDuBbbpvEOp3Hp0XW5jxUxYsLTixJmsOLmvvYOGvzlpGcw7v4
dginHzSIu03k3gTRjzkFAJiPPmAwKad9EmXyz0e4BRv9/sjxp5x8afVpnJLQpE1gV7IotGO278gJ
kLI+McPELJGUzaLLYXfnzupKg26hNzLNPO1cyq1lAV6pZjhFGeU2kdmC7mgVjRyPoSMTub4TXFLc
7XsACgnLmMMlSDe9EJ1Q2Z1x/qhbDc/hvEBi659l4bhWCTcgscoq76RMfkSX82KH2r9+HZSb0xiG
hSzi6AlCmeZnC2IKyLzpvIWu2nvelpLb/HzRxd6Al1FnbQb0ekpL9fAxGkBJEnGq0ZGBBOv1VnOf
aEHCvrcW/qUvhqix2jxy7cxDj+z07wzlWa+MxE2bfjxUUDCAKfVJlqCzTUAePyDVssQqHxfLZqwP
8FmNDiVbaDQsYOHAgGRDLaHX4p3yj+ep5vQT1iSqT/ERBQSU0qkOvDnmKJ0zYxq8/kHldLvR0eef
1w0xq6Jg6O+V7GNt9GVNLD+U8DuAl5gkp/W2D70aaMc4mTKXlCoeM5HicJeR/jRYRVTcA1XqFiam
8hWNof5kvbzxZYIElILacaEj/BlCTdm75FYvC077ovb2ZP8PLC00dK5TtP1z2y13HlW6P0tWYUE4
lPBrZKiyhPAC6zncKoltytylkSVkGN6Go43crdcvEHFLVewxMSamMrlh0TXd78xxbyOH9r82POUg
khFWS4F16Lbf/CaVOHeN9ufpFrGlquYivpmlppF+VmAzw2gFS6toNia8UOvgePcmwQF64/ojWUai
r/8IKke7Gxvhf4DQOaVSceXHjCLdGQLyaINHL4IMi7MHRfCOg/Q83LspVuNW2oPjvZQHJWiUd79S
qfvQfDnROq70/1GLgR2Yb6tw0qte02FbPQdtvPj3Zgfci1d+JGmB+OjEqZwCLUQMxaC5vSzLRyDJ
vs1zVWOYgiO3iw/lgDEPTkQlyXb6mSmQdoKTiRjlcqw7EzuFtas1JH1kGQlDLV60zsab7S4cAQmo
wWzcxNw4zz6ShpsV9xd5GlRHqGMHGt4/FTepb3vtM3W4GfD+NyrTf/BAQ62+mezOK7KpUGFXoMCU
rFQYVKnfmjGXl8S9GcPcP/Cr2h0heOZxN6+t73Oq5rrjb52A2r/O+PbSFvsZ0SC7dkkB94ZW19gX
MmprjP1xoaDUhfowyZam67ae7rmO1DCvDtUkq15HcvpvRAe9L+N7zePePZlLGDZMLhzfyrGBzX1G
4FG8FZEuggBKyzjZyGgBU7FlboXNmapciK7Y8FHPb176+EOQ1tSA3N0IOt0NebjQTwexATGESEV4
FOBufyO0oJlvFWwz/8sPkmjhU2nFfqmLDVd56BWL6BYZsN0sfX+EuzJRa8A22TKjxIHVOJyA2ceu
vOOjw6vdb7NRAj+/N05PqSQz71eh+Q/x7LQMHhqCjkpDF1V5a2xvM+AWmOgsRfo26Sur7sxuxqJk
ykLy/YKafn4FHAAqkBb2dlNetxtEA8gdaDvDWywMYE0OYNbVxoJ3mwIqBKH/8500j7TBB/CoeH4h
ceVqz54T+FAqRSU5K2vrqsckt9vFS5v1ZSB4qOn1V1PENJXS4s/bCFRGXK6NiuxRnEuC/OvVySiT
tn1zdM3XtC3zE0kPcYSrGkTnmWcmvgKW8u2p8X1CwNI76g5vLPpjCxHHBebce9k/FEySyhSxlPts
53XYHXbLNQ4wvt5L9bmCSMctyRHlceks5XdpkCHE0E5UGzBfug0tspOVkln445kgpMpjcaSUFZ0Y
QP6bsfHLmtU1paAyOmGIWf6uzTAUETQg/hZAGX6iIBnC7HFZTfNUhAas+SYfxurDF30NfUhgoJbI
GVV+FJZbxMdTUsRF++SbJxGpov9/PHmSQnqHsPGIPrMx+BcCo2Kf5QO3KavwHcAqG5vBwkw+DEGJ
NEvNA1N23lJdmxu/c8RrUdy6XL9/JJJC0S58fERCV1E4NNKWMP7NtlabKgq2PpmZ/u46J1V83zZ5
6RdvU6KnJM7QHqPkztp7UXWp0PMnMSLiadXRvGCbyCIcEfOdao/sQ6RFR9GANv+f0ENT74Y4gz1H
KfnUZXz2/lZ5hdPYj1DwRCNszI8Ht3qPQ0d/BBriA9JDbrMX2mPxG436gUWskRd0IjqmXcZkz3ug
3eYe9o67ovT4xTWyGiE/fis/04NEbe9XIq69pxIExhx+30L3K6B7zealIbGopAcAszmbhReJ+VrW
uoyy9OID+bk4JcyI156zKdAjchpOMcmeh86cPgGKe91o8E2iY+YNsjgseXHoLmR/VcfRYqppDGAG
K6tu6gUmhBa6uQ6KkaE0d3O63RDDILkMIRV/vi8R47PJXD8FsFwrGZ+n0af97Pt1mMVUbB/LIie3
iAfAgk3VkxqON4q9cO97vjLA9j4W1VZu6kUUPYIzxwZ6sZ+5+OMTJD7YskiM5KIk4iMIOo3yb8fW
cGR1yRxoKzzCwWyAA2DPKauesQWfDBcOn6OdzFJuolSZ1nNgA8NKV1aGYrUqdQeRUVObW0pma9/a
saxlZFkaK1Gq8XGHrtp8ILAn/MqGlflSqEjnBaw7xstCEjQ7mQRVdNAEii0RRKCTOtu2Gm4yO7kL
zCXhsiMKxaC0s7nRBmW5Hyl8zLPGgMDrAbOtnZqU6KB/TRbC3kZp22aZ1Y7wdJikFLIpU9A6KIqg
GF9sIroJxUdXoG4UbQMaJM7IT0utstMiyE5B6aV+VT7bGHdaJYGxsyLugV9vRKunFoI6z9i31gvv
l7l4EjAq1gYAbHDLESmHQulVX1Zf1GoWQRarTMu8e1nestnliFfbB2kUptJG5xW5eXSWz3Quk9UI
nduQksa9bp6okZZd5uxcnOzxXmZ3fmPrwv7fbCVu/rOJmxetF/HxfFffKKLEnliIcEiSzOTMc2D1
ZJwOeP1CrgQAMoCB1B6L126f+Y6D4rMufAlXqA5HVFhrikyTYKRtYDHA08jSnpEkdwhATaKE0SD6
AMtOswLlZD/8nRrczOnsotD8tpklfIBNKdG4NID0IKsrPgGXpWCqUBQ4Nyqm4pCtf4qbdfnxGkiD
HSNjElhZQvxt8g6u7QTZbFsNDj0VA6yhkEgfdztZ+XFg5XETN67t0f3N+NU8zCq2FbwHGPtYA+Oq
dRxELtqVhPtiDp5BRXymmYgWsjbqHIr2OuVHshy3i61d6c8ensBmVj1AhGBe5ON+FqxZhTYiJzF0
Ivi4IgKen38k3dbgNpXWZoA/xOgSnnR+uJLqWgAJlFp6ib1eGohYqDD9lcVvuSeMC/9P89hDZzHr
YbieYCCjRRxnv2yD8ncqyZTDmOBy4DasbXt/PmG4t2YlVW5PMUlDwWNp0/4t1TfFV/rIYQ207X0e
bvTtFyoiC9Rb5mvGqayPmw+NjmNx5JmgS07j5OzjUFWxtA8Xjri9bvZMN2duD3MXTCM9O7xmXJmY
GlBps/p5SNUaYLSRJyDJ96oMeRmzw69YnNmxmaU4f2W+yPbyigEH7oHbsg/JviFS9z7ycy3r/nm4
i6fLRtstBRUdtFxW3hwUe+hoJvOu56i04Jd8grn/ferKPai3Ov8vtTBFIZjfe6xxFGjVebS0q7co
AwLA+TpeXhAHCM3Dopk0Q9Jl0t9R9Kz6j2o4W2DIDnI+WimirWeBXpw8zlNRXpy1vQ1LcmZ5Gvxz
VlYKZA4/tBYf6xWPWFihUDMO5dMSiegd7Hn3DcasVff1rXeIteZ1UCXDGHqPmQIkcDUMyc2UYD2d
nCM6ZqdGtmmiJBIEmo0rsbjGKFNR4SIajL8DBn1GJd+uesHwPskr/R5q7pxLUb8QypZTnWHSURZr
kan7l0osYD7yi0E2lvEflt0Xi2IfVuEqFtCjJ4ti9WDBa8XmR/ij340RA2r4X/CDGiJjCJalb2lW
HgJfU38IFP+y9ew72HxkPk4r62CkXPT1RAj6qL6NrTUGJkXkHiTMIt2+SMCBVrZJGwHYwTY5tCSX
+DgQdnWHHCZ2Cy9N9M0LE747yl+lwUsQKH1aeGeYAasvofUf9NIuK5t90t+AVz2tgMBmFJ+S4Z/7
6eBm5WeIMi32qCp1G8NQbMHLDnwDuQon0QcdVtgNSf2e0feCKke4eaPMxhXahwUUHj5Ga53Oihli
jc3c39NHTQfop/gXzD3d4KBY8bxrwi8Al6dUQWZ2vMp9BMBDRzLB9m/fdjr6rj4O3sNbuhojboTx
773Whb7rrxSNzqRH23TDB7HAtZxFbBgv3ZVSU1FCwI58r5pOWZC1u35Lq0luToLZb1ewxoH4v6oH
Q9VdhdbLi8x/ov6t1ZiGDFK1uydYe/D0iYjsHoLGkF74dgALNFuZBVXmVu9v43vtMuIYixtxXwc8
3iMVdzQP/RuI9y7Z3igMGvKybkLS9C5xWGDWpmn6aWsUpqKduig+3YFwdmVi9rv3rVDh6yy1PLRm
k1tEmybrix/+tAiXglstugphL43VtHJj/of3F8XoFDUg3uOt89Nq2qMkAQOzwpAYbPJqbX+Ju6ym
e5wqTKWKp1PFDMNbBcbkJwg23L+vdC1NbnZFgjw6H83rpgM5yrmCdX5BGyUmXrAX4lVPx9S/M3Az
QJ2M7tC9Fm8STceUpnCTHvI9Qoc8ZLcAni5GGhdVEwO5eURdbCL9AMjFuUKbXHncWLqxyEfgvWGr
xW/3jHmeri60HAyCRe0RcwWw0mHzuWg4wKlUcswqv5+BTPXWbf3ATkMlMIwBhfaD6QyoQIbvGpsG
AOdfAdG87tsRhNh+LyN5JSkNW4FHvMvtcpkEwXrFQHJjkDNqv9hpmOw2wXKdCkMwBx0MtKXkGCzx
UjPAQZn1+48ZoQRx7yB1JpV8ANcG6CznMJaci4ncR6hMHUamYilBNzRreRl7o1OZMbIQze1p7Eh8
WIHQu/1yUqnbussLshSFobs1jkmKGAF33STK2SqyCuaW9CikfZbDPQTonMTAwxDXRuJ2zvrwv+B6
KQTco4Ivm6CjLFcFqszc7e8gL5EMyWRtn7iGSO/z/Hzfhescuyfj/6cB9yEN0AmkdX3I803OtdFu
EEo9xTZsk44/n+AoWBeK8eDp1iAvVMqd+Tg4ZSk4Gx1vs9Q7T9X8Pl3qiePiQzgK1P3JhD2atPdU
G822yW3Fm2VvNY245jJVg1msSSJHb5Fgz0nawmLLpF/28mpstvKfDb2eeMkb8m49QvAHUVlw68sR
WKn3Z2UbA5YlrvE35IfZ2xGekKDI1999dzKczsv3NunpwWpylrFRpQ7A78Ml5QkiFzoguaSlH7Tn
U/FARn5iPr9XkgcgOQwsHtS84qcEuWgsbjUNBzJEDVzKBmw9Vkr9jv5hOiSfGO4XUeECHBjTETCn
HpLuQO1UE5l1lkc3lmarjfqC0h/kh4mmvEpuGST6PZqiWTtuQ0ecLiNUmTcVK6NXOiqvvIv/kOF+
IZPopmfp0qgKlwc0xug36jtpZhRj5uKhh4/BeeASyBL6fDYr87WmgXsz8lKuzjW4YhYM88KlsRrA
h6UyZP2YcLIok5lhWO9789sur49UzgUJqYdqQxtFbwHKHXGPUuRHbFEXmYzEnGaIxMUdYMhR7ULn
8eFacn3loy7Q0rc/dYzsA1PZY2xKGF0IiV9OIdaJI7PL2/Bx2KwY+NuO3ORp6UlaUN0TxNrAYyMN
WwskiXP9DyOTdsxiC2ZFYRj0TKK5sK22CxxELJLY4QA/TIwJvCc9jo9gmnFZIKwATxt9SGy7Rj0d
XZUwwBChQ0LkqyHFO1BV9AuAG8A2nodq7slYKUIDnkz6c8ytbajlmUMiJLHLnnJ+Ybta2ybshi64
rKPjEyqcuJJSAQ44PoDhcbXoPmAperVXE/m/bFm7VpVgQ1Rj+bIIS5UCE/NMWKucD+DqvGD38vde
aYgeOiClWF6vg0NIMIEMe45Z87ckhojV7a8sr1gX1E7F+G2KzpaWp5CIr0au3Y4q0ph2r6KUxoYK
Jd17UsEZFTGux23JRhnWcwLrRMv04y5Jj8QvfjRpklnqNgLvwyy78PUo2uD3/jNBJldk1zcoM+ON
l70NttZ9mO9fEx/NcRta2OFKXHoNSutX/uK3kR/NhWvPhCoUuOHDmdjppdijVVkXB1zh+JUbeMWi
NLV5wub1RPuWrGHzH6Hj5la3E9CZcvw3eXH5mvZyzHqL+3P/l6gBXVf6BpkNz2iUDrnVEJxEJAzI
HQY5cj+icnj/KiEFLdRr9NQP+UUCuuYzDe3JlqXnbVns82g8ySiLxOltITmBiKK/6YDdJ9RDyd9H
FfV+4/UTVHMoWJKyP16hBS+9kyB9KW3s0octWkMJIw3N4PDKXqKRja64kuAJ7xuj0i2Z/CxZOJH5
LJhw65yd9HcKRblek2202Tx2OUbkVxqO4k562N+VP7BPNlYvAnmx5FtGLtFOT0Zj0cqMFTSJ9A8L
tH2wrIagFBLAYfbOdtZOCpUNNQ8JjHQnbOxnIwHZmcozJgA76HXPOW40hXMoZPtC08IFIK/rZ/iP
P0u9O34vudZeJdQZRKvw+PX8tJKn1BqOeKOe/WWUgVhZI9m0Pl4SYbC3AX5wfuKKGhqHwk3fveIl
t/hhF+/jzUwCyKluRDt1hFBde/o9EgBmpVLIRo6OJ3x4cANNge2oPvRZrqe98XXUyrufSEKFLogr
KogqJ6qSuwBTi9r8rOCkGjdqM4RMPw5ZWITL6nAkHe5U01GkDSSzOxi2vAh9yL1gMIoG24rpQH0p
3bdDQ+H81MPL9tdKnEt5MMJVT1AkrxEsanMqdvcvRAOa+Wsq+HpplSkyOT7V8/ygW5Pe+FHOGzZm
m8t+/xMmFEJA6Wn5TgSTHmzHhZai5/MEJ5Zt3ehn/xrUknwy8lQOVIRzxa1zjXajCVY3X8k0Z4Yq
vu0GNAWSfP+ueYB48NOpG6QXku5dFALIi9yYW7D/ULsN5+R/dIFBtTloqbFmJWJOZcjkAMpzkcyP
LACji7gCwDSy5ZdH3W2NO9tSJJgRjRMoNFj3CEgKTop5rzcjQ5iOITS8NSgDtcY17NgYLV5PWNAg
/O83XeRlcW+Iw7nfAtyNxQqqdmlRplq3WGqjgtRY9JyxTYAffeu/Ru6cyQ0zyZiM9BfvJaTFYcDD
xUrV4y4xsOtuZdBNgGOVI71uWrN07hXp+1tw234NR6cVmXh9P0pfvAjF6IwdV6cxITHsrOXpsNd4
XfPOBCwYLLv7VT4r3mZArmVnxlHyB+SdUUACoQ4GVh5n+2yMkFqUZMoK/mmCsVfeUzVcgdFz3S+h
Az29OUE9MP0xImXDqfv+pZldjYBaU0fwzAwrKV3+owFWZ6Cy92RNbAMRlbOvVekeQmx7UeRDQ5cM
OCSdH/+x7NC/HBJha0q7zCOsX+RcbqpA6/yKpeWNyi29qdxlXk0zQ3b9CLCB35FfWhmMiL+o2uQE
SbXbrub8+EMJavlDTIKa1n6Twms6ivZeTVMOY2xFosDHoBL2UNF95pnevjcA3KMtgy73Jr1jPems
UZcu9jyoUXvkUvn+u1CV6x6z/xx/zQilEWREsoItC82iaDK52xPzj85atC8F0XfVXbPnXarp4GvQ
vRozuz8sGqVueS+y2WvbGE86LEIqG9nGMqGbPb0tiN6B1CUCwgJnLHyRspOQ8jzB0s5e6zcsx9t+
Vc77JbW+WrB5112rPmnYxebqVPpAALiHysABeXwYKpuTsqta5KNBdQMKmzGqXr5UbR/Zj5VEyl7T
n44OoISbL3T8rENMm8PkhG0DmV5tFYUE1LfzO6lSSFbRS60glUtmVOvoM8qTdmebQ6szxnF2YSuh
NG59yBED4ln/IaWdBfdX9n2rY5dbWTaaVqyCNNkuptvpNgRRX9IsHI9AfEoM2/c3FrP0BATxdeIw
9a5SY/RFaBWhUtIf/D1kaQjLdR7YH08s3R0dkxH1DTr2ERt2znJnc8wyUhqIIgh0y2DU3ByuWcLl
SFOxjRoyWhoC88ycuKKBxCDyerBHflOxQX2UnxMlXLEXgysVh68X/mvMx08WpmDHHXiCFyB1dWNn
vbDHfbEFAs43ZrJNc7hMX9aSSCwditCq9iw4cA/12D5lDpaUsd8eWhSlCRmMJo2dyKBHVq5ZWBsx
jQsVcH3r+sB1vjjFn69E97Rr1jVYqmhnFpRmb4w6PLXbW9lNapHnPwOAGd87D0UtoKjsAnhHJhzM
ct50nbo1YuBXNjlw7ZG7vlSE3eKBN138D+PWYKYFcY0ecpKuaIdjT5bnXcLSj7IvcoJITUDJSHtp
v6FhcygprDNCTDcxjsKw9huyhBipI4SlD5y4367cLhWYHxO04lYPvBllrcMnda2b0ILJJ1/H7irP
bjsNjsmoTdPVRnSX2+rW9rkk54bR3DnBd/VtHowFXuoQDmSdk6Z3Sv6k2XZmU9Gq2unRiP4oTF3Y
1exYPe3Pi53wd9feFrb9rhxRflOW5znK4IojENXh3BWy7lf2QfCTeY5fqaQqxT8YMoasEh2PVfio
MT8N2g97+ZBnXadpxiRa3zNyuG7dXKOV6PbcMYjQgc7tQlmFONFlXrbzwkHFFAWytuDEwrlwdd1l
2RzVODnByKAz07wLH/VGjEtUr7vyNRVRHOTWKI79+FxiRGKZ67SpTMXlUZcCWnHlNINPwTGQfEee
ro/SD/qhamPqnf0O6R1LfE0uvxYvpQb6g7LsohIDk6+VaxV4d8XnF0tx4hPbxr+6VN69gTrSutw+
fLFPCvybJREBn0+8iXiwoLXNY0iGv2+hI2tpEGqKxe7ncLBIKR+fc85oqekCQySw83oQ08RX6aS7
eyuJngqCjeuulsY85AsseywMM5G3En7xEFlW9lNPnhPucwiiSWrvJGa2cn1X8uPoEatjboACVwj6
gMGxkJ9NayTbRtxwOry7nURzJdSxzozrywzbl3D9ITj9gKrN0Sgne0Rl44/oABBRVNwq6pYG2QOB
DiXhXr29Q2H9n5uKwPwMMold1db51MciiqvUMzDTlhjt6jdynbY7fmHoXtfjHHxLpKOPU3TeZ+4p
fW3EmtttjEtIubvRJsIi7rjxfrzaBauHmZQiklhSb4bz1VsltVGLkWIa3fswG33cqk1tR9tzB+a6
idU5PDUyJH5OjaG7U8FnS2U6WYs/fV0dkSyud2KXUuJ7sZYgWO7b+PZjhVoK9vTEsQ+440eSHAwM
lfNLi8qANyMy0M+D6OG38u621RVDpH7GWY6+q8PY3q3Om+Y55XxCXcGnYXMUafas//8HyZcEMGva
LNn7O1tIkl3PWB44vkj0tdanlq2sPkqagdWZak5A3LD1B2noPRVpkyyDRuvqLzi8lEXkarvJ9kcT
NFCJzmQ9GR1BgjEhw07D4LqH0P4coYOmlfDfsUc9r8QPVK8Qw6V18YjbiiOrR2MwWT+iY52KlkJn
pSNmlpU4iDCSxUEGn64to15D7WHjcUjBeHrCmx2fmdTeT83U5cko0/Y4uWESS/4mm03p19o5Foxn
QPx18hHiDZ8yboOw5bFWIzn2HtBR3zZM3FUJ2Be1c+0FiQm530vs0tAyiylWdB0P98rht/4Ls30Z
/e8U+vT8epDQJ8m7yC8uj+Qxtrh73lnsY/K0PM4veB50LcWaaBQJTBjrXv7YWvIp2mhYgF550eGe
nu3jLwl+5VnC5bKVIz+Ej8Dt2mxQLRWvdSsDFf6WOq20HN83TjvYfNVb4bD8rwQPcxaqMRNxvVzp
pLgytpZWNHHd9JN3NT6/lWqb5a1gg1LWZNBjvETqQgs4C+kjfToxPApo96U3kRl2GeArCH6lLHGy
iLf2pl1dKkwGCfkJjIuIt01MxOcxRf6wBgXTmj5issZEbGZjJgi+tydohQPGrk3+jFOomDqkAXV1
P5mtf/YozCL+NkOd9DuP8q6LzvsTxCOLzwbL2/dkbh5IyfLoCh++LMwZhtSltChO4feg0+D1Fbhn
OsTBz4hOXsHzI3H9arHehQ2GGXGk6Z6uZo5ETKKGITrbTWBMnZGyleh8O2rK4bALla9C8XMTH1nF
j0Jmw/+sR15+8Z6tCUQewiaxBeJFcvyBsim0EGbaaurf6TrjU0cMW6d49zzBJaHuEeTs/HdVsKq4
nrKBWFGfemzypKTySjio4CHckw0WCPF5Z0tLWcArVCsYoqDLe8vuM08K7rbRFHpxLX/OrjOrj3gJ
wdUtX0avNPlF0SkORRCLfk6onkJYsxDnqWgWS9W6FImd0jlDGKng9bPkcM+NmQZEUTdBbS1fLRBa
zom9/6MVy7uV0HAs/OkLl2jKLJWjd53Lwabbp8wR2JKbG/F67ueZo8Wv/nOShDvov6Xqv/dqSxbq
uOrZz2tk4QGmNstFW8vcamk1jlbJC0oxMbdA/UJuhRcYheFv4CUqDOaHniRoi6fTURpeHgG2tqXT
l2ldOx6xDyBNABMzepGcetsPrR6PseffQoegF+fkJKhYZ66gMiSabqGuzGGOvjVRm3mT3D23ze10
3PuxCVxOmpzE98tqbMS9AMjYKV7doaCan3hWds+QYslApaC6aQmucuEkLorL9LK6yAbYM3FBwKjO
qxDIHabOUrWyXluCPDTIIoBQfZpiojnyRzii1fJsYlhvRNe99bLl0vm2ousuDwc/7ENIu4cJUig6
KHMzyAx2X2xnbUwkjWIFOcSD5NCWxa5FGvj9mgfqU32qxWPb8BuKsSCaMurj1W51HkVroiHN/hIz
YOm9cUtTXsDdTY4WmQFOHdvsaMy+quKW2mRxCra2hvxxs1QFh8nEEf6u61qmjQ/OH8AkEamiWlb4
GZaZ80vAAHs03LbWt0YBiEUPIXBmL6sgXiXHB21SoUBeDqGkxlPqgV0X3W00WIanF45MBjbgV4lD
MFjwDchNSVKxmVsif35Owp8FXc6HXWHcUX3mfMxUn6P0WrwJ/3UtXELaJ7sKvhfrmbhNG3noeGEV
v+KvyW6xbBkex3pIoNVT+ozbV4x1BzJ9B5hCqoZ7h5WwtExi1Hp6Z6MAqegHrWGTMWZvqZjiFh5b
2NsEr2ZWSrqNZwAPDM28fync805k3kNY5FfGWPZnwCghaZ4tURB0YJSl3x0jSutBKadpf4nPgoJB
cXrApxy6C31ABWxCT7cLy/YaqFB4/jUhGRaXkZuBBTvELWmdJQIDP9NEdi9V+Iis09t8cdHLC6om
sJKlRdrtq4Gje9dzgHhYGSPdzgQxI/dEViXYk1AzZPcsYGrORq+weC3vu8Lesx1vcoWIz0otcQws
gq50KFHHuGX3uik8yU3FQpBCLGrjuYbT4AcjrdM71KLR0iTqrLNOond1gaEniItTJ+jgYN8HeeQJ
1nWaz9O6vPEY1UXGEXKoPBJ7jGYekizKn1xtbRkVlaC3e3ctolVwqwa9+I9f9cmP4gSptsoAPhvG
w6qwS4Hn9QoBU8nlwcBQ1Aqo5LytxIK1/2IA5oAaM6mqys4GoVavhFM9iDKowM4rotr/Wse8pw3j
gpYP5zH9He6dHyf/mPQH5+sxre8WhXx7N+QQJx0WSYCvUmGd+Yz+nuPipWAH62S9UV8h3QvQt1OM
M1uadbvmT33e40qix+GbHrtIzwXYVwCy0EZdTGnvMU/wK0hwDTtgDtodGSzKhHmpJOYbM1EG9RTT
kM+9l4115U2aclKoJUQCpOT3RB+7fC8fWIuFYF0odoBi/Kjk6ZQjp2Xdpa0+Xb6jLqBRc+Nodopd
CL6bbBKzWMCQ+8epXm2uHEtidriSjma2fDtQj0+Klg7LnGhN+5XTM0qBZD++169fH+zsqJzmpY1C
jJ9ONECXeYejzoc9qGbsGRKuk4z+3aVoiSoMxTAnN8pr0W6Oucf7j4B4Q09tFQHKB5cc7T4hZPiB
1f48uYY2Q+zBWgSwRo4zIJJx2UjgrVgOc5pOeTezDEGecJhe8r5zxk69Ib2Rcb796ueBF/7VKVQD
knS3UTs6G4UZ+crsVKju7OYTr2Sfax0fZ7NZpaAKXR6nLMfUPw3ztZ+kbYkpp1RIOTOyfACH8yGj
yZ5zE2CJD3n8uGKsqbOz4D2s+NWnvTe1HgwTeOh2JZ+rRqGoig7gOPOEkVW/mxVhKxqDTYxqwc1f
VxJFPNt/ykC4e7kiQUdGd1VUzKsz8xvqlsqATudLBb9kCWEnSVJyxSzk44nykBKqBLsB5PH4ddd7
zqDnTUF0MuxjBkm2SneMOEaqlXw8XCIHwft+4DMx8L6+pRDAlNqDUlcyYVWYyoGUFOq6RhVNEzlv
mcO4MIg9/ZaCQ4X/Kzuw+g8yAWGlmB7qIkjuJxBj9lKRmNhCGXlTP/Umd0lRIiUAbiHvpvNIOb2e
tXsTsrscmhsaZxWJbazc3AphbK80G7DL/7tQRkSEblho4X/Wti4t32apCRVeoENS33znfKyJa5a3
EbiKyqVzGBHAwn0CjFUVyDvkVl78mPrU20SssNnv/tYXvvA5RWwgg4aeqlKIzV4fFFJ65lMaNwEs
qyYvz4GPBikcm2ZIdDChIX1CNwaW8hADvaNiDkxbMyrFnosQX645xxYWT/8sVXC1ZJfYQOxGgcMs
H/3oDo0p0IUO5lYu6GTVwT8ppMmC9p3trs6upy+/jb4wTPNCBpr5V3Dsts74M7Cwv+wSxbECNiub
EUFYfAbYiFj0YX47FFDWVs2rWr6JVL3horgrpUfwH2KuX2fdOJaUIpJazk146AJhwseb+4UAL3/j
pNdGsCCy0tin/2eQExAgrLImqWizWLt/2H86657jmzH3XEbLlscYFa59nii7s584giHrGzL7cSSd
fA7Z8vQOxgk6dgyUbdYsaaNnNpYnuVYWXQeNT8gu2AYx/W9g90QI9yw2PzPQIPLcpnL3ALF4neBi
R3pNkvDlK4JJXrXW2WEcMh0TTUZHgYRr4WXaA8ZXaMFzje4dA6LJ4wsKq5UA9Bk7ne8mx4UiZHWZ
Miz4/hRuXoQXI2YnknG80TxE8ny7YqYU249VTBZyB/tecNoYRX1FlavjQqFqAwQKMQ57QeQEUei7
EkCS5CbqpHzsYEA1lo/SV0UwRpkpSv/n1nCV48RrLlhTzoJt8BFSg0nMdcm6Ec9KfhCQHfVhZAsy
GxWdCMMoEaoxT+s+4JlUj8jjLrsWdb81x2TJ/VxMocNid/UDroFXH5etc9OJ9Jqhbgo4XiFI9pI0
G8uXWQ0vdH72sfoADB9LG8rHTbpARxIm8po1oa/v2Q66rN6Uc2IXUhiRsPu8Sxg9c0Mtd52OkhR3
zcY0sbG7sr3pvLWAWj5EuLwE5AcUPY5iRNIc2mcqQWuvvq0zwJuqy+lag04/i/FYdrHNY64Cfg/8
+Sc/NW1hD0v1ZiYKw/DdJWAhBAUUtfz3BX67Xm4Jwo5HzBwOKn40Fy/xKiFXeHtuQ4cvOV29onJV
DEMAMljG6ffq/cBgDebzje5Ia3I0EET81L1D91P+//eNu21/45dk625Eh7trQ+9k3Dxa1wxBi0C2
BV2fkutjSX6u4/f9jSGB0SS8HCO7IzNhAA6S4l4YgmS9Y3z4Keps5/ATULpp3mFAi3YgPd8sdCrz
IldheyjrO3XRV7Tv4l/zVuocLWkUr1jq0xIGcCOUG4SzrLVrd6q9dqAKtQiyaNwyoW832CURMRgH
7yo1Wn/8jHtR9+oWhCVGFDq/uCTYi+IcsBvsk/m40VYnWUWM4kZPwhKysFPinqwNPxWSmippv317
vCKDG7kQTk0chWCZ4VUHzV59LKioQ2DILz1Rv6ZMvSWMfAGllFVj+8+vLKEZWqjUWmOjzvoueBeH
pdMjWjvHarRgvHAapS7QBn41tQIGKIm0IQON/iG1moB/9TuRaGGIl440GXlEXCKJTQNAsHRt2KXM
4uVzCqWvGVRUCPOROD/qA6L+SiRezen/82hcT598k4IUmyooV9y690zu2xtrC1C5/azwWuvMrjNp
GfXGcoSggqbDYz02YKcPY90HNq272ryz8YCfPAoAVNfSYeKxwP9lCXJsI79K7QRkZeDaCAc3lAj+
Ah+7cZaP7pVGJ+mU5K1wJOyr16eGSmGhPlS+Pkov8i0nABTu3NoDTtcgtNpVOE3hH7zlZUk8BTH2
pxtXTNuuR6j66rh7DGdorCu/gXIv/Xq1hhzNGbY44hXltrVe/kvpGd/mhtEpv6K9oj7JJPdrMtRo
oxaUWrMrO2vNlJLG8bllFBLKnc15dAX8RHlKV/TUmSayCPvRAkG96zZM6SS/ZZ3cODvSrh231sYi
eBFITRBKGjkA7fiysD/XlZoFc+5pP8W0KyMnnpyk9/5gfHje0mP3bd7AI9Hf4mmcDWYuekbf0MhA
HXRvkNPO0yPvMaNp0puNEJzK+nUg8B4uDp0dDDcJt44B3PYEKGRFcYzcVXuzHdRUz+vaRSCnThHb
2flb9Fw9IcyyWlDxOze1OcMIaJam1UKph8JdEawJjRGi5q4dy8x+S/vB6/2Yt+MmAPhd3IG40iN8
HxIdRQxxBdrfKDZyK3yoX9UTX3FPzJ4vlSrt8amU6D/LgFaMtwQwBXDIG3sGDpjuk6FvCAvUBN6X
GCZCC/jJ1/70DgJV/xQvkJ25gNgnMPT3bvHMUSDEHudg4Wl8S84fmkfPswZQm/YW5IvX/02YIx5u
k7UXdzBIpE472DvwaesMqPUTimk4r6Px0fi3nPYYcBjdqyEXouNb060tmoscDdr+DA59pYsy0Qv1
bBiq7CpwqgwckzZ2nbYlSA63eBY7TC3NERsWoRMD6pXPpFf9YUAf7dYLibPW1SKN+6O67+9RwL7y
A9+v4sat5A5UDzsZLpYRSx1rFI+FjCcZDRUgsgOyTUAKnPUlZBdjpsR5ZkQ7U0cQVfnbwxalsM50
KKqHgEVoBAwZlDAygf53aeNjgd+Iw976VWZYOSZprfvxwkQ4LJQ8wDh97TPaG4Py8XSOqa9SbwiM
an/l3utUC1H3ja2p6B3bFPjsxJFVsoluTA2gYw9qA8c5TZpkUkEQd2tbUfxX4CJuF+S7+Kh1sYJv
oFl9Jfygqri/9BtRRNWKxxKVWoiuBruf/YivVXM9/qHE5pNHEQt1qsLwkeDWQjCVbRN6R/h+A7EG
+/WjhVVJBYoeWY2OyW7uoxtCDVOOpcY3zQF5p0ZFtkN1LwgiGKngl3GSn1A5xLvzevAhOU0EH8sm
O+Dtv9vzAyvtxPBaDvKAw9VsV7CfsxwyS7eLzdO7EJSqrYwF+qKV7kFLjvq6T5ClNTNHOyymwjOU
iOY8RreYwZQWjpblxXQ8TcEcFUY36XAgos6Wnk3qhjZZPWPN4dtBT92eo+/8JkQicebP+VQ/6kg0
pVnWYnrVzvkcbQ+4fM1VegRqmef2QYD+dSeETq6TCs0CvAjJyUq0i6J5gYbtOR4NaO0nN2tY6MDl
xkkD6ctpM+D9neVDNlXF2tRVU7KxEnxnwIgAeKFflZj6Jo6RdgCQQRTHS+Tp/5J1sFoF21PdiFzl
KqGahwUaDJMZctKQ/nSYH8OCAq8PXWZkl12n7hIP291X9iP3ZY3xbKRo9d9qCOJPMXcosgcUO/jC
oKz+KbutSiODxBtDv/F0Bhk4NeWTMAA+QgwF3kzYee0YnD/DZQ3Dzc5GzOqBx1wNtzU6tBIjjCMj
NBynzNeAwicSZI2ogX1T43l21u6nia0b8E5TyMouu0x1z0O2baLFjqVHcUGzH2T2/jN4oyVJEVFT
RsyQqLUFE/A/BwXyRnSHEygZnpl2kU6IdR+00iK+xNtSIeiznIVOv5bgNeQ/IIBGqLHZIdDUzswE
4/11H5mv5Yd9TwrBMA0lADzDePdvNFoBKsyRf/FoddtqHk6WZNL3bqvlUZ/LAs3n8rne72L/XMjp
Oh81YasDDqSVT8JoiM09rHInZKjWFeZ2rCWUINVp3hsSFN994QOp8ufBkcdTrND1lucCiUsS4d0e
fDTTC9do4ErCxZhOCehXxOo9yoMluqHlVXdWAIFfixchCwBtszTqiEP5EFwrBfVvsS4WFegOAvs4
KQPjj2lzYv66n/AtWsonQfwfihwVWru7sMc7q6aueVM7LFe3nHES+Oz5PCFpdJsIPGUFV95GWMGP
dysvf3oOgQGDujIbvP8lkRLcQGVGJIY6A7srVhsvEszz1iYweIfC7KfGcWvA6QaSY8Kvf+n3iI4H
zcmoS5NY27eKEQVUzXVwWbB9mRtTtfQozNzfX/PSxopnFYGO3xoREC2YAI9obM3hM/gc4wOA5JFA
fjp/BEHpHk0dQO8RjnQ4XptO3Lt88vdYzrxOJaAoUuaTtk3mPihZ446cOGMy9QW1XMTiRQULBXyv
AjBxBxQ3L4JQyEYGhOpj+7WOGuGKrEkZlDLptvalzomqEcEolTKFZGXyzhy5ZTgK09eFCRMyVXqz
J12gRVf87eW/Pez1RlF37wg+vfLlNMoZ4Mh7xiKvV126rUDCUg9YoZTnyffQwh1UAtIByIKbKLXy
g7u0qafzcWVm3PMvDAW4zUzlVib0I3E/f6U072mUqlH8bJCJOPnzdS5KxAlIGOvt2zBSf/QKQeES
IFIw0YX8f3zWHP1Z6GiWPRFjWmmEk1zvCh86nh9Bpivn/xtQOjLNMjO5S193tgTV6mjj3c7DI0HN
ve2wrdxPgrdfqnGTSgXa31ixLVfVMt0W+I/FPcJcnQNDsMru8QxJY9By0UZNhq+Cq0iYzPS1+K5y
53t3q2XkojU4jhLn9o8OZKhPHszE5Rke1SpQlFH8xraVjbD8F6eRaq8T5+f2ScVuqBgQNtHvOCZr
zW3CPZg9/ReFBpQ4RnkGWbQrmDWQUZuBDKfs3sIUWT9XGwgCw8b7il/BoxvrlmnBKGjuvZT8kpeB
txGJq8y7u9MxA93jKb2t2tDkipzRZb7g8pN2DqY0t7vU1kKQwOO+CbNbG/AXJmLE5qWiLDSuCIux
+TQaALQ1JdWMEUTQnbEHwMT5M1RxspvHURuU7js52WXI8Q0bJA4uY3OTmJesHCHcoqz+IKxHeNwl
NYpVDnH3hINt9AW8y58JZAivDgSHuf+Zp89nkdsWe/OtKpwK4wVpwHepAM3rjEdW6RyYPPZntU34
bO9tRjbjvNYBajX2W1RZvgwyBzYrUrW1SkL48cOlXjDQLQmVlQCpqKY0c73oppAJNi9uzeK9MTyN
m1iRdAA8NG7Qo5Nd7JQ6gukmR/IOAXE7TQZzkonoPuuzvDJcoLb0S1HmgJnCWvDsI/NLSUTw5Iuo
flS85mGPIaWxMcYqJPnLNngDOqttM1ezIWm9KHpc2xsQfJvEg0zpvvWNZJf2XG3Ck9m4tadi4cC8
3gTguHdf/VNf+D9QF0TTIXYkAavy8oUP5z2ee5nAx7V4zlWANfdpJrgqZboAoHyEsZQdfg1bqbq6
MRGJb+k4b3mlRCEJ4+gFUgZL/NCkkm8s5aMBBh13OssFfO8N+ZfWrTcUUtfNw+3RzH1ga/7AP7zh
2NkyndafEU+xfydfPcNpQ08gVun9/awzqbacDztIRZfMJwECuMO8YGRWOS3fFaTKGnPZ/+SF/a4l
8sxP4M/oFovC5qRy49HwsoJpXgaUBpDJph49Asa1gp5bLhilPgA3yivZ5/JMUB005JBL3j0T6Hab
YoYe4MTYJi7V2JjISwIWOjz/TN3pyjx2785kKI/wdSysg2RT/yFV1dM/2Pmdiqkdw+K29HJx8Seo
zCpetZwquziYa5dbF+VAWip9Re96A/cOPjX+/IlHmHkRN8y6YCPoMMCNKHXWdW0/3OMJHwRjmPoD
6QtpyJFo0WWh03fKPx/taBGUhoDTNoDA2qRYZdv4lgp7q42StCGChHJlimXCeapnIchG4ctBOmQy
xDCOb/iVJ319ujOx9yUAern54vWYw3EH9u4OWaFnr6zXB4B8rbfmhWJKqbMXBm2O7GOPUt8+X/M+
ZwR2hUDfOUV4PIZNphPqGmTRqJ3nmLdXrd6y1iJoG0g7JTCkUo1A7sjKWvBTSG/ZHdrVMKlQeewA
4M0cBlJYZfD7km82Kzxwv40NmW1qF0j2Yq2eFy/1whoK2+NoYC1Yp45ETkqrn7Hcs9KIAeRzJydy
NXSlhwZ8DJ/eY321+Oq0nHWTxY7cEjNf4jopWQ4qOFSZtBwh+3OeicZTMiXy60qzHWhclCfe0Oe9
/ZxZmB9o4kUsVXySLmbQz8Kf222BQP6KIKDSukVul1J9kFqMFVkwNzCxA/D/CYQyE3vIs7TdIset
sDiwyRMutH+os9Ku+yjt4D9P9ciDJhfEe73nr7irfhCtRcnOg9OmHP61y958pEbRTD9y5kqgz497
B0IYTazJY2/7R5FhufODBd+dHhvwCW6MGuZl6LocjlDSO1n6YF2ekSUBlwMwhFiiTgO3Ap+POLoh
0C6MHAH//rp9RHxBDWOBCQcIRXIF6hFRmQwOoDrqh7rWUdyA7QePz0Gwp1SsrD3FUn7oGXjMrI8i
ZD/GSjRmY601ASua3BiqSfcdfYOPnQGxRW4ebvF42gsQPvwwI7hZcjV0Cmq2ERyl3tSbWTIAELeg
SnXVhDUnJAIJtI3VyJi8B+ORCnuceTW9eAxK37bEvxBieMfZkZWfUq08tXj9NmL9Rm6StPvDfQGB
ge3NnpEqC3l/jIlv2eBz83BaIX0jYfBQu0Tm8EbGVAuSfwUERMyfC6dggP7h0S9At+6S8RDv9xFq
WZ+oqkB9auxkdDXkEls4DY7+wrzqLzFsZSdAIHUxczxlG5M/DFcGTwqlVZBsZp+3r9J1tyw3NjwH
cXnD5hqDHBMazSSISAfkqgdDkarxskimqRd5byQKnVFDAiz5VLdsN1HqZ89BjiKY9k3gzal7OKVN
jg3hhO59X0PZexdjS7XBpXHcmgjaZFgMriiBh2HXSb3bqDVv0BVCyESIAB/Ird4RDxxJsQIFWroc
OfjfWHk8VjZOVsLFsoOBx1MRtt4059P+leiTLnoouCjfr6EW/jTcsfATNHSbmE6XWDEoI+rdki2g
zZeGLBymRoQGstTfX7QbfFgbbXDy6coWamqxy5OAv6LbdeUqAnJFnVDQqCQt0/mFRv1NxJZnYTOx
wmZkJC/ToOkZDiRjXy22dsaFpiextnsJy1TgMhNNBlugvSAlOrdAbCRIA1KDo66tZvFDaGgA2vDh
8UxKidxgCKGJumg4Ki25g89whBkI0iEAJBahztedY6qe/OGgQjhvDoTReT4boLDald6iWPRGgpR8
5l8zFwa1o+NxUnfoQAptuchb/2puwDjoEKTfqDtGptQWuwA8X6Wq7wsyIr79ArqOmfeMbmBOIgIM
W0p3puifne3Ob86qxaJ/Zdpg9XAQ5ByM/fqNPy/mCHrOBHuVz527THJsL76GzzdrTYruC+aN98W0
hDujJioBMvdsCvn0Pj1YBV5LzZ4LrA0PHQfqjcuf6nSmfYAM7uq5H5g8qI+FdTxYIn6j/lQ3zfuD
E0hVqAKendSztn9JeM8w3scqGGWYLsqneYP+Wy6vsURFvAM0FKbKpyeKyINryKRcmy6B7/Eq++x4
4cQBHiiMfAbKLGibae34VaGmq0HGWVYZ6eFy4mkrXiLndUDlv4uIjf9uPpbYaVgoC+8NzY8XMTwW
Ss6dTSTj7LQnuHUQ9+sn5qdlJcOyZZAc//dHc5fyTA79Mq5wpCIqhoPBkUtecN0dwqoGo6qQLTCz
TzYSbECVcKQIjKVifsX8t/HFSizZhZ/vmTkhzfajLF252X7+yq2ywpjF9VJ6j8VD7RkqmrurqM53
9G8/76BIgxuPdC9CrP0IM8qYLtZLM/cxcRIuRvSw7xASvuLu3Pi9JO9V7CYwg52xpF7SDpVcdnOQ
wowEPqLX8YU5nKEtLxZe2NBchPvTuqZahoOl2zsvoXAniOoaZSBOQdMoR02VAetIUAnlx56fFb8h
kxCgrG9kxTuc4RLUkOaPfZ4AxAh6EFgosSGX7cQFmqSj33bcLs6zHx/Eq2NeWY7eq89jhl1r9hLf
f9TorZhwq7XCI6rJAo06DJkFBUAzQNF8ZKTzL90kTRJmu4ViZejsMq9ZELqjiARx58Zc+i8AHcg1
u+42dY09ros1V55UG10OZ4nrUkXM3dnszYaXNIPnhMdH4nzb8bHCjBMZGgAPyzlgKIeOZhvOfl/v
txdUnib33BJHLNMrPTUJQ2XedeSQou6s4bY0DeaXjbv95IACrjrMRLoMdrDcWC/Kuv9nYIm0bTVR
0jhvrSR3WgUpLM7sxpRXKUZkeuB0IfVtFZobSRkm3h9sQWK9dOgFqc8VyMWcQ/OE3lis9VITowLA
/BWCKk4hIqxZOmf74iRpdNm0bO4oqT5JI5u8DLsqIbZinFtDO5tV3Y3CTE2y96QvOcUua95cMnOE
pAbz6AZGnfzWt8szVNYz9TPjZU544p4ZPlcYejvZamKlq9xXlvFc7kyZMJ8yK1CPajrtEoQQMFTB
GHIOhrbcnHf3y9kYi5TG3FNlHy+0kDeGQXpDQVu6DDLRpSF13fcR2hIX7IRyMxSfyeySaYM56sm/
3d4lk67JgdTM5duGbgMuIJIS2iVAS3J63DbKXFwxyZ+lypR+s6N32NcTYagLssUtZY4pKkAdf9Fk
OuDeX62z4ebUrqEtbUGm9NfAazGMCC8zuhBAl458bUFuP9Sr+tdM0Ja2HRoE9fmA1FFG8D0fjRnt
EkHXJJxUWtErV56zUrOglH7fTONdN21FFbiYVpGErSV6Wtf2T8+JS+oG2cJLYXK0U5f8bN4bkEhv
zejk9NqUq0jSCzcyXce/Iy7eQV/BPsSBpi8nSEXaaFcOLTm9ZYs5fTWN7a7ZX83xmyfGHWOsoQWo
BfMynC9BMr4PCKmY3c5w6IU9NbhPPl3926kOvWul3/dr0GDHWBRS2huh57QHKisJ1Ihxu1+Jo3YA
B3CWoG01W3qLzI539mOQOqFSYCX0nvxkC/wkEKRNHAI1iDk7x0aGeehwjLMgcSpoj03pKA8fCAuO
Et4YZzkq0jQWz4wqdkQEYHTKJrGvyeVla8oKQ0ot3Q1WgYSLB6tOFdzeXSYVuDLFAgy/qalGU+HV
smAWXfRtTPRQUEXhApN+Q07iT4vz+iWMIi5DeJ2d8X9B3G1NDttN79/E3+4Jja6/uYo+otWnL7+u
LrJmS+J5AEVSfTm2w7dJZmf/fbjWLXFh0HfriDEUITX7SLU4ijlxPcvsm+ny+eVOpQ+AtLBD6Sz0
nIUPcHCaYWsevTJSG4DWSrSwvluFvb3O/JM6ydzpmHrQf12tlhDHoP18rf3P94feXTunkvx34Xz7
Ed9FxFUWT+y6FTiL8EmujRIglCRpUih5cV1sBdWnI3jYHCw2R80V9sCfMYacZLKEgCyWZ9BeFpHb
NPsBwcoAzF41M8ZOaqGrs9lukIOuIUzbST5UgC9J1BZzU9LGHii6h9xJuP3uWOXpttV5W/AVHlby
PW9dDaC5VfgpJxXVg3cc8AciHUEFn+W+6nHrmtRNZ6JiP4fzq1SZTtE1N2/euTJz1EcXC4EXXaTc
YIabTSlyqwlexKQ1s0lwU0nBxwPuKvy8KiHL3XmpN4B6Ps8Dc4XhzzCbqzffV90MGsi9YZ4/ynaL
qQxFzHiGK0/QY+jSwVh3Y4iaSZx2iZHhL6eA4MfGpttUQ1OHHas1ia2xdwuH8xCXBrlDD19yu7g+
TW0SPGm9FB0BSGiKA+/8RFbJgecNbVvbl1XXuS6NL7sEp9nwgAiOISjidnSrAiJCSoo7bUw+WxuE
o/32YE27Luf94mQwT6glkh9PLigspwSkxSJtf76Bx0ef0OARe2PO+LByurTKOecTcAd6l69aw0JS
FT+Jh/Qsv+E2sFTAYnJzuSf6MGvEjrfIZFraRDuhUFahGE8dUqhAnJ9SlGhd4qXY6/SnFjpsnHLc
+ypSIjk6VnMRLrlhIk7fSs+vgojOxNcMNIdaJw2NLbtCNWsoH6RMxL1xTD62TzS/tbih5V5qonnL
vFzzjwMI5mnaDclnQecG3ToRYI76zndt6GgcJ6qOJ0ITfxl2RpE1qkH/cxfUVkD6RaWKM20TTFVD
3scz/Sr0JNAR0WBIGfXr0IAD8+7xKzmcOj3j5yzaHlPyWoLc4p1QV1BPRspoU/+CWvwqjBOr4aV6
OcpnMIgMNACNG/9RIxnpx62FeKAGNaPSfGnecj3n9B/lPCXffYginB87Eicwu/fY7wuB7JRj3fsk
2o9KUL01XCzqsix/nPy0tvrCu7C2Yyp/RpaIzPgxSylMjx2uZ6JAm4aBwiUMG0Tc+YYLuS/dPNde
ADw8k3PZoeGyuxB4nQMjSWa4QHI0ndAHCP/lDLbDkY7Rb5sIQ9h/+DdJnI9niQY4LxUmyYee0DAW
bV9Nd7lYhyRZfUPYFjc5dT2FCTh5VYwad2+dx54KMw/3CBy+2hVSfiqockx4heCLRS1DPK7irmPG
rbU4BYUZZvxDJGlv+MoL+yMfgFKeW51YOZfTRi8//oh7QDgLUbattwCt/73YrtiwZI/xj0W41KIP
DxcyiQX4bGJU5eoc2i2t4aUkPAvhH8bT2xVnwzy4lCyFq4rcQlhksn5pdefDd9S2vuzWvdOfA7zG
rX3B2vMQeZivuAHiUQKSOjHdSfU6EIMy6XcQqmOpfW32vV82gi8DIlFXgGxZC3xpMtVXPapUbTlr
flWI4TMEwL9fhKFrhRI0DpOMi1ywEBG1u5UTpWfnh6VP0h+Xpy6fGEs+K4IUxy9RhbohT5492GCl
6NPM4Mz9XvDKqUbFZGEvupi9e7f6p36q4y3+ZH5/rJv54zIZJ2uShau3tqU9SHmi8aoYEerzjPJt
066jJMINGDzKgE5jq+QlcSTBvfR9TeHwEBtYofKeHYNomjzm5FUyxA/0udWwQk8lSfFBjs2eTcnB
OkcI1u+cyHpv0YNS+Xw3Hzy/QxPBRh++7QANYFnzVTEf4hRK/EyMezQdYmnNhRbvVZDWIMQcFAvM
9ToxxeMnVzxCN0SS/vbZaHpzRaEmc3skR1s3gtwfu+AD5MvJHKc7+J04T3tyr1Orb5XGivtsuzME
cjYyKNyd2eLk4g3KEK3lvuApOFIcHm49lsuFwR8ZeyOpwnVd0qpDLnjgjyl0cxATYnTFR5TipkJA
qIHbFNDDX5l4HaVGabaBWZ4Pzm2nzUDKeYx9BiSUk36pLcGP4f5r5zmc3LJ1AlmjxOSyB9CQ599c
CkjHr6xGL5IOLEnvwH/mPDc7vtSEpljhl6m8mO/JJN+EXktGrmIN26leybNwOT5yLQEUGqxoQ6dh
Fq3MhWpQVTnDH5RvyFtloO/Jzs0MTjis32UYbjez1hqQJ1c3yvFyjSLGTE5ypzFjEpS/mvvdSosL
l8kIaQedIopw6ELT4KRnTL2NABots/RjwfmMDx0MiAGcV4mCEgvqHdR+QwnAwMXDjOXsSPxqNsiw
qXN5tcGflieCn5eY2L1EnrO69aXwUG1aKW+EAWxOi91JgO3UVs+Vsqa1o7DXwkF9xdb5dM9lGdeQ
U8mqtSaUIdFg/a+n5hUu/NjnqBc2edMbngSmmOf+o1RdeAIlHtD4qyREdkohUYKnaYIBpJzWqmmJ
4z5OrP7rZcRur0Z7moYL935vhaLFDHytgSQ4ECztxpD+ggbQD1VXqlph6gokfggqEKlqiEsTPAlE
wLTs+GAbOYxgz4s69oQvY9FY5tygVafeznmoBFQfUVebVotnHCFDFhE30lvSc/gdCTYG++mecEfq
PXxjOek7bwC710WlKZ9NH2eX12c8SnB5qIocEtuu3nKAW4EJQE89ZT2PnAtzOJhOEvlsZ1GM+dNd
TlhIMGYVl7LDOF0YykZ4IsEALb4WHp45QoPu0UOFNxvTtZIX18JzmGpIRbTvWz+17y5tOM6i2p51
hX7fHJVqG5KZ4E/hP/4spII8IGl0yLO6zFqNt69FnVao9fant0fxLMySimk60wD20awfJXPXb6Tc
/lhwaYN2IrDUJjGQI3fDi/CZTNN8yELPlPc/gO5JKtkn5MZIEBqolCrGqWysxE5lwSazvc7/Q4Oj
cDFOvwmooYeaYQBle2shaG0K/tv0pfafhtGvaoGOmSTYmPJO7/xFcAbvGTN2/euB6dKR+PQ28sK3
mnXcaTlbgTcwmCCQaJB835mR3DJpRpUHdIA1J+MZaYmjdiWzrtgwcj87R22ncQrpaaa4s8tkR1E+
2499Olpj1lhwpuCIvJHFYOaEFlapo5k1pqGon9cO3ZG9x616IkDpZtPUmHRzh30d2/jW39IgKwCN
b2htVm3QKUE08Q5mc2gFRVc1DCUh021QRvLVIHzd0s+IhHYIEUDGFlx2cmcrmfcW0YGLWNqOfFXx
zrMtmqdl2QWL99HLTQBUvNqY0oza1zbCpDgTUex+ngSwn3mgbgM0ecY17IK4I2HqGWV4touYcSum
hVjA0wOVIBI5CRqYtjKUqftgl8mu6zpW8ck0DrrdtU//t56mRTeHSJd5vmt7+BDAqhvvVAT5RSK5
TeYVDvQYHlppOWmDzzS4CBlES2/D8w6HQOPKWRRynhBOUTAMnYdKQs6YoJmp1UfFxMFMzd/j89cQ
aVKR+fnJcfbU3s8rFd+Fg4Csb3MI/8/LUbw1bwqarVNpyA/b2cDQesyMIu3bhFl+hwrTfVbKkar3
eBD8+mN7Ci+nYWhdyFzr5rQ/CUW+Z0aQ1Bz4Z3/lQtMNfWDQPZ2CAsa/2yO/zAoABx1e7dNcUsj7
iZ28+5kYYCH/d6Jmmu1CkfLkPjS7HeGVVQIkALfkkIHMIGNMG9pbTTnW9b+HoUSgZXzCA0Dhi92+
diudQGRKWxgzy+0OFigdTWTPJo7hVZcgG6or8FFYb8qUnMYzfOqo7LQWXjZO3Uzp4BORP6U9Mdqw
EtRhJZLJhrz683deSRKLGv9TaWRSA8DuRjsIwjLgCtHyAVXe+Pen8xYXqLmnlKRHJ+zQ580xv9w2
lrvl6HBTA4cquBb/pGHKvLo4F+pS4MpNvL3Dvk68hQLx8MYLU3+NBeeo+IOSu/Qrw2uPvqjcsFU3
LwUQmHNsTReUC7SnA3qvOtwuzlctqrWGs5NjfUnB9JUdUMA6V/4aXXY0pNqk5Ky4IVk1joCASPav
jIBOavhTXH1C9StWZKchXmtnOSYS67BF0STd4Ku6wtoHWEsW7n3tT8bVUb5DTkVeRFFTvu2S3pSB
LDlWQi+NILMak1QUxVDvFhet5w3qlA93gWzh6uU1ziFgBWhM42dvttxlQ0994Z0M1xHRyDew7GLy
bBlBpHec+63EEgF8vZ5phNH1RmMBM+TBsMFtFwbbhjqjSaKm4r1IO+AVBLKTNrG+lFzajatkeCQ3
inhVxIz7naEun88KZuIIgQZde+YUBKF4k3PFds43cba4g1j4kGC8C+iBj1vXnHJw1AWdHUxptgTO
M+xLp5Nco4nHBG2XDuamxNCsM262nKscxcVWhXXUcsZF3m5fZLbJqeLJtcVj5iSBZmf0M6w6H/9m
NG261MU2XmpBs8cx/L+w6jHQkez5dabC9/glhgC5Cl0Umev98PI9jM12jx5AW5F7eh5rFzcltWd6
Ns9Ts/bBFCrW4crWl6DUIqx4KFBWfF9s291gvQOx2/L/9F/PSXV8pEI+72M627ZgRwbMp+z6vKBR
nlWO9IW5/jDVdavcqlrui86yaLw3RB5KYewWKrNx/rA1VvOW17pCIH2QaoTUxJHRGKK+1341bzvm
oDJYOe9InnmDRE026m3wmDPnGAfMz6A1xKM3a8X1FwKQGrRgDuM3ZLWgp3uq9ZxwXjHJalXw/ZwR
JgsVLjh+7LU/7WHCsBCpVzq/5rK8LPFfs1nxtzoLe/6HGPEVUg6pDxn7SitlZZUS90bgqy/IbOg3
mi1AScZVHD7g9i1QnsuZwYST1hjH2g/apRH7bEfUP6dc0xyFvYy8g1dVXQ5wLfvLQH8e+zM0cTJb
Nb50SarUVL3vIT0VaQpyZHeXwVJF03nGi/Z/VKVUgAh322sOI9PVYavrrO92IfC5XIePvbnQASiA
gMwn29QbqJtj88cMjzmpgludZTWB21dDC1G/aqxBxmVow//Hem9CPLo/omEqtBHtWl1xlg7q8Uxr
AvwNcipIiqBGSieeR7wuYbiqnvtP3WcQ1Jclc/RZrA8TeDB8/6H98C7EpUPJnrUNJ/QIpMJGDJ92
kYx6GToPIZzlUUe7K3wGP/juI96sCSwzrs3VoP1FlOaiQdq5tYIMDkt/MQVWsfp8RXS98AE3IFDR
UaOmBR5hSLtQcTGrucXiKR5lQYAawNTI0luco+NgLfFPymHzjEp+wrrnyZCZPY2y04kYVqFUbqOl
d2U9irDtWjB2kuZzotrddx0Ao8VdoIel9vLpa/HNqsAR3oa6V0Xi8slz4kKKvSafE+cTSxlfY00m
ozrTTQLIYyMesb7KsWctT4aAqpbEKPKrWnTdckQdZTtiBgiZTOTRKvAtxwyVYD37nWacNfODrlJZ
KMomkMMJsskCxZyWfuAUWD0u3plv5HHtXl3LFuZ75OPG/WebNgGMjbtDnYHbl9cBOo62+6MMA33I
8qYZafHGnzzY2ieuOIjVhCF4/POxtXOMXyVpAYM95p0EibjipsZBGifVETBsugqsHPPSIwamS54G
+Ic3No2psEaQyskvGsy3v6rL/1HndPSwR8gZ2hdcQvS3Iw53m8SUKDm1aCZPiud8OVG1YT+2MLWI
obfLAzlDEaP+AINQd7mlb3U9t6TqiGzut8RQf0sAVvrGh2wcWSbArTR7lmu112v0F+BRyY0YlVIW
OEyle6hyYtaAEtePsH9T+eRYeEDFKB8Ovj4CoPZl97WkqE+GaC3zcjex0JQ2L1puCVAJtnhgv/yH
qa5ShQKZ+2SmL5l+KemtJDJLs5wDHSkf6h/PxjIYWkt5UFY5P7pzlXT/rlZoX8ONKvVYdZjM3GeA
Jkf8/weIvGVRARwxiVSlIvnTmmGms4bX/Iez7MGHxpSR/hXgiVyAb4ct9h12HWxk8Lhp74frArVL
MMAWbn2DR5e3UJue+B8P7aaURLxKl/LuFTQvoIEysCxNFqql09PYklNXKpt1OM7GMCFgPcb3sh8L
hrsujlVPSS1ubtCvnpLqk37rQggKNHTCJZTg75JNPsdJ+L10S0B4B70HhC2ZyyFhXtsWAy9Qdz0+
n8fXa1sj9iHIeA6ZKj7HjDkr9F79oZ+dTzbA1xiFeeM50A7BYzhkXXQPYrODlJhAkJLMoAyEFw5s
Fn4a4CEcu2XMrsAglHczViFYU4Y4gOIlGNW0y2osKM5k9MX5K4jISrHI+wClevl6tGE9JGTBxS/e
ljTy5SQkSipQlJxi1ldM5P1291u7B9QzLpkMR2JzeM9avBYTFSd3axoZwtoODOHJX/4cbl9uPxaz
vPU6MON5sQOZpjnKLANVVNFYO1fkMagQuCK4xe6NYmjE+zckTHF0bTUWiCHiIQqz3pro7yVHwl+C
m7KiewVtA8aQ5ur+kZuPekOtcLQfRPtbJ+d/wB9JsunWz1weOjrm/Vt0MkamR/jnE2h7jZqsa9vl
7XvXDInvhZZvnuOL0PJbxVeT76jRzvkw1LsMgI7JnBP7b8A3Stkw0c8sJUxxPSVMNTmYlXsf/bYY
HS96CwdNpF0HfGS7RStDmTyq625THuvstFXffgJ4zJkfYJjtZwvt/YGGB7a2Mi9naMU2AS+9IQCz
2y/YgtupB907bNVoaEZ4uNZ8gheBnGVQu+EZ05SRIN3jaq0s79E5YwPOxKl/sj4DDF6syQ+vInBB
lIiXMFgrYC+289naB/KGChgrp/RKvPemNMMCL7BvD+yNRS6/4NTEjVl6akTS8dYqd6Tmbuih8YsB
3DCkCEXsELOcjxSEcvL5qDnsfZeFL4eMXDtmj5Ra6DtD0D1KWIaZiF6FQZIFyAp90RoMaJpAxx6H
5ER1wEskxZC6lLhXMJuINBMWdCj6YLoALANs0L/WuCTlpY5vz8MBtN55vzGn5PZ8d4dG7I00SyTp
8GUntciRJ2fpY5bGauieDvvi7HAFv98BWSjdFd/GKtkzDpeCgUCfFgUrbVwufbBSR3FRyrzMK8dY
odWYM2rTyTYx/75et3hb0wf+NPAe5AmneBCjGORxo8zSQQwiS3E8xP2jsc8iQHANMjC1FnCGdwgp
MSDujI2gf4mRAGt3iPqzHlj0DsLTm3zl3ZZjaTSZydbsCReHgT33HlogbbeaTvJCgaQxuDj8jQ2A
jRdEoIUvgFQA0P8GDgEvjmY7K6annBXOZcy6GBdLPeapoCIbfx43VCk6bFfoQtTIvYUA8quvk+mt
+ZIFVzf7t8Zs/lvU24dOlNIXAytVw6m1+TF0VxJd7T5+wMbRCtjREsKvDJo2TJayz+97rVQ9Kf3B
v4aelzwiauk26sj8tSB0PCAP1ZW7Fee8SP1FuMXKkdT9n2PGAJUIeQLekinWQiij7R+ZUaKuxLAE
175+ag5xcuy/T7GcOOIzO0CbcnaJTRTQmRvPVkwhTfvCihTu44ndhfV0Y4qV+cVlXVf+8Jx5owCJ
iwuFgMmutRTn3bITn8NDBjmzDU/OI/EZZDIXR4wbQdx8YkuimBmkF5IWP3LTX3coNwhv+8g5LCMo
Il9I8+QHMb+MMs/MVlWPcslkcplGv30XicpxPbhrDCUPPqznleQzWKR2ZS0y/4IHcPalfDrg1J9e
iHI3lRdyR/Sda4Y+qtAKCxNC+1pwiCVpbpQataQlOc7Kzm6KH6YsrGi0EAaDQ3Ipy0+fXVk3X1Qx
7/i5pXCnKipUfjvG94odI5dqOZ7/rRlOqsGIleudwxp/x0uAxii/QRnrmpJbfks2nqxXI3zKl2HG
g5NLP7mjkgA/406iTRMqLPAmRf9OmxLK/ZLkfueS2x/gsvGyHlcrTofhHdQMEhRO7tjSWemMlMiW
CXviXCqyOxzZ/oEXkWn3cw4GsIjwh2wszEIf9+o6zkowHRUxDYnl6v3h8iQp2kRI6lRX4M7gmTA6
yyk7LrMGOf6VNccZvg/TqJDSLlw3j3UMSJO0IQrpJIHx8nHW/bNzN8BJWd6R0l6wVDf8mSxPZLmQ
Nf9rveBpqFE4Y+Fh8+UML1QcWudz3gEYpxEq6czmqLFxmQWnvBVIRGwwYl/ksjPaTywm2sHPNtQm
FTDQuv2tIukwrYwoOR0EHpAOwy4lKSZ3kO/3Fpdu056fl+kiPuSrTFdVr/pCxt5guBYCRodffq0z
411/AniafEfbVaHJ3bpWSJdcytAdjKCJDP6RJlS+emBmGUUEb4NQod9kgTH3f/T3XACny5dkUgWP
1I5GyvNsG0oW4tRZ27DahJtd71/n+o8DB3EcxAoYpQN28pfaBx87uDoZaFJMCxZTGHgBKD40PUOl
8MteN21KMfGLt8KfUsO5t6m72GWiBJEU+Y4Np7H+jj0DY2KtDvWzIrXLuIzeGk8pPIo4OgO/v2/t
vRRIuSsH22OHTy471Alo6mSBNcH2o/ANgjOexZpyPV7VIk6637qxCcLzk/rATv5KV+/HG44qgszB
A1MjyUxS9a8gQMrznTg6bPL47o1ma08lUzke+qQahpUAyzUO8rwZ1nYfSsC1rSJ1CzvSUWzOmaNT
avNQ0bMgiEapfXD40YtWHq1q8J8YWgwbEBJi5vLajwk5JE63Ns+mv9yGbBi72ycpUBkUk2hVm46o
tHVGN0LFUdiofJq8FkGOGZfPB9YyP/Se/AMkqntD1A/CgdvUyiGEqxt/Z/aK9o81e1LOuVyV+Iez
JAjXPOLT8nJQZz+PFjv1uwUcyoT1CUrMcaEPXcLgrINDct5eDIvzvx0oYp2dVMLX6DzsaPTL+ori
AoCQqmluR4gnR264QK7oQfCuNBgxjwFxJveWGHZivZ0aOaEFlr52YScqpW8lXKXZ1jyU4GdmxPyz
bbcSSiy6P0e22+fpjA2QlwgDqLH9sNGAH0xQKXFcES1t2bI5ZPVYU5gwNhkQlvaySTY9u62qIumI
gwa07mEaRjZTtR164CyDYsKLFhGR6zPJosPU/cM1SWizXCD2FtgZhjLCYo1UC2aBigbF3egFqpuk
SAuWw01TkkrzaY301+9X7SVJL4n9hN+YT504jnpnX4T5q9Nq8RzCzatrcZl5ByLyaNXafffL0g9t
ENDx9fx+VE4ZS2a8pNjCJFN7ihrGY/yTxei3EqZxYIfhxShU/likT04rOS3VD0OTXFEdHUreZN/q
zNhUisflzlqXGccQ/4hgiumhV2Gql81J0Vy0WhUxM8ihkHYxXn6YqwM1epzeIZTG9sOjaXRBJBP0
6n6fkf/sFZL8V8MW/3ox0RarfAv9cR+ZI9NI9yfyU4/E8BvfW3Zss2vZk4DFZzVmQX082VAgUCPV
cfDO8rLGkR70FPCXuAWggjV1on4rkw8OXBWZT1CNtnLFKG+SEDs8N9WnBLnCtxVy4fob2UlDYOXj
XmiXMOweWo8D1EgZITrhSdEDvA63Ni30/Amfky/Sfgmwd/LoLmWZ18ej47YOlD8a0NkjFQ8rydN1
o22Mt6o4eH4Om0Z2LZv+czP66Xbq4+xCVgZSeiBGYqGt7aspe4PcxmUCe9377PtQPp3nzqd7at4z
FS8kFWhrcKyzhYIvJhcaLwDpWs2goI29OnyXmmF2X9Acl9tf20bjuZEWggaoTSKDQV1SLesOQX26
UQCPCWG9Gc889VwUJFSIf/jUyK4r6xvFeZte3ZDycGBZkS0q8REoeI6JzYKB/l7eAIHzMKQG4Hrd
3Tw8J0hbiQwLGgXyEIVj0fmDybcxw17ROKC7FBzI7GER1tKoZSbPWU6bVAK0PkBKQgbqHIKizJ0G
KSZBGmuIWSeluKSWzIIGiKkX7gem9ehrE/0o3UnIjkOO60Z2nvWPtfhdNp5HIgJrqd8SKL3wgkw4
75NIP9s+jNNEmxhJuuTMDqosTv/Sq6OmJAQp+EB/Cq2FqCiEJH0uvoYt+AYZx+Pao+YzUGnuwcJF
nKx96mf9BJTpPPXCqCU1unOa/7oNb+9E3f2qQ0V7m3Ly6cOAq2qFHIacg2f6ZBLZU6Wy2dUUQ4YW
AmiMCqvfMqN+Vuvza3cQJuonfTNvPhwku+vgWE5nRfjnPpE2aHSkElDg53dkFXC/xQ3qzlbf+G0Z
WC9rErU5MICTUXsv0ZNiwxAH0LIxc39LoNJb45GfmFg0U9RT+u+QvFA/WcjPqw7c7GoQzmFOi/ek
vBYd0HKOYEnoPriNIZdEZCLRK1C9Pd9R3hFGV7J/RF/JpoJNXMe3ostU01r0UucBevdaJKyCLHQ1
Ekdjj0z0tQc1n3jPvaLXLf9vYZHjDOpSPbCgDebYIkPXfl3t71o/OvHADnhhJ8Y+QavByWmQpGaJ
tab79UXc9u4IPsZxbNVfVOj/iOF+4Wfrsf1lKhJGMZ5YPnHAh4X5g5O8re8EcoktZC4iY7/QOF4e
oFuBAdKSWOfTgEQQSN/NbzGwlpL9ZZZv1M6qUYPp4800A/BUT7yken0+kVlReyMFFOk79BGnZ+eD
ci1Qwto2Z3ZqFvzaYJGdi4xx6zd9ZBYBs6cxAY23aODg3rf25SeCL/Jp3dWKpxtxsSHVfiPzhioY
vYPd3SUFPejccRXQqfrlWJjfYxEgPeD73GH27cc2gRusZh8Epy9eT7yEScX0IdDoDif4HMgOX/P7
1gNNuY/VGuql4fDZRBqx04v/knddIO/yvjl3CgvfBwbutVi3i8pj9vtwzFpksbprK00io6hI7w3x
Ncq7nnjHF/i0IIUOazApt0WaBkJREzKRJJ7szF3F/RuxJ2VH9Y47FcBz67fZR9DhiMka5RBT13Br
jkzMgjj3/V0iBjIGihFvGyJGdoyY93jzPvZcYDzifJnV0qww082ONgiP2Kp8hvKqQbXov1E6WxRe
KFeEl1YEXWqjdJRMLXgdlY3ip7mia0cyRNhs1VQmujWi6rRVs5sBSHqlVc8KuW49LrWHe238N2gT
e4LWagO2EzdbQiOOHWnqQJ/SJJbRYDqa87M6vHzBib865h/Tv1woaxz8Uz+iTcZnHyj2wOnAMQ+f
5M5q0jWh0JLNog5K6TeOb9HnncINhdXMK1p9ZU+3ehp1MqySkarBOZSs0NzlKbhJ8ab7LyXX3pVl
bRO2jxh55+vd/pDa0fLJ1Nvkh9XGok0ryTJCcB0P/ABMOMR0aSTeB2J5iIK8fFxS5h43VIUkuhQj
lE4FhRwuKtC5+ZqQkTodSmWp/pErjTD0vO0xc+4FRqnA9jCMS0Qod8MNWu981yuQ/MEwItUfHW2S
3XxjoOiDB5B8+gi1a2Xmg08aYoyklysIK6C3y1rV1peng3DTfpvUqmoLGTX4qTxKeRprv5lv4OH1
Aw8tJjQDTDsl8lCll8RcpSCtOC2NRxQD3m7N2E7r4+6plU3by+1rAR6/oIWZnVVONYR3TaPXYI3p
33UYMtcG27guqoD4HSF0Pi2iSbq8QMIUP963mNAWW0MTVx0rgWCvj6O1HcbZTABR7zrW8kEW4m0b
uPE1/WLtc1idQaDlfouXk2jO4tLXl9xndLGYpPC15xAHNVZlI+ggjs1f3+FT1ZPNhzsh1fkQ0yz8
Q+TH3c2qezQZOqAzDm41PxTpGQPKNpKSUZMVLYgCoXCEiSXk7SPE8vg+Gy4BE2vISfo8dUnaUTp9
nm3JV6vNx/Fc5eiSh8c6FICpx1lhMLnXoSSyMKYd6IZcv/OeG/HEr/Kezy1BRspSvdGaiRRpEQZ8
981EkrVCILHhMFgF0yzkntwxfuPdaa1oIEpm0F3vy7F73E8RjfexIyZRq9vfXlobDAKg0lv7djDl
MR3/mijEPf3S1qz7BHxBXJhQ8CF1Uc5dSxa1oT36zpr4c+9R5JUWRdwtAM4KnJdStpLZ96tPyT1y
E+xijdT/CnIOMf/riqGf/mJXeSJkyHXn10qDj0VDhSiE9KsymYlISqY8djF1YbBrJwq6rB0gMKhX
UN2a/D+zB7ofXlrpKhWDGF6Jc3SvC/HWDOa8WR3K7HhFLeXfehHwNhkQy8HmYeq9Qgx9f8Nhn1T6
gY+Mq/qOVafq0ucOcQjrDjgPYQywX5HZSInuXbbTXFzlEAyVejBfYRF4XQKfyjdUNH1UFESqZ+ID
9U/w2KSbh6feLTkxppX5eBhBzmFn+9ZCQwmGwP3MtT94IsWd5SiemfbvISkQvRQ+DHBhbn4zHf50
An6wGlC6R5Q68Al6nss7nJZzUbo0OaZAqi4pEMC2rMk0xHLbVjjq/U6xAN7y1BG/BXrp8rd2DPlK
kEQpNOlk1YEfJVxpftDVFlKqkjO6PXwBaiEaFQ88JJBVsen3+rDridLkhWkU0xKlSid6Ru+rK54b
qQBNUoGuXpjLv/ql3pLAbwP4op2AJOBwGwE0GBL6cuuPe4C4uI+1Nq4R70P5skEnrTfA1b7kxrCc
cNSqbu18CB92+Ix99ILTQ7FRNlkMZXpzw5C+Bomn8NasFe6Q30C8Po4pHBxL2XiHVkSItEUhtZbQ
/LxnW7j/I1j2BPmCoey1k8lr8sgz5XShHmawxu99UW+d9gk3ETdbP891gNXZ/jeuPwtW+62hb9y2
Khf472RaOIt68JBT/yVAi/B7iN75pLV7qGGtYQoomOKhF2zAq/DQGy3xZf+yuI+iwM5DlZwfDZIh
7+nB5Lcssnf/8jMAlkJ3lenhxozywcfNuNzdEfA3lg26eu671QRVlaDuGN2Xa6Wbs90HAbq98/9q
dSiNZmhTO27hyHsjLswvlzsFlP6jTo5w2xszam56Vx05tqp15tuSJdzriRq9GeLIoN4PsHumkjN3
pT+tEx+iqOigyEba+ODcYrZM2bs5jkgPzm1WETwcqZWG6XV8GDFHXShvQB7ttZ+A6edP/eAhOeoo
eVttq0X/QMGtjR7viRtkp2a2vqemRL+c8DEa0I+tiRkcifo5GU272bqpEhc1v9lWZPIoEdX00V76
xb6u2gm2NahshN+DTXwdNbdGud16f6DF82Ix9g13rKdSur+O+OgR17WjpTjXLiRBiqQrADukt7fm
We1Zd/+zAZkhXrmDe/YEOBpngpqrX+tWzglkuGUdTsCeCSWHBsh/dZiIcZ6YDjATQz5k5qqYJAIj
7bVWY/Sa+vo5Fo1owve+dmnL5k0TBMKpsNiXeNNlbbCrWs6zY5f87hM59TUB8bNLZT5wxN5z5OKN
42ZKV9Y5HsLI0Hst/42CxcoMcYz1xIZL/Zzoe4aP6zTswW4r5rnS9iiwYJ9GRz0e0pNHgugPFNyI
GSBdwrXY0D3mhXmoUYHhCsi5VmyB/QL/aBAsctkg5Iqv63NVpdwgcfjinu+74ydtdv2jVpN28IUS
XkPh5S9CwVrCPm/EBVs2e6WyNc/mJjaHitNfVmQk+Dl5UD3t96EZd/aGN7xkPchYYyBNjXpFEUw1
Yq2ZKeEBHsjnIgaAwE8medm7DQ9WfRLUo1brKO4e5UHvdoATUjyexCk0zcpQc3ON41652lhpyGht
n/GV/KzynmMuFvtLKHlE+dsJ/Rove35cXqj8wV5jY/f4esPGXzv2hjFZAqOzUNO+WOTkGB8/AVNe
TZ8M+EivBmNs+B7XChbRPdUpxVBJcjyWpPWJ1qMci/cVQvABjA6tk1+UGYjtfxJwvrlz/Fpks5HW
rgK6SwtzWtSTIMWIF4y5GmVgkiJF8dqPfuUwHKY0Y0Smf1Z4uw1BonC4oyqUW9ZXofYwejTe6VKT
a16tJusHfiaBXnCpqS0/6MllNrhkYZlTmpGBZAUTv3X8l+7PuzdKO5EzuWnl4XtPX6G70uzI5POg
LbVxaAz9ngKe/I+ncwJf+FWi6LmPz8A22o+UMHTADMAeFMQ0pMKpzIBMRu+rq1ziaWgPrzpWM4KH
med9EEzKJpPq2x0QTzNDksNEOQBln4E11fxWvK7lJF992pIOdvfj4Th3CtsJ4owg1J4lfF0KqKlP
T+lhygii3GxFXODSyedrQPSCIMydXjdWBM+08G1DP6n7TefOlxIiH1p8PuYcjzQ96ylD6Y5Mk/JX
ZfvKiBphSE7B91uXl/FSfgGcQ0GoDAgKlhdaRzk0DA4SCl0H0ziDigNN2D9VQoRlkKvS3QEQ2OoA
FYJIXi4dlzX5hHamhiaROa7ygzoU6a3CwhBpNzbD2s7PzdoDbcRf/NypuuAPLhgChHmCCMskv4/f
bD3qw6rm58kLmfTBe2AiIJrIxQUusHYoYQOEO/BtNDE5YVJN2LVOah40xWBpA9htppC7LH67nOOc
Ygu/w6aeBJGNjsxJvNMmwdCOBCR7mF4lcArUOxVNLJlcro6exz8TAZtQfy3SJ4VdlfoFkevzdtvX
4PnOG8B327/vAkcLLlP8mxBbDReUMZMFShJSgDnIhdgUSojE1uiW1yVtoDcz9zBIerE+7cLJ+8UO
tn0/Y5nm7xmGs+2YnEIBH7wSACnmJLWUCvEJeXLWcd3vCRSHTUwOtr8nBW1e32kZW0VURpeWDMW0
bgmkikilMYnLt4Wq5rNM0nlBBsnggOu2NtG6pn4twJvIvh3BwfhS5LyrBhCWUu5h9bQ8Hnlmj1pp
YAKMirEb0F8Fnod0Jk2xwUvIqGBJ4aA77uv5rGN2qy96mr135hrNOJejBCLqLpBL+ATNMKpyMgIK
aWjJbcnpqV4K2oTVOGq4tZyQczSfFuThC/ccCiSsoG7bbz/hxJSr8GX3Oxl8VTGHSd7RcBGu/TBC
ne4MwLLHkxOpxxQRHG2Nuh+tAhNu09UIkYsZyeR4iYz9uSSV3MOwxqcN75VKmF39L0CqfFaUd8D+
fFtgyD1TR9bRnBwSl6V2cXlmwhAUO4a1LSfzLURIAsE578FENmdRq0Sv1+C405wR2UKa4cn3Vcds
p+nmyuXYB6r7dkx8vo/4tEtmZ05INLCyKsqmB/O67D5x8cCGJkC9XxvljflD8+Ok1AucHX8k0ZXn
mZXZKv5VmQFlsI4pxYmiMPzHL+utCzHOFJmNN9zpupeDr4bdQUbH7am+wGojn1zJ+ZxM3tVyWyOQ
vm2ZV+zmdeLWmTAd3ceFI0n2Cv5eRqj5YJFSnp+n4KlHwhOxFZXZxAoj8kVVwYwP3520OHVF6gev
CCIadLtF2h8kQEEsSnvNXrTAzAmC+SE0q3jBw1EweKS8JQN4BIhXnPrk2lPPfMsF6eiCpU7+TT1T
RGqo7Nfx/a8Cok1EwFlMG/iLUSK1HZAR14E4i7U1cn01TRYgGqn5HRAkOjjys6UDraofTYUTD9K0
43K/lE3JRFdbmQVL7rQWXGwT9vdeoc/ceFnKCo3mAxD9/BuTP5b+6Y/RJDUWHPzeQscE2eJp7e40
2aodcGpTLemz+2RqjBwWSyJtRmSFFRIjdHOBDHmBrxIQDMHsDsd4DmEuG5EYFlM2wzVro/kuW+0C
YH/us9225catP+I4SR48p3yWNaRAASVMKsgTKbzEfppxQMudEicyRnfkToJMWOKZz9bcz5sDDtie
KNRljdoBbxkGbGCr7HyC5rmcs/d1JiuqWVWOqX/CXJuIdkrjlv28GJuHb3yP5OuoTDt+23ETqVh2
0nLpLeMKbBOoKqgqdhy+kAW/ONLwvvuwe+XZPAgInVkhCL0cDtsu1gugbKSrQowrmXEauWzsNMgl
ytSTjAN+rF5BlpgSaoqFwTPB9GCVMiM2wV9+22Iufh4z3Fd8Bh95w9tpKUhO3Ca22w/wKUgOnbIk
G9Dt/fUi8LluFUQ3/y/ehWPUPx/AmCVpCjOYJCsI+CCJmglBhImL0FuOP/xZQIIEfiz6AgCFCubG
7BbFhrtG/Cw+tu3jY5Dt65riZMvysui3TMuUpiAo9AaBnz4b/VIjlHNRqLx930EeNzDrI70isrIv
JRhQbY3S59V+TDw7VnV5i/e82uQ0jh1sb7mzJDlJoufdKoRKH6MkChVCdlhTe06o7Yw4WBJgWI5h
LKUd9ykrFHDw3lzEnF/Pqwncb6Eh4p3sew7DBYYnm5MRHRLOX2MImq/5ez3L7JlO6YaB7hxBOQko
5mKfGatdFamXWxVIKRXNTcavqEENjVrUK0SQsCEibouMyy7d6y+G3bwqnYic64uGHhYQ4gfmqrAp
gAwMAxIuYe57LM+WbKoPrLnGUfwmzs/TrXSem6qGCDmDV6Jg3KGEPt1inwlCUxq57uehFEpNhixe
Dv5Z7J3lcawnAOJm8T6x6lqe1qaX01DLEAsMCxZ0l/yzknCFxHHJ7GNNfHjvuw6aoX3simPwLKPg
K2RD25SWKSqGxDisYxFlmc8W0Xf4r8IPAzJh9wr8rWqmgogXrUSwZN2YAzepb6nKG1/1vYsrqqbp
DGChbYC8+rstz8llbG7vt42symlWrwERYVBybwSYQAXacuNco7Anr5GLfZuL+B9gKhjScCwGgfQq
X7LNec9wfJfXGll7X9MkyFvk4Lz016O54zXtIxrt9wHz/vF6YnfYcfihFonDUHEMXwfKdDY8mvzO
hZVxTNvrZuA5AqJjB7PzO0Y01/y6l/HK8QbGYaET4F6waPGHf8N8kH/kVHvtiGoMCeZIWETIammr
o4oqACFieXo6z9kRRdrsyiHsRNkrTNGQlAT7hBm/ODosQ7nqKHA7Sk49Fu2EqbbrdX3trsGxWYA7
Fms2uKjF2UO9aF8CZhNQBlgid00Cp/bCT5+Qdqs3pbIhXxzsHMmTWNtcx9Ht+69+DGSJcdy4E+uz
D/DY83mQB917ceWJ/KuQfaaJJESreVEjsNRnM8zqJTjpQPZIQPZ1Q8xdMzoNA27AotXp/cw6J7rQ
XIdBpaGPclZ0Kz10Sf3uV4wMww0cTSkuEFsfFcnzU7QCTxEmOoIAv+n5ieUKbS98p8e6+d1eJJ0t
k5xtbubWUZceYfA58uoFadwxiAU9LcKdDgS25W+6+YZgeq+Zb4mn1YhGmYEnxCO70tOmUXZMbVJL
MKFtEwN+BZiSMggVjFogry7HgCN8Xp9ztSltKb7k6BtnPtr6ztQD8l1+HUL37I18XFl9rPbCQlEx
717ldc2uAoIM/3LKtWK5VFYBYL8dLzNICnE5l5d66AwTfAKtIocpm32lAQTReitH5ND0CMxdBaqy
uU6vqw20PDC8B8Bd+mBRqpnBc0Ml+lWA1HMFBkc2HfKx1GZuS/M8DyHKTAJ2cbTKm9PCLXGS+Sy6
FWKIvk5Avmmvh3zjTiUVm+vkx8stx/6jlvcSEhEhbB3zFAnPQSJDlWQD06KE/NKw5xtxN4I5Og5f
4jUivdujqLyTDjspjuLK40gMiL5sOs7w+1PPWUp33kh7qtWdnpSnNOjh60bLzuzEWufVqcL3tiWO
AvhwzebLSaw+n3M3JwdD+iQb9ySlGgRTpWzJYonbWZck8fkAfn6MoKm6yldj5v4ZlDWBoEwMhXk6
c5EQ6DsF9V/kRtJflhjlhFQU730ykcPKv/9ca0N5FS20VpmpBRJynUj3jxlMTnGeATKtC4m3gBPy
Xrt5UU8LVZy1kj8Re6qZnhTRhEDp8GunGneDreXVlHL2PJA0dOvs/sdGKoR1veDUoJvsKWu3np4f
w0EnsD4aW4WGNvdaB5voo+MM6+Vun7+QNMOj5GaArs4XkrGrLuC/FIJ3FD9TvIHecdzu8iSp25SD
LM2KjSAkUH7k70SKA9+3L57B8o8j5Mn0J1zL0pvoFZCTrG4to1nyb1KdEjHSggbXx6D9SSqdLPBS
hMUiIWKbnR70Wz2MjOkBqfru0QyoXGyEIXw0qodAX4WCbFF/vzEew2KnfIRhqW58+xke9X9mZ+Q6
kOKuWjjAoPkp0o7scqakbbvK9uRJCGB/pIoN9xMTsZl9FJRPv6VAojj8ojuLMfl935sUaVxpdLkL
YjwVgHT11VHSZs/941VYWMtmpqs+5Zv/0vEhs+pI88ikCXP4bNf6S/RaXh4qcAZZXv4DhDM9kB/a
8r7e2Mz83IdnggoEjvAX2Vat/H2E1DvJTBCgpiWvSnXQMPdoSc3Mg9iGN4/2stcZ8l9aDNvAQScy
2Fv3np7u79T03M2hLg9dBnrzs3xuXwq8y3Vmc51tlv+ZfBUSOFT3x6xlDp9VQC3cq4v9ui9HMwXS
a0+/6eNqb3PnP+Ro6uVj+pjkQEL3Gr8WLgdRp5LgxLOGINkgZ7QAstPROwGokzmfvPdZAuAI5PvV
vo+2epVfBToC98WIuM6hFCimvJ2X/bEXcwvV3wYswrJY0Q1KuMwunzvuLKJiInD8Fhratf5O2t5s
jhrXVZSJUGv1Ad0kzgFa0u5cQKRqNVB1EzrWm80fdw+223zYqrTU6ClP89+U2znEh54yfaE6wgam
eWoBt6G1OoolOgD205A5L41lAzO6mBEyyITaiETzepMn0NcZRPQWj6xzUZGRz5qbm6KeMFyxg5eu
UG1TFX/zRPW8DNdvYimu+zFEAAkWyzX62diSKfOdq3u2j0XclFG8T/JL2cnEuvPXtTUlgMsY1h3m
cJ7mRyV/Lbnqqte1k04dIUCVpN0gRp8uY8O8KbwPjEilDBqrjzUiFrXCHrpqJyC32g5AHs+gDkjw
xCL4QC5/W8bwLyI6AdyZiVT6ZySbDbzafR9AmJdE8W7ov3oHjdEux+vf2m3cEgoGUp3Hxegwf2K6
8z/bGrpDZXLE7ZOh+L6Y+C5YzgOiJ9oIITRuAQpUVj2VvU5X3zAIC3VUf87qMyzd1JJ1SxdZ285P
Jh2QMRyAnswE6e5M9WnFYgKhf+92Bp1xOyX5mZj5fZn9lJc3cwMVqihpwjwJA9t2SEckz2adgG2i
YWyPMKQWgnRD6LcYH5IcEcwZ+rGZTgNpuv0nh8dBjW0DrHciTZR4s2FUhmI1bB5vndbvGJs+DnEf
f1aQVlLQggC6yXL04YEVFAjSAcHBuEJf0+9xAQ/cYENzZVb/nXT/Y8CfAcwN3geoNFqCRqd77Tvm
Lfcexeo1dKnL5BMmj0+4poCFk1uuYsa8BoZMerth2BnS/JTIBaKhg6lZM0TIK3Jd9MPIYl3KLRD+
dAts54sDx19LAfHgPtP2ILOxFCZXsqTlIzwkYjxNlcwND05g/BZ8L9Tg+SrLelot2aMkdkvU/eIg
q8Tpm3wZCcjbrP3UI2vhI3CJqqHzp+vOXmkD+EtMkLRTCuRDTeKmkXOPS4YT+YNM+O5xzWUdAjoQ
1Bmcj5Ui0DjUTyfZ+liFW/iuBRnL5enG18CNW+aYnA3OKd/3MtyTAZ1z/qOkAlKhgijf+VHQFCBS
zYpgcmQfKuEtIF+9Ufp26iXv5nnF3VLdiPixpf2krlxwlajLHSCc8xsK6ceXBylBizMFOgLXp9TS
hedAq3gIZgsbc8gaZmOPU2vZF7GLv4w7TjAln4NPNm+FQSdJoL25+oFRLtHp7U+aTzzcukTATCRk
eKes1nurvyrqscJ5WUdH/kKod1S2bdMgherBYA3Cn/Y0nBlSxqnCLnujaQh4xARG1XMaDeDOwr6g
II4rNZssuXb8j3JNJVUBfDXEKWCdDf3M8Xi8zP+/pN0NxRLW0NE0badqzy/kwV1P7KVlsa7JiIBp
jLy28ksmD4NPoxxYRjFRpP/61S3o9unF/8ksm24DlqWqD/pBzKBjWnwGDpL8cnCgl0N/aNIJESYE
igv/rCygDdSik/B4WMAAUdxriT9trMxdxdmEJtF6ZaFlK+v2qsGSjUE8LpBRsN8dJinNBAmq2P/a
JvPfkbcbSCLpPZ1grDg9CubYSuwb4cMFx+iZjmXXzpq1ujoiwvX27AcS2WVplsydjr7DvEgB7vmh
Nqc3a3G4VBEovJleH/Mi8H0MxV3r1FGfzKWyBXyCsXWgMLdM3FA04LkTg1VLq7fHHhRjhQpkLK7B
1PVpPFhVSw8AQDowipRROqjOEv7+4dhSKoQFzTeO/pTurk3wT0dl5/16BPXr4Icr+X6IzRRX72wR
72xzKpHzHdqiooJ17vROF2yXQdv8kZo+dQe0mk6TiArFzTmEzsjRJkgbZuYS0fCiFLhPBFyMX0m7
0+RsIRFPrBlzrIm+WbDZ2TNiDptjXYyoXbU/YVTEwtgfBt0qmacusKDNUKHBWNeJ2qfNDXlrMCTs
lBQ57PBCr7lL7Gwn1xLd3yccNYi0DqlNluJD7krfoTC+G7lOeA86tHEPsMqPotfRbAh22LtzgwJ4
UydVpyHUuiNumog7zorKDlsOzNzca3IMMCH1QLLp1b0P9zM5Pmp7OvgfipMoy7dLeV8CELWmyaT9
G6PnMo/YXv+mS8nKk/kh43UnihhbbZDnIpXe+A9gPbG6NVQ66Z7iFBgXNX+3zsnSv1ux++QSCvoC
xGj94rBQazxQ53We3Rs7FV5p4gmOA4w96GZ8E9NnDHGmC4i4c9eo09SN8fL0uMEp2ZNbS8eT2020
BogUH+TQCngSLABbNiuXdaTJ5gKmmQDwNXiFCfTpGpm7MTn/Ah34qnPV2gqy6IqgwAZHdlHbv8cn
Kjw1ENnDel66Rn6YulOGWPdWbLj0eA3vSwtEiAtZFlHUT+kx4NovKEzfgxHiu6G6kST+ERW2PDK5
AaCjMcw+3XTiKVXBlP+KCpFXVnDXfMLHdh5DWXIqpGUKc7Bk6XrXmzl4iXvNzUzv6nl35ABlCIBK
bCxkhZapf9J4gCnanYRFiTHyqe5tDpAZQMgWf26d86ZyYBhhTPCpOleajSVPs2Fq6yiuv5XEfGCG
KBCPctPySDEb2hW5JNHPl0NwEM5o15+ScFokmvpGyvbpSjp0z+5z1Z9SeooWlQqqWM+8T03R1j2v
NCWwUchjQkYvxQnLnz0dTyGhzL8rkWVu/QmMuXLu75aewlzEtCKzghQTOloxgqE1urdZsWIG0gQg
PsGDrsuBn4/kA1zdeRLCYvakh23dtt15eclbhXBKAeQwEmzQLfhlntB1w09AXjUj7XXzj8zLWPaK
qSRRKNLVUuM7fgM0uxRkTLdLsHoD1ABAgcevL15pkLxK/Dl2ZUZngqRRGkOl3/xqriv+jWnp2tT7
UA0Mv2gXJuLWZgS0M34qOjJMeftujbXke1IAxF36HzsOMrNdHyLkLqVMIjG4w9NGYkFv5VBaieLs
bDqRMJ8tDI+qhgZUQ2VaQPliN//SYEWqRaXGAgCBMw2hjwh83a+YelRJmpzypCEkknHOa2n8iU/q
BTloG4rTCjYNIernkoxuCFKrd2CGkesGziiFYWy3ccw4qVshsa+QYLFo7F3KzwrjHhc0MYizUtxh
Zv/LnZw2SmrK0W5UulRvh02Z7hYd0aAYG9llGX+FWrlUCUeGfu6XBX4RyS4cMJ2BRR11AHR1TJjP
I3OYhR15GoxZqRfkPVJq7H356nJ+QoFi8qROV0hcme5FyXQEEHp8eIX93QC9tE9/0I91p/yKJIFg
QsjsX6ZhCepvFLWaFfcX6qHYEXEf9n//IFPM0ZqEuIvJd6kw7NTgKDTcYRiepjz2WAlIIBEgt1rV
QvwZSTubivlvnzCAvx/Nbr3fWk6anW8IyEhncUkqhiPBF8f7vVgNUc/nv1g21CF6HKOErJzAQn9Y
t3PZdTYZxXyCbqWPB2xDoo2OSACe/rygAd8Dtv8FGo6V9+dwHQXmFNtjS8KNNFjfoPkdOlZeq+/O
rpaLLJ0+9xbrLXYB6+YXd2TTPf3zwKENXpkXlxpt/8aIwVSYFwmHOQFT3ABNN7Q85SeI9jB+PDrC
fgip5H+PnKemKyDOolt71Qpa4OZ4xFJIGf6KjXXdHpIPTuSN5o9lTtyKAHeCB7GVQF+UbqdY7lLG
gD9NRKI1pwZwMVxYHI4YZXcWFeE52JLhGNeizdlghXP/hetsRpLeag1UAqhsgYpP3Gv23FgKGijl
SW+C6yUa9HRl2S0FP8SNCMRQ7iylfolWF2qWvprxHyNuTZkkn1BNQyWcKmUtFtsUfqQK0Xe5szVj
oM0YbSwtNcX2nA3au3JX+Dyl2c/AaBBIZMAc5aQY6HXuyOAOF3zn8ZJkKDK6lmriOzwBjn0SZV9w
iDj05ITMOb+sw4ZjhhA0FE3xxEiLoAijQCDRYWaENEJaCq9vCT+axYGF4Q5WAff4NOOGI9JCqqMk
lFljI9zrboRAyN/4KWLZ1lq6Jauhxutv4Ll5mGinJJJV8YXn2l6v3ldmh2t7Nrkga6kVmbEPkmD/
1jhAcsiCIxIeJbker5rznGxKIavAkHtaxNp/zk/mimXulSgP4ht7iZ3GUGgBjvSWL6iCTe8je4sV
/QOYqY9EQPM8aWJLv8oWgZJ32HpqEPvZA3hUOVD+K0GZ5o5ft3o5PXjhheTnm8Oo8SfIgGh0IDLB
xbvZ2BUUu3w3qbz8Xl4UrSS1rqav7IU1YrmbH/5IblCeBnzHnfaaW9BsdFiti//+RVVLg5g8HBqr
9mC1yxSanVO34Qq/nFjE22x1NY53Rjw+Syxjm7c3yNXMWb9A+WZPZfvEQVhuf5e0Hkq0zwBa0SGq
GVibQ2eC7eliooQB6EPfZAKkeLjgYLzbcUn63IzlCAnCoBF+jRlOjyYCrQvWMdpjSYgY5C5NIsP0
a5rXm97ZBEz2/i+HG9tC8uljE4sAOS9j9Y0DYYu1EIGpBntIiOlg2AVgE7DFFUrbt7OC7f4FD4FU
AYxWMXQBu2iLeYtPPwr7RG1N0jq7Ox//fKzNHAwS0o+4p+xhQDrLJpX20ubGRoW0UcbrXGMA48sx
A2EVsKSTFs5EndHa4BAi+Q7nymIbg20esytXAtIekXgfVR1Vvb4o098jGj95S2E872eChnNkHx8C
28z77ditdCaeJnwGwGdTi3USbH3d7M5A1kNMk4TUjhmVtIdhX42yVgGkB00HjLO1bZ44erowMkSv
IrpcF9jB5Q7LmNdIuFHFpoYUA2Zi0ishR2Ee2MCXpJU7rOuq6RUpvQ9gmBQkfd4dPkpOcSwP63a9
NddiXURaSOItHErgM7VOxKqSNT3CfiVA/bZ6BbgzrGkf1oYYbz2nlSDeeCUPDcd4oA4kKTp0Tk/9
/LB/Grhd/uSjct0jAUWP+8L0lDdUG9SkiRZg8nvrDWJYVteiNC2SpRJcQEUK/6+rmuY44cET7/do
Xu9sFpRp/WuUF4S6NATJhQP8J92FKOq6EYh5EyPdnnYgP5q3Z3jviewrXFU6EidTJg3jDaPyUsr7
Wb/qqLx1iKhDDJ5EQvRaglyeuvYbA0M5wIJ6q/37Sc63P3hu4eIAZMzwjzQhsaiPOaTrg44L0o3J
vjSVJ30HT8vFiIBte+yztGtETbBcDlUHgE6BtRkzFn3Y/hIAhShjCo/4Q7vyDgU6/QUaC6JUqwPd
IJ2t6tIbZfbHDwHRPVJThWtji7mf1r5vowqZvM09lj8zQO0Fpwk/kfXHUXGBflnONYcaxDpIlYL0
SKWc91z8xNUeC1VJbxxtQi3bM0eznBSo1OO9KNXeyXwX4Yy+6r4UAgM9JQlv3Qy+B+pgMan8PPuC
2/sCOGIU6mdv2XJ3DFCi9cxPaL4Y7g9Bv451PG9lscjP3d2pcEOXDI/Yamj30CMNhz7GT04fwizv
Apcfxg0+HcraipT+tjcBXzyhLvFpsEJ7egZtW1WmlZaunIK4WFnPzrtmSfg4312EM3eiqrWfGrZ9
1f8JcTpvuwUS/dk9dVLYtEQf7LazTHO975A3bWC7rxmVSApnoIIRTettX+39fitNCvBoX9z8ub+K
iMg9hz0S4bi4Tm4/a/eBxS/fIelxlJ1foqpkg8bW//Z/tYbdXYLbkCRkIKBiHbN2LibdvnmzZpRE
iex/lcECB2OftP+ZrTZjWQnc9QIi/rHLYJnGzu/JR/T9r00NlXyee86oEdeyLlMLwilb1VoFwDCR
6NjK/g075WUffnj+UEgqYSlbtxzZ26CN3eoeSIn4EFMeZI7eNFAOgGRvSSFzIeTLKbjKJhQjHTP3
mUo6Djg7k8e1VT0Mms4wW1aKYQmoNZw/yzL/I2wGTHFgx5XVyEy8VJfQoolOilD/AlZrzILQBGam
RafPtc++ECTYO82UwIkb0UmOU05BgMxOkFN+xb6OCSFrVzz3/lyi/ijYT+emC+wZfa6c4RUKd4Ex
MZeZifS5uyg8H4tWWSkWlMbI/XDqzqcELaZy5qlen6rE1tqIUPpy6+8dcZSU39WCn5D8F8uknrjE
ZHckle66s2QALPKbq+ktendTAeNIsFyqbr4v0LRjcRaXyTAE/Csf+TZCO4XyQQ5sg2w9wzMnOmUf
+rXongvCn2fjzgPl5DYgP+qBfaufhcqmNffo5q5cwmrv5XvTTAK9NcQhu79fdB9/nhMEQAPhhusK
G8FxcGwbrWNSQxoA1UA+xwhH8w/aZobkk9PfjG0oX/IAuvUAQXGluB+2mRl6u9HWNI76fNFxpLt0
dzD4nr1+44J+x1Z7PaFEYO1jX/zdgXTKT692prErguH9YqKI1eSFJpuQ0S4gp9vCRUvG0V/Cz+rj
iT+0TOk6Wzqp/xiKq8TjVqSNCRWJQUPrLW0rXVYE6GuK+Fvj88IIqhQSBtWDq6gO7QR2h7oloNSS
cPrt8HZdRR/7mHxhHXoeLeUO7hAE89E/yaKluT9kkPT9gVy+qZ/xjb7L8jEk0cu429VOkYhRyl5R
bXTIlyRRjRwC3U5e6b5a7kskDIFDx5Cp98X3Vfp8D9L0hDyizhOKFFldoYNLGhIA2wwEGtE/wuq3
Crs6pJOY3u4u/eRDvnnTS8kZog5LJ3rXNG+Gn10IFYlqYzUMKv0LYJQwyhftKq1EoxnbgDoJe1U4
skWbnC3X5dataYXQCKW7f0sV05zgzD6smvQlGhfWShN5Ndj/imomyTOzA6dSIGzfxaGjjdlZ6oWp
57cHeFPlVL1BgygRpEbqFoZf56NjuaVRnimPyJgB/1oGnzu5ejBMuc2LAUxz2IczqXMv9UtLsxAA
IKOPs5KatuMO4TyBdFiDVCdZoM+ceHmXW5tnmqALfB6N7qVo06+o2QeOfmh9ciTbQo3irB5a5f3w
waLhUu9H44qrPvvXzi1hKSQQh1/URwd8ILnN0Uf/CvIPpCdHVUE7tVIzHzzGF7mucJP9sGblDvhb
GQtemPgUytki2SAi+K758JGpdpKmgBHG7aa4FgXEPdO2AkJC+M5TxsSemd5DTv9QLXzsUg8q056D
2QkCzCmsn2UPNTNEv7EvjEqvu5heEs/ypMKbb5Y7Q75k3jHAPqFvCZ9BgHbKM3A5IYf6Si/aMCEh
0KvwBLhP9f2bocFheOlm6bSRAUys71ULURp+YvISs2vMCnWEdF7BA99IkWX54kFXRut3hwzyK1Au
8Mix1R7J7u5hy+vuJ0bqArbE144eoQaDfWMj5+UBsmMNtL6wYTu1vsPIjPlE72BGHdwLO2pHDYG3
MAo1wbTYLXUX+XIwfqHUIcO4HSC1p4R7DZSSjDn3CRaxRiNTi5vLsj3PmI8ZE+uDtlH8yeq0iaEH
AAs4Iyqj9TXdnbsFPtlMvi9zt9EHU3kpeLvFSHkeVS9C7tkNp347J6Xxz2ndPibAjj92CT4Q5N1d
iA1PrGiO2WvFMNW58WqruPJHogd9R93g0vfOjK5SaZuSFLxx53S31o4Z1/5HYdStOWSaO0EMJpHH
4fkWb1jEGcwhXJjjUNJDxD0XfuV+vhRxELBeWUSSteqPOlZGsLSC+LGFBRABQUJIhKrt58Udmv53
Lm7iTEfYdRtCXBApQUyngs8hvQlPiXx/f1jJN9k4XD8KkjAnCCXkaO2x+6nSXRhIrzm0Ip00ZQjv
RCFBDY0fTwRushuR3f/j7H4u7hC/0t9WwVvWFk8k8wOmEqpWDJVuwHbmnw34RXdiKgWCrOWvm5c+
zjPZqTISJo7djus6BRTcNI7TnAqg0JBddN9Edjsb6nYCKmmHqWnB5P9ckAcDxrdfHJUmuoc3C5jb
4+FH/L/w8AMGeqNFSbIDdjjZ0XuveDjZEkD/YlnxIjL55OCW9ii6uZ23vMJsG5g06RWZCFROn24n
84DTyMlmN5tT5VyO0uHy3Qisl5mhaV8V/WhTsimT1aW4hD8rt+dyc+UVe8BeWFf//1HdcjYlx413
ycrcWE7Jcrmq1VjjLeAPocvIVclRs8P4zEplFPf0l91CPms6IWtlwqgknqjgG28mrbzqSOq8wTSc
NrHHHEUvISw27v+WROpexi4k2wKGJYfd2R134xsJoGPFBfKfMT6Y4U0JxfjUACzZuCCtShDvmroJ
WUHXrDXD4SJ2ZQDN/PXt1HLeQSxjYhvQMTlj54ppnCv2TQ28plsdwmxCYTBCNOgPV+7HFIrqwdf+
OSM9Hl7llOhubsspcee+hym+9e4ZqJoF+NCJqCbdbqgvxtR/2QTzHf1vtVCDJk8P8qdFMumNEtWf
kukdr8LJ20mHwCD3tDArzI4Q6ScbjbYBw5S+kuMPOCqJxHAIo+1xV6EWemr+L8I3IcsuvxNJDaNZ
R+/SZH9nFaOtBbR3ckcAAoUkcqSrMUC3eVQj1NcH17LF8YJNyR6MPc07bOl1gKBeYwQ+fZt0UqG+
ovFeB9/O72LNGWlhTYDEdGW74fPpKbnn7LXwa6YmlLzdqYDy6VbXfmBx7K5CQzwLx8dd6KoNw0Ch
7beXl19C1YxnNcx+LI2BZKjUzBoaAVKwxY50Mu1rqFDx8O4UpM81lDzXcJexMH0q7fTvRxjWoBhk
Q541B+d57iuP1knYsHkCo2UBk6bRVMtLfgyohm7gPOe2i/xI+WTkCa7+iWyAEaKhqaKIwD3pf6WS
X5EBgHQ07bRIxBxk9XyCPGQPS+cF3TL1yZRHlrDbQDXIY2XJu96yNK1eBPGHbS1zOnlOQLux5N2n
Y7eo6SXS4LPv6bj7Hq2ioMxQ0z0xxvpEyC38fGC8DV8f2MtcsuujHUiiejoqIS0nHEQFm02ZkkSA
Zd0QvizYyIDhHN/MqGxqdBTIKNAxhP3wjP910Qr+E4DppxfgOWF7AlrYon9PIlBVzez6SkY9Gzbz
Cl/oKFb3sV8Q55nVAaThRtTpPlFFTTmwefpK8ijla12vox3fhEzONnLXnhM99Wc1b+RPyzfUX6Iu
wPdcCnw1OFZLtMUKPutXIKL1o9bkTkIuCyypCbZEnBI1CAZRbX1BrzEObxinG5/DYT+4zrFVXlhl
vMea8IYuBZPqvLaD1vFNbFd/YXMBZS1nl3DdeX5hG+WmIwQl5NLB2RVZZKNcunVUEEHdmbfEwaDp
dHdzxrwHJrAzwWYOCRu4aY0MVn5WyckdhlucThNMHJtJaP/7ajdwww5seok9E6JHzPfkzXzyjlEk
/pA/7+AOnFFXMa7lAUC9P1sEJf4w0EVmKbJAGmn221th4Kx4qYxxhU0IMt3LtZQFLtgH7/CTzz35
IaxGLzErneNd7q3KIiHjbKIZQthkRe6GOEEJWhbmlmnKZ05Osy4ZI2UTjc4RJ1BrUjClv3Re2uXU
/4MGieEB+xhg6qMT+K9deAJP3DqAZQjzgEiwBi1SdKQrDXNoUi3ahoHPbVaersachczx+zcRDk9O
2gMVIWdUtFrCmKLj8z0FdNiItRclbnsa6xAxy9VUn0kh60FOBXsMO8Uvq0Ow1XkGJUFWc6qlB3xU
wLCls/w0Skk1IvPzo4APJsvKwSGIy8RGtkbVseBPJe/nte5iVMk5XZ5E93O3uUQ551TkiJDt6pF2
s1zPTj5Zq3IpzrbhBNQAguISXRX171oi2OFnulc+j4j8+iekOsxvGUMqMjMg0LDvsIoQeM1zJ446
wdMxYD7IDbQU0Mo1VETp7zI/iFJ0oXCkKopMtB33b8c9f7hSTwAavPHy9pB1d4L7noG0yVO/JSy3
vrmAOs8bOQTrPQ4/mr3gHmybYgunObjfbBBkzNLB6eTDdAtGHkK5orZ7UrdQ4Ec+o9MUetX/Vh5v
gZbVNf8BvGQmS0LEFIom2s/ByNqhmwWtMjH4Pvkkq3ehOPwgapz0BctDQ3WfMFEKXbrz9+sfOg+Y
GUCyoJz8w7Fw5onj0ReQhLjMCIIbEKOkRwzp1lWywMPypun6grXk1PwImg77WyslHLqQyY6IgMZu
TnjAXCkq5ZpPeZbZHsIQlhjr5IQHCSeYpFDMs1LLH1MDwJfES8WKN8W9aOlIVEKbIe/jdCuZKjBz
fjgbzOZ1TzHLYYFzs/zrpSETWf9Cbyqq4+Nde5o6RFaljp7vlf5RPYt9LPS1lFf/uSIdpbqQ81/y
DKmvzOPdWwsxNpF6/Zsw/xXyd03CFJuV5Ac7/AW5Mv8SUHflHlFO+L13x9PDfUdEG/g3uzwMEufc
dIDvCAc734sEWiwY7rKNuWmv4vvpcfmHk/pQYf80437+0QHM8vHF5afKJBKk0MlA/UFDikQ5g7ox
WWJ4AT1txdFRo6IEQNvnmpLV/nmlDXx5eusQIcYy+j/JBILngH2LdLiBeeXotNcukHQNhEamL/ok
gSo/Ip2xUj26RV4sGmOFQPOhCBR0swMuJS9Bj/6pMOaNUGeOXxd1WE/OxNJGXmlUudBd9jzYCIXz
0CEauo0bUOd8KFytD2aPdmoLfnsZA/W/LCqoRHJ4JUDhjkLcV5BIbTvNuAV9JjVrY2f5nYaEMSlr
wRJBaGqPpEp0Zx1cR1GeE89l45jqzQTfxh75RMpQLJqOySvwgpu7InOdREUu6tvKwpW0NpiIo9lr
EI2ERjH8O6h/7zIe5h684D1jY8VcGlP5LanhO1Cxdj2gMj7maiWp0mg/9J/0fP/tNechllJQ5sMn
FFffl/85qGzyMfAab4x/icaGb31vrIg2+Cf/vwH4lAe3ZsPA+20mDHDGWIj7oduebFcQ/WRSNHUe
7jQ1pHxwCLakeNS0wWJqlhN+tGjAwqEQLN4B/QfZkIAS6VtwSBI26LuebPOKVFUkZwt2lVt9iFT4
iUH8SDlLuWMlQarjj34sKESXMXiIvZgi0p9E8qmx+ZtCCYJ2IGE/w4ydZ9yC19PFJeley1yS3NGg
wMlS3215Uir/JwUEy22sExq3wkMXZzTjSL6h7NQJHUoLUoR25Dc3jKz316IQDTyn/0Bl3jgly9Rx
xkyPyPCGHJdEkeL67IVa06f0VrIrcYmngVeLGNi4K8NIOVNRY5Bkqm99l1Cml+j12/rZrzCTk9H+
rPmNWvEaqMd1pnaNIJRycKp01vdvAODf1B4sy5MrtX+hFcrG5OIGSz2NL+uf/T1anQwsh4HOFZqt
7BLcUfbI87E+w1yAqiZ3dTGLfOqAbsFICthHqFgnEMgRcb8qY2tbBX81bBs8i60URKT6FWfeqYY4
dPtbiio7taX9KUwiZdZMSvIlCGaWY/4xsYNBRVndh/F/x7aav6z9qi/meJuNYJJZOVvJPoriEy9K
rvkqC+ptWgwxJKorisUc86y+vcwjD3f8e8mUs3+9I8MrIatAGY1k1nN8JCIsdONTOHSPAcwQSEaN
2a6tRRWub/jZ7y/XCY+Bz/SQZGILsXvJzR3nUO2phSWV5gnz/zQ82uVtcmLK0cRrCVUWeWD4gWBQ
hd/Dkp1X+1YW19dqriDL0XNSMoz8XbcKySbAeLsSL7hPTW1209Yc8dmkJCGh3Xiip+h2v87Z0cH9
lFghZfa6jzTx9SIQlWlgnW7lY13KFo+mDH1qfyPJjYiDkAd/yZ5Y94/wyuGdHVxIJckheXffRsoA
8OroA+C6Pwrwkav6IO/f0C7NbGV3k3ArrrlWQSSu4PRL5fnm3bWVHlQBOjRx/qBeMEOvuVo55eJB
o8UzBCCRICSI4AYtTojdtpTdTjXBGjYKI092OGabd4zW2Y1oc1HAeTrPc8xkwfp4BqiO9NDF7tMr
CRjX/pPfY5sqmJoOqjoQYHN3djbWocJftSWLP2XkumItyWV9FfbvsmjKP7uJAa5nl8wCbwxlYB7c
R901QGntQLmFginwL+n1WS5Aqi2wdA3oqO/C2AR+zH2ovgW6iUYbKTCRwrgPxOwwt97ZvzA07bQt
CeALMbju2l0yVXFZED7ORLOzRcUdO9cFKW5aSQSX1onC4jz1XOxpj0er6Mvpl1RXwS+58yszbzon
hPVAVb9DlVU7ZARyFt5tuWBfohVMUVi2EvzuiCmnAKxPwcYW79MtHQMWTmRy3r4IvQznz+uz5ppm
LJi0juSE0f22Wfys67boNviKnq4TtX4DKf/axzvA4O4C3x5PeJtsZiLroI2ID/7kLkxzqpq5e1Fc
QrhiUpLHlMQ33DtfHCrCOpz0P4JJU4y2gjsBtwV9CyimWx8Ws15D8euBjiisub0duy71/t9rZ0N7
aZWfqRi4+R19MlQ1O8UtyySkyNLyGsqT8zP/LmlPTKGJyZzU3PtzntgVw7vnPFP0rE+r2impFUSg
R4TVQ0P+gNtmw9ahzIpFToJgmwSUoFtkgdlcYzyyYzR5I71bcQOYczC+Il0yOyYqlS8hVLGYAWbA
TpEvn/4RAe9poLNL75a3esRFMJwtsCSswnJSYf7Lx9dSyjkGv6glvVD0VIAUX2x95WIX7HxMKWPi
mOERW9B5TWFIjzGLrEdZAHG4kZjeGvLNKodr6k16+tKUH7bMt7Iz2MuVDMbxcBZRKczECbL2udBk
/JyxAjinRyAA02uSV4VoRPqvd3w4JnEdMmycmOhn0dOp6N02TYUSbhCKAZA14KpigKLF1SB7HgJS
cPgv7UQM1LwA49yRj+f0v4BC51uchWm+KrP1xvPj5tZJMd/w+sburO39Lus7cOLXbwjwn0VJkzrL
XqKK4yxGY97E4zROqjsIaa6YBLyOnmLuA40g5yKrg5CdCtD+VlBKOE1k7mFggzt152Yz3Oc1BdPD
DHYwKmoSCNUMWvdIjbybnuqyhol0EpMWLWr020raHpByMay604bXa6UrVvmjulEJkiHsO346QbB/
iqK6ipKn2Q0c9w3f3zG0NIl2bvpDxPzN5rCXQXM9JxcTH66nxDFku7VQdkXtG90XKrdhfcug+WjM
VppCfur40SVpifFWAxa0rxa/fCRDZmA2WUzhWcDBzqFJMTyE9gP2FetODwhE+H/ORqSTkaBGjzVY
c9LVqXzCC7ZBoRqIGDd2HfsorVmuVBzbXdIgdAMOGP9iy5yl24BTz/Dah/9LiBPfn+Nd3Ct75Gb5
ZkB9FZGxs9/bpyJCE3kEelFP6dOsXkqosJzp7qQiwsXt3oHrX8FmZg3xwr7Md5rU5gNB0jFGcqlN
UlnmfLF0k+mlJ8fcXA6ue4jww12LWUyYaas/GcS1FVT2SrjRvQT6pXsBhBhhi9TwQ6TqG3A7y/j/
c9WJaWz4TB+oe+b6dZqHSkY3M8TCNs0Ff8A8Fk9lnsay7WOWJNPIf+JpK/QRveekpJwWR4nU6Vj/
HTJ2KTC7T8atj1gvJ7ySZ8RlYeC+9N6Uxy6L8em6cDErecCfMw0ezulBFqo+wtxLl1lWoNMMp6WT
AuwFsjqI70m/svzAp58OqqBkqzQeq3EeOmPGYBD0fu2bq/QKbufoNLVI9nDuMIu74BBAqwGhKUal
jQSJSubtjN5VbCIv6vOI8id/FQxaM4IIbQPYHPK1eooLQUfM6tx2BTW50F3b48UZ447jWfEda5OX
TiPdIh+vMR2I4m1IRyr5oKkGj3Ot7o6n1r5ppasrimD8qcbBsC0ZvW6aTNjmtGMG8oHU+VXwD1pZ
CXEbgJgL0EodfZ6UE0JstHn8/uEQ/WKObWaMMKzWgEKR3W3/GcWN9DabvS0OwmER3XdKa8TW7SDZ
RKrp5yKO567FnKurHbN/QdyG5OXWcNLW1eJyGTA81AknGT4/8rgs3uHUSMzXo58e4yo/lVdfsWOa
5hbofnsBDdDpgfzzOSbG0fmdJZ1TYjDR52uQwqkJ5dMhsjp4u3spJTwiLZC22EA9BmY43eux+djS
gUM7PH4rNEmt6JUnNFSA22z3pZ9kT3GMesXNRZBTPO0HAl3N5wy76JUgjn5yw2094QA0m3qlJIkw
x2f/EGipuKLS844pkQvKlh39mSwgWHZEYnqjcCAJQhn7+g0JyOQLJ7LJXloMcb+3ndPsoshb502r
O8CSAKIGYBV80licfcsVl8LUgSXE1PO9EdzUPLNpsXgJRnc+P9sOMjlEPOhODmMDZOOhLGCfzLE9
GXjn50boqeCpvpfS/wTkNHd7uT2c5MEdiO3wbKFsjy25ITOXknM/w/ndkGVvhWz2IVW9Mfnjp0ci
tivX78AQ2uPGpkTJgCar7KginXmRrj3NVjdQahtHmw/uV8Y5X6/2EA+0nng4SrWnMbcyV/Il2GqU
Fns/Kel5ijUGj5Gk78U32jeP+5nTj3+Lui/OomnPaFftNFuPgp5rvCdYsds8cKQDgE4uVJCamueY
JX7nME08r9hH1Xb1iW7+Kd0T2X1x+HXoVR3EnI19g9GksPne4HQa8dWToeUDafE2OOY5I72paepZ
1bTy0ZUAy6ELh2ZWLVtUSHEeTqHrUy2H6x8Wvl5Z3fa40vrxKwueluyMf92Gzo4sG+bosUuqrHlk
WFjH07bWl9LwZ6jtq9vFQqvOai0aooZsl74Gssa3BtnVO9SL8RtYMifwaYEIcpufAUFDc1Ma+/8C
5tsCEYuMLAuHrLGxvBiCSORgYc0Ekg9XqV/9gH4rBndL5CIMFG068N1ArLXSL3vAcFAP1M11Q4+c
gj2pK/P0nSKbldHQPWNRGkPZZ1v9VwWjY8hYJFhFB3+RF80H1h9lptfBGKnbW/cLt32nvvTuZHx7
ioUR0RcKE1fr+8XXkUxTKNDgz6FsaoBhK7DQ9WgTa7WIMefFGdBtmcH8Sd92I97YPqQlKNqwfvcD
107qfL7Nno/n2NxZCJiUoRKs4TeUWDNMW9eP6x9AJjA1IhNI18FKYsP3FXroPkedR41TpQfAfA87
VUZk9kMo2I6v1pd/4iMHGuFDvsERUDgh2NGnWH3X5xySsxrK/luIFnWeOLdmXLRB8WdOCORWqdiH
dJU4/uLyKXRyBzO+DjW6XCa+DtmelNcDSWdeq3i/VoBrTA+TscBIFZ6476XhLSQIHjR0TqTJiU2d
LJ6HFwzB1ZaNCGLHSpcaX1goV4r5YZELTknv8L6nHQ26vFKmvp5WiyBMsD7pKpcS/5/LhQcleEuQ
66xPGaKQV2BE5KZwxE8jFcIP5pCwkAR1SpuNNxJMKuB8fsnowgMTTUtstZ6YcN0HsJftEghMBnTJ
0Nyd+paur6oR3B9UProcVpLRmY48whfsMlsIpyvjb4QG8uKyxvs1MX8dIhayqsCF2Cggsu1z80hW
ln8CzIaFHNtiUzgZr2anvN0Igc5ijlJZDJj5rw5Qsp4zZ6SYtfuZJGT6fcn1xwvk6kmSPrPpKIlS
BWcDP7K6y85X0sw3JYkyqiog7TJHzcw6tu4aCs0OGXdrJDFMfIjFotc+IB1rFsx8ZuysF3DgRxlx
6Pb4pqw68VAcsUODaOkUTeekkrEVppLocjMs4ZfNfC4NTjb0T9F38lWfGTRbtORZ4M9ELzXMXMIc
f9YDss2TaCt4lqNu9hJZWXY8x47DDyAdSeJvknm08smKzT8LvchF19pw9ygpDyLbjxN5lmTVKYDM
VHktTlfPowskpgWFWNunuUmxcASUZQ49c9r/GUbtt1E0nduzvguPFd95VRgNmlSe4L8ZFUjmMiI3
58PBMNc5zenIZU9Z/vevbMKL+crOu9XX32lhXhjoRJk+bt88WX28x41cIKM6eLR9F1chjVFEXGJI
tU9viKMUdgmkBcUGsGNO29eiHgMpmKWsHt3V48JD1HxSjsiUyEiczYgLKslW9cyms6sECweHfBcE
+slLb8rChJw/+iwJwthCw63wSse5UhTt7NGs1vZQuqcTNqB0JHcQePGcLNrCOTDFfS5TCcjElXts
N7xJVbj6YMwrYyzGnwFYfedxjLblqkWWBRDHrJ3nhFypqyxmIabY84EZzw1Bzp0DqBx7lSY4EBm7
Ck8jfCwHuoVBkRRBz7brSj4Uobq3Ear63vEWiHw3Vi7Zlzv3SKs1/+R6FGnEYA7TdASuq6vK82Ps
dLn6VGmmhG+KkF33BSp6r98gVP8SnWLT3lqbSqNdkrUfg/TziBSR/bT314VXR/KAMHtfWQa9R/0X
gVu0HORaEBaPkewzD1HWhQxJ8G81U/318Pqv7yx9mwv9SkWKmEsKb/w+WAWEYCWAzYohGzyY2228
goKk55w1ViycJx0p3etsSr4zHbxFCL/vYpN1WN35JrRYDkLnEkhfK6wo+1lc2bCb0GU6w/nG7ozk
JcpsHeXCdcxPV0+8yEUCZw/qMH0Fn6s36pn8Pg6XNQMR6N/tS1P//wxfk0Xt+9gAA5PAJeSoWUXW
zzZTKZ1dNm3wO6iDdb7ZnpB46c89V2A/rFJeZlMcrY/f7n0KfFfbWBAbA1+IhDXtcQ6jh/V3Nufw
YbYh8+rTIQIsp9i4wLsViuau/gspKKN+3w0b7KoxBashPekqjcnZ/T/ojRqSb6fFM5iC/lUoGcYU
RmgTuLbv2vt1j0t00vIh10JyORVlhrXuUnRqlON08YBuAgcBDBfJKMl265P61RE6KIDsbOlvpLyN
VriyUbxZY0WHfCryeMXvmd0CY3FB5Xq/GGQe0z+4l0XfZPJdJqGBX5A6mI2SiZ3P7PsTdmHsdZMa
CnmAQmIhcWGQBB/MuOX6PQ2+aoXfdxDNlmERanP3uCUiU6yB4MPfIJ8gzPRv/bWp37bbp0l6FZ3Z
YaWL/gt2348IPeu4c9uuF+GTTwIAJ9UvRqYYbUkyDHAVp1l2QGU603sDQXUxsXFqthhXD6ZPTsOw
FprpOxhCwVQSxw0Rg9gS9//OdZCwBKixHdvtFOqcM7tFIRWpQwfa4K5DV56F/UyFKsOjjvBBB17d
9KDAxvXihFwFNvr9TjyS8J2KHn6/0YW/Lyjd5JS1ib7uJiW1lnsGEs63spFeWy4zilZR9+pYahA9
1ekJ986mmQhh3MAmW24A+2CHKusrqFcZxmpX5eg34tb2JCz5Ep+vrXoh7GT3/6WRiJ0ZjRtmZmMJ
AYpfCGJ0qmUiGO4JLUjK8yqsZGmhBFY/BDAcFak/Jx/Z/sdQAVid4jW82eOlhF5555wRjF1JWq6o
PBoEBbsWiTGubEgg/11hcqg5co/Xd9l5dEZT9x8+WNSMKzmdo5ogtojupH+lXt//wrZfClYxoWPC
eeHq5tmFhFFHS0vWGTouotLhkSsR2wPTNI6kciAwnir/lAQynYNcnpgwqATMSrDp47qFa370Wq/9
vfBUw89wPsNVwllyXArNzurXDMYMujkJW5bNkYcuv34tZC3hc2bukQ87x41cJomWGK5W4Si4JfRl
ConCzBaxBIyafK4G3C5zTJHpS1LG/xk6xRdOBVidbTgdZHMhgW7iZpP+rkP+UJysyKdKgA6aP/lA
GzynFjUs2FBXfCO+W96E4Z5ZBIE11sfapPzjO1BlIeGafWyPQrAgaYlV7rE92t26l/xz5VuZXvbl
40ao/WgyIzbZNus5z4cs1cM5zQZF0nXymKk5vEJx+NjcJVz9VPubeCh6fO3ouVKzzBlFEYC3vtlM
yvWkJuJWVBYZCY78zAaXhX8UtT3C7wepI+oMBtZ5tuj/90717forxlZzUXWs/u8SOeMREiq8zpaB
G4ivknKhLAHuts+e3MiMa+Fg3YmiGdXCSgdBv45YYcNg5KzXv5JkCAUsQ7o7E3FFsyfrvDU0E/C7
zzMPpFkSomYXZeL/dmOXoMaZsv7qi6le0tr/3eUQz7YkEcmQFvbCpkHSG/qhwQnjxtP5BFWCXRo0
sF3UiS+mvtSYq3j/MqfLKanBq4bmE1LP7NKL6brjDZobBw+Pjy2ih4hGoRMInlKT1cNMxpAPezNE
lw4Xqdg0eY6scO3fWbWNuh/oL/iPtfFejJ+ovcHdc6DDMsWDxjC0aMb1Bp7LmYZcTYaYUzJ+6FSE
235U8HQeY4X7G0iDvNfpHu2/FtwbtRrAV+/C8d13PMvhtE1rVKayWreSGcXyCeAUlcR6muoFNCU5
mCACAUVnsdTz22q8fbSfcF4VvBF22nX2kpxQ0Rvq/ggP1FbKOt9CFFA4QnRCw5buagCxn+Xz0A2l
2YCxhF2K97GTW8TWbweNix7QJ7wtShMu2iuDiRGpaC0pexJdwNmpIaUdWaXtnlCvoFtln88KO0gG
Iqyj37PeDlFvC52dQ6DmLyF5B43LmHJ6pouFxBzsS6nFmj+dG0KQc3xepk8FfVzRfTLai2Gn+cnd
Ex93X0NSvf0swHemsLTG3MGHTIb+jUlhuKismf1BbPmNVcrkmhrpF+v3gzdOVA55ZPyxVZPMxAxN
LmBqMRkiA1nlQDYk5/KR4vsOBSC5CIVrAa7IrPU2YJa3yVmHK5Pzt97HdjxSJO0AC8fAm6EV+fsT
Pil1NHk+yVal6UwRD1H3/PAfkwuxtNCOLK1XU/AGHPEnTGgM1m7CfdIX7alNlPTrsjgrZlB7J9n4
EotnEmtMDB82U1KQA+SPKPWEueBWk5aiUGfc7/wG4knh1grJ4uVHZ7rSHWqQ2DzrQ6gbNKCxrFFK
0MIv3cniD6pa5Vn2FeELlmv589XOwjOswWuPjgmFlSdzt6ZBdqA7Z0U0z2JZj6d4OM/hFj7KWcNf
k7qv7DIg1kRowoxQ6VBWwsvtXsJEbSzoyyfRRbkj17GOXc1m3dFwSNJy9i4gR7bceHLkU1srxt3N
6pnAoUgu8hcfUvia1MsFu6Er5m2cZtJBlyb6VhbwRJJ2DL+zFWssmCqlVMVE1SLrRaH+70iWujG4
5iBqSfgpEkh5C5JvqqAe3N8vmE7xaSeefzaa/dOPBLe34GcYn+HXeI7FZ4bS6+DNlmiWK2RCcm90
kcUBBMQ/TKUNx63StbKPWNYa2Se4kO22N5JP3zmhAaAy96cPFljdTiyQaGtnC5UxkB8SQqxK4etj
qkiaumODy192HkqycAGux90VdmK6NoWhDYy6tb0hkBzPRxnMUTokV9+iREQxQ3L8ot4S7IJwu7Ds
vcLH+wdW925mZgdH7d1hD3DEFoSHRGF4RdA2EUCggrL6ffGLx3y3OjKH32GWDR1r2dTGCiOtQXnN
2Dq+zr8yRQ07sRiVhG/YQ1WLttwehJqKQV2NzKfDQwSaLZacnClOan23EdwqnLuNIRADt0ueXZ3x
UxC99ztWTRO8KFig2HjowKxNLKh63E+L2dxwaxWqGCm9vLIwFVQUTRo0LDln+kzNpOIkGiVOW7td
5xISK9/EVvntMQmzHT/UUUBvAuOxdtVCly5DewVzO2QuzOYvtEkqCOhRYpcBUfbPDnNk7xSrZXKx
3wKm4QUd9jfVGTOtGfKy3lizkmaiYRrRd7Ub8K5dyb69yQOCFut38SvtC1wTNACCjx6EevqJD5kN
xKPtZtB2K28pwdWSe5vvHH3X7gDwvyNSV3tmklqMjNejD2Soqgf7wzVtydP5evfB3wX2a5yedU8D
W6Ht9qu1dtjkh6HETFd5fBAyKGN4ZlWc5GLBoqDY3raOUkl+5nNRd9XJEPnJyMjxyT3Azs9shFpy
Ukm6m8OLBKD4DNfX0C+v0KHEqr0WzH2JYii2b2WuM2IA0zB1GQwq+yHRsI3CuIBVeKdzqnr622Kh
XBSb8IhMFa+L5OZQEsbJj9f5qfAXhduUl4p13inTbj72jdMAjb/aONj/LOdQ1wrRTv+cXIYiNrot
WdZ/i1+KE6ZDBf0pEZQwjJLqFAKwFAq1lmkKer5MzxpwOeofEAmL0/PdS2mg6N96pf3TjIP0M+PK
a5WXzbnZ/WR5xhl7N5mD9yHdwQD8dRFxp0zFkOcd9iehECehCU3diV03xVev9HIxMmIeKhb8RAsI
tD4gzMCaLw50H+xgh2IdiPXFJ3120WIQdMqLbTEfnEDd/RQsRIqa+Y+EIETETJV51PJJU3KIOtoI
OynAmmr6mBMCxq2Z/B/eayeILBYfPe4dgyhqwH9WjwwKpbchRCZE/jAMunPFD5k4zAg010snigmb
yDOGEKX+8NLEFMnTb/mGBChxmJZi6wteCZNPDbgkWQdaeT4nzW6WxwsMiRwTkKKB+sVTaDZ1365Q
8/tga3HbLp+2n9bBCONvy1WUiWlv6spBZ6FH2yLYkrN4qAVb6LB7L82orkkoqVsC0PB/wGhGHl5i
rGACMc+BmYCh24qf/jM+vit2jEYF1ECn8yWMYEBgqcjLWUMdtxDB5XSjWaR+4g7GL87Bw2wRO4tT
E5LEQ+7GZ/l0kR9Q99oqGE6up4NFU0UartK0m1/abaWCmCp/tThiXlUnFNQJ/iqr7IfIAmD188lB
BqghRjwHTkaEWvGUzQJXKiGkkISmSaByu3Hk4CMGsJXhdx9QLXgyk6pjPG9qv1ZkUc1Gz0sd8+Qr
Il6VGFDzKtaa31HQNUMUpZ6/CeXxRi+XUwCVoKHQVjweKn0QgBWXgULnte9b7/ze8kcIGfPtwPqh
ODUAsgdcsrtRDDXukIO7wd5ce6u27h9gngLiL6yo78NTnMCxDOryoAZLQf7wY//F5PjwvyOd60kx
B/D4cy+u3uqzMxXkCgr96VeJOPy/ErMJK6GnNXBzDzpzE2TfyKsnuz3+CCd689zNXoOuqbL2COJA
lbuoed2LavA1XmO8iUDZzo93UUmaxZ/j+wl16/w2qGI3nJ22K7w8HEy1KW+j94U+eXoYgVItJCb/
yhJ6cpHtM/JYmdRavlHDjEDGYAWOZRvzZAzv2CqEYfMwLpwkFLswlO0Bjtnozhz1aC5H0Xl+HxuX
gPn0HEnBXx6m3ibgJvyvpjZ2VjSxeMjGVviu4De78Rr1/ECOleZheJowTzqBYX4QggU6OJeG5aeD
Qu/GfMRWi8q8/iGi0KBilX7f7k2zmhudiCw2NJttBsu21pBDUxigd3hKZ3acQraUpLqOpoeyZVao
7YgPsmXiDuMOqRuD0qcfu8icUma6rEYJZv1bbXAkD+PUxjzCGvNkfS2FeFXkqm9y4VX/i4CiP8Dg
JYz7FrX5iycrri17J3gclJSW1ppoVwXiECEKe0PAcb1ej3ATfoM6eeBSP+age73RJ2WcoFHbEuqz
rJTE3qkuHKC7Cu+CuJ3rjfglBeKECOmKjXurTec0zU9hcIl89KifFtbkiq6c5UUuhz3rjsekWRFa
8OtLuN+XSVhAybg+ISCWSJgXtkogn4Enb4dAuBRqCUUl5GmOANElVWi3eZZHXlzOAKmmU5kXfvTi
mqlXdtgpVOr3IWG5dg5k5VokzeLupYiZqiwr9GyEV/wJLbRMZN0Si7yMc8sBHXZJXJwJFcoDpCth
nlGkdBttLuGxl/E82E+Ul7bNtIDdSAsl1gA7FXE1wW4FQun8w8LMZCghQOewXuy0Vfl1eBYYW8TS
8Z+GerkxVxmMse/eelUC5WdwyrZpjzbYPUl3p2HDo4CvuP+wLD0W9MEq/nDFDThYCEXo9olCBjL2
scIooIPW75x0GgP1tjzKzkb1QGYRUEe/SlsilfntbvxyqiAtrhu7FspJfj+bwe9tIZ2wjTdIyvBN
+RSU5dYwkgdtwEMB9LdV2JlCHN17UH70HjLzTLKLmhyT1RD9K9p0tkhbRS9HkDsFHzo0tST6sXSo
Kzw3y3cP56A+tNKJLYWzZtNKTeZb7iZ0FuZG7eFTjhdBJilX3ws36vqwiPJowzlyF+439bTVh+kA
BVaojomk2a6fWznzRsp/KGo4NZaJGvF4RE0m+rHCEQH3hI310D5CRgqj8DFB680Kuq9MrJijmXFH
/20Lc8LpJ7D3vSsuCdkzVytRNYccaFe86uVN+aATE2+WkBPCCoo4u14FNUNATxbjyMlOknj1687Q
eilKO2OtUoA97XlSwriAdz5fKYVcHbWOo/owG4GxUoQLdoL+OieVrLCyBdxQ3dooq0ypYha4dZkp
MuprETx3FecQXd7e+or/Z+TIxX0uL4AM00Lh1xFpkAlR7G9CrJKZ3+p+gnkdLUdBOUt5O17E77+G
1v0vxDDompEk7Y5G6/1Pk/60WdmM6vicLgc/MR9Cgv0Gf3ci0PrgHo//9npFpHWwsctgVMuVr2Xo
0SymEfQyfKUL7GyrVtSxzTLVr9p1j3ocMCJR5AhEBzv9PYsrczEuoEgSlsEpNt/PINREyYCQsl1X
ptWckIbiGYHkKbF7VWZCQwXXCB7vhHnIaHTNN5CvpeBUJyoYwvmX6GnIUGXKLBSZJ43rOFmyxpJj
w9DeiGyhENXrvEfEmNUD00/GtDX5WSVOZZxH31TaZbgEivh2pt4U110fJ9FJ5pOOMhWenfiJXH+q
bNrAaIfLu1aTlo8y4cW+GB48R6+L7WtYNjbJCwSWmVOrWX6sUwSLwae32O+1XfxrZI7C4vp7Z0EY
BQkz9K6z3NviTYltWFWPLXJsC3rn4EqSMCF6p0+IRbCtFncWZKoqmLr440Pn/2qcValtduvi24J5
mgL8KaoYdbpA9keEY/70gF76xMQZrhHSg2ZRVeQZjdLs2T6hdXAv8p9xyqdQGbQtOrKlzQHmixCf
9v3UiAIIqcksqiNMQF6o+FMn1vUB6LY/YTSrzJ6Od6gR9AeY7eB8I36DcjqR/utCLU8YWO0dX7LF
PteA3QjXN78b/6DvMvdmkRGlXD2HCu3VUps+x4y0eX2qYifgRmiC7z8DG1/puYIaIAzcYKSqFqWC
wGW5R/iwezXU5CULSMEJMNfRP+HN5v39GRK2ws7Goa63iraGGiNrmmky/3+a0/h/j6rxXILjZQCE
Df5JwX5ZpBs0G4DkttEY4vyR0YBX0x6YYo9wQzIgwCg30ujPi9l1NFe6H2VPDACkBEY7lQlV8ycU
pHqzeCXoofph8jk1MjzxLRPOZcF9zFeY3CS+gXa5w0GR7UrertqB0DHb5LleUL6ognOihTjmNafW
qt3fO+TQbgl9DtHzMqUVf7BRfUp7Da4KKFfLSw/GVfOn9jIobWZQSP+BHzD9czhZKXKp3/jvJ10r
tXbLhNNNwt1hxphog9SRPpG2ONgQqT7cpPETkBaE4VYx72ZpM8HOMWi/umbgkZAYLDMVmioPTCTb
XxqhD1ucqQYuPedTuTP9W6VUhG7m3vMdJu843KCkBTNbn0/Oqz69WYADxeWAssH7kirB4YN8f5Te
z84vTbYa1RVDFtJBevcOSOrrgDIpoEVvNTcUbw1uvA4myPe8BVWMphnIWq7+CLfHW+ZzvP39MdG8
c/VlNPls1hIQc5IyXiVj5ts4rLLUErwGWbn6uN5ZRwyDC/hBIVeIGBFTj+1Y0IjgfSYY0++UF0ic
it62QjindLK9lM9VIOqzmcYqdExSqzzRJVBHrjpA/T/ZWjiCOmkb4E7qUOyyOyhT7lmHOFeCCbht
fCKehh3GMayQI6vyemaIS9j0pJUbLkL2rwpJX8FdK/XiCRKLNMcYk64V6VLtzsC2scKMDtm6E8Xw
zFM1NGJUMxJp3U/vTq36MJLz/Q878cTdEUWUEBYEefo/HD3bIi2gUjPoiTh5cS3Y3VtJhgNFwkuY
3rxB3JuvFwbZ7XPjxb8EFTzxNh2aTX1G17AjUGGGlvRWaA7bhAl9abu4Zz0OxyMr5jnWElSTn+ym
sP2i4nCbbYKShy2tQ5vQhDJlzDbeENkM5teCVFKsatqJmR2fLW4dKtZx6f2R110plX4+oVdFfuXL
zdOXL7GmnS9BGLxJKp+nTecTGuHyOUFGU/MCjAcl5WHjGBPPxkPdb7udw3M0i3xue1/4AUZ+Cuup
eaOeBKsrmsMwPsRS0KbnnXTA8ywyywzpfv4YSV603mMYOW3tLFLqQqgyfu45+aviCf2nwMgcVeKW
Gwq+igYqG8OepIqLWCXa5Ed9zFN0VpZO+0CNML+mFWTmA6gj1NwSkvPBKICUKqYq2eCZX7EeYuW+
Ju2JHoaBzM4n0CJzHeuIngbHq7H31BZVXat163XAfAmLthq1T/W4VpLRTF45c/WTsvFbG5j5ae+i
BAbUUSxT0paWHiSinrK8WL9uhf8tr78Ab+JKfTvTq/MrSYGKBfw/CzOBddI18ToOS8IwyekAqIgN
FlzFv+XVZ5xMEixuXSGAWeiGR5+W041/xKxykrkpqV58yPgL+5ZhXodIq/6+RrgeoHAUxLzuXJo4
iKlxrlZ6zX5lYm6Yxk+zHxkXuJHDl+oKGce9OJjIEqGNNu4YTW4QUIx/XF4kTMnnYTCHZWpywhNP
u79fKkiTW6UfzfUXMYdbzY9NB9mQ0jq01XBzQSySA6RVa5kGZCdFxaRMgJYGAmwEDBxNH7v+mAD2
i7jymtAKy8eiJCpXQiD02gRU2s0uE5O73rVW0CLR3qdq+CY1cKg8kvCdMKEftCUaCC+MLRM6Z1Ya
cRxTiK7su1hBg0PFP9BSJCsjA1jw7tCUMQcRWRQluK+51LQxMgSaYDHXY8Y1b7O2ONwL3fqwnbtL
L8LH04vsQOG528elIEnGgo3C3jaPdAvc8NXj0xTI6XLDs0PSxpW4oYWHmYlFoAk97qm+tft/nh2z
CdPXpi9iIUKmPNtlBZufgdv2iDMZb0f0QQvouNiw7kWOV35wDSkESsK5uFYay+scuSaDTTOPuZo4
+MVU4cIgCN7NHdRTcLXWEa//vn74XmFOa1nUvWCJH6rihMO03Y9H16eLU0AJfgDQp/nU6iSCkpy+
eauf2zPeBdSbYcFU+oPv+hQGVCDClbR3H/X0DXFx7RlAGbjo3MhEezcSEgP8YRuyZ+XALKPFfk/y
2DVAiIUTDnJ+uCFQ8ScitaLtzVgKkpIjnrgPY4C1bPdm2VFKIeu8fq8t1qrduspvuoUouHeUgbim
xE3LZtPiUOiciD9nl78UaOR8bx8HVCwaaA3Ia54K3qcATk+UZLfnXcWPI3AIE3W79lYq6t9OjXXC
qRJLLlyFDeAl3pbWgrnPudqzUP/0zRzcbuZ6FVWxFs+Ld09HMQ+t40KWpwqIQqi8sXKjAuraPU2O
QwZ8C3NYcd+f22vklQ4m2A+C3wXWRyKeykba3jU1b7fxpsXch2JRY+NkIyWkwT/HVM/c2rxQyFtb
vE3/41MATj9bRXnpTN1/eMYeEdrxHY6yaAN5qyockKFApWfu1r10D8hJe/UbTg0WvQjOvGK5MoYg
Rd6bOg7cHaJ7DU2i+5h3DxrI2k9JFTdm9bWMhkoIHQXrW8Tpemf8mhWK6sC/N5KMbnuMtSmTkFVA
P8uLBPP2NvPTTE1YRtohS/O0axFgaxuVjnhXMuF677GC65IF5LN+s0/vdE5UAoBVa7tBvV4ixpqG
o3FQGZ+yEtZv1LriJO0RisbFkCHXYvlYSS1ifiYp7AiZ/q56xLsPuip6Zzc3G7Z/3wjKvtYvaYay
MVE0dXcCaA6lhQRVfPbIUQS6I9kyuktjvvlb4VQOHTXVDqsqLZb8ozH1e5WkURNx8v8ktTZjf0lE
wz4vG3WJV0BJ9LXsXldvEwoMqK8RCVictiYdzzQ3tO9FVvGiDQ6XR7/X2eUpcNGq9NDd9FwLmIUv
ohoyshy+8ix3V/ySIR5IFfTdtK2fSdWwj6CuFRQp9MF95TJTbjTfOAHkP1YkITrML6ckppAaGoyf
HM4ODDas1NthGpW1xsGITQWMN3kVy8p+0AcHUC2YiAdMn3UYAR5kho89WoOWURW2jZ63xRVXTtS3
Vfu9Xno2rtiBR5VrjYVXhyO4uTYvnqg5jvSW5KGIGZIp79/SErzLTp/lCVBvlJX42OzGdjJrBIaG
K0MAkhkigdoRqootHHvlg9K+X59xmR62JzChgCHtaGRqv4lw6vNmr6t83xwg+mt3XhdGZ2RzPRpC
HeoVRm6dDDCZnGSe3EegKHdA8afAVdihp/9vR24+y3ONP8ai4vewiy6qmynas7rAW111dFPeWljJ
3df7mZXkReVkQlTGBJaj1/JnMmEa6STtC7ThCpeXzaIisjxirqdP6vP8eWu0oswesA4jtjIWpDeG
7lu8lNq2sT37yoyALWvcpk0hdpiH0z7R7oLga1gJNQol+2MDo8wT97JrQ+ylqPtSxtI3Wu2py+4a
PBi6SrAUIJUI6U0NW89aiaGPfEs6NDjC14OH5aGD2ulvHLRGujMc3hjX04HujsThHY8Gct8SVZ7A
iOZmNYzC3wGuE3lUPCylRkr1laMVAImwQmNwcVx0tVVgPe2X4pHcpTJx7MwzrcbIek8dQSG0pYJP
cvi+6+hFMni8meJB0pTR1RTWYvY2bCGSa9Ek+zk9K47oeMc9uQqgqQkyJ2oVJJY5kcg4cwqa8OlX
8yQlYtqA/Zht9ugnmAowGpqN/2kipJy/ABBexa7ahxUEqLl8CWDLk2lx+WAe2qM8/9ZjrZ+tAAPE
zGcIk/IW8WUIbOdtzi0Y4NTx0E7hHFvOHKgqIs1/66oTtfFQ8zg76VidNa2L0KVmUxG3t2PjK317
+vC/VwW3KHKRyGSw3HeqIJrTcfdNs6Zilx9b//CjGkD1nB+3TcY/xR6gq5VJbhHB0qNE9Znr6oT5
M93B4N+/WCvrj/F0k3dw0IQbgvL58EDWOsIED/rs8TtfiOTb7zL2a8+wfIxdrAMXuZxcEKL039vk
pVMh4VbI2h+r2rNX2U/am5peWP/C0Ch7ZIk7QGGDHR78rCuvn+9S9w0R8emIZx1x1a/KH7fZi4kf
Q7C+YE7Fa5vd4ulO6w+bygX13mslUWJ+bZVuCvj5KNdkkF2t4yhqDteqKm9AEirZPVmxBi2DeNmG
iN2DdN7v+tJE8+ojqQTKIcG+9nGSvyCzG2hVvq75Ce51oQSYMTI1HZ5lLahPC1e+jbDGnVFejUFh
iaJEHjSERJXphRX7LeJ7hg4xyGMZa4QLnIVi/jQJFsr8mcOwpJSvH/gAwOUmBrVqI6McWiSr56t+
ajXIiuxyyLzM+RG4RpDPvfNSckZLAtDvYahbO3Dv6Kg4bUOt28MYB9+MSEIKmUy/2T1p0GedMs2+
uOJ1anoQzbIHt7PEgd/56A0QV2D/lEaBtv9OQQH/Uiy+saK+tluz4vSrQjOTz5/XA6E+0qt8F59L
+Xz4L6ROMJ6HUPfEVp0jWBtrkMgAoUxD9c6ad2D/1wtDYd7sRYljQbpTbE12ieEYQIHIQtm6ZMcs
brVj8L8qUVNSrewvtxG7UUOGUnM4/d6XKbn60kW6ZYo0DZ4uOjwxlTKkq3Uo5ffrglt4QHXas+l+
h3l/FjT9x/KXGJSYX0z8bePIG674DxrdNAkTPCALxlDh9/dfQYgnt0FaBMfBeowvxWFi4WUIJU4y
5Us0x+O7cGYk9ANT5son29wOupb1dNCRXuT4YcRQ5m07fxl/9GIVU4vQVMy+E9wug6hDrStvtI7f
0oRtae3yyuYjEUaD5i0/XfAuERe+atTr0RWml/cICIl/ywmoat/1DrQrE/1RHO0W9n/H45c0B6mu
ziNJ72q7GNKiluBB2+0kAnQ8cpzHFJFOUXOZNJoIzWAaz8H/KYBiPo8buM5inwehQv5/RL40594a
k/If1BLlJJ5q6CdWSTKehRqnwzkEw/9Eefz5NUra8iiEs/Nysmd+DHifolxGUwqCNQKS3zCuo4rF
+Sggph4Dx37vxZ5cpx5BA6qQZo0ChQRdDyGGz+SFtHh+qDYBFGjM0+ZIQPnx8F8bkMbhPHl2+jDj
OugWS72Qt6Xebx0eW4J1qzxgbn3PkE1AgNhorvoAoOulGc6ZGSrdeXMM7QX1UGz30rxX3yN//Iq/
GdAvGDvfCvyIghC/9+lybl/Bh2Re1mKTMbBbBf563CRyXvmJhOF323vVabFnp+0rJqeXodA/RDs1
BbqN6gQ0/FPY7pYVfDklEmxtnKuDgHbc+6qY4THY6VjnJLWWClZWbXGFgZMtKyjiQwdd1x3rfr4z
p5Ln5fT/5r3kL8u7Si4ZJAgKMwy4NGnw3iU2TjjRXY+gKyrmJWmmA95tm/egJ03uDdIDE2EVK1Rl
WaZy7t/p5F6d8hJPKMtQMHjq86JYAjac+CgbbA6bipUgpJ6qcZlY9Kg9yVZZC4m1lwoE4cb0SN/b
HQsyqRBWv2bC0nJDSoIeh2bfGL1L5MGLm+sloLNivLJp0fVRuD3CrVgBwHVtKDk4rMf5LFvTpS0o
53Q5jUngNQgSkPvV7vyvmwiH7msIgStVbzFk2xEIEBuuIqIocT7dwHO4rjypT9ygkYlGO/RM89t6
Rj21gFIHzExyRt0RSCJR33v98MgLKXEIU+2HA/oqKHR7HoyC/VM56aOtVlUxF80w3goH5OXYvZMp
uCKlw7M++Tq9Nc4yhBRYxjNmJlxE/WIFMpGbTEe2V7Vg8k86GM9UfO+Pp9R04qmTZkrftXEVHel4
95NaJqkC8gKNE/aHg/s0JgMPIYfla5wn9ft69QRd7wzBjPyWwSOHVE08ryhZK6GTU/Htq5i/+DEx
sn1ZMs1yWLNRY3h5pGnGEdxpvIFc5Y4U7oCpj68KzmnHZcAkWekxIk2hHE/1s4HED48TPWPmc6gQ
7jvNzXNXEcRDt3jJfSchzkf/G96S6sB8fo5aHw3Ff28ZYImnk2ln0r9cgib9zXuAs9YJabGoeShY
h08b8grhAHAVXs4tqyvxHU5R0J7pdpqFqBF7OFjDLdc810T7+NiUIXmsLdBKqbBGRMcr5fTF3rKj
wP6cdiBBv+gYdGyVeLjvQsIpxmYB6EdZulwuziupywwaZXb8aZ/lhRj0HRXkP+xpOBjB8UQiVZfC
ZQnWUQcREuWc4RE331iyLfp5Cl/y/jPUlL5w/VtvZ/a+GzIV7/1DmRtO3GOVExj4MFVKqbOHmjXH
cvDORhrlxxHkBMutbjub4ELl5ReI9UOejKtki8f3T8t8qwilI02GozZGTxNrohWHspi8KXR811Qw
SUIo5bTo+Qu/x3g9OsfNKDYfrvwBtp2atyzFl0GIRdesXW8Gpob7scUy9XRGB6P4Z8KWsVm01Z+M
8okg5IN6Sm+NyHqQa15o54fCUEMS3ACZHO9/OLe1936R1PFqbLU6LFhVNwcq2hp5o1MNcJit/gfX
V6JS81C7tY+oRQ88grGnqJFVYAkc78jZQeJTy7Lobiqy33Ft/jnRmbx0PIm2rti9/FdEQbPe5VU1
0X9RrJ9bHWgo4h1NZccSSUo16Qj4P4f9a1Iqfbfn8XeZf6bDXu3gLUFkekMw803zm3Prz2PviJyn
W24oTIzk9yOX1gnaDRVf/Yjonn1cr/SZlSDC7caKFlKgSSbvTqhayOAE9YRXtO8eNnzXVfDVvamL
2FNNbQNG4gNUnv63qKRP0iUSVnpK/t4RSQkDwe9YO1ZSd1meZOvoWXqdDu9zK3susDpKVHaL9ueW
KIC1JtY7Y/PcdwfVlJZs5xV62V2bzveJvkfYgnVee/h0ydV8XrcM06gOlP3aqn/lmsIn/vUYVDAY
/Yz5W4U0GYaC0QfHGKdBggupTzqcIW9q328I0LDrvtTA63zksjHVzDsvSpvJnxmYsJNwc00jh2JE
tfkZpTm1XSfFdslfxTxnKGiXuqLpzOCzvHvMAJjQGTJeqwsKNPpJo2SZDh71qZG8j0AE0oM/Wso+
Zb00JQ7vqPha8CfrKwIEaldS7RQeGSA5YccjocIHqR+3yx/9xiYg62yURxRc/npeL+VMWBZHhtnH
dXebUhKHEMXQraKsmvP/wXt9lPl3zYUTxNFr8ZHZHCmO4twccR87c+Q5ZaCAjtwAlaiEKC8q/E31
ByagedXJgic2/xQlEII2yLqidcrTx9MF4wqKy7WjkzdQJXksAl4GXBjuITiucJ9sFB9DKpH5wsbn
mTl5BtsMYUqY5z8/eTQ4Q/qSEvoMMfk7n84nfAEWjqtyouZphDiTqK/cnJmWNHXSYmAA0S1yDsM/
4r9E+buE2FPsCnlP/1yWwajZXGWVgj59iLux8/wdLwZPOQHkq3/6IZbh0n2bK4OhVTagca7lVzvD
nZ3j5FKecQ1Ixd/Yd8DnAVTREkoMC4JvjKls5a5lzUAadhPWXsq8g1A23hpMrJZHEBibquv9t6Fg
HaHFndJubFFIQMiYZ3QBuPefqYA6M4Oy7YoOEHPdi9/jVBXLuDBR+RBTSb6QOtzLsjRyXwGXJib4
9aXFpBRUu/8/vw1YGHy+1rhifPfoitWNLPb2CiDKvmbSSl84HtnwNl3SkgbYepEuJWi1eQnccNju
Zm1Du4yvxX7XBrD1FvS3axuoiYv2xumEZ7ARQnBnw99mucFfZnzF7Ur07x36ZoqFdgfFEEs9VO/V
kVb42ybyr36YUCZ1lpLuW/dEITTLuaDsOJuqnThpgTY7OG/Xj14OAQ0a2UTiN98nyLvAEem9+45Z
5mVia5TV/hYioTpGK2EwBiSPWoca603W9hMBTrNmeRmGM3aVGCff9ABThPsujKtR+8xSfZqLgnoE
j3lojPWhJtgfMk7NbMJGxgwYkczJegQW4ReXtZTQWF6X0axchE2aku7p+ec1pO91XCpXW5OHJQB5
Hu7BkV+VKd4q1XZAOdmBYm7NzYWRsO41O1G3dcMzCLrhUqwXntW8s79G+uMC/Y4iHlPpJ1TbC7k4
p1SEkMVqtVXCT9fgZsjhZJTvC6nOxYyKlqSvarRH4uinCbpjx3cWWx2NYGltGH8OfLaB8aDCEta4
FlLaVwxfwshhrxnhTOSx7AKonFbGow6/Nz+qxo69vmUnupFcO9J+APGDuGDK9BF2OFMnhcCDaZFk
HzpMsE5SZgOXPBTPU+WVY6gwvfY9KvzhnfNNuufhAJJch7Ht1d5a+6MBynTEjz5gnndd7fZhIZtm
oJ/ccR9tXFi22oNN1gns6Xj2byzi9ydTDTr7DjiuH7vJTVqNsdzzfQiXrQI6YtJCEOb9rUEO/ZjC
OQjR4qFZOYfFQM/vIQtnnQT/Q1lCdsNKyh1l1JdLxnsjL/gdG9t7xrkHhJ34lmM4CxVZqHF7r1mG
V7HBvYNT8ma++BNl7l6SoBXWrscqF/kh7yoGYFzgwN0wmPYuQIEvYF9dkHL++/YGMEruEVvTjwL8
rq19als+QCUBeHQsbK59B+MDJsuaqOviweD37TNX1GZPmXgUa+vWjHtNtFhOmiRtfjoi/fjj5MZA
jj10HE3GPPHBKl3vDQEhlcjtg+PBOE+h4o2qtSzylwJsLYc4BfVFS/BAWouB0/TrbeZx1xWPpw0L
v8vTl9v0cvgkFrbEdkyKnKSAWb6gYdqrRRCUsBFLmuiJpdX1uwavrwAnmQyLZVY0gCmnAAUZw7ow
AqTBr2Tg9hy4rojd5ijappXCy6cuP01jw4GluI9jhcVv2QOiUqkIeT2r24SdxRurEvak4D3pAaB9
RYYxjfzGlewku5Am1H9cFPnw11y0uLMG+hZ5YL7sMgnezRT+t0oFQVDMtlFRXzZxAtoolEeJ0PUE
mVbpp4NBEwhXI8C5vMwU6fX3VfGpAvdaQ5+wqYSQh3UToOzwf0YJlEAjUPEsefR1rQ35Jiy7e6Vt
h9q+4fgeQA5NQidcstdi1MHDVgG0uihaixGpUGvzixx7uEJON9RZ4qEZYKGVQFZpkTZFI0mU8rsd
0v9DtC6d1snqbjAz9Hk2HSvixupLjUAPMpCbo7lxtk/oyGj36PGykiOZPMhqh6X6TCmGceCjWYkx
5dz4DJcTDD8NZ7MqLj4jnxVx4sTIk8hfzeFitSAZt9A6t4QuVQNlsYWJ4A71ksRfYeYr28nozt62
7c6MOF9vq+qMIbFM2AXPMN9Xsw196rvJ1WWRNiMnmTU7sPuUI74hp9icmnAGExb1Q6Tx3rlcSbt8
Sb+KZYz17Q0YX25ewf8MWrQT3N4bi6xWcoCubcVudCE2enDK6/L5M+lwExqhtPjxrXUhLTClhDZK
ZktESt01zqYkkHwnr9sB85hPOxfE++FTTrPwssMyN/1ClmP5NNh51aiagIVvHU4KY/oBSycEYjGe
P6s/7oHWpE784mIhiBavIGNu8zY/Zgz/+Jiz9EqY4kL6FIb2b7T+TVpx+8P7duXkRsbtNTZthn2N
WzrrJ40k60NX3X+XKBk13A6VBSyQdE/UaVCWoqij79P5buB0P5nWoJ6LTW/y3+JCX7ycq48XEIzn
gZ6hY9U0SnfhTUZLG1FR2MWMl9iGiX3TihWCxHRXBibqoyPfoRw+XS1U7cy51MvZ5PRhuxoelSZP
dkigPI5sUvzvbQKij5jwsZ0cuW7vGjvbM2EEHFZuIH5bcyaamkd5rDhbZQxCjeWho8v2FJVlItoE
Am9IOn3Gk1RqGe6LcgflwFRL7bbKg4od3lCgD237ECeSQUDldjLJ8bjlp+9Dm7w4zBsQXRpRBf+C
26PVDnXKT38apCX1HSZXXVImGB1FSUeS3fxGCrFIjJjs3BVtYnrx7P8s5RJ1SsdB8QPR7JOnNSrR
wm3hfTC49wS7D3rhpS2GsX+JQVI5Ch+NIaciBkS53mTuYOtw2tEQR1v6zBtL9m+K7vQrcmbu1TlD
baN+DtiC017/fHge59ggxwFb+MDN1CVeMLXeMNDClrHXs537ahslR6UWjNnQKTrIUj2I3n8zuY40
DTNBwAWLaY/mgk4FAUaukU1q4t98MZ95nesnfZmrdQOGLtgduLIaZNhxfVBCRm3qC7smQhryGhZA
Z8EIjM5RnrkqsDn1BNWma6fbzRV8QqFnyfXBAPyT79NRcDyuz1oJ1Og+KTrRjHwZlre3UJfaqhWy
HnGOlfcXLMfqsd1WyhYvZekTEMtcS83IF3HBA/Ru5A2Il0llyCyrBLs85U++M/BgBfjXQ7Qp548n
zfht7EWgjarp3TENMYWpdlOsfyNAZgGohz2XBaUvIsgQF9Ga9y7h9ZpAImODA9iuyHiWigFEvl5E
llF1A94lDTqGUPX7j68KUjpk0uRoPlfNxaI4EU9ZiSTFQaN7SchbFVZSBhstllDO3eVif5jRugtN
lH55Y5VpRtxCF+BEGF0Vk0GZATOKdmET9tjRYvTdRikjoDW24JWZzOevD9lvWq48fkuH13zpGv3l
+OPE2Kt7E2aYXOho2K+rHSeo84r1ESHKeI6Yh3ra5cvooIfl6LJRYU7J4soYrqcZ9gsm/i5XTZcN
vxviXVAxuJnnaAwlmkjYRNkdFrIh6YLmzDSIP7Va0ot1g7nwbfivCEcjdun4PxYLG4IcTgMv1Nzj
rGruhPtOg8pFaFpM2BVVnsuY+Z63e/N4icAQP0p4ovdPJ80Sn359V/XpZqPFb/PU1FvFWnrbqqO4
BOkdRg+KigF7F+JcAFEFRM6aY+Y2EGPqBRiWwOC7IuU/gv+Cawcj/oN+oygqrkuBCAlEMnVhmR4o
g9DakaJzsafQvDbXxgojsmwyH/7eskNKFKtCbqXPYCJyWipDwShdsDJSnY7yTaN63x9tDuNeOOdq
Q9Hf1t330+Kt7rEoMdj4Etz4JADdk0TsaSCYmoQTfTKdjleXYRA1u5JLEINfJfXFPKEFJ9BYaV0B
EPs7crwMZl/S5gcXN5YtdVLQ2xvHSnJ1JFRHxB8Slac3/5yUi/fOnij7HOQ//0FFkvAa+ppp3vS+
Rl0V0omMjMAX4q8LE6clHzdMBOVtUQrE7BmJz0kNKfnMQ7MjWkh5dAykSSaH9OTaPX1RnmTga4Mk
y2DkvAqtDoNjzqBN8PLkm5GBDxvJG3zM3eZeF1XMiURaYmf0Dbx5ESy6xOWd6863R+9BoqPGTeeT
DBHf+YAnTzJx8aMTwvHKpjmctFv0vmUCAoiuo99eNjZfe2Vb8GSJYahHnRFOvxnSFEpzDFSdk+rx
ltnHyQlpaOS8CxJMw/wU5AQ+0c+mCOgGks8jXtG/xE9OswH9p26j8SuhkVJL4eoTqveVbRXUqQWf
OJGt7ULoY4i/o4VLpeiY/cVDODyEnLbahftx+hK3owAM3G7sbTQCHYZpscODt/YUgxHCAQc8YKIt
ij2bWmMfBAdqJc++LK8fSE5+eda69JqVtQCymIkzVNYIFY6I4ZnETPLe/c3NRRArJ8XJgBmyWrDT
VOKZxakz4M7c2N20/9udEJDiw0ykDR3YpgqOIS6rAQ32G0MYUsgB3eB9tA0Esi8yoiNrPxv7rdrH
kXhvbWk7D2EMoXFvx1FAmH06b5ObMyD0Q6qNPWjckO5cwBql7vNnPC/ksjZIZBoSUUk7QAiPnvPA
4EXDCQCAAPyvNlPeZNqlb8lrSDb9YKazNl/2CReu8XlM6s73o3pN2zHe10Ff1n2sATHnJ3uzkkB4
nPNTY5wPUpG26O3dMOCGoJZr7gbbLfwTcPcazNBTbZv5IQ5AcjOjnqwUdHtyyT3xQZ2Bjg9Rf/1C
F+zXuee4NLWXxJ64uVBcP5kHlyGuGsxavkPg3yinwiizu19omFPcvyGcyBpuDFXDMImpaHqMrGg4
cINz4MX4PmsEWyiL4OgycU093XbFl33wpsVTVN2ct/PJsuC2rVjV6abhxPz5yEANK8Py1PuTxIer
m9vRKcRcfpn8EwQQxH94Po7746gzjyoJkgz/kMT8VtKJe+DkdsDRrmLwZq5LZ4qgUmDxdj2agwPU
vBEGkEYTfG1oeZYtF41N/RzRk5WQyrykfQetP0BVpqcdZEtXKRxXipVUDEqZ5dH0MiLLaVXsWJMk
boWzSTm2gFtuedHaJ2FsMnxFT+caXVdRqCDQbr3zONCZ4y7ARqKzZVp2hgBbHxclc79eKdbG4ux1
nqUtpTVbl52QsiaShIYZzznbneGgG9aIxLjb5npBINVUn83V6pOqCS+8UVVhk6wq2bEyUUiG7ZPX
gh/TiAhvC1EPbLZF5H3wgFucCncDdYOUhTk3G4zSzACnhETTLS3Je7/Y5WzjhYJd93L9CcCPuKbp
UcKxa+wQDvlvMsp2ymLuM3W7HgW/NySmVUg84swkafu5DrXGytSgUN4+oIZcH3wV+AMdkacaKoX7
hd9MGbyofmn7yudcLXCXRjWOf6j8HjfA17jvrVkPyy9uBhgAR+AYBJEJVopdf4nxaMj5iqo+a71s
dmCsECo5JPmKVqPYxCJ6vQirRhZEDUs9rb/o0swNtuFzQEQCW5be6ac7fybX/TDEteqMWZYVleHz
NQp2GmOGzRt6qicyvf8LuO+pGA+nbv0s44B5Dk9fkiIFab8nT3JF4UohWF2ERftnlk9JMtqN2YsZ
6L0W/OxBUOzG87t/nmhNzp9COFEJrKbNYoO0qrw7L1xlyjWG4fU8FS0sBeWfqQVB6BH/BfYwkF2H
xuZ/gCscWar7QvDz15012dDGOpWizAN3GpSZqT8eBZmp/fAuRsgs69YWJo59bVSgwsghRUeECnBF
nEVU+wovZsyV6ukXqq3jOedpAcowz3LBc5+ntCL4qgoMU5qUkL+XmjFWre84IwuZ6JybkV9FA9g+
/unwXB5apn4fXB2qw/jcB0Qy87LKm32MkghXNszPd9LAa2y+s0OMBbKSwg8z15etD7RmuxqasfCB
k0X7TGEWoQcITSAMSSahKzIdXEwsh81S5uUIOCWtwzh31cZNmeMXmUjvuJGbYX9hM62zqSA2zou6
vYCesIvNfVpOhPP01WHPXqWQ8vsYFzQJwtm1iYF1oOfwGgVpdIgSwNCMhe4Nc6ouCeYZh2R3vuFV
TYkfS8o8hnrOBvLEXamW3xdsjSUytXEEz4EwRLzejdqVZgDl881MjB6GS6PtnXfgWx0J6HCV+fY/
LpD5k1E5DJ87QOVKrcHZTmGOoxk3zdLzxcOY7I/emGLIIyNhVnrpCoTYXjtXn38z0IGjAeGzEQLx
8Edc/ccWRHYIe4CyH4KVzM0r6AVuGDm71bMbSCxd4GbFKna8u2cHN+jCpTFeW4zbtBx//U6PV0Za
f/3plYQ1gRDHBhVpFoNd/PqIAlmKtl0sozEm0EfcNGAVJnODD+b2zH3NNN3YyQu4rqkHPD0lmcg/
iu4aYbWAJjaQos5pYMlREkQtnHVLS3K8OgrYvZTbSk+R+4J83eSLvioI9Vd8jjQR4GDulAuQ2sW1
FD1U8JP0MK0q39hmUcIVPytNv5G4zRqocBD/CqIBrV8FWUYk7NfLPGqZQzYpXc8H00sElYSp9Dsm
AvY2plCOhbZKCbULh8Ifu4ltoNEi9THHD32mtzQgJZ00purzFecHYJSldl0kjpwvwowA2ASB+v8z
jsrrShgRoIHFS5yZWZNzgOPc/2ZOxc/+thb1KogVEXh/s7GF1jDJWnlBObDwTs/9BnGA8n+qX37Y
jPrhpZpzs9FhMjaG2PPLakiTWjfpvCl9qh93GwedJ6q0SkXAqHYxDna87Q06IHxlpLdMmL2tSkAi
4IdTKt4FdwpCNwfM3Zu72bFDXw0MAFFUv19/37oOC0Cn4YZ5UnSFR02zFIvE4eVneuAiwD0nHmuG
H8jIq4twbIWywIc77VyEpJ8uwODxrqSrujPXICmKzn7xDlgUYUY75DzNK1mu23ZwqwIxwM6fJ6PF
xRfRDcpziT2RNfOw4Ayi8YH2BxCbObfp5Bfl4+yVtVau74wGFtegYY0zbE7xU+/NTbfi9tsJ1i3m
S6O2PENKEempB8RsPlUUsBTBaaFcl7im3bYRS/wDk6zMqzg01RIad6O94QbAABSIAtzNsiTsr4FG
oMMLDZP8mvRoNCXuSFopiLbWtGZpAlAVQ0u+8PhozUk2Bh1VdagJvq56lIs+ZH4W/s3dbluwcDe2
JvMu4jVPG6rZPH9KlI/cNDrReV65NQvfTixOSczFXG+w6aQ2SbqxiIMa9GvMbnfCOCmz3RYSplNY
F96r+P0Z6Cv8MCEvEBCGwgDXFJ4MRkL5Tjfp+vGbuBncyOCIsQdpkt1Lh51YTSoBIJMUI6X5zGAu
RPiJLyv7yMa6I+S3xNiBF45SHl3qTtIBi65POvuugLGnUQvGT1y0oeAV97+qcfUKJvFmcijBBrLw
yUcs3v1E1upb/B/5vMJq/yTGh4amxMhEJRoyqmW+cHc0/WkJRJNln3GLTa6U9dHXuy/r7S4QITG6
MHJ9mqRjgN+iT9UHsM7Un+ji9NpL5/XrQsN/Rzzi3NeZAMeB+oiuG7QfwTbbFomqSd6raUoYvmsp
kyO6MCqrcu7ceuP2MS0utZTnN7ymCtTRIqxmoRiU9YW5DUk5+6btK0Mi4aTJmi/P487S0eUdM8JH
jNuK0NzOv9iVOPJMsQi9IRTWZ8yl3zQTujhUAnoGB78+7IrcsP8ium0n8pUt909aBD4Ngyxrvkyy
VEutOkeCL4jy6dBkpRZ7CDrjLKaSDOU596fM7Ysf9cTT9DkrauC1n2/VHYC4L66kTSmUMd7aFc3c
1D4vbDlrzclFLDfEPSvUxnpB/DIPzjLdNKvcEBrmxnNfzda9iruDCowybJ3HQbeXsIpWRoweOe3+
3hE0L5MbUMHEnGOSa0dWPXQcoRJ/PYfG14wxVmQ3EZ+VIFmzFmhATsKNHict3R4cnvFCehDalvdg
d1p0iYQxghiWmEKaH6yaUn5d1uELW9g32dpPm7t2uYHHF9FzhCqOK55OErBEZ8J/LZ9Q4aat0HYg
tR0mDd+XBdSwX4gsfxd9D8RuP4heUvzKgtsNngXScd8bGXzycH56XV/h/5F2qt85zb1z8l4diMb9
JERbTfQK1jNSdW+v26EtRwCKelHmTODyTibFh9ACHfLYsGdNHf7DYEW+aQoSa5Do3LWNiNAUJamb
kgMuAFIhrxOf6UlMmfbemXdf3g79aKa0gZFL1dk5R8tzwzdh3hcQCksEcN/mN6ZK7+4KUCx67c/e
FEmYJlyjwmLTHuBGt+bhhZHuw5ByMvXIYV0x9DZEoTEuIRFS6ykLmUaZQyA5Q3tI2jiC1wh1ZKM0
22J3JZ9YSMFn91hxFDgHu16uITFqVBmB0cCz9b25rjLdEICS9ISmrB5Bq+BWegSDkuPnEDIbM/mi
MHZzBkXeIpWe9p+5q5oHpiuv7SosgiF7mb2PdxCNeTTK+DZYJC5Pph1/XMxu+LwAsOtx3BK0p0K2
84qBiFBF6UrRqfS2qmolLGxaeaU3bdG6KxZCTrz7I8iKAY7UcFLSpSXj/2AGPFP5VM1aPWOq8i1c
8SZvVzzjMJGc/jjYBcFcYKkJAQijFLs1B5eOjCrB4M9mmrMtm8OS6LXadsOR940qNxzsYX/weBKg
qskzA8PsTlF4RX/1IzL1HzLSIdFmhvHjbb/1G9uc6NHNglacOT6+cUZifHu185udiTgsVeHzmNge
ZXF8nMdcP1Qzm6fI3O9w0QKoDIhF5jSZ7ZKwC5GOrUciJr9kp6/nv+ShUwwaEhixhYxiU5oEiCgN
xXwdatv1RQsxFTxMnmGTe+hBK79EAWyimhBtAL5ht/wMUCt9HnNYTOPFj+8pA90jdBs5QV2jIbZ1
lWKHJmN3/chYVz1UkwnUXVEMyPKmaxPhQx/iVpJlW8bZsQXybbbXUuNEoWwgCWsgpP7elfPdzRmU
iQzimh05LC4pHIoqWEIW30LiFn3vScLDp04MKaysZ7cV7JWC13ma/wLO7U1K8Hf1DGFlAtAmUZNh
vWKLmjJ5Sya18Jyvkr05LkgoX6IcY75bGKwTZ0HQJBzDHSdNWEmsJ5QnYDWScuZS9tSEudkHmwAz
l2nvxGC9alhsFBZo5lEiBQuCiM5A24hCe1ubEYueVbtVwvQRShRTBTXBcx6CWTtPYUug63dX1oCq
ckL5iE4Vz1bY/0oYPgbS5LTReSuTcmkGszvUAXmlCxQm5EVh5IItj+lPFg4zzC12UqQJtejWYrri
ZiI6hmGoU3HwHaTDFapDX+jX0aFvT6W5Al8XXH9PkFM1xj7G/ykcdP7qGxRgi8bSQrb1tXYNq7TY
s2hAItnLeg7y87/uNsmpvZlBfTRttzdeXcbU1drcsEs7efgnJy7FMXdXJFgwt+bjL2mAQZFqQmZd
HfmRxzq0ZOgV+92a0Zn0OLWzCNhtPPXvalj/VQ7d3x3hCXqNxkPIwECN1v8jjn09PlLLGavLlbLG
z9wu7hGSRgjEiENUPeRl1eJhv/h28kvHmsjMfbPA4wnuLM3zCTkYjahAjUK2BRS16EY+4Fg04FNb
mOLIttLx4qRuFT9fkNp8B1A5oG8SoBwRcw5RhYbsXqNYBfvX3lFNGSGOHRYAw0qQmwm0RBeVJsJX
UonPOhZ0o4wjy5rG9fQWa1+px6/FqVF94POZSXsnINCA19UP8n6tByQ05ZvHVwNAiqDrkt7WCW+3
nEzBkYf1bUqCDOmHZMWN0ofgOTLZyPYOMwnt4cc6+LYrOOKHZEKk1DLpU1T8sGHkRkS1EBqOsbto
SIUn1UCzS/v47lR/72ocaYuwLLIRgBlxSFThmUJ3noI7xdcNrwv4vcO/wFt0soZjLSCCYrSbdG02
6eCJr3Vhhof+q7OyyWInNCl9FEyTXyqxf6jbzLoQTkcDypNsNQ7GsJdQ57ys+mfv/w2so3WBYQ/J
H3vC4ubyE2TqXSBdhXqAI9735ciGD1ZrzZQJKOmNcPR4aTp7cQAwqy1nKaL8gHR2MaSuoWO34pdA
92POWsc9krZTaqR21ksPrzPQHDx1PRZ6kALKx+0EnhEIuFjKrOHOTx4NshAd3VbdAScM/ECDMWLJ
V0g4Q7L8PBltZ+E44w1Tq+/MPDWrlptOrllSMDnWsn2jQfBOosb3V0aVMjQao2mU/VXCXOMXE+Xv
g1axCGccfZ5f2Pzd2fODGeZotqSvzBbEvthOWlhQxltMUZ7BmjdKvVBdj6JybwRbplVbdWfrp3eD
PyK62KcnMP7Twg4IOoY5nBuZQgZSx7RLlHO2RAaivkg3nsvoAEbzt0S07S/DURldRz0Fwq8w5iMb
00ZOem6LyMRqvapH0EoFrCmhD8qckDHnnd/8i4mqWWd+cTBAFXzqmvI8bTxDk+E57p2OgjxDXyrQ
l7NZXnLGfaNgjdWxnSWgRZ2qGmYCLY6mAmy5dQh2WznPTHCfSGZKjcucAG2H7vJaGmCsVe8qMVXl
2okH3ooaBRWdqzgSyUJX63dS995YMNOQ/AJIOElcIRNtnal0dIi4OFXHvTWfBmCKkyDZMTmQtKk2
uSypKJP4nvqkHkbl4sOtqGUGvYOV94LiW6dELLyJXIzvFmEtJZQ0v1aBMRDggWHYd4h+z3Owe1d0
1Xi1ng3uDn28TboMawKPhoYKI2P7duwhH1ENy9rWF2DrP8E2OcOFNR1a+8mr/n3BOtwGTal4bjOM
+PEw/c6kFxMwa2+uIujZztALrJfpofaoUW94s1n2P+iyKlOQfU+X9GOMyVdsVNTngu1mxrhKhHLR
ftDbWK1uUk6sCGGZilLbN/vcK8o7e4FT5Q5aCvGIfQwlt3/7CmaQF7+A/se5QISXT0xVZs3oq63W
/mJsAC+y0aIo/+RlVswkZHo31rxpOxSfWE+ADa8TlbbJtbNQenxgaw/Kl/RU1K0PH2eOSFZFqgCU
hxQzLUBnhjISjEH/U4e88lXPMtWO5ePGMH6VQ95QDTiIXMQ4lVXMuUxV/8S9qZ7H+KxLY2rFWgpM
GxZe51vpsLnaCAIZCaYM5YrekHOFRj9gjvqVcehfUob6F6XlQmm7+x7XJIovlz0ygGjAHbAHBSvb
YIS235rf1XFw61XESSNuwAiEtP3khFc+HCHto/bkLOuO6qNgyARN87UXktBTmrPpNFmdnFOORIwY
M5YqqgKCrMu0lAdcdhyPH/GMe10a18CGOVFDljMnV1YKj4PdLTcl1cTtw+ShJF5QtX9b3qDCwobe
CWDKY8TmzDnu/saxk1VmItyTiBV2vTzl9NTM4BvSAPoWUG8Vo4NbQFEq6TTxcTnTbTfG1daXaGi3
5kgi8Tr63Nx6ACp2xw88iCV76H4idbQpek+0F3OL4mT1vpUfI5hHQ4Lt1qHjRL+hPReQDiELRFci
3gwzcX6HmP+h20V+0zFTB1ZBhEkONU+cBLI1R8YnLpYiuvsXf7YY8c3IybFzm/t3JU3h0G6S4/Cz
ds6BrHr2M9IXJj9q52qfevtZ9fShW8r3RKDKyLz0wYZXcdxvocorsypizpS5+LsEyLjl1kCnUaKq
y9T+nnV66/9HJ0Yn34T3hrcpODBqT1GC6YGuh/TR2rCGvTDvywEzJDQ0p2N/O5hGc5DJeVkz6xkr
MmjfuFQ/0wq0nDUc+bs+LXf1dpznI+wwElEgVrMXUejQXGcxnhODgmk0BAL8wL8p1smo9RRUV7DA
TfIwOVxBQt2zuLBlxpHQMf8IWMeNkkN3ahoH3ggu6hcmOVsTtUlF+/kXtGd6ikJyXo4Kgy3br7yh
/j8tQFPe28wG6Td5gfhS68RPbhNBfDKO3uV7OJXTGCoh/KXE54hEpxHcQnnbWoNweHvNSAtSJ3LB
tIAPODkZFTzhULKuBz/8NjjQwgQfQDY5Kfby5Eg8MMbmKtWnt5CbWYUhPj6x2jdWEJBLWL39U5xb
hACTPVA1laA9KpMv/JjESblcQ3ISLDdzhx6MRT6qncqDzFKWoDyUtNzEHbqJmvQAQ6FAy4TNauf0
uJVFQ974RdKQ2/extply1B4tsfTRT7HWKCML8TUpky3/R+D/UWnWnPsum9tq60ocBBBy58TxUJHT
fsrdtXew5Tbx1RVEaSjrsgGEgmYye8DFWj2XQIccFQNtpuCXQCqsfhtLkufM5Vgz+PEovYLOX0t/
1gv4V/3PBA6kgrPQBYCvLCitJc/+YHmXZTU823DgvKzxqncXiTXDxgCFnhqJbrpUPOjuaN8E5dhz
ZPOYgxZHq7KHMFHNVLkDOmYcDR7VH8Kq8B8ZsfqEKDvBqDsnls4N7YHxinKYyS2SIN25NtJ3DUkI
+NFF0jDQJ9weyjBKKB6CDbz6pvImjHRPdaTRZWCV6sYrUKMDUOKD6u9Ek9cthqqAxjEKnQEfdvej
eM00DDKqQ/XtSd91i1FOGIydSx4hbiffc6jvviH0GNRAQ4d2w30rxyAq2pkO2GQ6ZuQ4cd9Q1Aiq
OnhxQ8aFU1sHsw2z8Ohf9EpvTuyXa4TBA/CUjJWa72pviILLvDAxXaJgUEAyfuPU0ndUvGW1enTZ
Fhx+4gtIhQFuXeBMIqTcZNxG87Z4oe840eXR6T0S9zq/fYyhcf7VhxJUwcROPL3OxYrd9ZnwKMhq
qxYt7+GuAjoxvCE6hrjiRC1dHwP3GEultDF6EKXGKRUt2Yl6S7/ZolsqiiHuPD2MvaaF9Q/IB+vZ
7+XAGX4FeXeY8/3O9URDo5w1rcuJYrcR4qY9StsBjsLzXpFyl2TR4sSY1f8ofWTI+MvJ7wJXB4ne
KaPhwQ6M7fnZA0b129/VdygsCXBT33/jac0luZR2xLZ4DguTy2zB7omtnHkP5e7BI520F5+xydzc
3nvRnC2r4iOiqMPm+wTKXAF00I9pj9oc25AoR1mF8lcUkmrnGcsbiMdcuqHsekWFWgBiDSHKg+g/
QsW+2yXvZ10GqcI512rn0kg9kbOtKvHWfINgDwtq8nkOnMe762sLUJM6FawVYC6f0eUvjnz3R4DR
/lwC/jgLPz4hnuu+hHh2KDe0Uz+cTtkPfLpcA/s6iMtrhLgu6OPQg5eAegV3PuiPcIXH8zaHiZAT
HNgkbKnOI7c1h+ttQRr1KMV/BpyJR6MpeQBJsHUZKHhlWAB6qrxsVeReHDxQ9tzw24PCxKwiHoyy
100Bf651mAEQZ/2TEXY0Yvdp+M0A0bDfV6h9o5eI898Y9yWhv6y32gw74qfrkdEXF3e4gXM8rCSk
AvvZ7bfmIAF0FYsEgBnttF8Yabkn7Dr0VH4ZrZ6yCfHyca8KlDcKG0JX1/JPW+y1nJTydJW0jAIs
/gOTpRvh50D8OyTn06GMoG8YQ95Hc5ub8VSW25Q+iVKnU3TQSqezOY6XHSCxNXEYdnYgxWqDu62r
wELHwRLvsHvU36yRvOgkwwEaooKiIXJ+XFUJTPHKEvsRQeVc/ENNbfaDCFNd98DUs3GZ+PzVu/Uc
nw4HjdxH0OGrV0je36OmO+1KynNmGxmSiSAYT5KlPOkkmqa+c6zrT+5dvDBmTo4rpNrKL0cFxV7P
P/1Ad2/QYRWHsZi6Z8FQLPh1vOtm71oM6Lo+OsmXZf/3m4WD57SrWaH/8skFneZzu5ak6kIBcQ8M
faad6MilE44aGKj0CCroqG1U/U//rF8I9lGrUJ8/75w936G6uj/VeXsDBU1K4k0KNTwiAclJ73nS
APs19pGS46TEUYw5gTO7ahYPDhodFpCDH3fuuo3e6864w632+yR01MGqxibgo2aGGGFUtLbqHHFI
aFsbyWK8mtq2TBP0fgmeQMS1JrwoLGTRU74bJQKoGq08nmSw7gIGnqb2eLP6niuhCPcuX1G2dclP
hFuo+cYgNxVTX8qOTUer22BBpOX1Q/a4sYTN8wYkmlye94jQ3apc8KKkZpiGIbUeZdFF88dqNeJP
8e6L35eNHFbx5cyls5h88PsPQ9HIkuz5/S2j8/iwUd6avCxiee94Tlopnr+k8fQziFTey1Ibf+H2
Fj0ed4NZ1/l3S/+WmuUZR6+XS7+0M1TQ0G2+RAh5Dcec0X/3Khxp5x9V5bnZ2DIW9M4a3PZ0uJlj
O3FObLtc/ctdwlGQH42XWMYIGZyesi/UwU3VQYd5Ii3j0YVB1qdijadyLafv9KfUTlTthBKxYBbH
6wsYt1g4KPhcSz8q59cTiwyEFTIjug6zTJEikjo6l0cWf+SqUHPcM/F7Dml0i85NL0cBYVjmkl08
p1IA74ON4N/FiR4weACgummsEYP/ia109yR5kdk631F/D1UI+dSZyytTTwgMFq8JVcVprtEd854F
YFCklXQVCKGOjcCYNez6UES9lBlHxbLMwYQ6r5x3MepJI++/v6MO1nj03sdXyI5xF1EswgxSJqg1
iPeyJ2yudJsbpenjjCBWyY+UoJBWwuUvpnP3FMQHQz3NtCjROUoxB7xgBVvJBg9mBU+hHeXHEwI0
0N9k+v0OBWJS0qX0nhgV2ROgt0F8suv4Op8+7XXOK4qM/dc5dMEA8y7v1EEjfXKqMWA4xWdpwlYi
gsajPqe7CGpRSZ17sKilrp/oblOHauJCNpq3jjDfRa73fuVLEDWVMBR5xW1RiP+FpUmZ0MYZuUvw
ZhUFOVDccGp6BlXD5QovcZjGDXCdW47Rb9/PtB0hF0FpkFPC12PI0LTbAmUASE8Iw0YGFhcS102F
Rkr3MxQHd7oDgDk6r1UfXqAwrryYMsYbv2Mt1NsTOuPT9gm5GDWapyAxn86CugEK0rl9VKheAonK
+0Ztgb5J4OXMqFYQyRdOFX2DIfK6N2dY2PZ52Oa1NAqLz5Kps8oZsGVvRQqr7RCIL7iTRmUnqtFf
+ewdWlTGLvluEKe6PmEgGNoNsYHp7i97g6HvcuOByZYbcr3kAv37BlKC+ucPdyFbkxzTIkXma1XM
CNmRTArHxmIV0vGNDboeuZnynF0YK/4L9rW5DwsIKKfTVAViVUmLf0fdWciI6HGekF4GxZsSbetU
7cCp156Kg9zeJbwopPzam7eycA4mxcSm7CVBZy190Xde2VkTwy/Ya/SYtaGaOuIIc78gF+PjCV0M
RsgzQaahveNNtKxdqyUEHO9Ab2AKPKD7/A5mMVvjLsnSwl9DzOoimHR0+Bcqt88XbMC+W1b82E92
s0m3QdSutBPYMPEUxMdlN8EzrylLo8kOQn82Zhtn8XYeuwoYPm0z64/hoKZF+uzJ6ReJJ5yz7bWR
zZQsGdKE+jA8c2GSpGrYHR2+z5Jdnm3mx3f80784pDPW+loo85SqRynq5mraNbPJk3/VukAd+7Mg
1qEoLKkmg1JGoybSbhGjD+Rm7m3aCSO3FK4lndL5bnxFD7X1NJiJffu38tPKpJpmgPpvrjFzKNZ2
kgeVb0177ItZ+xT32W2r04UEXZ0HJWAHyb9W5JS3hWqPzhrSxoYpCj5AjnrhdzEKtvcgaEAR09Eh
LePSaD3i6nQMrdTUz9s6oKFwmnt73J1N/nkPTvgPp3ztTaXSqzgV8QmOZSKEKyWz9QJbAcf+sKRk
5wgk2Ve3yiU3bqNRo2gt+6gaxuP9nrrsntdGZQEHSJEWocBdog/UsF9VMqltqaFUiNuoaA+aigtv
e+Ja1sc6LfUNfrC0O+t5e2tE0HT54R66OCvjjA+5P242h/CBM7Og0GQOtvNM0ITjm/xJ/RykaTTe
Rtk6iK6yGXdLT2Fawyp3hcIwjb5QNmdkvIBjf95dsylTByByNPJ+2VbpHjDCf/pOYTTz7BPSMct9
LG06gxDLpuKZN9mu4I28KuG9pXapaiIQRrVAvBrZz0K8JglMXrMckngJAPVtbK373IerHUVkvDm9
TONjNxiBt6kIErD/oJEwwLYsRSqrKcAi742hWpKSINlaqKZKF7NAn0KpLfn5j2iaLLzqWv+/TayN
0n9AVNpFJCCCN8NElUOJATjS8MZg+S5UKs9A2VO6GI8VoW9kKYaULiyEaBfAqIgdNwaOx3AaBiLx
kZpYal/krPdqgCGYFYkVPy3/YkwAXuASGPqRbxBsEp41wA3d6lCzjz41nRht71SI6IIf7tf5kOpE
QjBx4GbcN73pt9vJw/fLQN9PIL7gn1um3cv9jVGnWd3jdrZdgOUfCUsQux48l5xqEBZlpVPhvwEe
liPznz8POBOC0VyVkbBZROIUOTRfLdkKbBiEMU/cakQxLGasLzquU79T8leG71NfuJLzgQoApCVR
/AcN1UDpHAb1DhCRZa+ljyeW1qb2aDHgqYWEfUnDrwId7AQFmfTm5/ngX03Dirm2zOIjHlt0RnW5
RcUQfG+cncLUyobwcojqm5DvJSyPzCBxy3WfrXqVEZU5vIVDb+gojOBIThJnZ3U9KgxNHyht9M4c
dIYmcsDgb67wqLzdATugLEvkuXq5H1TqnY4s5frq2QNbeK79LusK3BUxV2aRA1U2LbBUMVN8z2IJ
gegW0XcEzL1bhQjW/M6kzO6K6QOcBZdQ4nPg9UqzexxIcjAV1mnkIVwFIQ7y0i172JvAe1QmZl3P
htEPfncFuIAdbFEK840/5bFIeV8I2qlM9odrpGAIWTxlE77RpiQWfdY1bUHwoLEQIZpHfXZYNAk+
OoqYKaWA2xIYmw9IvGl9SkHslizxPMGPWRYDatEMiXi0sPGQZrw12CgDIeuL1gr2UveASgMPe0MW
fGkVwgGzMdQ7B0helSEp1/w0gJnYjoaIcwfAHoCiRT592kG+sRs1JBCLGegxL+mJFisXIxfR90Oz
rA074cs0fIrwGye0EBQYzmDIYjLldqx7L2WWesd2UYEPUGcer/SFeTfO+HqFjW1XNfH9Dwv3UGp5
aYEv6gMI2GwDbhWl1Y44ilQsXwC4QjecSSakwJSO7Iu6V3IEZzEyDfpL1tQ2/hKKz8YwjqxuKjcA
upBLlwF4BDz65PZy5FY5PztMurRCzdQAfn/odakwZFLTzw/MGFs2RGmAoQOXPueyJXAJ8gb5vFoU
zA+6mxZhnhsSXN0t7OB+3m/mnMhyYDEkVXg+NiPYTiD1A5VEzX5RcPdtP1mWo8AOfQCTAJ2SX8Dx
UqyrY1npsUgYAZ1wF5NcAoDx5uibr9horyi37AWvRSPi4m58G8r3lJUaqYEtu9jPibwvkYPefxLw
I6OnGlCkpLd1q+FfHwcGxB2JtWRmYSAmzDLt270yxFpAsUF30r5r0oasa+Lq9TuICdgVLSJUg64L
K5CcYv4IZX3DvIe0pUDwmuab/hoJAK2RblnthskqdGxzD7QRFRaZ3ZfuTl6ViV7DjLYdJCxiRSaz
lTryplDb8n5PytYm3KMbHu44wVL/Hl54OVIsG6Nuy0HD+wv8ijyz0tLM8BkCxkbvubwTpvaQjcjS
FpQz9KCTImFdNSf9Jmw7PJHqLO5yxOGPv2BBBqvmOC64u828yw4VfixjIHOHCtKSBhF1FuGVtTSj
7nSPgMITXA9G2ySPrL8RHXZH0gdXCbh0410EXcUhGQA8aB3y+UQ1Aq32oy8ziopavT3GYBI/QD5Z
Maqg1OAgpDbrQfpxkphBgw3zcfFtaKSefoQaIzxRaL9TpYWqG0V6kA0NgHauBKX9vhrHVnNGPSpc
qIBQK3pAJ2jnJWSet7FRaOU6aGFk1FNSj8MfTHDfEJLEHSHCUx4ENr2V6xabOV3ykowBlslsErEe
X1K83xrOlXYtkq1xC3O+scTTOpWmB+oq9IqeS09LBx/da5r2cWmuC4YNSGUmVKwhKABSoW3GoZhh
9uwxQPwrzQJ0ncIoYFoRm+8UghTVUD3ZCMs7IfkNrd1Ded/3BVkjTfLcv7usskQ34mwDE3cInpUq
gZGmLbVRON8pRjBjiVybjiYZkvuShfMUWziCh3kd5hT/YekBe3UnUGX6SbeBUHC21KnSskjq49R3
3ZJS+8UgmmV6wa/iBl18jZ4GB7XazzfYfc7S15WBSvgqMCOEUgyje7DRBzplg+Ik/WcsY561fKgn
ZeMuW/RA3fo2UQndWJSpUVgLz+TIwetseoOIY3XExXn57/kXcX1PKAPu85qJwpRlgF95LgUynkhw
hlgEAzbQtQ6/UIk4UZen/D+jvS0p6u1ExU016vIqYXRzv6lfkQd1nlnGckpMjL8Fts3H3JRSzIAL
uwlxEPKaPYQAb2lAh/taXTi9S1zWj1+qd1p4PxiDKk386Hqblu1l1N3w8jxumCwNvZgW9OHe3Vfg
7dyg6CuuvziXuXhXDg4wD90MYbhVjlfWQWauV9ubJsUiI+DSZMr0JOd/VzYy/zn3e1GGcelQkyHK
4ehBhXmHKzw9Ii0ElvSlHuzT7hkK42o8gxCIzUYNXgu/+p5nDntoz/vcWjDOYDMs26pVRK8LI8d4
GwrPvOELBp79Zr5BfI6EDq0t1hZ8T0wZhGp8u0AaOW653D+Q6v+DFBfgRBucWFLbsTfXmNSl4D5H
Kodd8Xrjy7DkAbSxC6uNBbYsZVB8QEOUD1AHxtUTV1CtlG2knHzNmPmd4KnJ9XZENz+6Mgvoz9tL
/SETK1Vky4SOBB5eMF3h5PQfQEMzplKmtfWWXRFc26MZ5cchsUGn0/zGqt7UJ6xQdHQd4lkgNWFc
hj7pP8/GVlSPL0eF4uvyt2+Mi6d5PhBrg9iKFShOiA3jz8kp7igBnrs1kqcwf53XPvrjWfShlDTk
9TWIwB2r8fJpAAaM1Qufzwgoyv6aS3+IoZvgt9gbsadfM3njxv5hrGrftkOULx495+eUEp99k+wk
Tm9J4UFSJJ2lsYNdF2vt3kbYy+oE4jXhhFTrmCzqjLnmgKu1gqT/l1q3pUxVf3Jk6hKf/aoTvMXk
tcN9GJHFUIfAIYzl+X2aXuCcs9v+xXX2qEOKo0SulC0KqwHcVfjpDCt5E2UsHqqJjCNUaIOL7LqH
sbyYvx6xu52w9l3fsG+PQT6rhekx5X7jfmGGHKSizBDua+vaSfPWe5U9oE73I+6aEj9D+TUWxKPa
Bu7lKXkGZoWfguUKwkk6mzLHm4G0CnPNYt5eHWsumTVx6BFh5i/7U+ght7Gu+K+fZphBAfmk1AK4
bMjLHolFwhWW052+KVGksYPtSwW7o7jf0XJIizsZ6rj2U7KT4ialTiQ/3mbzoAGkcj1STa/GFZwb
I1n/x+izvSAW+LVvZBL14hYgvbkWVrRh+/lnCnBO/nP05lousMdcWu4as1WuR8QEt/zvRNt4uKUg
ydUdXag2P0WDQuBQRINjh9oEBv4OmEGm4hhhe8YfQt6WvAmneIIz37jTY0Nb0oRu/xZCNMK4P9Bb
aFrx2JgqHh1UTnQ8lT6VVFB3bzARgSjVW2/GtlbI/Q4M45JZ1Vesm3SrhWeJm5FcaKiUVb7D8zuO
D/W5gaUm7L5zKUk7H/6RkDazbihNQqQov99AnVO3rBccKbMHreNawMtTZD80aEilGWMkaOUBvAa0
I0eYYyQM0AL+PQffy879LHA+UgPwWJ1758/Dz5iH422kp8kANP1WXuTIhMgO0tihRXM5ErI8+f/V
Jn1bLbEfXhH6EM95EL4H+V+RRohj+YDO3Qncp5qUHaM875jDHUp+QTPelSn6vVfZS4pe11OcFUgr
k65mi3uHwcJkx6nXvmuewaC5g1BaKeFsKs41jDun2wb6sr8Lp0ykLZsqdKJR7XVaaug30aMEzaGO
abSAY1NApznzAxYZax6aUcGoaYsS7Q8cuXyqavwXuh+SJjpHaGJJxvl6k/1D0Mzoge66M7FKjL0W
9f7alGQ0YddX8Rt/Vo8iXzpRU9W2RwF/3duf0O14Vn7bn0JuzU40b+aSnWkW9JXSzLoHEKrMuF9S
NN84ARunmGU5kCcCxG17nBV1QvANmKUJHz9nJklFQXEvPKG2FvHYWVkbT9bZiEDSJSJeE/aGSCO+
iuVdYcyVPK6sI4dbYMP1fvHCXppxxDM7numxpYw3VFZ6cUb9XnlnvjhhU8iMmMcVCw1Cwe8wzd2K
YnX4RAQkCCnoqRf8rAHHftB0nlbXdXFfF0SN097c0zHgbH1/T+e04lG7sV1eOPtVY4YDTjInrzB8
+c1fsAj5olueLmCea+Ktqb0jTYX6Z4+TIxRAytR8l/o0soGFVN2WOWp6OiXFdLRXD97yQkkhCei0
lBQtWUhd+bb0wdEOJ2Gl1npRNomy6XEllMANo3UGWPNQF4TqSI1l+FOyPAZTbFvyuGYTlUI5wfVJ
oHqOdAiS5uyrQI7SiyJokuQ6UUdCGM83BZTlMFtwMoVUTnUUqQc5lKYoYvIhWUKrbOdyv64Yg95d
CXmSpX5VEoVLy0yLyYxJc5p5YzT4UADEqqF4nelextjRJjFvfu3VZ9Z5Nclih8rgh+fGoBNGBCs/
FsA22UrtlUVxBKTztIdszGqTQqfQcjaW+T/0SAJyKtnUbTFsOuFesqGB7w8i1i3KhnobyrJ4KAuW
1rIonJlviuCiEcqXRadJAFGWW0+AZgwTazcr/+ksHsyw94Eda6Zyr/e2N9Ni83mj+2rp5RIYTxzq
iuSoFMtAHwOx8WfBRP7eIb1kUIXJpErzwkjwBIiQTn87C8m9pXwNla+cpKM5VMmYF1i7vBYj6zl/
+QepA16urqZxDp0J197vLtjjdFKZSce62418ZOfg3BCMStxiEqh9bGHoFMlV8vLJG9QaWwSQo/II
wo595fw1dMhPJ41B5s1ZC4eXnTMrEHAFbo9sZZ8LvNjoG1oWT9CfhE1WnuTWMpNulFOIZ/PHvObc
H8wZ2WZMsZsfd9+ihF/LMFFdoXyCvJygyqybv1ZKhWC5V6sCC9VuoG+nbKxNsuY4uMTp/bDK3pFZ
uwGCSf26iKhPMP9hr4XABCF47UJtQ08xDBkPGjAZNeEtScWu1dd/e6La5mrBf8midkmzov6mV5s+
0cUXo6+yyqsJgurrI51kGKVTNzZNVL/Hv9at4EG43UOznsgcIBxwl8B9VyO7YRzS22Grk+EoMYfN
JXWnEIiGJRpBRDEP7JV/wpKq8TlO7k184g95lxCoEYIVx8kJJpaF7wuA7ns7Zgrs8HEludCGc5Qj
SyDpTdJjbocKL7dTwG/lGBGaqKxF1sgVhz77oTWYItUouZoRXBIQvgW9D0BhkCOrsNV48L/SOSPv
tdeVLaL6NFHoE0gvstKjax73iQjjSA1RlKYmxdRDhCu0soL1onGdhbOL9wtrgaLzpVgMOYZ+fQUT
nAapskU48rRAnJIcDEcW7lCGMqbiN9T22Vvv/qXmKHT3JA0SAfUU/NuCO3ZT7D7l2XtaS+Az1MS7
G82xRj1ZmPp4YLynE7WbBcArQ9O/Fx8RAPSr9ECYL4wacbySp/0wSydbIrlsxkfUoPPVLKw/37LG
vfkgQP8pcAOkgbhDtCprf/Gqg6WETb1OtQrzLWKQHxcz3EzU2NmE1E89F9qmdir/RoQZU4nKt1Mb
OLKcWALtEYIT0VL2YGxB6qoqRcQJCbDNLXo656gbBzTTbXgnShFAVdCGFN2SGcSIMiOtr08UNFhl
ZOe69uWZmdAhtK8+QjywR0O0H5KQWSB/MLVsUqw4G8DsC1N0wN9OtBLkCoFoOmzI6/B50aZI1h/p
m8Qd+0R83Bjt9z4awkSZALaNsCpSMmoEbNxUD+wuXXJWGowkLGxqj8g1BRxLzcEhJsUf2W/csrVE
hicn0DMHtFh71X6BeJ5tQY+zeY/ENzVJ88jWH5lh0z/8LvKKwJgpo50D8/Ot1ML88LGgIzrytK7T
YmHcmlzMfZcqtPnwlt09vy3r/UqjKrXEeoMm4yGW9mj+iSupiSdYXbLvX3aso6iJIVmVZbIPNiJ3
T04/gJ1CJ42uRMiXCoVKRy9BR5JztY7dxj+QDI1CUGgyuonjjQDUWToOkqeJ70/1tXTdsHaBF4zW
QmOSJDaq24wvOCuANMfGfgp7qW+rBVD2AQoL8BgtqFqHL7bViTk53rq2l5/pSbfjRoOk3xFBEPz3
dX5A2lyUZONIN+9AVQ4zIUHeiL3iN90Edp59SVCmahkMyfBrkIcf4YOR5x4q63KtxDPQWBMnjPk7
UgbbRel+a8RwgPbTT0/Tr4s3mLVXphX35DoF2XkR2lV0s2qhurMjzeqF0HaJ3w43W+UI/CySBaLE
zQKuOrmsuUgX43eX9HHnpOBy2uXOTtOWJx8+mcrnuDANn4wJfspWrCuP8eO2HUPG+D02pGqA9cgq
ndEx/TbCFMfZXDl6uMZt5fecQzojmU4xXDA22t0SveMx7Iq/uVQwDavbwnwEYjIsg9UvHdnV9ARf
r/IakRK2cpupWx+DLFuFsA0mXn5Yc2RxU1544Ryawn/Z88/ynMOiyZ/htxDDSY7Ixf4J1PgJFvXq
qy83MGstjwBhmqIKol+IiC5ysgvOP0+cRUj6EPd5SKkwXf+xSE/Ecqa+HLD5F388dzQHG/jPPDVw
LcpiCpXxR7KpyK7EqkUPLHZHKC/vYk8qWRDqEwkr+X3y8TE3ZAJhglTzWz7LH4Om4tOcHlCWfda+
fCwEHyp05tD2lTRZ1icl7PBI6hi8adnoyW/u0zlJMig3FdCJrBuEgCR/jPgZRmfGJ/mIWaM2o2+5
MSUPtnJURBrcVy9VjScT/Dul1oKUwOlwb302r15IatBP0c9OMa0xA74WAma3GM/IOO8gBIKWfyy6
ZPXU0FPfl5hJn6ZkK9VmhNHoMBCzB3Fg9qoUwvnbAeA4VgDRUJQR49ciZW+MyYWURolzu5/mDrLZ
nkKuv72NBgIHkjD1O6pwdLues69H5En2Jx5Ll+2SKF0JH37DRpYWv9BJnF4Grz3p34p5Sb0qlwCr
bL8rljGDNBPV9gKRrXMJg5xzVJ5ue+3p8z4UAN6Wt94/245s3/QU4GVM1btPDugLulI0fwyzg4Mk
kdJ7cpBgTo5EeVG6cHyLChrcGbsuZDLud4r2m4zki3sZkIB/I64skRDrfp0Y/EBP9Smyb4+F8Q7m
oPpaGiDIdQvGm0LIiiCRfPFW6tm5qBJogd2HoxjVf5A0NjCUpnywUJJONKEv/3VlYlnkI3o8tmc4
g1oRg3Q4R078NTwlIA+K5i2dmKgR3//0g3SrMsd/WaXiUlQTTOeygIXDBHj/pYtdpGN//GXJR5xI
4AbL79c2MGTEW9UZuZsqyZPLI1bQ/0djEZDXHT/JsEKIqDTbVnWF7dAk5AQcr+z/S8NsW4Is9iCS
jsDXJdcXqu8IPM8i/BpgBkIYJpOv8dIJssUv/a0qnhr+I7T4QVzTAch2lexWGriFH0lJ2J1oL16m
7uTKmlVHKExMsKUonm/ZQ6bUk536XO7mmXw9hhUpE8pCskt76vRBG0icK2CUPcSvIutuy/39UOj5
Eb1GOMZ/c8K0emXAahmlTgu5bruxebqSTfm+aogzB5QnBqoT9H6qqe133BPWPbOFE3U964T2zhJs
uE+FvoAL9UhX0s3Ez4W4ccLcXD+rVLgwFmR1ZlKxz0SnrGRSkvqDRuI5QPisPrRuR7H2ipeU6NrZ
HuzovgAY1VLGRjpV4BoLNQeZ7OtwsJZhOBPPGc/HGMp4PTLba/pEp9m4fHl42YQyjGNXGa1hqpD/
SetrxUu5aUv8wvWEZFmsK4Oqf3lV0vJynQay5LLBTu43cER56MtJhZLl6Wk7XB1NjcMVdcJPiuna
WQbjSijMunFGBgj2iIvPtCcXb1pFrZfbGuC8ufoklXmS7hn24BHvAroTVH2Eq1eEyL/nKpZK0sYw
ZbdAy9PFYR5j8V2JDikCOURO8AMj24xxHlfEb1wpj7OHwMx+x3C55XNr2Pbu7XFqJogeIMLhztyN
fvKYjWeuchauZXWt8kLqFn4WTImTfzRRroZRK/nYrLYK29kDaj6LzUMjcuZb/132Tef9/Tj9yAJK
p6gxNjVUY/O+t7wCd/iLm4GMgwWfXP3MO4oCHH04TSdJhBY2NTN58qCUt7Tcca3zOFSKBo0E2S+0
wqBY3Is/J9bSirQtN7MJgw+EYx6ouzhZdEqmuyPMSlpD+gybYHksnKlGTbGj/gODow5Q/y+SC5x3
Xkc0CTpZoXkTKLNBTDurjmYSGVTrXh3zDmf748lpoUfSvjYiWhFt9XTwWQL9PxARNFoGHuhQmWkU
/htCQynbcyrXL5onUiciRZywUa4Ona+lhyqaX0OZSo89PFZRrj1Yjg/a3vLq9oauKH/uxw89c4oL
suMcKW3eN+UN8odhI0UokBI26EEF8QMWFphWdBZqvKn4t+tqFguY1zA7LL7FAMMAjHAsOFejvNEp
WpEf29eCJ6hTRlz3zfm0FODOfsbB+iGltr5Qi4LRZh4pzNBn08hxSbPHYacYLyagTbJywvy15w/k
OZLw6KUeUEW1MDSMR3ntMIi3F40nHix1Ns/olMZ97hShZSzZbNDHXeCivqfhq4JYt/mT2ff5+1zz
diICe60RG3YwBMbeXD+UNay3hsCQ5QIMOPsroC4wbSP/jpRt2a8RXTaonp5u8ttAlUQXInImugVR
tL+N5BZ2qx9r8z0Ex4PGoVFqj/hfS8WNUkZeimJHipjsoPukC7fCVfXk2b5YFdHyegcgC94cHDct
2unbmzVO/AXWvjqybHV2JZaVG0cbIxx3lwzC6/UwU8CLkKYxzLyKjNyFH8zXhc1bxSV9nC56dvAu
ChMWF+zMlxDFjmNtBucCvi0h0Vo2XqooiqO+8fvIc33S0/Ak2rvdYqir1LX/FIWNcmw+tsT+IUBQ
8qXxZ2bYj6T1edcFxu7HegzhtkEjD6Ub1RINOP8JnNBEr2NMDqoQhcyJa8pfp6zVNKy+CAyfFV1Q
1KvPH0aC2pcoLe0/M/Dvbf9YNnA+J0qarBDao6BBEGgdMJggfDGr5UVF54WYGEsqDoijhjLzeQ28
0MJa6EU02j2kzouLqdGjLdJhY0nQaJOE3D0D2G28ugvB7D5lPWYKBN/HJEn5B2m6ih87Ne6M9clf
VVYcmetqS491KLDYObBUr6dVUwWqW5sfQT4zYxJUoNYgpxDNfPIwSTMiawJKShEJoyOlm9IGa+1l
9kEtXqiTlD1WDnE3UkWFyDqc6UIKI1o+35ytjSYRiMyqASHVxYacYdHTDr1E1b8r+4DuSHcpBckI
SvhHavjuY3gNFMZMMXdHN8qp9X4VI3W1zNTf7b2AGMr9DUmA3m8zgIhxAu7/RJJ3aJQfgsMbTu/y
Tr+lueh2LREjrRamH9FVGSb5ysn4xdH9+rroxkPfgmPI0+ie9X3GtghursDeVfHWzQAALjpzL79s
YFiL20sigMlO6qnMCCK4FC00VdH6YlTyQVOMx/cV0uDW7ET2wuVKJx8TN0iH3RanYT/R2we0+YH9
SZA4p3cXLlv6tmOBQ9+rpRlwMrCdnnlinHeKJWIEpJ+vdICfBrjdHDGHG9oyJlIgm9GAeqiO9C5h
ZQwPID0HkafMXwxUiC+VfEULOPJKiV/95sbV+dLs13WjYOMLOsV2lTiR5JM7ZT2e9p5szJ527NR7
QrPCLVd3usO0rbAf9lt0gRqYhWNcmjQH6E9kNmkspItt7bV8g3xCDrnktUr1/dhEVf27x2dQ4YKS
A7YT4fGWYNBsYL/SJtsyPeOz3rxpFhDdubjyzMcj/GCmBeltZ/VzW48cZBB20gkabZ1V1H7NzAJP
/6Yf3KqG+gjgr2s3cG5K3bCdUhvhgktCyWqfIxLiT8dF0jjx1DZLpi8YpE3ae0HET6J0owlQhXdI
03e7QaQoJPT9zd1jzpTjbekqPg7Xjeoy1lFl/w9ON2ZYHU8YhsxXSbWlF6ROLlcAqlOS0VQ5B7BG
ZU/T7tHmX02Qh8nOt5jMlmQisStxMWlQVPPWGvxRXXpdtvZAZEaZRRLSCXjXwMlQ2M5wQV/PkI2I
v3C4RiRB4ArHfmXHoQmqhMMTD1ATe5HtSEaWDAHqI1d0O/+/efr7JkRs1kfh7i2jAC99b07KrKNJ
SbZixcED4gdeg6TIpdTKsePDwg3MEtgZUkQVOziLBxDSaM+b+KK/2nrrvCtkvlgmfuKlRCWF8bT4
KPzs2oqdl0fKBBWuElq7K7H8W4qi6DxQA7TjtBsqNlR7zbns/zKDKPLgQT4Ac5neoxLy0EV/op4A
nTzsEs6lfMburU6p0X61KROZ5Qah3f3YIPCJe4N+niElFNRuk6htf04/1ILRmD9WuKsDrb5qyikm
M5cec8x255UrPNkVAAlpg0O+MabscLxXRu+7HefD8RUDNR8R570IOlBNK28lVanceYUCAMPXtFsR
rO1xTc96qUrzg7LqW0dCpUSLNWe28bnTKw8HEDxj7iR5QiE7vAAQgOnK0xkp/7QMu/OKgh7LMiet
cW36n77c0OZVe3TVmvC9MX8lWt6WvfjV03HYJ+BfwtPcQzXBs9+1uOo3izF9CmgDgRymI/Hzk81s
KpMYyVn4yWKO+D7bcSRuPYezHdbu+C+QAX/1bu6fSqcDl/CG2V5I+6zAbKzC+vwT6QhpOlmIEfMf
1ZV/HB+gQKfOl7mgrqnzo3LldceUNuSFRpKh0gcGzXSECxDnzXnrsgoa6/xBEVU4PLNauQ7JWKyP
9DPMIZiyh5Xg1qLTRL0v4Urdz1KEvQlf7XVTvRcTLA1IJzJjYvFcXfwUpLkmB/52WH9vD5eoNo91
UHw8uIDX1Wca80mBtfLl0b9gBdO64xnnQprZK0ZJpLWJWOqmdR/gDeEj6e9vclV5FyTMvVVjIW2k
A2N0SxiwWuHCPfd2qAuo5snHQOjiKksl+BkQhQKo4FfaI+e/QgR/13pCgzOiRp6C7k8qN0+6wdfZ
Xke5Jogz4PFuzNuYLjzsKH6qVUzpJrMo0lZklR8ufiyOBn28Gkro9CBC5EBRtuI6meQR8uDR5z2b
RuH3fmwDr64M7JShnk2OWJz2JrrcPGy3lOynXcKtup9ZLmcgmhx0BZ8YhKTIj82u/Ntu8pZ40J5U
70CesIpP7NiGHLTDFxmmWTtgCF9x8ZhNuHvpEoPHJnG7gwCGq2jW6BRWSf4FsaMAVChst3iQuJC4
lJLggLRM8trB8i6sN5WdYysHXjR81qK1loK6YbfJQYrEh6uTq6cqunlxDANN0pFZrg/23qPV1/kb
eFK8CcDkW/n7yLCykZl+mpqsK0+wWfNZQ4P6qoX4Ttec++TXLaTtUxFshevYhTyVMJJxroqfVtyx
iZrdhMOsWDC+yey4fa65fGk3M/llJXWPfXS3UIwNI8sukDU/CWthav78OgRxzh0wx3AIrlbCVG7l
G5Xiv6RdSrRX42KFW8A9u0EhmP8MyC6C2UTY1QxX1xX/X8snWONWd5eBS3S/jiKvisAoJKYwlFTm
LyScFLkRVVU9z1u4ZoCNwQquE8bnEiqE0orECR32HosADdvOgf6PIo0W8NQQHznEWRKwJ3fL9BSx
wgO2MaMIf6pi+85EvPJDq0k9NPMu4Bo6KKkjzBtgamrWUoMFBobxdNOUYkEpOwRd1XpSRT4n+a/T
DW4e/WBB4Nh+WNQEAzfpMwW5ceabwereAkrOu8OGRtUClyRR2FOXKJuHh3pgYoB8ea167uDQCvah
yKRrafOMwFtXO58xCPaDztaNLjsuMNsy7wlVUHVzeqzSpg7UN2UHGsBtfgVQ3/zkzQC5vzLGULk9
2fuwfvRZ4tNG0o1ZtKr/bETdsh6YD2RyQCF0or045zCTEiIumF35/G1nyVd7MPyl2xwls1wod0ph
zlcR/is5HtyeM4Y0StHw5UHG4CYPr1I9Ev8+7f5q5AG9F8XpnG7ow1TZGkPl4BE1LEtctdOU2Ohl
SveIZGSrsU3/at2N7ZyFqX7qj+ugGMr/1QzlL+Y9Ad90jIpfPdFI92IE4vjSMkoW0qtxyg/w+jPu
q1qatkcna0TFnjv0BkYztB53Xd4aj1D4MtynpCx9AgaodtRJWi1zQVk6NduJtM50AGLap55xykmo
5QriQGztLBXF/mhH7ADrmm829j46AVEUen/69zWJ3X6DDMzPJ1xG+Htk8X7acnuvXUA18OFGJFnd
s+le3skbjQUd8EqJxuLlHNcUxtjR8J8a9rloPTaBa1RtowYROwxemumHXvyTBIgTk3+u8r9rDimL
Xt19SuQZ4jfe7/SmggLO2Kybux0u5EeYbpG9R2yR8alrVn8N+2Nn9ctb206itrZJ+/MxgIye/58J
jahs9QcV58hv8cFCeiEg0+8a18srOGgvoH63UivTj5sNjsSVZUs2cyMCG4BPO2Czq/QF/kYLAQg1
knGp3pWLshzVHt6T0STgQ7hnWkEQltKMTm3NUj9IOXnTcoiVTXWeD0xYRjKNue0lymJSstJSwgpw
BoRcJZfi4lBDN86w7ojTqWrhTwSSP4+0Dd66etHmiyuVe5atn6VsTYI9Vb8CIeeXQEzwT8ezrOcV
hobkjrHknnYSRonFrYL9BFu0T8g8eUOVJJ20os6LOWTBrDiDo0QIpgE/G+jVa2jjNQTHSHAf16GA
Q/Y3bYDKxVUSA6ex+itfcd0UKekcxp6X6N4+n2STc2G2XWSQvM885ogkD25EolPIz3hZIniWQ6R+
Gs6aPo0y+Bw/HTT9COmBEfxzkY10I/nI+w7ej5zjE6q7zv4/E9h8MWN1zerSxaVAo1a5BhRli89Y
p3Ah3YJluyy7dN81w0yEjc5etRwk270kQ3oHYgwJL9qS/uNsgj+cjB85BoLaQHgQ08MyXVg491w5
u3tkyT8JFmsXOdhKzOZpu9u7hGwy4oTL+S9Kwt4ibNVS1fl1FnqCFPURjuCkHX2nt433MIby5cee
yW3gp3cNAHvrG72joqLarn4c6OlNBnV+0Tq4XLPkf7j3M7rzA6rSIT5chXEgG1dHztHPOyV60F9B
l+Pf0qSrFeYrO5zIdX154CaLXOLY+zko94jBJozmyfJBG2fiqwAz5DZy79qcL53UhLnISBRq6eh8
DojV+xswUu6lPpw7wK4C5c4cc9w7JkAdf6BrWPQbd35eyjaaMpWaCk2Kf9OHlNezZpGnQfDPEud6
JblMlTd3Rtg8y4RjFjnvTiALpYt3oOESGotW+Uddw9AptW9VwB66ff7IquE1iG/3s6f/EzgdipxV
WyDQVXeapzpj/adqryCQozJdInJitxqazptb8rHjza5eAqXJo1E8qj6Ku91PZNPT7o8ojgvzq2+K
83u45aZiZT6o8E/fZOqVSDiLNHuZaXVmIKnlVNazy7x5tWIX2TdFxG7a1zbMQL7uD2ODX/HM9Bqz
M8rYQVjfCd/7r4ISnAKIzdIYsrvT0B9ECXXkddynY3pGY0ffJoJGznNRSNlAkH6jNVhNLv7+yTQE
u3pY703Zj/ATtza6e4/rZJTTY2TFf1+VazBAAfCrazFzYSDMmt7j2iSUgUCid7V8dYBPiQtKY9kO
Vp7wBBkHvUSP7tkbKUhsRDME3Zf+9qcQDk8RtrZVHJLMVrFZ+ySM58ZtAp/G0B/iHmr9CzbD8gDV
XMPPY4hDlZ8AmXI5PGQNQ4PhD386orsm9zpU1rr6sMXsmvJ+lW1LMjMQfBnnUiAlo+JR5F8HH3iH
l6PfwktGd29DZ2Bqe99fSYmmYcH6GmuU1F9NNbDzTW9MbuaSJNPjfu8Z+Hlx3SVkVnpBfzSrTQjj
zUn+O/kmyfRobfLtvyJtPx0sOPdgMn7J2e1JVMQHiXO5PURY/uewf945AwW8U9+lBxxoPtzygPlL
yLLg7QFQrhWtFHjA3EyTUdholPYE2xBtBKTLQnQCDkvaf+sxHPjbmIjdEJMlZFgY6JhdeuE5GZJH
XrHYPjSZKrNkDAS8Xt0Sadx+x8VTLfbiGJ1iST4EEpH5qEtOsvKTP3Ryp9ro4s4irHBnpGEDNFLC
5WU59z9RhsuHO1ZRnzVH21TKWqijjqA+/2xAbY0/fGJd3djGv5Wm910Iaw2UiWtEcTDplYJCzS5y
6HjKkkLoZj02Y7n6enyFjgp9oE/nDXIA1MtKhKwCEjTuOB/cKlXhEKZO4UYdr7pdz+oSBQj4tko7
mvQr3Gb/spTwVZ08i/Zx2F0JD7f5og+lLDwqtny2HewkmxSHJ24jDUsmvsveUVymvG5dIYz/ig0L
2rKsybV7zxopR1BegBmVfZMHb4s1cj00LkZSo0WX9fLLNyKeU9MaxDtXaUSGTv2saT47x8H0vcmn
pssYHZ+TNJ8yEfmJ1JPbvF3Ii+8VCmY0LmcocIFWJQCCIRHyyDNTCtnP/R6dVSOQZOev0grnoAoJ
c9j2Diz6AGejn5GHjJxdrAu/mo3nsaAbWx1aggv2uHYyEo3i9s500mAwufVe1nRFS0BqAHeI875j
krklxpFcxjZoUVPPgrXbJUFoiNT98PBx+VZYkiYvVF3Gvs9vmH9uJF121Jw02uVACmcX5xxNLy69
z8zo9TntfyWR/a5AkvKZ67QaPebxzF05xcU6YAPr4G2NsHMB2FhfaXFShwy2uK7hznSLdj1rv1zT
grw+CHuvQKuk68rVUtQD99oVw2+Lbl8/Ya8+tQM/nS4HN6Hpgxn72RLU+s9tUDVKcovFlhTpgg1C
WYrLC81vfh+sFzcdJGyLTKoHCGvdU6L01fGVVhQUeUXyVqzIfwWvBUvHar3Nn472i5t8m3VdnP/a
RIDLKZM91leilasnIgb1MdincRjrQyyb18fsBLc7/roUl6N28aR+cmbQpKnVuhAxhIknyCv46B+I
30I7HJoOdl+zQvSXUku2ePEkZ78w3BVv3SQVWAX4yD7Aop19giANEtGm/xMV0XBVFhrBOEUTya10
g6z15dnYFtn1Oox8X0HG3dvu0orDezkjlVZzrin5gFV26ggYn0yu/5j39vnbVoM0IwAY8hBuFQbn
WLgr1NHkLVcsm7KoOurxZNh0ylQcXoM4yVL9FiVreeJoirQKJFq0ZxxX9D7BTS813LhYCGRA0ul7
wbn8awvipP3xG4RagMucH4LkSIoiIAYe4tph0ixDLh5GV9jJ7UfOzbqL68JHtorkjxypNAbCclhG
bTaqKxcxpwkWq6pB3ZwljELJ80eXlB3R8N28NxxKUCzSAcOKR5MzXOq2F6Zv2a3yucMBgW3tiFQE
yYM3i/UljEMjmk78XrAeFqal6kYDd4ybkwXxI7cX2WbFlfUitr2bjCecHnDGgq+oXfEBO2iA5m7y
C9Cr6W/3PMHc8GCG0TOdAMJRTaAIsBSuD8sEpQqdVh3PQDZ9015S0DVJBDjAlgma7NJcoVjD6n/R
6p3KcGKQu82/5DWRNTSNMKDEq3zDTv+aBJgKCT2MWlBCDjXSiZaj/DS14E28HA6jwqwEFPMf23LW
CQrF0KIvd8VoFTs5ALQ3dHl4ITVCsKYf2BTtmByIm3HL6B9VjLJ01s2uxqp3+p4ajDRRTtJlNIdg
n5SjOj5G16NpPj1WstD/JmwEe3XFYcmcYvW9QysBHUupb4J200aYzb78qqLNQjpuuolbwazwKkI1
Jg3enSfUPltxDpQZVWmiYMyWhZEqG7R8NGO+z8SubKCWk0ker5/XNQk3kIUQg/pEWJM8YcvRMZQw
2pKjUyOFZCE8e9ZfRnitflxMGXPR2OvgpedcO5j2mcsz1WbYGBHlsZYUW6jaYujyZsGXP2VG9Gxk
lW7UTpXyHwB3EDqdUKaQ4eEFjGPGsjV7zgst7iawcLuWd9bb3ydhoAegBTd+EtNIXpK0xRDQOZmg
d3Lic4oyqmTLJBgOXH++a7bzrHy5S6MI7PqvSLR8lqyKtA3OVZjMSFkubuY4A+AWjKFgUdK1SMlF
GBsQujEWcKHkEjTdcyCw67ELBkpsTa+UpnZu1pFB36M4iAR0Tr6rVDfzljTQz6Hxa6W7GtnApqJC
+bNfulntXKsBv8FTlQo2/kJTSe5qqSN1ZZdGaQBQzVg+bhcXTXUndaltn//ojzBfjVD7LQgPjXfu
m4U7ilqiFK6Xn9sdFEaRegJPqBw31K/gO57TRxe7GfAWKY7CCv668hYoEe/PUxkhB/YhS0fXow4z
7Iq4OsMgMzZRRfUEOOyARHc1weJNtOsj33+P0RsEMU/pIMpFETcSaF72NecfW5NdSdSfzfxNdgQ5
iPoj88FipNpQGNNM19PZXPDA1wz9QZe6ErH5GYsTtla/lRIoMDA9FsI8RMvNEM+9OYbZ3/J4qFii
gNVNW3qQm8Wr+NawjnCf9pcjhEydrCmfAbp1Gj+b9/hQhAxFChRMTcUyRyPLEq6cx46+2uasOPdN
8R3t45aSy/37FsiIMzuvaiCWp7uQCmQgpp8IEjFAnQBdY74FDzN7CoMKkrjnM5S9cug0noFESTog
+Qgor0dxjU9FwhRelx5QJYBq0PxsryEJ0kglR2kU+vOkRK+m0kFs0DkdGNNTq+itdDwVb2RFZ9Ic
dRydX7PWoaa8adQDNBKyEUNiXpWu8jY41Ony8MwZv7CbL91R9Txyb/mJqhbiYjLfri0X2PmPy7Ss
sW2yNJqWQ6kROgfYNSQkDOifyPG2gfCRAPyIRCy9cEOVoBAjbj69l73MZOXV6F3mC5cCeiTOqJo4
9ny8lUXH8XzI0HK9euX5zQf3lcKDvORCeK1C63pNbymxrIQCdTU+5QUt/3g/OJ/MNVirtL0w94oh
7/aYPsqaPcyfGFOSml4gwv+MjlpJmXXlcg6VESWg0snZ0eGxOl9VXO67b/yYck33S3piyrYLDG/Q
i42J+jo4u2tmtn7i2FgRmFeP0hBoFsrUaW/hg8B0+MbIEjKRLxeKBbVDZSty4Fxiw5B7DaIOHBWx
jHY6RQj/GyKyV5H63s/NhxSYJuilR0azfOGkAHvjnuViQaubQ/VgXWODfbxhLAx0XpKx3PVXMgZH
MBeBVkBjyIp42E+hEs03BPGXDcTrmcX3LetW/WJO3BZx0hqkFfwqJJtG1M1ykRadsk/nhG5AeXzl
OboSut9Mf1KAlNWs9XF6s/rtxSHfCZBYnjbPyhqrhrjxsyPeytYS1PfvbPQ7haHbv4AJQ9HzKlp+
ghfN3KMjq35kiWZuuLSMzXKonXnsVI4JbtC6l8pOoZjvwJbr1Ug94V1FJlqsrP2EgODE3fJSOGJi
EJ/HKzKbaVRBQGrsJCzfmUnZuFwlnOEPoliTgsy8OCaA4aqTAFNcMfgt0cURfnieQcyiLZK1fuST
j81pR6VSw+iWH/xEHSuJxc6DHM3PEB1X5zc34ZBGMBx8dbE4VAJCJ1UWfSPP3C1niTG2uMBXzPDR
nd1diCTbdGXpRI/QmDFZXG2dh90E3sw4jnalaCcS54bMmvhpdEZhMoDPfwnNHHeuinIY0bWHqzzq
VcO1gyK2IWdY/pdR36fxBfuHRoAIFrWVj8uDGyn4butiFj15nNkV8rf2Q0hP9WLwnJbVahI/R9A/
hT1Bmp3iC4wc+FWoD9LyZUrCiqv6fKQDRZjpqBqUsJ3YhYyAzJ+BmEqS52SefSbhgfkqdRX2Vsu9
fjcgOinyx63JtbEBoqoidGGBr8S2/yYvOVTZgV6iMy1HUKVBgIuw+V7oLIZDYGygE321zNotLYXX
zarjgCp7dM8YNdc9KIdxECLnnn/XzCsh7Vez7nDnpNsRic+jWCQgsZJQVuejJErOPN1yNsXMEaQt
SkzrJEsMtrDeNVcmuIYi/fa4xMHc8MJEc7jdXsWXs+nSyFBMwJmU0uvE/85cnAxHm1S0GwXBRrka
8s6Z2vAtJF7/sapEzoH/Ec3KkfV4Hp4ET/9vj/dlmEJAbCdhgL1wSyojzkWGRAZIa60TTvowhPMd
WkSmK/r9E5TAw0y/XVt8Y2m1V+iSExRyM+h837mA8ZoOXAgnItl5yEPc5EsizIlE9ElkrJJQwcxl
D8cYcMdxToDgKTUNl7UpA67YrpafiAeY/bEzRyWFe/lffnEGI7j5lEj/1QSqr9uFr9mUBh3Yo16X
Kfjtf532LiaaGZMjF1hB5TfZNQzuEMSyxb385GxqtJzT3tjeYHEVNkWpnWFxnuQ+jzGVmwJtRoCG
K+FBtANEUjwPn8ItJEBgXpKjegmSZ8zFoHsIbf6fsp5ujOpyUr2yTo20RcQ33bz2QqbQlbaexmpl
cKu5Lt3ShEFjT1KNaAQz+kk9I8VObsQj25B+RpSFQD5mlXoGNtua0pG0FMCRVcp+79++lqKVdkff
9qz3ggZJOC1MtUajJW9sBwX/Se78Aqs53kUv/GDT8/Zfg5S9D9LWNKuVBvBPRGw94oPbEcECyjls
oqmII2/5n//E0DXiMP1qc5gwRYOFMb3TLeLN1cNcZ4fdaxEZ0ZTB1q9irYD5R8CFO83LFuuvHV0d
d8LZSQMCui8xfRMJV/qct3dp/Hauv73EO0SxiEsj6TQoATb6XqmOGW6NakQRkjXs59ky/CQTJOKa
wVjAQ4aDNERXRPzdscTJpDkYE0Jae/hGVG0e6X3DXBLKuK49QAxd21yG3NoPUjO73mMwvPuaFmMd
M0XB2KlA89y1UF63X6rHNgiGjTh0vF8ImZ12ykt84ThK+xaz9GWakMkZ9gdfXCWnsw77RO1+fD+v
w1t7Kgd1fxG4USFa/c7j71BSDffeFt2NzfM1CbDnWVh7wEUc44jGL8yHAha2dK/pgNanEyRG/2t6
ug+5KKmflpX5PUtsFsdAanSX5F5v+94vCs5r9s6hWpU2pgkpPNEa1E3bMfs98ZOZItrV6Vtx5KuX
pscd2DL2xU62p3r4Obb6MHK3q/bo9iWKgvk8NyXxbuuGfRMOW2KdFwlt+/TWAVA3HItq3iiDxxBg
xVueC3RirCnE+XBhwzUA3q2AjTLvG+K/OQ/CyyJqZZCVcxapvvWU5B/P8Y2L1QzKoDY1k+8js1u5
w/hV2F8iW9WqVCwpVXk+PdvcZiqaycJs+QLO77wN6LbMGFlLpJ0Aur9qKd4Rs/jXrHFBY9qhOToP
ijCwJ++85dPwOJc1GR3/OzSAwx7TA1bpxy5XBPgKgWXgkENU6PRjA0r4oZ/MtR9XPdh+ppKW3m0i
+TPuQcjgt/YEdqQBPJMZn8aIZi677OXNtVrRb2AuR9etOXflXJUVs5f+FdJAsvv2M+zaaV4iBkes
sO6dFfKpD26tL7ZJkji9ED49WIkd2LFVYGUHHxoKaQ5ZqnKzN1epQ/F0C4SUavccuBkkHqkkaJqx
OYjRUSN+YGVaf57yT3cWnACcLd7DaNanoY/l2PyOmB6PvXtXtCAif0oqmmK4Ho4R8p5+aHV7oFx3
n4uFseaiEIJBjpsnApr7QY7x1+Xm587RweZtNpAxaervIIbFwrmTUrUzEUqeeWfaU3oAgKByejy+
R+N/jlxTM4D+70XBAyz2Ei22Z4Xvf1pSmMOpZ7/lUnAu5gN1toWyJ5AF80mKucjAa/vt+ss5DGmn
EXl11biy9JP2UBUbqHkMDKgsiuPYnj5q8m4yjf65eqZoaR4+xScRiO3j7z+DYLFn5r4NxljEStY2
gV/PEJvgsCOEXoqO4dxCg5waC0PsY1ekMb2OfpgPfOg4AxvSiVyIoyixE7Zzr3O3kRVyo5SdnYqw
Dt3oZLdlOC4ZHVD1yJp/fG2Qjx9qqFtdiYke7xDEuBQpVw9KTz8Rvo8/cbWGzQDrlbDvk+qLhWvu
8iCGKq+lVx19759mjtMj1IYTjuhVOf2yAancgSx2X0aR06pM37siC+v69fI/c++d7wx1wm4BMWnL
TORN6k43FP9pRyI7Ako/6wwNw5Ky14wrevqiz87RmbR3lci8fJiK4xS6pS1bsJSzghy2KhEMFVr6
fttw16MPByYnKCaGyz5CBw9rpwxxTNdc9F8dzE3Cl6QwSG0nvTr8bR9OO/PRtWN0RgtyjH13/80P
CBYPF9qUDDW0Mo312b4ngSXt5zk/hUz3C1B5tup0erQGL7pEyj1ujF4EY6HMSSSL2Iennn4kdq4o
CKAxZwIis49kNdR+hioxSOlj6TyBq6mV4dY08swJ/DWU7KU1+0GCI/zgZH7sTww5O/8hoctSScDj
f9FocsVPXwB/xI/86S7denAkLIdHwWXl7nbWryMRcwqdZ2hoTx9K5bHgyGK0JPL3etgDwJbpGW8K
SHmvb1h7xr0DEXKevpkIUBi46V/fuXbECVUrcJlBNcC+W3Khi5qVNWxUF7UTor0SgNixVaBB/GNW
qRcqZMvlAfI8GDAEBe+GnIBFMH6zV5NrI9/uJbNo726vgfms6/k+ccaWIBh7Y4H/PSj5vxD2e8qM
7mOvAo67HZH13rp4QkniEdIuZ2161449C9q5KbfLm9Ne3Bx9dGii4uAfWpI2euFTfpNFtCak3Pa9
TG9wkkrU+13iC1pB26czLxPO997Mb74fy1VogSWL7dlOIV9KJtDms9sq/0djjqpVczGD2psXa4Ol
xb7Y9ZSZeIP2x6VUfM1xiDcAzpwGccuJVS7C6bxO/5/uztVEiuFpA/Sa0KEkLGGtufmNgg+uAept
vHCKx1Xf7BQ0hU45jGKcWA3Oqm/N96KLcLrVSy0z3SWcgdKM3+M9incb+JQfPw+xK1hYW9uB8TsA
Geytq9WWvwWkYGfxj2S8T/JQ790KHIfTbIjKoOZrxxwxlV1qaXU+bdiH6tZEJlGx9GTlp+QulUsS
RfOFVae2PqbOMnXpIuZDgYcy0NNyCN2bCgqBhmq28mxkOcM2fvcLUqSylSoh4nQaCSqKIAm+ozoa
4I+Iipu/G7tgKjzFRcfuEdBAGrzWi9sS2jF32oUZJC1tlZ7jOKyexn3P+0lCtNCOfh/Hku/yHfPB
35+qrU/xZxUEp+bKbicXJFb3EEnkqh+7pBRD6b9H6FroZhqL/OPS01a4oVz9FEoN7AJH/UXVzld+
Nj8N1I9q9e/HI77aet9abjO7pINglmlnMpDjUrG8+atj64cIRQHDP08ixzQ5vbDl158p8sgPC1pG
DYbPbugsKcYuD5LdEeKBnJH9CuGg/8s59waiCukOVowSFwFCFqyCwIWjk6tkuYLzfU3J8Vfshyuh
qydTvzLd5BiMECXZsMeHufybROoM2the23uYC771XeGm2ku3aaP+Q30af2j/wFo5dBlPfvWQOfbf
+mXeNusXP07vzUIh3dxxOmha4vua46Svq977g123cRH79A0Rbo5e5qY6YjQWIvGZsWecozReojiy
qx7VkzOVSxFjEZ+z9yyqHmPv10zMVvvwSwvTgBhPU+bJk5GaHtJGPFHxD8dnN6ryprwavDViyj/p
yVXSTJqD0wxdT7WaCIDdww7Po8VarNV+JhcZWM8YGRfFBzuQetfUeBynlzOVxzeFWIapZiot5v8Y
1qPm3eE8VAlFLK9UJFy64SprtY8R1lvL+QPjhAW0vQvucLEw6x9uUyL5IphUJhVPl+N3LiuFBVTd
ja+kpaI/xDV0PoMvIeKFYu8iddp6eylwM6bfEnSVjoQqwNi+NA+zTidyuftn4UOuKA+K1tTj399A
qZgffygoPXz9a9RWCfW7qOmS4HPxJU9Vuz55yp7zLe1ea865xlu9BCv7fQZLMqvdbSmTofdRG+Ws
+34n/1s2I9jVyCGi48CNmPG3SLF+I319Cril5ChlwKjg3hPC7tFJuNtGtAv7fK4JNbo3aaOP8Bem
pUslG9nnn+oD6OBtOlxSgqefidfmIWiUm1N/y/2wV+fdDHOPFDmABICBczWdcjd3j+YB3QdSoEhN
nOQTKIlkA7mi4KbCzwA+uOiZyxilvjJ343yb6uBVstJiVlCpiDcU/bTlnQjZW6mMIYCPn9qoyh3l
RRNs7gx6paP8yrUMc4pkZr5o87W5qaQiJyqfx9d+DKyu6Tp5Hw3KmfwyG3PH2DbRmqMUoBURxdJh
qJWRwv7GU9i1hTT2TwSoA4dpU+MipjxOVStHhzJ7DFwoXQ/AzdXNDrpgTqNgYq+fiZQ3xOUYzmr/
9XDFmp1Dc9T3x3p7fTIwMYNoZsJg49cnXWrdrzvUQjYz4sqL8xasjwBJErVGUcS/yvSHd6Ztky5x
rArfXeNWMWCEMwN+BZj+oLgDXjoWZ3DIVYCaIjuy7p3oONvRCt/339d4attpwJIb16dFG3PqB3yN
/KiFeK6ENlQt9ZhZRAVhsId8xwmdAq/Rs5zdMrztpNs5wtkx5da/NBR/M2dGGlIICEyqGiIiG8f+
G1/iKgrQC/LJBX6JnPTdrK8UIHym+L41/klvlwa24RnUEO80D1cLY3JGe832YaaAt9R5y0KXrgET
eItiN48zOCZlLRwpygdC79qDLFeJj5jNn0Vm81VQisCOJSmX2z0IZe+iFm513XxUQkn7/YQZIiLH
pR7Nd4nmLQzeBv8Oy0fJQARW7mW//IGbA6hb9Cmy0XbdooEW8/9R9pR3v4+zqaQSIlQ1PME/FVRE
Hz3MrMAliY3JPBJC3SXwCQyVOpwl6iaoudDo6/6iU+lAzQbLkRYObXxFqL6NQDwz+N8u9Q8MjnMD
0M23tUFgtCErpIuEnFd5b8RBLo8v12lpzYxgZYvpqkR3LIsQX5m7Q+ihcaIO026NrBaS8YmmwEtG
1mVtcVJKwtRrPXxgOZC65/2NuDzuaDkYppJJAcclw7ETlKAriJOTfQGRrfcWrCIihizrDk6Zn0A3
t38SetK38J/qsFby0wnIIiQnLIzKV6lbr81JFkzIQPfR/6rJadF7rO7YHpcQlaTUkVICKCKd3NxM
vioILv9QTO1O4Qq6MPx53rD4kaerH3tLlzZFS2wH74MF4KP7BqICX0ISqq+ToGdFmQyJ+wJGp6UE
uoArTuBpalGiE3GU55GrMSq2eyB15xn2NLW9LBOXDGcmuf2S2S9RcDrDYQoGPGM9Nc4sHfuB2jkT
0zY3Ml70OCnhnGlLEYpknzrbYMGDWtr31VHAVSpsJYmY9g9wojSFF7eC6Pj9mH21qPYFk4eEV5w+
vngnJloR2sb2kUzl7s5cvJnIqR3inSrAvcu1MLJTVQ6t7N9yIJLyWg/e5Z074/6MlbrFib06h0SP
bNqlOEslzlxNvTNIhL5rtPgalEOtZK7eis7x5GeKtdeyposq0LcBi/M9vgnCxZD5Y42WgBTt/0bp
z8ej5AmQOpy/Tlq10xyREuBFUWTsYZyRiB+ZZbsRf5NUy8/ggshyvFxxtZ6lVrzzGn5a2dMZvsUn
B1p/mHVEFTnN/g7unqyXTfGDWfMqNs1UvCzNzFqMY5zdwejHT0stmXFWZr1NzSi8OzrzgSKPQXtb
T/KYXkPTrez1fAUzo+zrzFEAuA/EYp1WJHYPVpzRA232hBQcad3hQHsAGArggq9qBDPpvjaGjznv
zNK8omMQrBYWhQJWeuIq4KTKI0uIHmX5e40AVxRV8MvpuQzO5vm/Whl85QcV07f8VJ1Z+PThASP1
KAoCQM+S0jWOrv96uwz6cjIt/5KbSauOlFYUZPuewE5e5iSGX0YWyC9/htFHwDeF2VixJhMAlO3z
ChpHJBXGVjjFpKtb4H0C8vrItk4JMxVPAsKJePZFqnxAYe5XtiuvF08Jgm6tfIGltMQ2Q7Kct//2
O+dy5sJa/GO7H86/6inb4yF/DnZBgHTvr0ulko4juMb0cKYkEwEHJCNzqJ25EmP7K7mLfmIFmb9a
WanpIFtFMi1FFbfqjIMSxZSFDKWTVC1EpKY/vepBpxy5f0Wi4tP92mVYxvJvD76cp26z0GApchJ8
nlCidB69FtCwuac+No6KjrkrWIjVycHkkvR6440zlf5UC4LnJ9nzEPbqE558AsFQOZZbua0TnFke
gZC3D4ywU6rr/7jTRGK3ZGHW883qRgehfscD2mIb9K0HRjG6YBHa05Ze3+z6pewQkrgpZ6KT7a0U
UtqtkF0zPmFy/ejRKjHkCVoaKW61+oMfvz8pGtOVgvExt9OVAboD3S0bAUFpkZgaxz8nK2S7LTYu
+5fQ1xK7DKYeJ01Fs8sFZRQYeZxJXa1uET841/3W+Ir3ZRnjfkiegpILfle/Wh6sTdDrMieER0o2
0YFh2H/5oEXRnG05Yy0CRb8z3HMSy05FmWecjxWlgndnySH6J8f9k++06paHsoHFP7lg1s0Oelkg
M2X+HPUbZDTT9jsh/9BleInHBmLF7t0lZKPVwVJJ6zI4FnbHYWnnur+9uBdjKooS+ystgXA//LtA
8xIA9SXnYqlxBehgh8H2Gb5xjUM/IZmO6rfgDLOd0gIt5iss7hwl64q07RYUe3YhvvQHbWZiGiiP
rROOfrTZTmYJP336uZPqMVCKfBIbmG1n+LrJBCkslHfMWGQV83dHOhnFCTbYytPkm+Y2Heget63o
tpTI+AkQT/qp5bT45kqlXcrJRJjhBOLiRCaMPOpMXTfwldFDtNRAT+pPBR+DFU74Y79B/3ey519D
AL5oCLf6+VJok/eBEjueXgCU2yQpEqGZfxqSdIMaPVACc4n058RaSSdpni3+QnzzjjPbB+MpEoAt
DAlpedSFAtmoMb4o9HoMRcqAcBRY3JKrMJEDaSznqbwryK5uOqBeEQF78HhvOe6CxAH4v4tvp3yO
AuVFFk2a0ilQkvQgqFJVR38+Xa6ghPnJ4pMzOhxS2jXJZVI3MzPMXWTNcas+taNr2+AWz1kMey0S
oNDgrC4Ov63IUTDJEAT3ND0xt3oE3mZ4NADOLRX1oWDucp5VdSKByuKQJHBBErLipRaj4IQD1zcf
C8cvb1jtmDQO3dc6w9SkbU5kKnp7untl8+2jbdVZQ7y+JHM2lkKmdt65N4RxLGyDK/BSjcBpipUV
o5ZfyUwmGR5Ek3PLyX5fbp+KqX+nhQrAeIVhNp7MzuPomPpRXcnVIIBFzDzySWc/W6535oiBitPZ
04JQaRaTi4/eP5p/i89Isb28B6ilO48Vb/Sr+852BpDeJsIMKM826XSgQJ4WewI3zA65Zmizrsz8
GvMKtgbhCGoBD3OmRYWbyxcMyKjrKRj+wlzRB3oNcplUUhH5cGZn6wGY+BKPQ7MDXU4cuqkBi82R
ghgCi1JYOrTvmmcvgzHujkIaQJpdihzUi0F8eV12ZnWkw+Hj+1rl+RG6DqhJzThk9wLkCplyFpFf
Pnln7UB5DjgpdhDxXZj4YCA4+i2e7XvGxJhvYIshE8xv3TFPp80E/DixDzdrihn84DSmJ4JE/ZOx
yzs5xE2KWWdYES3Sz8isfLinAA5x8ajDcJxnCEHWtyVv5hW8VVSxcdsf4RG2AD71QTKNkPBh9p1F
JV4BjxMDvtC4hVbBw/j4NWQUlwIjURlqG99V4lZE2UZvzxhFhDaJLYgU4FoLfxXoXkY9AiVISlVa
yu2tfpI7jYCD3tPMz8xswjo4W2+AbZFLTF8kLvJqh5tVoNskx7hmw57lr45WVSaneblMZsQRVhkB
ToI1Tqna9gOQPicD7k3I6W4G/rI0rml+CkXmzQNlIDumvuaCJ17PhDrX/boSa4ntBSeBlu9RXmCq
XWpX9EDpBQtfx4U0E5g9n0S+SOFI3S+DKWVEdLglnXdW9x+5vYcmi9hn1PG9ZyQ741QG5GM++y0w
sJquHwvGM5EI09qH85ejq9HCadpd/HMXWmaOIscEdNhVPdDMqn1/AsPdRV5DMgTETnYFupM4cFeP
uYmBkBzwcKGXx7pY1IaYs1tp8XTyR8d4vNeUCsSvYFbPSX/v52sdRcTLgDYcWCHtAau9JfaVaPPT
bWJHnGB7QijdGgK5wv9FAtYcJ+8ds2MYcDmrzSv6rkvohMHtT5u41wRSMmReVHYoHx6KCvoii2ON
YKlK+mcxcKqYguykYSMvWUhTNRf7/9o4aD4Ex4fulWYHRIQXJNtC7JnDFEj4TK7WDN/b6H9fd9xD
TSGbidLotFrMu0UVfYGTMYzelxl9/CTNQby2bEynLbFkkluToeB+trld38LPn5ds1KejPGkPJ969
RV8zYHBnQVPXybq9YEoedMKqOvFRaJK4Z1K0po1OEty4XG6ItfzKhMy6E2sQ1hXz0x1ez7iya9SI
foEfUB5h8/F1BrcRpdgH0IM1buGpDX8i/+w7Cy0YmnV6yichADH0r60n+RCX+pXzvqFmSYo9p0p1
xBfnCQ0ubw10B2FA1vq/QYoSyuTapkIRkbSLbliRRJ+Fw9IIiBSPtz++DKGVM1/ta5/PXESmpHbJ
JXHXuvo8qatZmJclwF45wQQmFiP4MZq3lz58NA2/ZOLOPj2OLKtRodB3LXaCiBi+ZOCMD0WG9Hqv
sX3RPP5809MlX75OqJ2gtrDJPB25diDDYbOrXzBAATW4XtO2dO4t259xmrW1gjN1XWTinLHOmYp9
h2bFDBlbX2aFMYTThzhLgXIBbj0/vNG30qJ//kgj+sbi0UDfUSo3Ln1lX1GDghL3aP3sVhBHPn+M
7V4ttVxM86ORYLL/jy5fW9D424CVrNkARlOVcxI1eD6glhHo0AGjab0ItwuNunqfEbNEg8ovWj2L
bkiVRDAzsayYLKvt369GxFOS3tqDQ63sPFYxKdow52S2mJRgZ7yP4/cVlgAPexBorVTLfs9rhoxR
BuGZXyryqxjntR9Pte2OdykVG16XsUsoGvD+hO42YMXraOi1S8SqtLIrkosvpKZhMOBZmnycxQJ0
FqKb8xwfe6TtytJmjSg8dUFvGnBRQCVFqkYC0+eneY65xkoLlDpu4lJIIxDfpBUegNYWWhVUa7Pp
baqm3PKNaM+Wa7txjRzvYBEtnnLnM64/hRs6E0U1nx6qwg4wfskuD2Sb3Yd6TRJavWBFxbEiX+h3
C0wj1AF1rl+Y5IWKCJ+/gXv6eeCQ96bXiYdDtjvCRFY00NFBS6ovItpKSk6ZHogCdbh5Tg6tlhh8
re2YItHAO5Ar5H2UwO/oEjxiKnTBbzn+vzeLD8HiQFfxK/pPrAXTvPzMQQp4Vie2+s28Y+l6x8xz
vzlchnofD+gSMyOnRveYDKPblhlWmDbD/XXu+Y8nvpQFlV195yBveeDcJzALyfDYe02nRl8I10re
B7sE5Os88MC1ApArPdQgkGm5E8OZbMiXLpKpYp+h2NqNOMvdFrc2fA1rAPDQ0ptzCBZYitVrXfuZ
2jjWwiK4Gv+s6+LrbOdIwn5FK78nEhWLcSt119V58VKLEAVlyZ74G6tIiF7DSv8OTb6TXvhlrIVM
7q5fAZZImv/S8LDz+z+N0wcrz7InAfaquBdMkmQB78gO8nsM0TyVFyfoMyUhmOGiD/j0g2wIRmSz
kUvloivdQ1/L51JQNFimy12D50k6wGhToZ943end8YMzCFSZH+iPmRhfmUuwGQ+GunjZlF0ldXVk
HK8G3DkKpe9b2tKZ89jvk3swwAhnN9ntRCbdSOGsBPtjP8LQZ0Rpbg1lxtsjLav7qvd6j8bOAyER
YpkLkawYNsYMlSOALdM4bHtWqlj/bNwRwbB13jfliKr/xr0GVbF6VO5Zhx7R0EczRNjj2zBkB2Fu
gJAVVRR19lS2yKzuGKTa7Z+r/qPYl3Di8rwV6IUrPLMdBSTeg2JME12lpXkcnVbJ3PaDrL+psSy/
BmxRZp7dddMw3YZNz0rasVyGWS67WrN9xFJTxLsY052Bka2yNV4E7qtyEWeJKsXIzlpDtw+alxKh
l0/wtyaPKNIrz2D2JFHva7HijdyePtnzhH7lRA85fiLUnBuNEOyrtKm1VB1lvdGUu3dVw3Qx4pSe
wShK/afm3YJDhKZBST/gjoOxe+LpGfFCbplfKUXBS2J0P2vwsrWhZ9/yfYPJDuGpDX6Flfm2jnD+
C7GjWH4ijVMaSrFLQpt/vHo6HM60KYGIrbBJ6lHr8eVjpEGUQwxqZq1YSS199SiAGOZaqKbyHb/B
/Yq+/l2D+56NeINA/8D2GG2L+Orj0d0Nk+GvSGdNVt8r9gMqDGMqeTQUzUwS9+AH4bvPC+lIaUzn
7UX5t2tnYMKGB0QHZqWwD0CxMr9WKL9UBqAxfLRTfY7MCLqKazTmJc2j+R1nFQ3sGyUH3KQ9Iik6
+ztepCRbbrnTf13KG8xVHIFOyCYVsx/fdcGwLvoxBD+usZ7CCM45xpsElBKC6nZKzkqqWTF6XFzK
DPR2CoBi+eGx6k6B0eYwS8eX7KtZYzfHNvh7isRXIHKsOooin+fqvRurgTql42Xeh+R1kbhZqU/2
7dgGci1nB3sEffcJFviuTviCYd7IajVR+D7R3atX6J1WaxTE/ofPI84sFoy43+YiJHXpSgY5lyS/
qhA8Syca24Exqd+VTSa61Lzevj9ovTCUOwq2WHCwiZSrz8cSo1PWjb+Wo3kvI8ZY/kteiv0j9ICJ
8xxMRt1jSnQBkbSKVxMy+6E7PLd1wpKhL2B/7AhQBg/W+BOP4tAjsRJcqoWKNddicS1jfkmQGV4L
eR/l+AswUlEmvzuveiuH75XwaYMI379ErOjZVeqT4HkuGsH4kKm+47DYNlr4fmOCERXK+tUz6yjj
tYTjcKxUfx4JLvlY87yiUdWPwO2wlsSyiBHDdQea+HzTho8oHbCQ7M47+dw+wTE1vbBCbX0TD+bt
sebynOTmsRh6pjLSGRpohVY6MIWMIjm51EXKJOsYDgM3uDnlbkZPR0aaNQ14qXqlnWNdtpeXvEKr
zx6cm3NB+VRyKCol4EmRKtbVnkRxdx2pKHQvzmx0esSZy7abcB52AEfFJAqOmpN41KIV9nPMI1xE
TzSKFYDa28QFadolus4fAAIXkLzbl+C79ui6q2BUNzkaWLV0O3OKMJSkUkbMAVsIBMXmm1GBBSAO
s+K5SKOCpreb+cPOd7kReTWq39flhYyxj2QWxlrvK8EDZe9SvmG7jQbE6T30L6RWqW9Tof3auJ5x
Nmo994k9WGvZnfWhcZ+jvKNU501vpI0K2yaGSBAM03CTzIHdi0h5eToKjbpellHLlEZ9NjHo8n1K
eXEeYfXqTjLmthvY+Lw2mkFOmdSwSSETCEaIwkso0sDM/jUMTx/3xRs63gse9tO+xUpZv8JHJ+mt
8YhnMfGxGyy52RuhpOWxieVJohB5as4I3S6ghTu4RFArh54GxHnKDGfMsEuxflabFSa/4mmd7KnX
u4zKSJvagth+OXzgabIfz1EXCsElxU5ObU37zBurOiAlwcC94fQZZv1fI/Joh2UML66SC2qYnjpo
zbCA9DUFDoSnMXf0zpFyZdjXPDh0+u7Lak1OftNrLNbXMx0dtCHQrMIFzx3D0SBSQ2Unh6mqKb6P
UjIAPv+NpOLwWYAvyPQWjI6uBadiRXiJufO9rINyxY5cOcMcNsbmdkQsJBAAcnbVQSW6e2gzzdVc
gCWC0asPGoSeA8LraJO52CFB9mp7yiuqfsTcsQwbJKvLNchLVT346iew8b3XCLO5KIx+g20K4sKv
BG/oorL01dOSaozd5lDz7aEZMb6mMW96PPFlQN5eTJJadyO0bOIgzJZ0GXdpVPvSJbtTbPRVIKl3
/Z13CIo+orE/8I9K0myNemPmL8q9Os3oxw+z7eRL0INPa2gwkT0XZQ/9DTcQipYiIrxB2vPbXYcf
F+iAUfMEE35VVYlaV2FAwzx57bMR8HYxTRewggcP4UyKj4Cbi83PFwUeORoJbpj589JljH5QsETj
s+j6qBQxw63tIWXPjk2alnqM6y+4nyIXA6Fz4qjkDnmc6J843t8GfXDpMm/7a+SrBAobZwTRLqvY
T5kUVG7kRJlLFz5zM+JltPJdcVOwA2QCjhBGUdlEgxXioQS0gwQ3z4CGUEgn5/nuwtpvx6yQOkrD
bjTrzEyeo1t3iyCd/OTj487pS3D/CPBVqQBgVNKw9/kkM4xDbYKjOvjn29A3WTshs2bx7mvVZ/cE
u8UBoGT1wwEoLi8zLifbI1BDTiv/NqYguE86+LobJUxP8tPcde/X4e9g3r15af1RBlMgiixttsyQ
609QuhJVx0l7bPdbsDTx8NcnTIfmrpJCOpaxp3inO7Wir7C5Qz6QFDmZSauMz5sXR+mZvhGq4B4C
NBlVu3T9+sulyhgoedWt+ZiaZHRNYt7hPf783J3tGLudSUYjPnqcEvls9nS7HJXpvnzuhY8o2nvS
szNAxOUMx3JmePS787WPUq5wxSXeti1X8t3Xr/R2qkfL4sOP30eZcr68gsDk+CkykXRL0PH49WgW
KGwWF0vi3zZO7ZAIQquy3M2aNQ9RZBpx2RMCcTLhS/cAI9kTlw8ueTMd1alg+35Tclpwsuz+/taD
zW+0iqqw7tTYbMFkrwq1BaiWZDBdMg6Z5N9WBdwd2KKmdp+LJ9k6usOkwDGDidjYgfvet8ORw5mk
xZKaJhN2sxFcvQD9YqWojR9NcduVRLJrSfcKsbDNf648O/AXPgBDDVMNnYYAefUHeVr/cZjZzqCG
qQVtoFih+Ibv2OB63Sw22fTmc06Q6zF/HSygVj+afuOQZNP78IfBhpUgwoyGt7hbPJi70aLpEk6s
V2p203KUw8uJN03OJIv4GvSUOHkriomwcRsy8tqh77makKutDEulMQ9vuM1SnUVgfFcLVPmvG8Un
Sh/F6FyfX8F+FU7XnJYeK5rgUShQwZmAOTAYZkGMBDqhghD6voEVP82dZrgfBKWIjBKQfmgXtKLO
C/6d5a60wWkCSHf2OiVSi9wGPo6Q1rlxzFZ3c8RauQEs736qPc3KXpYacrIfAopABiUmFl2zmrd8
zykM2AZ6amKrkb/qo/YEbzlLKgGxfBelwYP3Vdg0diZcwh3T+br+h4+HaIoRN0BU0vIFxlrJjZVN
rgiNGqYo0AdM2WHhoo3KfZY+blRGipU3nBmshJY+MFRgu2hozaVr8Ue1geJv2zKw02tEynkNdfln
u2/bNld8Zpr9tPHv2BtyP0AHpmd/NMeExxv0SZehWOFPeSUt7Lgc7DMGIWauljLwRAoHzQfaM+Je
2iqIg4o/M8GDhfGMNeCMCln3oCx1VHEh44FZMnCh6MMJ5MOyiuk/a4oWWpDCyWxps3MJK1kMLmt8
f5x5oXPvFXpFfgDckkxZyY4PfczQaeY7lQhthfMaKu+EKSz/WveaKykNX7OS1CCaYumCjWi1xnz0
R/EphSNQfeKDZ4yvM2TM6U/bSET2e9GYzIQ33YBQwwPwa/kzV8wPYtBg6j+4NzbvfYDVS0QMCO/H
Hu3rbzLCv/XNphJs5Qta8C6AqprYRyJsh1A9R5VArVYYdgDqbFNHwaoekp4he6tZldIPhFaLdwGE
xeqMDMzOvlesFodOQxMM+UaZsWmZGMpnVbpjv5Rtyseyjsu5l8nCcVq0eoslMTA6A1mry8iaIk9y
A7PA36zQI7AUWVIhexi0WWv4LdHsmqz9js3XahiEF1Cu+X5ElU4TBUvuiziCRQNe5rkyU1oTD7ex
9z7IdDPLTTvPdC6xWYqa/k/p0ygGdhCXzZmehlLOR2+tVF1gvl1/+FLzD2eOloSchPNMVcphFybt
mr+ECFljzxnLpxMr5ixbwLkacTy+3lbvduIacBE6s1xYv6C7E4irGvkJJAJFw9/3QVDvfpoL9g1c
uMTtAtygizOrcZrevio7YkG9JLwzteXeEjlNuQfyGMUS7/KURhxQEznaVEO+XSjx1ITayxKlCmiN
6KJlPoJAUfYGUg/cQMzE11okKU7FbDC5YYpzZidFBG7HFwLwQDtprOcY8ub3A5KInDMcAOqbVXlL
L9gTV+fGeAWieX2D+1J71fvimXQsRwQ+Mqw/5q0J9GUCJkIzIzrZkJ3rlzNw+l2Zky0P+DRAF07J
98daeoSrWTML8aKJNLFdJf+0zWxVKLtgNtH2GTp3HpeBPmlbNR8LIN7q/ixTWjyUzwY7Agmy0IhH
HYmakiMRkVAPXg88p7p29Yi8EI64yvFj5iMYflRnoqfdJaLQwNIlWJ3PmaKdj3GhEGy546rGTkpN
vnTUSH66ibJUxTFjyjnN9b+EUO0afbi5RrF559EYsMlIqV39msngIS2xgiaNRLtMZnddsoKai8Qs
S+nhJDs4TztKNkq2vk1szXXdbcYD/78IBHd68qbklVt/97lr4Y5qIdojPXKlNWJhHK1o63FYExFE
QCEU4Alo0YTKm/iXTmY5KMMHUtR49EOUr/GERjTUsfu3GxGuZyQhGqH+Tg9BflkHknjud7cjW4bg
/HGQkszhle7eQX+++/jIprUCRXEUtmDoy2J5Snq7T7gEIawt6+o36A9TppXtrBAJbtlRPk0ZGVW0
ZEVkPz0H3PkFWDTyBt4HQcdRJWbDdb4AWmk2TyPV/tEPSyJtaCPpW3t6Iwt+WuduyBKhAkB5ZpXs
TcwL1F+vfvfISx5c+MkrZaL4bgNU1rXcezLwzf9y+pr7Io6QjNNTtxlPR6UrHGTrd9ba78vXlg85
mJmmn0AyJKZfYszl5EGqeAhwa3F6/+hsWJ7k6K/AqVUEZWn+C5P5JAPA2QCwNM9Fl+1XdqNE6v55
PKs5bdfiWkKWmR3gKooc6CJh5vCxstRm8hzD7jIHpDVhc3MjjzxdZstkj4rCLnviySec1qT60qvw
IwqiP1Wb8fTp1KGSXJ6UW1ACOYjc7qzsd4wTbX4FKSE9DR0y8JCFbVNMuafJLIe1JgCcpl5T35YS
8n8j+LD2yl+SaxDe5go58fr3/oLUHQ4XRRJRATjhKg6dwYLHx4cIf5IPbyA6KcuH0nY/OuSeGfAQ
D09scVkgyDMZBVETDWXPJ4JMcjWblMDtJIji44HGMWUHDuikE1FTkRQTuJAxMwo4oCI73rTwb5Az
x60gvBsKFio8L8IhWWnKsbdWePBkPGzdl7Bl352WXkdJ5oMZzg3NaNI7YFYaD0Lc2cVbnYGNMLs9
y9snSbaDVS3wydK/gDN65nMWZJejKZ8AOzjg9kQioZSkiroYzesroalMCqTJmwlPM0GCwaPNUEAh
iCwDip6dOBI15WSXVZDaB8nSPpB4w93OwkhwUMcFvWFh6qsb2gu4Rzd8JiqipmWijOqXtd3xvAjs
AKBsL1yafItdZDak1DfbrWOkdlqZx5R66VPrwsL4QhDZd2kigi285s84qmUTDEgYOfS9Wi+F7hK1
0uzpEGzoQrolfq4dAl+S8v3LHa2UuytlJbuGbibVdgglLEqfwYRFa6THH+Q6bLZWFJ73CTEWdzyN
8DiWy9vSECwyASliuQDJRyXVHkgOCCIYbuS4GC77thAvFyjxAULusM5bPKwjYlVdvVnIK3n4T57R
jO2/iCUxtzKphn7UujzJMnfHEhN2B+CPep0hEycd1BfF1YRGnFY6P18mWaDr2BQO92AF5EIj9rV0
lWoBC2+EZCdsuaC8qQaMq9EMvljsHBSEti1Zx4+qvTN6npwZsLl8TZ+Oa8cVJQLDrypHU5BeFVzw
BopJ/7mBHOK6Uio+YbC6uA2CjYDtOAIPAMyRaEHxMOvW52X8ofqsVSDJjSD9vZfU6EUZ/l+AoLjC
ZNoBhG0JpYZ+ro5m3lGyLoWSngrx6imXsqdcAz60/a/AqDIVWd2x6sotwK2r+3G6bgozPFN4R1pe
uCVjsCWqTfK5S6W7i4kkFmMoQ/UpRyqVYvXxateQRF0FUoGGy+E6Lq4UQ2Pxez6fqrJ5FuILm/+K
5/N/uidiWopaUeU2jp97E1EagvtVh28OlKozAzzfgoVOIniUBsaKXbEnXfUaVAJ3d6whCYPYaCDU
L2c6GzUtszXzao2IJ6WozWnY6PKYfTGeBhdEfuZ9OHZRfFG6EmxisFoXL0HILvKN5UJsmBsChzcQ
6iwOWd2rHZIUWKUC1AHqiCHQ4saQeBbKkho5GmRpJNmPeZl7T8B5smrghGkFA5inT9ZwL24ArBVv
RPsOba6vPEvRx98NXEN82Feq7IZtaxBc90Bhp22TRro3IjGdC8pPN8K+srCgBizf0Q8p7Do6WHDG
FIWk7QajEpwS1gpZRYnlI9GR9OkzIoPX3CVkPksp8byKBv74BFK5KmgiEDKAlRpNrlviiIDOmzCU
LupVo5m6drhiLOffBNI1JHGql7QgSdlJ0opm8EoFNnbuV5o8OG1bw7k8+WEH6kb74EzpYiTUBouf
U6E0CtdzuhpcYkWnRyPk1S2K1Q73/b/VbOKM0e441uoEo2iSku/4HrEmK9N9wjQQC9JWVGyeNIX7
onLql5nra1Q8jqncv+xQwz6/PM+bXo3voDEG01qc7ONymejiJfhLeXCJ6o85iPvr/Ed1hgF1e43e
U2adD9bYRFo93kf4Xsdav3vQXzvolu+ryzG5qRHxcKd6EFXMCdL6ncy07TELOZX3HyC885OD1jGP
zQjqum+S6/DPMMH1mfa8W0+pcjX862umnV0nrAkiFKe+mbOI/pbc+uD6vDszXaSDk729I1QREB1h
SGHWOq75lfxx8et1mVr9coV16xzsQ7/3/1/LgkQ5hbyejOAzUPq4YqPUDdqpMWjs2OS+x3pT9ah4
obSlqdJZGHeoQ971YwVy/bIblMZgaYEVEeowQHiFzPpymae5K7nxt6r8+LdidXm4jArR2GDJ+uEg
Yffk/51RiFJU4IFMNl+ep+Cspg+o86A43O59LwmGHSmmoygGWsVuf+7Iuk93VNQg0OJg6QgjxBN6
LIuPAqsr7bTGXKhMhmg4D2O//LPHgXbGtELFG6ZhoDPuIF1Ddc6dFQIBRWoEs00WPoTjkam/MDFo
OMmJGxItRRowAY0WsSoUgFkggknmBjAcmIhBiHQQhCnj+x/zgiZ4DTP+pQ7Q6Jqo7Csssp42DBjT
4/MRDOhKB/TfH1RDEljhKffbyxPjf5aYqMDjTTpWNab6oFkrDsNz+ATLeSrMfzhE9VMp6ZFWMKP4
6PbxUxaFgOJVbnczbydvu9B5jbPE0ms2ivrcVKpPQasHkkWyZfOe/fBcKZVHdaIICy4+oBF82E9f
CUq/zT8h/iefmQ4wTkvHmmx5SjCqcQRdzx27N310IFvG3MjpuUBNFqWKVdr2MzobiDu1Yrt7hfo1
bPdy6bwMen4vbuitT3Rrg4WthVSdDQL0zoZdmhkm97faXnqTeRh7/qcsbz6q+1/56qVJ9FvHX9pf
N6/CN728h9c+e+mNDAIgENwJB6pxiSbnnf/JdRe+n2454RW7bCCwJljuAgjJIOS9m+m5sFs0Qsta
oj+Db9IEPxZ1PaWhZfe0j0dDORNR7PLEF6p1H5nq3WtLbMavq1TTehqavu+eWfouLWV5xq8+PJjd
ZNrVKieo/tZGDZSAaHkSRPf7QepjjQed8tXCLfk1q8qpZG8GORS1Uvky/mCXREz7XEsla8XyOslF
VCvmIfPoEGTOwomjQhluOZs4g4zSi5/GMyTyGpdNAUgt9X/EN7Huqzv0+rn4OuecwXzovbqXk9Cg
SLXT+AuW6VH5lmFyWeQG2NshMx/ZGdeQ0I9BBdBQkZDNm+t8SNvSQaImqttub/yUQl4LBzqQrIyk
bsg5bWpNn2J7C4CQVXQ7m3ox117d+eTQoInYlIFx5hlCCdEInEEBFQEaPrkRRILEf8Tx6MC3H/Cn
V9HdUsLTe311wEG5maDmN4ll1pXKKoohGQ0MsNp3WwFrHITXKEwE7nDcbtgyL2yszYbCmrE0Nw9t
gcNI9Sdqb3Y52TU1UINBYv3ilCXHvPhFyhi2xkrE13mjRS9ONzIqobZm4Z4HZKHncoBjMjQLxcJS
DQ7jgLViswPR1zt7FZBndB8oaJ+CavUo4LIgboA3OPjFuhAMPEFVAR8gPEJZKbvZktY7srHUXtBf
h3ya+37ESVGcwc81u94rGApbk2AsCw4zGxglb2Jt1+8rdmWIaqHp4pmgqefj96OkYQ9Fx/yhjEX5
LSwgi2XBS6gW1bidT2mE6/xS6jv1qxF62/FRjIqyfMgeyRb2oPEQulxmlhy00hpfiEpbK8gIWTBE
ESWE54+1uFdcf/9c6h0jjSS8GL4c0LMc3+LDQ+rvZISyAELFiIeauD6kTwsG9rlZVvDyATvlw5pU
uoflnKOJ2YX4ZouqQtlKGF5LWVurItrRrBb2mB7byAdXRTHXPzTP0SzW+KEicMKF3/fMEhilXX59
Se8EvzBPA2OTYQvx8aFCQmwUkwFM4JPWy1G+bzlje0TcQhlClfvURmIvZ/FW7AO4Cq7wuLdyCwMo
fmX09mlwBRiNHS3nS5GEFZjTMlq8yN/rQeWQx8h21ufuUeO3wrc33CNN1+S7rxaYi0jnr6qFG8cF
gBq2gV1Birdb3aUFtLDpuRRQNicJs8xtUjLGc4VdZI8uQShwPTSJdOWlvD0wV7T8nOU+rA5OvvGS
sUHfWP2tiG7hhxnlrETOPq7jpLRAMuGLs4bPAyocS0XfqHaecgnK7VOckblhWwdFtnz7PGEYiV5/
qfZBCAluHJ5ArWWgJhyAWEdfQL4EQmQ85m8eHQBRsNzogF9gh/BLs6gs3zWDLMaU5KBMQah4gOT9
Uda/ai/H1eh26Tt85baHyz8E/I3B/RcFIqFgRkkbu8ysvRGE9spSrluMiCMFHNpKnXm1FSdc/t/1
angOWcFNf/5VJrNkxk4byeNqosp15EvpzaloxFmUC7V43wr6auLRdhNtk43t5mAftCmQRAxCF7U7
HsfF6novBhN2r5gqFV9KVTRZMPkUxfP+lrcaddvMuKPZj2RPExB7mBLob5bNZeNvXBHYV2Kph+43
tE6VMhjWwVwSwat1UhD/OjaK022XhMR+BXgtBrBiYx62gGVTpNHV4JQVgb8auFAeH/zVXXqjbJyB
5tuh3aXX1avbOJbdtVt5DgnRa41mz8LizHDoLjVighDQfclN2dLupW+ofdvhJe0jhx8NOfDj+bxw
qtes2whtjHOfNZO47S2oq3PLEIhXG/f3g1imMsd5x9PQULfG0Kc2jXn9WmTTqlYv47/5L+sN1XHF
N7pPOhzvccaLBSlH+sN3A7PTd78MO8kGZM0vGu60YYmEmPX/cQiqKWbJuiXrEM6ppVfL7BW41I+V
QyCuzj7jQvftWalgpR441UvG6Q8Vo0S+EbeC3H+rguTT4aGG6HvDEVYzpn2tswuYusmEt3uzkdDw
NdJ+FkzpGk5lLmNQ7pOnwB7tVKyE89beVDIGrNaW/kCXI8Gl7lzQULYYRw+cW8ue6LeNR1sCyahq
tDTzpFVH+NtCyzh6rBBvn72b+y9n74kmYkHkuXaM07aJNw6WbaOnl1/V/GBi3RbrRgHYiPcvVJ4i
XONG/8Rshz/yT+6Iy85YXU3PWzfE6xcsHGqFz3qGBNLoA8jvjhMCZ64mNqIcsrp3QF+zloTs93Bj
taUFoiD23FzZUt100+WFrU6Apz6ytT4xGZg9XMxpyt+NtQMg+1YDw/Xhpg3GQYtFkw1yNPVJmW7g
JhFwfXfH6U2mlVARsu84mVlTny60cMJjkVeTwK4fkDH+C0DG4ETAUJlGk3DbnBDwRbmdXbuQ4EFR
85apstrhQm2cZcPXKzKvAkxbYkqHHMsOWezEKJ0781WVMCMrvWrOhZug4DZU6hKYeAUYkaJoE4Ix
38jWIrXOpRmnkrQBj6kZQWHzkZIraT6KaoWZBzuUXq6qNbRllxFTJIPSbY3IQ1xCFdbHmI1RUQXo
eV1ov4IzQ/T6AVY8lpZJoTlzrmNM7uWsTtin3P4OiQf435+e6iPvLVFGsXICmAjMwECm8kM5d1WT
skdPy/bfhkj9l+MytYpXiUXGQBpMwMAeGD0sb7TThrQtxYNecqcZjUPlUISSooXkSIUKY2cXiAFc
H6HkAK0uOyIS0k9h8nMRHHVCuG07xd9fluxtotwSPic1tvI5QqQhlPaJdbEBnPRG0Kgoi5GQRZDy
Vgi647PtsLE3Q7s44g87dtnoPTI6HRKB5jS7GrTVNTYAOYQMTHv9N1mnEyOT+zCOVOE3UZhcYjvI
WChCDPF5b7AOWXZo5C5NuzXqGhNVjjmx5gFSqRd4mJJBVO0nEeebGbIJqY83YQgeBfLxfoRWrKQm
nCJljllTXtv919529TslH7cWAXBzW9p5YLdYxPKB7bTSNEcdSlwvccyrieY0U7+CdtnZFeDfu8N/
bofQ0RibaupZfVhXC6aSrPnPn5xQvK31hE+glO3CUI5SCM1zP9H4kwZZih4jZOv9VUjHtslltLGd
Xa4kkJ+UQCAJ6PuKPjr+20jZ1UGItjszN3W2LDPwkc0kxmeGVMFM9jvbX9YEYo14G4smx7khjI39
mvTXGjT1O50nUu/2dJsTlf8aCijWKCyCVPrw5J7N63ps6fz0MU0vkA9TFcFCw67cTp6XiTjIFfTf
6NMhidsE2ArGKqGDq4lk7S4OfSdxvcCK8xM72F38zWopXyTZgWqkOZwoLuAn53jrLn2RhC0AK/zs
sVLKxIVaIUTrwOUCN/kzsm+DjivHb6lUl125Xrh6NU2Bnw+m2Tqv+BWFyeXkyys1+jvPPQzx0hgg
1naf4mXnTgoD15Q9g+mFSJbOB+PDu4s94NZwX7Z5KxuETdxp9HJ+6b5M8v0u1lfbcOd4S9SvHZgt
u6z+znZYXWO4YDIErCIITAyj42Vk67kn0PIxZYOVPfBzRL3d3L+L58l8EGFWi7G5VwlJ2tvPm39C
u3M7NftdgTZdleHxD5oXzXV16JJJwehPYvyIPoJElkF035uHbIzNl0Tu+QRDsU47KmL9TpuZ9grz
jpYkbzbBF6osak7kUX+s634hN9O7YRpMHlB2t/zNHt7VCnffUP2Rpb7sQA+ka8up7bdAvnSUtfO1
C5Ku73zyLm3pJ1fPbYgWdGo+y3iEnzl9WVy1u5cIYK95rzYCvtG3FeUXkj9g66uQKCexv9E+vV5p
zZhjuswoMqN4VbeioHNFTpcRJymXKwQxiMteybPwVbodZCp3AZI7CdUc5OqFtA/3WpPV9Ror3NVP
m4Gb5LElAVqjuJVM1yCGiDQSvug8hlKlCUTtYtsD6Hm+Uj39IzhlIk3ntOWq4myObOyjjGWtfSn3
hVsQ1Q2uRwDheSpd0nsbBDq7GTJAe7y4EL3Wevh2om0ElqoGmO7PYaDjMk+9b37mvJ11S+mlQv97
CokNRp6IOYCBPSYqFTUjF6viA32vzZFzSggDpzG+nxww4Mqkigv6XgicdAD0HKOuP+LKqmVeO3LR
ImiuKljCVh7pTNB5pA9UpoHtm090HEc7TrbsHo1xOVxvHReV0Kkyxo+o92M2anMF2jwVNByaWQDh
mbDLgjomJGvX74mB6nHvhm2Znsvo4dvionGrOXdkZksMngHaY6MzTt/z+Y5/YE+ewjoWNchfKfAm
kQA9d4SkZbskwQt+uDKMhjT9et2GejTvkuHPovO4dccnIGTxe4OZPaFmUsYBLEe5BUCPHPzVz+sq
os+Bdb1DSsA00iltOm333BRny/qBP/JEj5gwE4k1qYYsMISV3aGXPVMKR3PJrj4jtOKxTF0jtBzw
KB8HD5jN+av6/yWNZyVB9ftaUYpN3ClRSNX3WTucxc5r65EJmfdheD2LRAPrJ2+y4upEPBzMLE18
FLZAC92p6bngeg50boR7snsnnAUEaG5GGvZ1BoEPtxgdofRzP/4Ylit0Mm7Bty8i69ONI61wjbrd
/qWd9S4vvESuVJ+fsXDeU7lK2wsHU7Xol4wfRcXuW9aNba+ROpVOKXGSSFhmQYDQTX5Yaj0H4ChC
PrfuP077HBLn/tpxdymGImm9VxPkd/GG0gm21FynI/mTY3szLLGjJs6oArx9rP5scXZNBPM+So1W
Kc0AIWB1ZTfJI3BF3bp85DMMYTG1z3w7Qg5f7lo6yj/jlvqgGYe0xYCMjQUE+q41GLFoOyVVyhLY
+HJZ1hNT6T9noocOWu7wNZwNC3OvSsdCSVS19syKRYAZ7p15QPpcnlw5ZeKoa+nipHCOO0nlC1xa
UFHNH1jujx5nRJ8TA7MeGB1TsyX74en5k7A1chX+wYqBLvEyNZFMadNTD+dDs+VrZR0BCGm2QEJZ
mtvWlU6ejXeFedief7IH6eTgmYWaJFULSgPUolDWvdWxKbtX0cHcqsLJ8PNivCcufpzzmvWQVcGh
/bwM3pTxMkQj6Kxk0kZnc9ElILHWg/rzXtqEj7TBw17w1AgP+efYnqOJYqvlXkkeqrYXONO8nmsT
S1fQs6hj9vVjcbCyX6FzuWCG8EMMMmPSpV+HekFN3og0UhpjTaeCYkYxALr10jY7spRW4FlNIvz6
tWX7805kz2YocWePzoK3ffjDR0IdM7TC5T5VeVxN76LrLJ6pPigP30RgvjulMjjDwR4Rfbx/mO8r
T9KHgGaw5+Knf7LTb8hoWaPVcxQ7WVJtrfWCOEZCKSLVO3Dov+RtGAMsEZMvR1u8//0OhoAcd+cT
jkZZenC1anX3ld8DOrP0dyktbWh+S26BuDbfajnUqfP2EIK5cnXTEsRgf7gjhFREDQ1Yjg28SNKl
mObW90OzIAKJC6Q1O4ZHTyEzEfMOXwdf5bDIbOnYGDugzUOdQLnwHey3FO27h3tAkHZUHqRNVBsi
oJ0pGrdEDmcSUB+mc9/zoVUiYhmJ+VjHwVuVlezHZClbDwn5rhsn9+GgeGipxafGSvn7AVbXvKf2
Ibrqld0KFm2gAw2lWWkUnKfWN4G0sgrshmxPVw4H0AVJwcpncnFn3sn4zYDuWuPByBza48btJZI3
Dg18sy06Md7+rr2NiYVYvg4mw3EustpLccmMFkfNKHgnU6tXzRBeXesUYXJp7BPm7uUvp81rfZxg
dwbnSSoL1uHM9qjMDVA/UsbxT7XdbPtwLsGpc5rA/1x4vbRq1Dgk26iysB9iNgrJdx1Tts+mYtyG
bKWLiaZ7gRLkdDKc03J8VZtyGaNhg7sdz3Jz5L07vtSsJ1sbsxWnHbv04PlGVd3CA+2wrW7GQGQN
0FD/nDbLS1hYz0YIIKiUbi1HDV/X0dSOn8aeATXv51UFU+IAEs8kcWeg3KRRcnGbMHR6BNoEdGYe
WqJIr+J7nQWRrzEyXwuccZvMsQTybBlU3wTvYm9IxTSb5m8qvGz1kYvkk302mLuRPPS40ftu5FU+
r0dc7QIehoMjIiZsACR8ZfSxUt7/AMf21KUDSj61lXpky+xiYwdcAgy+9uvsvFzomVd6VKzkjAxa
qkeTybctyWSd07Ye5D3uAXWG2GhzKuzpJNfz+InCEZ1oXPByKqwrMoo6rCx6+HLDTBot92QvM7J7
RuD4qb7jpWOjasZ4SBheQFrffZIKW0BxQgfyYw2tOEsazMzmlIkwXw5eNtB5vRXOfaurXCUJOS87
LuNr/g7z1Hv63A4to7SaPqAFhfO2E3BOMHBMQ2OQ1iED7wG0d6/YcqJNp8P5t5rbGizc1/shaCcM
e/QEmdAwe4z78dbx4rdJsfa2H7IRkEug9n+PciLsKYTf9rZvadpq+yFwqO05Uq545ZaBJd4jrLwE
RHJBoMfKgCLByyTgJeBv9B/kpNvvU/TQ4S423jfU0o2lK7fD9l2CqkbE7zcUSim9uoVCLXHSLphC
Mp1oNAIHMy3DwUo4Fp3Q9l48jkjFJzNl10Y0OFDyX7dSl1r36bqgyNN4cJm/3nEMWlPAKMHREmHF
FOxtuwL6L+gSvKJt7Es+7q9dpOZTxBTzKj6EsmSa9u2aKj7G+ZSiCMKLBEFAy9JmD5XPALnYutZV
dbfFGEwRoQUeu80tOPf4PZxANJxsrUAL8Xng1HnEpodWN4ogzIgrZ0WVlfbAuEywmnPx/VPgMrq8
jsHtrrlU0d9N4+Q70VPkNs2ZSHJ4p5zenZPAdcRZrSlO4Iqvddu3H2AgGEBwwCuvGMLBkEDyNT+q
68K59wcjLj9FY5lJWWpKOvSJ6cw98nqT1cdrb9+ONWUKRTgFMmD4X97bp3ALqtT+cM0EXE4pVfg4
QWhWoo1wYMmWJOaPYH2M/eyFivIbW7YbT16Zbt/lZPSanUMTjmugzpz1mYeXGFYTC2A8fMBlxM3o
53XPTDiQ7S1eGguhyf4LfpniV/chlBo70Sklez09mN23qFaQZ0DkEgavibaUIyEwEWrdwAUi3iyn
rADaQyHAI60t4IjjViXPWmYEohlBHjLQEJ9s9DHytdkd+bw8KsqowNbKoOy0rLWejtsVCKE+gI2v
BsaH/uhtJZgYzlOCXXZDGIkJIEQoPygthB3tQ8y5MH5g3VnJLkMRxR2sCURRn7CeXsScOf59r7sp
eusZQyoxa2xadxUUohzbEwPaaFsyNYfO57o0lwIA4+n/BWyST+B8i7tnE1ORfg+l45vNZrK4LuxI
kMk3kCTHJaxE6fcI9KM8Ai2TQP1mhnGlRLa29gYghrjmTD9BvxgghzsmAbltTQP5Oz0iGmFpn+Cq
YFNr+B4+pQsqQJ/km6M/PfmfNvNo+0EmT+XXv0zwtrheRBJOuwn0xUkXhaSDizAHm1bmUm/4kf5t
ah1Iij02RwW/80SOpi0b7KUgkvbhNR/k5kA23BpBOrs/yInCzmMzgavNi7sLiFkN3P6bmk/cNjdz
6uTubeZl4128rAqD0WS4yXoasEN+wwwG5o/FMz8xe+vx8i2z4L0E8cMQXaIDm3qX+sFilOdDz5nl
oJki98CJOS9f8U8j9kZ1zQDthrzasKP1FBJHKacLd/uauKy+OtKugCf3VH6HWnaNUUtxpZgqCvl8
KEDv/FS4Yv9g3YwrIBMNSSrWwFP3sdGQS0wuz9u3F7WiarWzBNCuYPrFbZcFWZXURMwLgVS1TBjm
OkeP7RMecMFA3Wjlmr2f4HYPIjWeg4Jg/OigO3zLsKBmDxNcmMkvw4GSexSqS0GBlFAgnP5ReQ+6
/W86Rjy8l2ik2aJFrYewaYfCc5T7vFMLmEJw26NXxfLo180XBwNelKZXkIuwK0ZIN9f4L+SrduNo
qqcGoxRrIEDGlpfzoDhwwtnhy74lpV+zBSgyZoJwoYSdEhzTyxxgEEOqbG+fmL1ks9ZIOaaTzt3I
yStbonx/rcu8wmZbOQfYow7OF2erqAURQeLd/D56hvvvcskfg1cBeeXmpTpfUa6n9ae0OxsqsATo
ZUxmrBUl/JYFFDwuOlAO3O04F79RFYo4Mt11amBSXBkQU/So8OjLp+pTzgZNdP53FBfAMa+WYA84
yqjY1EetNGtVOkdiWNMxQmJqQ4hLWcZeH7ldBL05pqRd3bx9FuLG/gA9tj5bs9+OKbbVr5aOOHsZ
np2JwIjP7syGPDtaiPKJsUTklp2Bb0hcrVS1SYYtoN866EMa3EmUarrLV4c84mspqaOSKcziyGNB
fXp6KknjoGlwZmAtDBsazuB/PEbNtKmjxSGZJYGxDZoxao9hLxFcoQTW+PupHRBvBw0565zEEsP8
mCNTKDRnjor+knSQNSRlI1ndxMceQx6lD1R/xTC8bxZQVWlhjUxVgYSxr6C+gCT0Hg/n+/sZn1Nv
ceUur9wIg4LpC7pZ0XnFYKTBL4ucumG0lBKne/dFjq6C6uP5AEIZi7Ruw51D+XoYJN6qVDHKgnnm
A7wyvK7idumEPBs2iLbZxbP6n0ygkb6MX7/z8jmQsS6a9P1fOG78hNTXicqSV91oKhEXKi8Ey+9J
OP2ycX2oK+ookyo/Bw0PfI0jL9dbm/9vj72v4BicJr1wLfaM48TJ+0gmTCnzuYCQxyruo2FhFpN+
GUT4hNntQ+93drw/a3iYVctNJyLEj/89TaiDixXznxkC5U2JHDeGi6bCUgDEbsQleSgQahk5Aee6
SwPKLD0pSKwPIYy0+qyolAHK4PR2y+YmN1WxWswLALn6dmQP8oZ/jNlYMj1YzUS14OcvBk2TH6It
YPiGs+wtSduLDYThKHt8uptV2h88gkCKXEg6o08d+OmwPM/q4fCMiN1yBLQpdMdLXZGeeDQEeLA/
okqgDiQRYqCDqAZzGX8A1td72wkmo3oVL4G3cMpWhCSVXQaDJo+y2aZxM+371eEuQT0+1dNbHrnm
unjs3x4hh1XTpYXJ1e+G1HbXPJP2cp3R+l6EP2FEDcv9PpE+deqLAgTdkZ7FDskqkLl4sH6UogKc
FLD3PEDHohwhRTg/5dfvzEan3f3a7foDjjJK/ikffNrDJSseMDeeHOOI+ZFYzgxTwM6RNJWH2JvM
8ZMB9SrHGMCiECM9MP0vTzt3aIzOOrxGhJimke+i6jBBGFwoU37xNwKT/zA7olWHmoVGOWfr6FoJ
RxKfnb9S1QUHZpgmU0X+MppvIeu75QqV2v/8PWVVicyYeMDyVZRB25rafoHa2rObIagzn7T/U4lw
IVhQ0gZv4arjd47Mq6P4IMUBVDiuY7SzfpV2NqE/qKy9Y+X5RkQ6/308aL2qfBfgpdGo4YKQJiOo
iBEcWhByy+b3CoIq84gI4qvlneR/B6QmxHev2RU3gDVFWR9YeV1G0GrBXtOFw+BwZD2MQZL8tWGU
rxUX8uXblM4fzmC7yRLcVcaakDb+FTDKCVPhLzy3sxfxULCZNE/lmmrGkR485zHGq89lTJ38ra3g
zuU/o8KQfkrfDcoy9hkX8StwSLq5RR/e8+zS3l06BgQABdW0STEWd+6ffBHSMaAsu+ZyDD+jkMFq
M7t1nHCxuLQK+paHVQvvsiXfbrviuekUOV/J+Z00jYkm396PPNsfZZNUKGs+tZN96B9tuBpzuYdS
IAmn54orGyLwQKfF2alLmEwYCsd07GukCApIMXPlhIoboaA1TCxoPcx9Fv9H82ndaJq2Ru/pim36
DVs8wvoU1p44TejL4hCre9t5PU6++Us5I+0eCISsDA/AmojWCJM95IPbmtV2DgdsRQRqjjTlaPeT
wtp69gktbcfsvJnlu69I4rjyfF/3SonUuCxSfw9LeLx6knIZsx7ObTNd/bYWoL9D8JTIzMyW46zk
yPGp8zd5yLb2icmJKb7QGU7MkB8lFLAlbFfBOPmIzztPtZyvAEoqvMCmWXHV2OCNcgRFMLwRpK+T
166/NcQQ5ZvIP2qaRmQtO/CJRzgQEGPkGcoLKkKkxGbqlMm1/RSF2V/abyjgRSgvufLlRQfU3BZH
DU27YYiT8Y/XBbwGYELDWBS8O184BTJQvf6HMl3XEynwkqH6PQSsQfuJVxDIG8OCcsw3dUS9n8r0
eZk9CgmyJrsPrEVzGgNfXgbro47f/xvTS0xkEhU/2b3ZGcqJiBDc3LBjalgfPg4chlzCDEiyFCr/
CLh0+36PctWL7htktb8VxoDhzN1bhOXxugfDv3xp7fyHf2F86w5C8sr3JG367Qhv/78IqnUZgBg2
eN1zGFyPhDwSCcWv35vvDbUL6LIv38xiw8p6FoDH3I6OWUd5u5cslrIj+HKOe+ZsgdX2lB89oqg7
LnaFTW/zJRdv6shUQM5flkwugyRQNjMJzn1Ioe/z6mC0N8sTHsjgzha5KREu6bzVvxHca5W/zO8s
32LRV75oYR16f4qwzvPxXTR0cFwoXFpOP/2Sf4shlggRe1szmvTRCsAkDg5B6FoL3WseENyiEsNV
ptUfSvyXkOF9kT3ZoMuohpP6ih/pUdTiam+kpsEIORI1AITqyZJZ5kw8Hv1r0DgY3pj9MdJtKz4A
J7WhNzakrGvkeCnYUb+ArL4LqvW0N+3JXScUGVfGBJ34yqPnOqAUQvhmPUb6cI5Q1fUPtMvxeawN
4K/PIFR81SxW7dXhZqkQTIdJ3MSBzH1A4E2dNcIuo+HqLd7TaLZGa0G7Vrlf3/PpGtX/KF/t8b/e
BCGE9CJAkk3Bkd7TJ7amkt/nJ7bEwGXjqbodCmIdEBD9HHA4sATZ8QHmPcCHZIJsG1I+BKckCerc
ZT1LqTmDUPtY0+fTTq7l7B1Z1/mj3TmzH0KZqxnWV+RV5y6h52AxSb9Zhe4PhevgY3xuRNvi686Z
sFUPvbpEz0JvK4QLXANryVncTbAmL/Mw0dnhE90qs/lHLYiNJNllSanwEIPd2JryAqsUdsii+jBn
kt71fl1n59LuNZqqd8S6vQnur3nQLNq4qHfufcZ8oY1PPb4DjlqeyvC1w03Xesif4aqJpJou7UZ5
xC39zNi7VJ+zlzXvqP9UaWgup7QvxWXAKvrOA45FTlveyL8Wacsyd98t7LNSBt6bBSZt+VHteLRM
46lI0Vkvn42yl7vF115gvkh6bEqe58GD4rl/3nnyCgNZsA0WrIGgq8nppCNKV3+8MnkzlgHsb6KU
G9yRFKOQl80hUKTtnDRjkAdgLiWDcaPbQq1HeKKf8EETcHlCBOU++LO7OK7biA57NGF9pvw0zSUX
kMC7s1F7ImvnLTO/cVDZeeAt9OyHA0cO/GjHmZgOJSLiLykH/Hux+ZBuuEPp2egwiEy2d9dIgTka
r8QcZrQBGMxEF3+/3PE2XGgOFAXtEQqwT9+9Y0Swlaq05+Ol7t1BKx9Bb91K7D3kc8d2kQb2Ni2b
4eG7A1y4T7rqnCOFAgeVuyYkJdWAHP+ydwshhjfq1i2tTPt5gglZsJUAaFuPKomMUBJx6B52m9Jg
YZ63Djz4V7cdgZh9GTGN9rMzyFx2KCrLwSUkKQkDGwGF77Cfecwl+REB6dItFeQjKRUPlVKSeDL2
k8vTKtmmfewlcYZn2omDS/PZtlegO33qNbIWKMXj0Q4QBpXmG4SIg4aObuk76wyDylKuPtn9Vbu7
IL92a/jVkeonGL/j98C5Qa2vXDL9Rej4ngXwDUJxs8XBh2yTDWiXis+8yyFgbI5y/kI3JDtx68WB
pRboc9Nkx/rjAju97zAa7aJqj51DZp8FZKoMjNaUxBdAd0GOpwu+73/mCUwPMLkAW20qAG4DTTpr
FHTwmvv0u9ERB0Hy24JQlwaOl+8XXrWne8rQcoxfOanQL7E/RUxiQ3s3NK3TPCmUM0tuB3MnbUq7
ROJ+tOUzMXALQLa04wSUmo0Tp5AlO3BDcBVYEmEix7Rhi6tdVz5dZXtcPqom2FgnwZoTeJJf7b+4
+rqwZKjYk5uDhrVpt0ggTzu6GpYm8w28DIiPsrZfuvuHFMUY2fJCkCD2Y+4iFDgYn1GmqwPfZVL2
pvZmAZIRlMOhwBeUV8m+I55ojwzxvLbcLQOSRByYJaQl8tOtJqWXwzYabbKGmH4LQqqpjdaJ7Wqn
u0r3DEzhAl7uC1p9Xf/NUdjFcRptj6UHQxoJAp4/JAIUtXvVVyDIbzyA4P5/+bOqQBBiGXra+UHQ
HoJ/U+MGYj7Rc4F974Stz3oLNcOCeofrxuVoSw/brSIRi7ED7PiLwZ5tqh16/SkYbE8ntKa+456Q
GTTxYJUP3T4LIMJC7DFpT5fd1gZLHMykG02NTpPGUxZU9K5KkaufwTG7HmbtsvfITTOcYpMJDepx
bLN57xPdeqhY3VkfLVmRUBI5Aleq9fUaWEA49znYRylTBIxOFhQgxqV7/1HtTlwl+i5qNezli6cW
NjGCQGbalbAxAZT9uh9RoiFVP4KFXsmOb9AzZQpnfb2sb1ip6Zrg7R5fljPsa9WzepZX/vpbUkR3
wtyRdBsbIbWU883nbIhpuq/DrB2sMaRxIAIirUtgqbxRsa812i5Wze8BwFgDiJqQ99HPaSnKjjEL
apjs5n82oBBNzuq22E7t1VRTaxOQfNzkZVhv6VLczXodD3pVPBu1J97+4przV97Ssv01v2fI15Wk
2LBBHDMGL6Xq3ywsmujIQZf0yexjaEa4z+u43FZQU6larHAWiKrVEGyLbTJ/9+QZ7PegRIEr+KYx
VWLUSlJ/SIjH/7F81ZMMSf9eD7TmIf0TTRCjbMYI46wVy0xE1VInci1N26tQ3eXncYVFGaHrV++1
gUMTnzgQTTL05y5PIQn7ybxNrKO15JjJHQiJfiP7HxhKzjMtDsqxpdf6aEsAs8jFrhSqk6sBn7E3
j+PF66jaELCEe/1nXNqmFU1KlfYadiUXXiPViSXvbs8+jNr1ieeTzDKFJ2mCYB4v9MVaoGebLBR3
UL5aF1gqRQJClmiG04rgQqf76oT0z/jptMYS34riKCIEiX6xGKcRaLaXX4MplcM08x4WYALnIHIv
9D6FU5tDSc+lw+velPAho0IxPLqJEW+JSopgrSlw/ShwfNraZJ881995HW0kQnPYtycZNqw6q3lP
MsMJGVJRAmxejlEECWdS1DNSgI1oegIyHYtUjrWNj++dT2ZuHXSCJeuzhU29l0es/TZ689BIKAUQ
Oqyec9PHUvgsI6voXVSNiZ1fOg+2ykvwXPq/ITqyC4aEGx8CO98j5xHUVl7sUI5aa2Ya2ydXuO6v
oppGEF5QI2Nqmewl/x3Qgto5yQHJW3ND90qrqpPzO0GBmMMCiktmxoxvTyWRoJnxqS/FDVelJf5Y
Jn2Uyy87Eui+tDtSJRZBHdebgbiSQ4QeG1D6LRY2q83m/I56uobtwOE8Q7RgvejmSOXGmPz7zZk4
W3PlpAbpRVlN9xmVRPvc0JXaDekjd1CkL9PHIlRu4G2mVEPVf6cBcXOYPGE79k2WCaVStVjyNYRo
HbWTi7HrxjO0ktkQ6EoS9+agfW5Vzy4vHePDOkF+NU3dccZuX5j9e8C/uxkOF57KwABEIp9KJeDn
tojoKx5PK3y3TzE7n3tien6qivvaA0VZpzgkeicga6bK3Y6oDCGsr8VqJSz4yFGCCTWpdnVfVhem
WUVmrrkoc/HPiZ0uySoFFoeYx3EAiTqGKUcZVaqIiHov3HyRTlnSLPjlvxnqPk6d4qFMNhakd0o0
CaU2IDDvt+sxpehEz+Z0IInwVPJdzGavFFSb956CFzoPvJ0hlI8XPaK0vyMkdeijtgL/7GNnmSq3
f4Wr9nXyhiD9iHilZ/Ufsf895SIhi0rSY5pniNDhRGGRrxKfqhT0xHMlY5CUYJLMOBJUr48sBZ8s
yW7rzDU+LkvPx04VROME6nHW4v0qVP9wOhvMueioY1/GftFO7geOS/H1UeCREXco6/lRSaxPmB+m
3gPTdm9MZEmR/2qpO5FrAKMwQBmmFOKGVF1LZ9ZOqq0TiNC71MJowx3DEquSfjqBtRFO5p258W3P
qWQehJGkyx1bMyKEAK4axzogyTBLOfY1czTdD+NgCJw2f+X72PVZHh/+qEsOW5zNJUAGb/mx8zo4
r2fsht2N1SUJxkgA9dsglBe4+UaZjCGCRVLtblFWcXxNRt1l8tClE1HOHZ53cKcfbP2kd9IJRLNE
ad/MNa+j9hjSfU4dfx9vNi9oPXj6wYzl3aHYEJreDbQPVOsSMumDaCNG1DHv/XCeVDk1Fe838uKX
jy2gc699GN2BPuMkn/cqc9ycPOti5UFau51PHSKvvsEHLpbYa7o2RjVkRstSZfLK+vyFzEiMN0Gg
bLwZTxyAPdefQyfnm75YGpP5wijjChulmmXy4NepKB76xFKuguswL/ONUzFIGODJAwmqvZdGZjiP
nHOKDNr8XczXjkyHUgUPs9TrF8CyJMqtTerRAn3q19/c3P3ubmHUsVOVwR42G6/jKy7ThmGmPMai
ywOI25b2+CIOoc0bhnxCUhh1x4ttlSu9ccJACDFPPXY9iMbxzzsco4teRz/j5At/kyOjL3BARjGo
t2u7H+MtBC5plMWZaDNWJ0Vu2NOmfvvIllwScQMnqqrXN6OSdAn7wTHK7k33fAxQvM4pyxul0EyH
bRrjsnxR5hh2vZQalXxyl7aSIYVBOepmz21G99hzcnbU9LLfHLHe/sZ18KgPzIIUjcJ9DtT7o0Yv
A/OYefeiszA63C9NzYe36Y2M/TtUK6jgbVHcxiFsm0bfNIyU5dEFn2Gz8SbfKJp1bZ8DLAewi5eC
4Bqs+DQjbObIEFTYJ1i/BCEhmU3qIS1WgSaK7rIRqqLOCswgPOT8B6NPDuJR/ouiaW4SgxkfEybB
SuULaTozpa7H6+KR2R1Z0Xz6nXY3BZsi2zFm99wdZh9mg5NpcaAA/xueexhZZ+QBbY+qaTFyc6V3
F4j4uIV8LOr8db+UR00g+/CtqbHG1r2DeiT6dxF68BO84bLMvw8+1K3KESjcyBDjvEMRdBHeOnVh
oRuGHw7fQbfS2Hf1nesWKfMpjzy3Je98YTZA25gE15rScO+WdBwu4srMvSulH/cr5g9zMNd9n0ET
SRA6WE1ruftNYLDtpkeFcYg4ydkrvCgyE4oka6Grzx6dk9limvIGaBubAZaBlmIKH/oIaIgMddFb
6763K8/4UkS7t+/nE1EdPuO4hWiYWq694RTMjT8dsweit858tuA1MGtstkBZYi8wCRifkLqOKts/
xTktZJe3FIHaze8W5w4umF6vTWwf9bNVND6GEq34d8PrQ05ju8SieptRrpbkDOxm20Y+TYz7xXaC
R9c5HX276ozIkA6NSPlIR2xIoaxItpB1WSKwBtMrPn30psIUi2IhmsXGG519bTPuUi8LvP4KlOAq
rSPTYoXIh6jmh/iMS5UzteQKPn7w2UdGQ9oRazfbB/EN5exHWZJfIo6hvXD4gyMeaNU0BH1WGri/
f6eG/uH++sf2ot70Ba7hAi0kFeGrFab/SMMGYySSchBkZe2NE4a3pY3OvNRjw75IU3DujzYLS0km
B1INu791Zhzib0RZmOM01VFXUnaPqBjHxQvCA1X60w6wWm6F7DRyNrSHyAc5Yd+PySXs5S4yeqJs
1WLNdcWSbJlVFH/NfzFNj6tLJQ5VUz9ogsgU7Eoyqk2LOTw9DyIxb4Vsmkk8vSzt5NLSWBhoXI74
u21rpxE9iCQicZgrTH0f1rFNB11ZTh2m/4U52ddr4gi5e/NkZRjtBDovv69E4HqiSGgsWuhTiuWM
PPNrWnn+FME20I2/WU52l4SkUaHVm4KUrJ5PHBRRxFknGwXhu9uXH4Sf3noIrrH1kaFDuCcvyv/E
6qhbGDaFumnxJpaBqDN4+Yv8wGb3nnYpH4Nzgs/IyHYta3JOcARYfDPE2kgNSiGxFDmstQPPtjGQ
etziCzVW2baSHmweAjRTF3VwFWBNHn6vg44EjgARfR+l/vJB0x9ID0KbVD8kMCBInBso6AIWK8Mb
xVMZDDG8kx2oSO83cy0OZfj6auVVg7jAIk6qUM0Sp6tkxq9ZRioiO1J7b5/WYgBvOjIOPSu9eu6Y
03/LHDIpwcNV477UrX2dQm1k5OPE7l/FoG/mkHGVRM2A7F5YWoeYxwDUDk8O69QZ6T+JE0m/WlvY
0gsbW2CvIT2RpGdd2c+4KRdj0yzXW5ZTJGGREUJMfzSKrTgzP6CuCTNi+G0KLNhJx+0mIS7cdO2y
DbfZMDocTJaHP8MzPLSyno+Rezj7LWJqLAouki358/UPhaPEAeDUYoFcxoCpzzmHR8RIEI4Csj6f
pI58wXmGto5xO3jZ+Sid04juZnyAehjsWJzaIWWqO/RaGI0y5e/J8rOqn7dS7dqPlouZLCh98bea
a3eswHAlDD4hSsT7kCGfFTmZopsHbm6IQHR6vcuSTByI6VzlyeGZgN6TWw3Rg7qYWx4Su/FOrkhm
2+itAPqhUyie1mccW3fZ5CPRX1TVEBlCzI+i9bDU1GL5rUIp8eeMcZ1tfrOP0Mht0Wq4qF7dveZT
rj1NKflbA4ULsh3DXQFjW3x1c2DQDWqQlrssozkQ9ug9MdUiaeqJdWfZ562Tk+DwHQIk6hpH1d1a
297w9Vt9LhldLsOJsobwaF/eMUuaCpMS3z5+Yw6MlGWEAzWiwc5KOWsOOSm4EF5YN/Ht0030eZoz
bWk5FBGBfTddccWOkiVc9619hSsEKUKjujbxKyt66LaoHygrayfLZ2dTpuGf3n2DjhLMyDAXRgNB
Jh7OZU4b/rPjlyOH6oDOTzqXPRnZfCU2FPFcK6Hpn6k495aGg6QJOXc8heNWRw4E8W9Rk5WcVs93
WpsY9d+OudKBP7GQJZ1BSMccJUbd0/MvEf2KxenUEmuGVPYby51Y557yV1Iy5pbBUtM6mxuJc+2r
a9E/PTqn9YrcjBpHpt48mOoCcNihEFfGZGVVSdelQWfJ1+ac1kM36oyZMjrFD6dUt279W9Q6Yy3R
f4lDuLNZBXnVDz5smsWDcrN60B0e0J1YrmFbJK8IecyP0PDcWVLhCmsmn38Z1pnzdP/fL/WYZGet
XW4spYCkwqrl5R21ZA89oU6+G/uRdXY6hjYAEfV+F+biYgQwIbqgw1YZwLK8h0LgKCOmSA1Cccy4
Q92dBNKbkqA1KJk/BNYwFfZfyBZG+1BtVGosEp6qVjRh3Ip+Zg4QkENc2xGvPRCQEML5WoBXk/2g
La15mOKuyAfos5R8Kl114ML0aUbMfC7dSgcfVxGZL+Eg8dxFSuQ4M2G6odX8VdT3g00obQ39hc97
ZV71SjFmNht2khxJ2GpoBOw0QJLrswRVd/hL4hDBJY5IAJCdYt5KcXoCvY32fWamK9mCfAtzTGIK
67r2SQKDdJrnSUVhVFyj2hfpD7MJALHY5FaXJDEV5gqWIKlboKFrVEolMTaNYVeujuZW7WfVf5He
UOMSDz+slEtGhPzEZBx2Q0etRaNJ5hBSGGQdgqfrlQ1Z23M+BXYNOxAcFD3S6zoWPQUmTAbheO6n
muxyOZRjCoXHjkyNso//c2qKdOObvpQVtC+zOPeylt/8U91UDMKOgnWdTE2Mu+U9CgOxOxJeLHib
NPkLZAgyC2v7RsX03OHpwTmXQcwMr7nNWI46l2dReHJdAUfeGtbP8jxLq9EC1V6IxpCmBHAIOYYQ
3p6+LlBEJavAOYR1NiGCiXXurGwpG0ism2+PGbHVc27evHAXUvFGZ0rPYYk/t9h9m5kYS6cqOzxy
qxrV9oONif4s863Lure3FtQoLy7NTHrlHCTxb8mcaZZZEw2+gpzvZ72hxQQpw4B/52xwMY9J6y+O
QTBSKP3RmV7fJfkZaTUMjK3z0NMBPelRZBuHbRBhvM0QosGyXCv9IkEFLAcDB9jnsOTlLGoue/fZ
GvKoQREQ+LzxwqKdZZxyhXHzrvB7fTFmb1Ex3GW6+lLU5s6Tv0NpqKVirYeLXjQZxmHM8P7+R0/F
fYpXx+bQ6JjeBLynGodIjBIjfSob9bDQxdIzawbtCI71FozgolQAnloaMMS9WS452SMVpy8qaeLw
/RtHV3cMsxzK3p5t5Kl/ZNFopE9fPK6hpvVHfycyfgSKgmp/WvMElBCLeR6GWBkxgPvqXOe1K4sb
+xTsRK5iyZ/8q9vRKtEe5Vch1mz4WawNWFlaTBDevC/un04SdzzArEAPiYrawN22oN7ukMgqIMEf
xDEuo41SdvuIoQg70WEZjJW9XZTTalnYvwJ+alvLjkWCGSs0u9wLU7OlGdbp3TnppZWIKxODxq5o
NV7nxV3zBXMaGuq3FNwZ3cdVsk0H2Md6RHkYiqOChOc/hLv+mFSAUZtGmTIdP9urveSImB8hP6y8
daQiwBqQ/fDpOMsw3HwYlHMqmz1R/A0ypZsRM1CcYA3e5740YfpGxa5RqUw92zOAOuOCvbiIUrq4
fnqxqwD1KPI2ksMZHAELQ6/wrhKrlHt4m/eGrIA6La4IkpJVtq7daSFna8xcxceC0laz4ZoDZjJ+
aP1c1wsZeHZAkqZ4X7x8gdAdVktM+YXm12qxMRKiIIfUu/FRr4SIR/v3lKlrPBpx9ZrJ0W4Mir93
zEIgs5F5gpt1mntXTcIpZdrN3prSmLyjUlVWTmjrdJmuUcGOPJ4SrCbtna+hO7htVRExV/LAPIiR
4A0rnJRcWx1yvK9hqm7RdaY4wADR1yc9rOOIVEXBBHj3gjZTpnowH7cLryyfZH760bDsCN+YXGXx
w05dX2tSCHetqEGHqwZ5h4fBucPu49YxxSFC2ePIyIHxPwQDPknTaAxKaCU+CDp1Qwvtmliv2Ar/
V1eP5vkrAUfePFTOIwNqUOFXq8c+6Q3ZHhWeKHwWnsX4qt3MTBrIpQ5uCXcbF1OgMzwnIGVSZ6mg
kziD04e9CW4YoLWVQ2M6Hjn9BQFiihT2ETR3ZOcVcYtuOFgmqUDhWPjSgSxFTKmbrFaZ+pUZEEsd
uZljUsdDN4NitIdSYV/atuIX7fs/NcVaJmq00sd7DnAiaudN46IW4sAJN+nkXTMIn4gJzngq+eGy
l9h5CZ0fWfgBUk6W3MxMKBRvr9LepXhkKMcc9tYCX4qu+BceofrihtaGpxuB0yKpvaO34/0vSn0+
jb5QkeCtw7+iQw08ucZyEJzj0VhipLJjleIuYVy1SVkNDMyVm7OhEjMUJQ7xiUW6c1ojNGHO+s8S
TlN6qZJoXBTYJcuNbTCMx4nnA/JumOuidxpPrfaiSvkHPdArr8wHHi5OlkhGVVQ85ZZGhIMrGrvF
qOtVsYZETnAWJ2t+M85aUFWoqpfZg6KLjks09M71oX5WJ6TEe/Hw8vDB4TqSJufwdrHSm0d681LC
cljA3i2aONkqafbUD9Dr99rC9Fmfy8bvPUUehLbukJbZZX7k+JemAvZVfH/evEbiG39DlqptLkxr
sqAQR/w/FdD2H5Eklj5fMcRWiftQtDT9uGoFkvx0XSiF6ddvFfFVl4fjZqBLYPJUGXb5ZRykoOyx
bnDU+zUVRCmaHnDFEGYLisR7CBysUOIp44GOt0EG/Ss51xVtioqQqH6DEzADfzuAwRVMoZH9sWyl
BRlrVH4phcmyly3UY0Bq3vn4AfDMufSJboasCa4+33dxRIc+cUvW8U4u2li4W1TKrCjcYpKqaVdE
KVx22ycu9J59ANjo9NrWGD6Fal2zcZgq5sln0EGj020kz3QeL5prchL0z8AkWKZXxdoMBH10aY9X
1C2nFhTK0We/KHAYfaeK4Ry6XXo+BuSRee0xzZKNofJgxKDGfwTNNU2sa/fQTweeBTSVLJ5Nj4H8
mNm60e1IgC0B9nnCBuKLFhh3CbEC2IbXqreTeqGEUDMZDyzc4dVJVnhzHM/ZU/1vUVkr4EI9mDOT
UEsTybPMmJAxShk2RMklLvVI99GBOh6HKHZ45xuYhSpnYp9VqCNRhZHEI25daLMJGi0IRsCiQXyg
9RI+sGHIAZT0Z/ifE+5SPLykOh5cKLZkaOBcZ7ikXC+1/Eo1riTvpO86Ut2ELirMbGktLG/aOu+h
kqI+y0OXGVZxaaJmHunv0gcO8d2ByH9sj/HJor/ecgdPyCkPHjBgGOv687tJfjMnxeb5+ZgT8mhD
m8zwM64MTbrcoJeOxF4w1NVd8J9Qgawp4NufAiEw0e0oYoVg+hLAdkGdWfwW7yi8xH5ltdfihQDl
nKiHEiap1vo7WS3OWAzKRqW8gqMN6fkZ2xYKv0BEsmbRWRWn90xe2nZLRPNP1A7xO/25lJ1pV1Ab
stoeDHSQnNONV7d4QIek2qa9khadmI9Whd4Sgub+8Z8o1y8JI8t2Eg7yJ8FTnpeum/93VymL2kRI
Cv8MQTVPf59J/sPPaYQqqfS509OruL5VqTDjfZ2ItuOisKpo2HQq5OUL2fLFyHiN3yhVGZS5l9ie
RX0Bx0efH0j5sFVv0lweaXhNu8IWO41ZYSp6j5IoJ+3ikFGfhSAIBid6OQZoNOuQOWXjMMgfFYVk
R7BhxhqhPvihlJXnRpAgGRMX4lxNpjQxoAVI/K+SHqXVhoDydGrXbsbwLiD9xhi7mO7zt4GJmNne
yUTzzRcha3DS1EKAt9mR4xbg/FE8pRBIpB0hsBo4aAGx8igDw9cZcla6Q3lnoDLVv8i5ZqnwnGc/
VPkGY7ZTmYX4zOp6AlxVOsHW0m1EIfSDyguvBXaPUJvOWZc/XP2ZkUgo4ZCqhzeOc0MyrlMnagIp
yjzZngjrz1Ai2WzuVs7DOoo8XepuyHDB3nm64YCjZh0qmuQ1wjZy5eo+VjoByr2DIG965Ktisn4i
xh5YO2Ve2+dJQBQ2p9cLV3Fq0lTsrzyP3cNs42MAF6nXOBIZs2UqAm90Z/8AZ3YD/qwb+NTv0Myi
U/byw6QmH4Rty1uO/I9fkt5BZZyQotb5w9PLGymF3jAEcisYFrraAfd+kAlJ3aL1QiKVcQRp14GC
0FMtzkdpgHaKEAZrZQ7MCSkl310bUcyc6etoq5e+9+5Oc190AmmHv//W4d9yJOeRVK27uqJxiQ/n
X3CMVNASL9cSrzEFoR9BEd//zStf/DB7Sikjyb0z+uEYOJqPw0pW/BLy3ICd655Qwq9IIQwT+MNL
vwZ1b3Pyln9ydIRIeR5kaVkew1FxcoQ21Hc2CHNdc4tUwTyoPl+EzL5JTG/4S3LTv+hgYoFNNgy1
60gs+B/MMoCsLC0K8tNphcLck52n2SDT85IB0cOmeMqyvmqhQciVgII5R0EMIwotz2T1dX4z0Aby
OxSDEsjv4YlmAXpg312AEc0IXEfDmSBX/CHv8anUSCnAFBxgUN6mtfzBH+eqX0rTFZgEIsixO8bS
yt1Vc9IfCt+keywxelB4L5SUOYTi/xO5W1f13UJATh5I0Hfr90lbfYdVrMqJG7VUdbE6GvK2PePS
7IqWepbdXfFs8KSXeCcN7oK+Ss/fEGAEBxLluL4z6Ajsv3OB9Fw/z++QrUBWvffcW+6TFFpH3XvR
gSR/rXg5OK5AKbF2O4B6R7Xohs4OOBMYcswKF1xPiy8pqTv+axoTe6qBEdwY13HmAc21pTIRf9tv
/0KdkP1B/dB4lUc1Gb3evu+uMMPpdZHdfdj9+HgG5DRWUDZyUkAEm6Re3yRTitZ3yLXXujXGfwDi
ndmuKSQFk2WqAgQNokSgX1sRiUINx5fPrRnMVg/FdwDrpDdCI8fra+S9h7sAfad57PpSPT9egyYg
ymEtjsqx1vD3o9qeucC9M51eUalhzgp3+O1W6T3MGdJTjJxKw05FEurCvf3RdNmEoWzFH3xmtfkR
CQEWDKB/YlF2qF4fW48Ap1S5XZEutTTPXSzxIRMNlBciCx7VSiitx5oEJmWE+MOaelvt5I0n/efv
p3YMJViKr0AwoH95J1KT1HcuwMpvk9d9B5ExF/DmzQgPSJ+bL1cIkuHLgAfB9M4Ifabe9WRBg3Uw
gNIv6RDTkGlwtqGDaFTS0R/ysWi4JC9OMqs4mW8mAchADR/mTuwt4D3g/SAnrmzaD4NZ70q2JpKd
lAIt1F8gC+5tzIcxL3QVEJ8ZQ3kHa4nZ2HMylRDWmOGp0MQkyF2lC/yUQ0IjIREdxGKyxVmnSBok
2cH9fuh0jTeQwCteL91iyqSKlE+Dxx4QdFcPI26XylrffaD+sV1pKJA4e3REZf01+nUcE7Kkx+zg
7+Pdx4oJZkCv68lrUch78EklB+OjDE0J10mKpjuPDdBlc19sjXlLTA59S2kUz24fQjk2LsrbllD0
ir6R2BTqrsmVXceprDFBGbiSATKizBlH4Ur44tLnIxOD23scnJLsm0DspyQCRsTi7cr3DQGJif/i
fLmB7ufx9nrw4OMrpWEroGKJT38hymyjWLwoicrM7uq6ZCU+DCjWQWCzdIbcwLCgcJdBJMsMpEGI
bCTrj2gvYOQyvOkaMFaOeBP9aChg2cF3FeqdJxYIsJVbVrzt5znL6alTlBokTbyXoe/MHVSx6Kis
rIZVqUQDabBsKySc9Ttlvydsx5YeIidwNKqZtl7nHHcf26MholqVTd86mMpSz6R4wQCVJPy6rXLa
sD+3XiSldOu0IaOOc77BRZjqpcf32qc7h5y2xz7Tde1TaYN4e6FRYC9hNZ0vbTEIpBp3NI1vMOw7
xQh9slfKecHJtonqxOokBEMicM04uvnO1uahyQOEUgVCLSDxSEDszEMBh7fHwZtiIE5VzN9VLbXH
L5MvJGRrpqe+u5Hm7V8m0QbraAtoBHqGktAc29kvSseRdP05LOvkVLah1AduVDHFnyhZkjicDZcV
o/f4NgUVSLnBWjWe33tNVbR19lKRp69S/qFM3kS8aBEGIdl8xgFHdXya5UdamnmbK/+M1p2FQJ5e
GKlDdlnL1C9loqKTlL5VcLORNiFKjcA4CzTJhq6AFQ+Qo9KzAPnaKlsAi9LCRA4MAcEqBq8Be5KS
2nGpODmo0I2iTZzKkxdqwcIo1QfhYbLqOLulqtehPZvk445y15RQkwinrifzwFEKO5kEo/PsPBMU
B3xkuWijvOst3WUrjHf5JBQIRFTJ1OaIxGOelN8V8StIsZHNhHl1bNZSmCM6jvnex9pMzXA8zIkP
Arbzn8mfO0L40uqhACeRF4uc/gSUEKYc6OnxBuejnepC5Qc+blbOzIaPhCaX79CjhHu2TBj8C2UO
d/kurwi3HrLjcJTQn+FZZR4qfAVIdPsfXWhSh/XkkoyBbBqMc6wQeeNqPlTUSuwRs758waSLq9Hw
bcjvdWrbMmsSW2xvF9u3Ql+4vp2p/MjZALFDdeqduF1d2hhOyLMMLJahNG/dfhpzN2GpPYieXWWU
cmM2WebQdzZMHkmLMBThZhoN8Rx5wXoOipcBB7VhrK3E/CdiXtpfZ6HY/osDQYVz0/Y93hrcX3YU
l6R0PZoYfWwbBHdYPhTZg7+KeBVn7MRZmwROby9o76fIVO6tueuzW4kT8WfLahUkKpZ3ctswLQJM
1uYKg9fxTLiGnrSS4MhW+ds39d9mm1YLyoKBIlJ1IxjicWUmrnil1mnSrP9M2nAiCoAjQInQ+8jH
5iTj+T8XV+nRVkNn0lRDij2UBXzH4nd+4mbBrGbQqdEX6Be65yjWgnBt4Er3vP6KGlkwr1pH+Inu
KF4fcuTeozj3YCxU5ytm2FNw2SCLCHWygyo4GjL8lS8H5LtlWBf3yyCLdYugEcJdWL++WjDJVp0v
lXhP3juLU+9Z5/2oOPgA9ik70f3mHyoYONT4VKVHuDTVSnwYEBkRterotFLevhhn0SfoEs8sviA/
MnLSZm024Ma0gqcN2RlgTpK/yWAKg+K2DmBhxBPc9QZ5kAowGHrCEkjAK5baw//3mrd86Pkg1/b1
yVYUGC9ZFsISj1ddTSKJZn0mkgNpuSifupSCh8L5IZn5vetuYIlN0jdArM6V5A/DvRTnhKWqC1wU
YH5BegeiMkNXFEDDzVvj0LHKhXXVlW2Mc2MZ2idKE4OjSvNmYLg7DV4QjpWj0oQ4a6oWSBloZmOD
iLZme5kGUYZHw6K8ij96nayDLp3LsVc+aL8mTGfWG6XuUVYnSvRhs0oFK1HFS5Sh+fE5Lx0gja7o
bqZMTkoRJqKswqqN++NLIyB1pn2YR5VsPoWXotdeFAzHUk6blymdZds3xWQBCXc7E3Y3cuDIMevE
3h0HwNG/ez8S1toQEALxTiehQwvOxuwd4fqr3cNmqE0ANFg2tr8EhtOVT3IEYKxCogXvn6qbta3m
QcTXux7QMN2DGFmPvFZriI96CHuPIZeSxpQmA2NKZOUjsVyhOdD2rJJYo0mg7J/UxcVEzkRpK13t
FRkICzDnuOEh3hvui/WdFAu274q/roRKZat+tZ0osNsYFmQlORULoau+aQikoVZdA8WwpG97EbFn
w1vNiGAP2dJyX9qGKrKQuJxpnnaLDCCLfEwmtYiN6+a2WJwIEnp9btjExaFAcNb0GHbTZiicr6b3
VxeNOrDbY9e/auZWGFUyV20eOuEFkTxkcqIcv8jF8mm+oXTyLRWxqCj/v3xQnb/JYBdJQDXrCErk
vqHyhaiqBhFRQ8TC911woiO4YalO6hfXtCcFl27qKoWv648jvjfopD+IHBT8mRpq+gNhPmFWulPN
fNvRhmBd9jNbsrXI7xeUVc3RWelHD4BGMrMBeGGTMBt+oeGZE2RV+EaNYgskHivbDSvk2DStaf+w
n1jnIVyRwXViqrqz0WFqySuYHryCk4LjutncPR9B7VOrYGppzLNfZrmFHEqKtKQVV2pAdnh5PrAr
9/oyn0L0HpGBZfIV8hZYs7sMkBU2V7Cfr3Y3rBOvhgMinUVGoC3L/ElgMvhv/50u15J+ybhIbNCK
hvcudqjtv4NlqYKFrQ+cm++XT95/v35naooXYbqe/WosUeZSSYFeAffhdJthg5iLJqb33zWJ/dS/
RcYvPNKrVrK6+9w1U7DI0kV4h2VeZOWX+yWaJLg1RELdJRxLHoZqhEKxtZqQM6FnaEvw+dqNsw//
qqFB3kYUt2eulhhrAOIMtnRR7ZFPOtMtaU1YTFqhVIAjgxdtyIbZSG+emGIfV2NWHBqX/Hyhh+Ct
tJK6H9cYxvFbV16DMC9x+YgvhhHNVc9Rs0nETz1lhJ0j1czENqoTyvRyM/peHsin9AF7CKiB2P6s
uqFrpBdag0IfJytQLl7vmSyqmuMLe7eIgl11xPFUhCIYhFN4sF6o+VNuB7rJ+DFWePeeZvHH96ss
Ev5fs3jEetMwyd39Cgz3nU5R3r6LzYfvktndGDFBuTqakQyt5OtTABTWsRIQq3abFNL2ckIrveKz
KlOW0pI233b+62IYs18AaRTjtPgId1xjP+CCxl++SBBZOhUKqJlrj7FHBvka7/giHmpQhAWNKETP
nH9lwEd+nFCq7hl02Xcs+jBstznIdoIRk+gvynrZpRTaVhY8YRl4F9PqKfjgC7+awjxO1ooy5NO1
e6XQX8zbJgxMU/U96qY8VvJ4w+iIirmvscSTQ0qyS6fxHZv3xdGGlHumdXEeDkZlTujeiM4Wi+tE
cUtTpEmYDCSGPve4hVoqNODVehNvj5ZfxbOlX5QxR19oinLEcS6M4/E5JIHwAugVyeRHWqLl70AR
MiPnJpYCHeXZAYzsjxLUAth6wimHQwpQ1Qf1rSFhoFrtN/CEiplmVTe1qM+JqV9Mw+3bmnWoi43B
G6YrZuKP1rh2d37GEwiAwk5XKpLpEsiZDqdgpRUX8o6+zEgezte3JamX7SH0/o60zP4pSHj/JGm8
UHzObya3z3cMzxjrxGh8l36qO5yOBpdap7SthYLFxW/8KxIbttQ/klKTD2lerm4obBExGBUnA/KB
FKHiitQ6PpoEpvax5iF9OzU28YqAsTCFWENhU2Rk/WVDTiW0e4Ow8LE2BaqTnql+eiAGIdnIZOSH
oPmQOY+haKP8aEu1EEhc1Ik/mEscE/cNDgebHXfn4OcTCcx0eCruAUhxPSH5RyqtJwFjqL9tnTQ2
/2Nt7DeW9vFR5sgsKP4tnodkNY/mAUedaHd4n8v4YN1ZWrrB1pWAPdmnAMSTWkPYVBm7rrQ81bba
E0l22/CxkdBM970hoRsKu8seZhqNuvTRLGIFtdSeOrkgkCCkwFEZcRd2xC3RP3/o3njK1G/8E94H
Hfk6wKfg3mW/Deg3VyDmfyAS4QxkcjkZ5cWzoy2yzfyKaffH8CjGaG/N3nXnE2RoWdFBMa60RYV9
Kr0TmFgrvWrbmy3mGaGzEgUW7iv3Hy96tWRHDJO3k1vE5AfuquajOeaT32ISnHiDEu4n5YM2Q6Fg
WeXdADd5GmvuvidC6SIMEENrGEA/nrVob3kcQpz68h6D5cAV8ByRMoZQfvKv4GECZTvd+WWQDkOW
oNjWcT4E5LBt2O4hmoJUzF26olXTjh+BemXozZwa0dwAjaksXhJfCD4jjWUuVQ5jX5UCVCHhLDSd
LukMoRd5wN2a4+vN5YHpmoPx/6aJKDrpjbuJIOPJp9ak2Qg6FBr15lXcG/qwANWPYWRRbBRtGRIw
IpKECPKoO1knw99/VGYJwurvs7iMJn1Vxo4685Aj7Y5/EqN/GpOfx/XK0ZEpDHPts2aspfOMPRUZ
vUxPb1yqruUzswoNeIkMxxg4+m3w/Mv8R3lPXTGhO1/qC1Tncsc6XMwDgEENDpk66RWGz8eqgN/D
rfr7OewjOukXQJCzJHCcRH5xaZiiXF0EpXWNavWafT7CrNhcz3tOIfUFHinzrqWS9bdB/HcLIERZ
hfV3iC50so3ZdCS4xNOevl7NGVCixwoyjIT8lsl97kokDbnvgWTjHv9nyhNVUJzm5oy00xlw6TVY
cuMTqbEDHvoHmrKTlsOGvF8foYhk4+JjVww5kM5z277LaYGnLR/+ivKD4dxaDfslCtw5Kvg4M5u+
0fP3tXZ1ydjobbVVzX8SU9JXnSIKPpbSxKrZBYlB0jb6VU6mp/bcF4cXernwI3aiWk7xfBLZ/DoW
ArrGJLiSz5GRr+YwS72361uNZofVkM6UtejxJBAPvkobKxD4tXMQH44aEKTav//JYH53yYulLaB0
qbHo5X7F2JMmgjO1Equgdr5wA0ir9WlUANDpYXONHRmIL0oOBydns4V4MeGLrLPKjjZS0mNWsfSi
3SHf2Mz7VCXtbqB33A0Rf0maKSXtzqy2lxmlGsYzTRVKkjEUFB5orXsxMpCJpu2e994/4QUNKhDD
9jYsnTo7VP2yViVWLGQ//9+GRanILLQscl28OCf+F/PY8/TzGS1D2/NjnacCIm6OBkIJn5qwYpQ/
k+v//PYC+mfYIIE1EcfV4lRHXEkPlvEFtvFGU0snwTwGrzEzzm7dJcPVYveKDJq+KeWP/F3RUTrN
YyGpdRZjwGYHws31iPNrzQDpDSl+STIxLNCuOZy8DOWBpckMB7pa5jLy4yd+tiHuOJI8l3SNDr7q
6jL0rBJAhP20PN3KhGBp8XgPjiQ1GBPi+kZXOk7MRWQdBmEV9Dlr4g59vHT1V4tgyIOP8Qjd2Ylm
w5esl2HLEap2fFkCwpDpsuj2RiRktBgQR8mQAQh/0w1HWhSutu8uFdJpLf68PpS1tEX+GgbwVlZS
GvOXaqa4RiShSonKFYjNTjWJhPHGb+4puNT4cuhKKGRfUXVxPsX+z1m1Ba82hDQXX4+NCuPG/p4G
Ii9AlUYHvusMnmbWiHhIkNRREeoKxi1Rzzf7j4QVSrSoF2kWqIk1lndI2PcdjzxdiIADVB4eCTfA
2Yp31IqPFHAr3EzuDRs5ZiFVof4mtcwuuY6VdkHK7WsKlS9fK0cher60IqPjU8rxqv+TDPFoGT8Q
pYrydIjMTPiRiSd4t4mjaETcxzVeZtTlzV3D4bAFM+Pt9bg+lywIumTO99zRu4yS1ygaHjngOjdq
vLKyfJwR3LiJOwvIJYX55pcUD/MEVB8Un7zW2UCSPJSAh6sOsvnNFkkua8aaiy+41KWdgvHNH++N
NPLNbi0MBEpKFOwBnsZW2sk4Fcc/9cygajEg5cM7qZTLSuHKtGcXaTG0Y47RepqPm13/ACgea7Im
Michoq/rASuZuW/hRfs7ammCRBwZdzkelfwXRAqCQ8nWj5Z6gEg7viRDCb+5OvAF4IUA9sxD/AKy
V+DMGC76QWdGpC6ibGcuCLWH4nEWSYio8NPd36gyfcFq7TB8nBwm5WT7IaxzxmsiPN88BvBy9GGU
SzYlGtKmIc/59XTd/qaJ/YrsyqCfLSqUUveQNBbwUPhs63lw2UZZXDjLF5iJxCrC3L/euQLkjWMZ
OTihOKM2ydsgrINnNjhPTySyMy/jhY/XahWbJZwCd7JvxifFiU6yXRy9ZfT8cvyEEgmLA5Kv89KX
LA69HFPX3rMSn2K+q/cC8ww23EuikMm7CH2g2BfcBpkqJh+qkXlliuO/f1UJhQNDCZfOCed7Y1IU
ourSzVIjipjOGeko4+d8DfvdGvT3i/Hbw/ma9br5LqEdG6QJAqNLp6mzuavJ4QXboqglJzyPAhhK
iyTdsFfLi7DJmmD5imMXcPiYAmao2zw25DptKRRCYGJRPkS5luKpuKA4KQWy5mnmsLEApFqGSZRj
TnXGcFoC+H0s3CG5VPJCbirgw9Wb5HtJDs7efNtDt8tfPkpB2BVmvQiw8FWics3Nq6fCBHzhw+1P
YzDsDh3omQwTo+V9c4jVyiypKrJNHsJm0i9YUQsmlUO8HkMdCZDkH6jtj/YtWEP6QZkBJaVkyZMd
NgBoDPuxKrSOyWsQShRGAPWpM4uW5vn6WOEs5eyw1glXrTx5GlLK4pCFha4AOdPIOWcTEUoI5lxx
J0lNdNfxMxPkZBZmpZR+4zxxTBANYdlAF+X+pht+W0GucmylP1g4A43KNKZk7MG+y331eanQCNSp
+iVuDEX6AlqsHsgYxtrX8qGpJv0nXq6ejKk+enpxzGl60OZ13PEkwgtHi3UQ5VIPFUrQmpHPUSCD
MJW0ARcD5P8sPfJ98p+xYpqNfMbO6ld0v6OpnwIGYoCB2a3wjJxz0h9ppXg0JgVAsGd+RRuNlVI1
j7h/hR3WmAUZX/pOAd/bzdhRYM1Qw09dxNMT0aKLv1X4OBiHfBSy89dPyPDJEnKTYlKxh2Pp3qCX
f4shL6Z2aPSKcU+DolPPuZk7thO808879XerVecasf7cCZxgUp2tRLZ6+3hI8UyUMGanNaX/mrWH
8OUnUn94km9iLjPoXTrWlzPPN4faDkxCMdLf6H9mNn5M+EIKqijTzkOh6NNrLn3AdFpvG21H43rj
NupzpdPbvsVhoGQbnzV4sD+xD0OWUwiV9CwE9DXlkgOZYCVl3mSonwbfHF0WbQBshOWZcYPbBgX6
Q2FNl/BfXW1C+NqblvuPdULFzNMuVRTP4+WrF5m3SHIOJ3JEUg73NMGziVp3PkeNpLQuzRbicYc2
ZHMDp1oSoNQTzB0gcZI+YAlcUdNCLEy8zUJr6YrGamQbmejLtjQPNeQ6HNw7RyAboxisUoY+uqGr
QqK6owOKtaX/5E22tv5mfKuJfIk7mqEUMA6ANGxxJoGPahGxMK1x7cJHo4sFr8dn1F/OsBBc+Wcj
FNa7WYWa3braHttQ3syoXx0nz9eupjcPhkpVgUwrju03cNly11dhCbccsAymAKK5guDWKohHNp6k
TUHiDaTRCnYrOGwsGu5qlnTqSoN7FVXBvcopD2UBaBLhfzyeSpB0Ecz/XGK19KjC4M/SrUjYdagK
Mi67nORvzTXMMlD0q+UCLi/hUi44Vu0kNJh7iFF6b47yIipK+Cw14Zv05XUv1Alr9MRS7VZg1a6d
Bfg07W3U7dpIcVhpvbIpuTH2hdyf5mu0Ajt4hudQFGVDQ9DIAjGbkbb/6S3flvifqYRqrWvrnHRP
nthNJIYm7eCmZwC8JNXW9/DGOm+V3n+39AsUnMcXFmR7X0MDZyPu9a7wSnDOQR86nLv/y/rKo8OO
RG34LU6JBMLqFfddh3hKE1DhWHCzKaqbhB5vfjX2MKgsNkAprpWEXCdTINc6DcLfWp2DkeCrWl0P
UIuA8Kt+g1b8rU/nsJnSYmZ1MHdQkYIRxvH490rdSCFq7cfS4kYoRvZa7lLNmfVSc9bKfliYPwsP
orVbG6PL2KPLczy93CJy9nyj3UxUzho49OUoKqeKrtpU0kZj5bh9vb6l5CUh0vkWtMPgM5LxrpfU
E4LJURC46AJiOBy9r1sZlkwh1gbp4zYVsJBUSIg7Oz6NzziTkO1pWX/uYI9IF/H4YUzVQXbtOX+M
CiyxBv7xg2ZRPbLFiwRrPk0KqHCCXeKayVv5EY1CC69DgR/m0QpB6hV3UoPQEnB4LMiiSPeKX/VO
Ft61fRMbFEKJj1E7tGJxyhNnnQHjfvXETTAvxUEcX4MjkoDlyjABUixfWksEwPK6uM1D4aaQCSn6
VEEFJJ7/vyOmJZqyDx7DSk5lKfVb+m6bKopqfONQmuRGgY/D2A2qDU7yyI1aQwDnBXqzzQJKPoxu
boO5X9o60mQ4/D/RH4IWZ48t4v92XfVWf9oY20AYKuEhVvILuNfmpPyihJsLfgn1lEtayzWppx8q
a4GGJI0zJbQdaiKq2LSNzgoFFar/2zUhYE1zVkYUMJ4LNkW8sLAhIpBTr7N1Tn8/zkLMb22OMByT
8V1iM0sXUo7fXHqDrc345/gKhwi6aDmyYZzTbQRc6EcMes0eoDCKofW6SPzKZuSRjWJj1i7Xe6+6
riy1scXoMBpxKUhQRmQ7n1sSvUM0+qf16bUHv66IOA53nGrad0NY5h3ZkRMJKiJyVYOr23Gd2aFi
M/NdGCBKu/UIrj9CX2i38zYp6TCMtgavz91uP+BtfCc+45GWqj2lOLFlS4QGW7aNz8f3ytRgHIN8
paI4Ta4DKxF8vyz/OmnYUrn8IqLAOwcxqDmtEvqS70f/kd6rqOhuvMmdo0OEhXXo5dpVTjLkKX84
MP66z3SyJLccs8B1nbo3aV91J+gik5/FkeQkU3D+2OruDsP/gcvBnqqOpHnW2xFvjJJfdpwImAQ9
bbNtir9F37V31F1ezdaHoxgMhGH9WWAPqSN+bx3ncXaTLVYTBdsd6R+T3c59Pum4zvm1GKrNPpUF
cMH9Fkf33jVweFCeFfnSRaO7TOGQT5iibveBv7WakxJOyYAvLAyB/P3Vglir1WyvEuQCkQiT/AyP
38qhXXp1F7JrfnAlV9eSj38T4sYP04h3OmJab59HoBfBwlY6D43QChPcNJzpms6Q2kGrCH2KuoLs
xrG8rMBmONcMuhuykDrz4EforYpkvXojK2Ak2raYAzZ1kH/pq826Xq+7IHq8q/+FRYlD1t78Sxbl
foOMDUeUw7qaxlZ5IR+WZ5OXHVVK/GNpBAFNEk15zbNG15dnQ6PUuUZCUoMvWHS51l4gCEJsnyfy
5QENE6oZDy9T9N/GIi8Gf/c8mNM+EZfxhG0Hp1ehbJ+/Q9SVNmyILe1Yg8ApCmQE/FF6ilnpYkh6
CKbO7a2KpmDCIihinSll+R1vTg7DLx/81WfpN7y4hvVftJtELIzHvY1FJtdVk/n4q1IILMhN1ymH
cT7fr3ZG6DEmQAoY1kndD4XKnk99pmq5k+KFEwbCshK07REweiUl6dcjJNkQsrpti8MTjGbJlL9R
f6GrWIh7qkqFhk6MWFTEZ5H+Yg9yTLEGz8TzUeY6CivgHc1HnxQIKtyAvu7xnP236C9dHE23YhVY
eNYtAeJ2F2i4ass95ihLCmUI1GdA5oEMuoybqKorjp84ZF2/2Ey+dzMQIDxOoLAmvjB85MOzvYUK
D6GSf1RQ8CKvFqNm70M39Ju91SGSDq22vMq8yQ73TBLCRK/r+jtzZcNlHK5Gb7tO/Sg1NkT8Lc7j
bJTugMKXy/jMLHo9utC/PJzSOeLBnYEe3s7UScZWPN+oLENbDXde190G0vGPsDJJOAq2NmOPZ9Qk
egUN487esS69VuWrnOI3DqGp3HXU+ybnqt5Sg3lbEDpkKpWOf29zT3QzlfeyUs3A7rpBvCuC6Gnl
labVM8zx/KeCKtGpED5Uu9FK3UnuiUzXTdYMZrTZOvGJKvHK8+IiEDVzIPyfM4Shu+yK6UHdaYsL
uAFKREpxEwebmwJR85M/4LNlOY/bGhxgHkS/uz9ZGvuOPkaRiwVc0LHYA8/OSMLGQsQbbEH/Atzo
TnBaHu978Q2i0LZuA+ZHduxdmQPyFy/RmyZYeHy04cirMbK7qNdbj69vBjNPuuMzoGjydcIUAMov
l1DsXYLsISDnw/pmrO3/2341qD0VklttDxVBCLPXcEkZYcIZLUbjR531TmR3fZZ3T427NWS91np8
/StMbJP1C5QO0zUnI72Whct4u64dz+jrki9hsNwGq7jYJd1GgINsnIcfBHz3jqkJFsR4CCWIatMl
ZfqQJy9VNGcH+RS48/axOrmClnpcf1O8Fd3JqasFR1zjU2atTZMTo49rBEeWs3tWuXhhXowqQoHT
Gw6OyA+Cz34vIz6CtNEnGkXPWPJYiBc2Qk8JcsdcDzQCaP9qm3vj75Tg8Y5cTcOIbs75lq4VnyeA
hjyA1AU1iZ4sS+Wxk2LNtErTAVzGsqNsKmCRQ5Tyc3K4JWvTRP0ZeOa0OfAbdMy7A3R5BBKx/40o
XFd7+sQ0QW9oCXSy6SWBiupwEuCd39yEhB+hJ0RYU/d82lpp1zwS7FLh9Svtqr8HgH7d+3o9FXoX
+7yYZmpTtor/khi5SWvvIAmbCTcHTkX2OYIn3EUcGas+LWiPvbacDtOfF7treFtiUlNYp+1Rt7ks
/t3cXBgrQ6EfOmE2lo9rmv4Af8ApOiQJivHE1umZmuIqbXSQtRM06PRoQM0DwJPcGXT/iwalvqDs
AaRxG8LWAKUbrq2s8s1HGB6pSS9UGJxI2bx+wqj3YXf73QMKJ2ApcS2Q+kppJ/oyoAlP5CuMMnXe
r2w3F+UfrcIHkuflSj/5vg2f60C9zmrNyc4OvW8VrM6WQtmQQGNDnG7bOq3AYl3PNna02nTLAeZg
95NyNn8AzRgL86d5PGO0XvYdKb3zJ5WGBAzAfukeIPoiBE9lNWbENYGFqcm1jUQtrTVI5v93vdDy
XCNbwcTGvF/R4xzAEsN4CZ6TR7Amxu0dezhyjIJ9r1kIbpo0XHdyGf0VvTL3lNKJAbqLBq3rMdFV
2avTKi3aBIWddiLA+LXgaupSFQkvSU/oVdS2lFsanb1rJZNmDptGj4h+Wqu9EzkDF62SRlLfja96
9D1Q96Tx0vT8z9PEjm9axF1SH5KIdJdKe+AowvuIoMRO5IMxHLfnm1yygPldGkqX4jqzmDtUed+X
qemYrAjdTJG0xxEJ9TGigo6r/FAaNMRJP9PFU0lGPR6ET01y1Z2DyaLkxGP4K7CXX37jXGGNw6DD
3UnKLqVC56o3ZrZXng+FcCmWeenZGKyn1JS12gHIAJBkceza+IU+LtVLHhvxVSuGDDtyKsCACxoU
3i9IHZ4GGBtXs/5tYFxj36i9qOe+kxHhCqtOrDYTESh8bN0MbU5D6vs4g9ioAFWAPYC2+KFZ5THD
UDnF/fOvFwutkr88IAVQsrELXA2VjtSRfKfHmL6qjgueLsxsldp6aiL+kgNKW2qOP4PIHHRRPiuS
L7Hc1DHqiEhnKz7LlxhagmgfjishtC/EKmD46nq7raBRyPT5JMUsLipVgjrVGLrvadBucsNvenTJ
fbojDumieYYVIt01PZc72xhlUdlOseZuemiEqyFoEqZKZ0JFPQ+RjeNEXSwa7pTGBR7lbUHrV+EM
+WFrVV75CrkIybEGUy7Z+LJeE/rz8MYh82rexPYqlDaP6MSF8TLKrkGRxQqR9HAOGfarjDpLm7Vj
ziPt0xwS3pSzUHzC62l262FN6N+cDfzUhrvNKMftzPUHR4i+cRAN3I5An9rW1L60qXcUwiwTwkJi
LDYv95RnAXLywNfhjhAcRshKpYS0WVFVZ3b7o6l4mq63zXBKqjkRJQfV09aLegp+JPtTRVJOPrZj
vndcfDdMLwY4qiyQi9IMg9QpKPRVKPCnkTvB9siH1gx53xnfchPgkzFg/c0Sroo2h3h+pW9W9kHu
BjKNIX3yRjt9St1kci/pMfL2HeH4lY4/5o3doI9fHadhPWIx7Jv2lnMt+vaKaMs3bH+C0SYilFsk
O9UQRUoreChIOpjA5VYr7i8kkZLhZHFH/PsrmvL6yF329DqofwqD9gNPayWrXMtiNPUs2jtGc9TM
ORCfcIecfrLQShDOj1mNyA6wuPretpZsuK0XROw3CkY3magi8DfgcjojDXzM2KQp4brFuQFEBRBU
1og2irwpnneteUQaF+EBDsnKmctTXGk3tUi1zOuOf4dkdPc52Q2irGr+7d3kPJ7zJvLyEvmyVlra
LqQLDItq3PEE9gnap//rDnfLiTCZf+bQKUdD3sgXaKAqeG60FRSRlaliYdrGcKknm+E5kNC6hZvK
vsocqcfL/QYv6oBCoDCkjLDmZSZlYg4OsSsajaOgaiBGZ/X8c2klKX0qNHgp9wrBGlU9Khg8mc8D
9GYChENvlS/WaFgM72cHjwObDPzyLJGNwpZA7IloE0CkFCU1cEeawNg5ECDjw7qVTNWMW61J6sji
NRejZwtlA/7pkUA3tjZiuNioTWcLPrvkf1qACB7VAJ4lggTzHnLl1t6D3Bt+dex19ySiUVDeSoZL
8DK51cUXP7hDArV9NVXHGf+wsKJV6Sc3O3Itp7j2bqsLSv6mkaDSaijEsC/gLY3bi/LbLx3shkFk
h40LyIKnRQBDPrLunpTFHepc13vHSEnplegvl5HNcVzPiGybS6cIZcbKs5rqfoqMkgG17BRopf8b
iJE+rKTZQrfTWQXSaPAYsfTyjSlMSXS5rRJWSvOdgDojxFkVNkf4r5Ig/WS6V4A6JsGoeCLRt0q+
bmDua4tNTaXi5qU8x/r039oHiFEF1eTjlLTSiHNwoPSVHhpTnClqwAqD5okYCtjt0JfdQWjkGYnH
Oq9zSRXrUW/qWvRXxwWTN2KgWbfYu5tJBfL8rwckefKWKtL24WGaDyQ1ztnjEO37mIcIxtu9xLyF
QhHZNpUHIb+uFrAgajwZicI1IguZp8qSUpYQjcSeQNtU63rHa2RT3KA2O1F+v2Iw8aVhO/7CnlqA
+fm6k9/e2vK+8kSIv7oQ3GvXbVP9njynmKMFJquwWjgc/HHuz7VpWPkQmyArmFNLO4W1dqc2aVMr
uCywTbF+zliK82lqA0rXYtphYEuvOKTvoIPpLw3fvhtzOtb554DmgRP5qiNeTu6OKxX/eDB7fMqg
jxt1txbm0QIG02BrVpyoKZr/qoidSHbz866PpyBjWy2xi+rPGvuSpmxVt8XMuxkMLI5a2a4gSyhz
FF4LRbVaH6DUnf8r1ZA8WJQD5EZ6RZw6Pj6gDJpgWzFNvIfpFgsWQxJt3j/15PJbcYRgbFX/0jMy
lt9ObIKz2z48ok+GzCRudjWeawwJyneGWlLt35ybnsKHNv2H0cMFDoWEIh4g68sUoQkjhZdnq87a
CAdEEwqtltTIJip7fMuIUQw7A0lnu4iKW2dmQraeuNg0AnkMZTBFWCRI7mea1BOxlW5oK9GhTPYf
pvTkAYAMP4NsSldW0AJjy+5j3EKXMUJiANUW0hkSk3T5uh5xtjIUbYVH98prm9wwz9sIsw7C8+k5
S8XsWp9vxgpd05fcLNh5QwaPLY4zqDSDeW103t6n08Wa7iMT/BTrqbrJHE3hVNq7Ld+qg81kEi+c
7iqH+RbBjY7M2gpPrzbPn+fa0ovdHwps2N/WfsfnuM5cWeKp1re3zaZfYJVVoD9AG+KyLkZYivjn
5vLfkQCaG1pXuBEg2KV2fpeag4+ZlB+F793XvsqxRtMwlf+a9muNknBfDkpiuFhpl/rsa+QRjJRb
+Vw+FSxX0IopyYyEjbHdRsFtCWiVSv/A8p+QsmAKAyItvD85j6u09RXCaMQ1frwOTO6WP9FRc/cT
4h3Sfo1diWPAtgwKTKe9mvYnB7xDO8juQaRHCpJ9H9qUbpgSUDBnmr0RYOYRwi9+G3JC2hPdbgjM
DsEQs/zvdVOoNUcrvCh8mKql8I4JTwQtmDnVoST9qN2l762E5TpOObaFycToNoJG18tjNGS+lW74
DeroPAAy9/AXTE/zQ7hsgpiwBtQecw81S23+nefGq5PKDLoCCA1eoI9k1FgtgM7dXEx0N8nl/Bbd
/aDszA2h08YZMC67Lk9p831LsOLqqwKS5MQkTwsxlE1J8HhLG6mgYlKRDT2F3ZnHhBePrSHj70cL
Flo35e6liehfafxZiQBwAv9mgvbPqj9eQuBqITIqEc0dVfO3WelHBSQihEgTLaomVV+3zHHajopx
bJESnqlBLZsa0Vs8apanhu+6fOMQu2JL+QhKgegrpq2lgAB+U9P5kPWeENE6PLw8Hgy0FfGl4Kwx
n0JkXc/9saFJ3BMw3AhSpWomEpNLnTMfIq5P/DpMBEcrT0cRuEe0ypJ6yA5a0unugskXx5dNpxPE
PQXKNx3RLm3xOL9lDNe6YbSsH97b/zaY4RcuI2cOMvioyuFzp+EOwE0oTyhIxQAibLTJ05z3QqzD
IS35YHya/p0epxd9MFcXspTwBxyz0NijFqbP7X5hnqm5jn+kogjQYkXIDxD5b7n1qCpkvDjfSKz2
OPCn5v4TcIB3062UFS1gTQ9Y6kS01DVE74ywp/3ghrlOThvFlQ4LrbGdQX4VoADkXoHBsamq7kUE
2Dzv/CleBN9hagtNOcs3fDCnYUZIvyYidCb4ouC5PxXelhLw1U0YKm0vxnVP31ESwCTp1CFB7icH
CERg27LQ2MaG5CmlRAzYIW9815hqaCZt1Y5I2yMYPeYmxzBndg1SoI9vn/+Vmf51xQF344ZNcBue
iuHsMFLg8BYpMiI3TH9Wz2mjQEQFUv6eTd1YXTm2av6gACt4HSgzFiLWS1oNzCPTXk2+WD2NB6RX
qWTAvXgYCEUOM6xWI/JDC8rBusBkajzgUOZxFuCFeAeknzdS1IXhnizXHjaN3An/jXhrbQyVhU8g
8mmRyv1BuVbtdcNn1+wzsKVK8Dudkm7vCLU9NaI08FbwB/Hc3qAUMW2BDKGQQKw49DBafC+fbrDx
n4b+vTdp1gSBIgHhofk3kkZRFoP3thuj3XyIbURv5Ubud/01uiR6QOxW9NUE2987bExSGL/gLEUL
s/lT9L6XA1tpyzciOEI75cUvczm6RpaYbiECEKiWEBWjj5tJju3MQE4NTsNKMvsXsvUO/9XgWLFs
OJzwlLk9i5G9wb1iVs09MIQxhbvA/Y7MqArAZbki/gRBREdouMfqurutgVjtScbhjWjcgV1KrD3l
kmL9ZrkxmqnFPrrE+TTN9eKYIzs7B55oDGdCTAFgBazEDni6vtcgMfE3BH6G6SR/wrICT3VnGR40
Ytb/3YRPTfytslqmgBK4Fkyb9St1pSYRGQqScgntiOY7rDI7/fhuGP5ofhlbFh/PTPLIdBWBnxsB
Jzcvus6oAJVIRxrQGXWa9LBUFwmqURX7T1nuAiwVBeNnCe5JZMFrZ2Wq4kaIZvjrGfNyOPFWRNXY
iWG/BRe3cw1lIOTAors65wiuC8AsTssG/xrtQ4mORpqDFvYuO3/yfvYF5uB/tbPuWtdKEyxhGaUO
atDnnOFVB1idaTIbUAtCpYYhdM6DXd+5X6kn9m2/mc0wpJ+iI6xpyo6TXoL2yUex2tzxtq5okwoE
FuW4QuDgF85BG4MGM64XT4Wmt1WYSNwBoaez/YVdOWqcP15jeT50XFglr7/7Fw2CM0P1n5GGa3qo
ig8PibavIClQGK6oiERXsAGwDL4JfKPfwUHF6aa2NQLVXxBhLJR/mv/JcD3yNyueWpe7AVrqBOGs
7KC8PqjvewqhvGmkn8NAb3vdKGzeR2JNesGETFj3p0IsmMmSTeOb1J5JyPscXvQxTqheGYQQ1ykR
4Zn7fOf6xFajdfzVENI4t1fT0KNloIRfA4QFnI7d+YA9PCRPlG+2dDKMkYiZ4i1klfqHddqNQKCD
JoX9MtU7DzOYHw+2gxiSAN1DWW981QY0LK/u+G117RcDJzlcQxdp6gXFk3D0GTltR2YqSQBhnUtm
pqd43IgEjeswmsefrsB/fi9njccf9U0XdF3WHV0a2xz5IWP544d6sl7l6GSkBRLXLkFyFXdLB+Nw
a/LkSOmWL3ICiB5GMzX3zv1+Tttvp+d4Yd4vfrsosXH9ZJq0oTZIj0TTVNlwjgwnvFiPZeGOvOfL
X1bfSwEDcB38Uyc5LnNH+JFqYehcmnagEkL83FxCJhVzrC7BnYPhE6mt7Yj/WbDa6Jq7qVRPBOCP
JNx30LyYQeOJYNcGiKb1EkDImon0WZUPzQXJV8db1QfwWw0wGRbqSUqlhiXoEFFQ5atTkKLf9t86
g0nGVGz2JXVxw2lBcUATOoas2RWopX+9rLrmwuEMrOsGFfhrfeOzw9QQSczroW7mhIfcVMG7QYJJ
dZIB/NwoZWfmF5C0xjRJSSO/q1ccZE3ZDPjcM2jcNlj+8FnUGiHLOzLxLLImOpTUJBFFDmID7tcL
PoOXQHJbelhQ8GC9CdHhmV6istc/ZWUrHgtcFD9mfHrMOu9VWrWwGsU9t6Z6qXFCHLS3DEY50hC3
Osq0F7X5Y/Vl07k30B3C5cxEuWNf1cHhWUaF1itIDujnu8g++rZqyLtIcZwRad8gfpzeAsksS96a
e9SwrkfIa7hf9iqS81q6112sLElVqi+S8/DuT0hROxHQQPJYIKDsgOgXfg4YpwdFUuTB7WcAeUR3
vdiZ/B9MCfh+s1YbmrUG8TVZGvhr80lNa6j30PkjhZz+iA4lTjdACKso/leUU+b39a/N51MMBq4J
tkuhXsx9aruy8S9cR8RAX3Gki5fLBIrUDG9QPEqwb+P7XboKT3AJHAgUffGQ/4H+TrGNCLKJ1Ccy
uOILspHNhzZxlW8RnnZGCxpYv6Y30vOWx3WprEMYP5vZqWrpAAzM/R5xr9bXT0eIsZTMEEBpEAZe
89iaLEnCYzqeNUHRITcnn9kxGKLoCf//9T9pXRmI6aWBhhCW71vpWS/eAH884vhMM8Ck7t6cmv1S
oCLr++nlceBI/IioSTdL1uivcwAu4usn7zl2ZTJEKi42Yt7rmghn9ILVnv5FcBvsw7dcFxSoO9fD
s0SxEx4D5e1C7/qY+jf6U1g2C57tb+Hg0MLR3XB5wadEIRxau07JOB9nuZoglrMSVzijynsLjH0C
zK9Htq9r7yMhpbBgkFABTPaXeTyTUl3J20ezLpMvj3rITACwPWmftVP5twhRFPPqyOO0eT1OipEh
MmMW0F9Q3XUWjN4AUtTYK+qLZLWczcVau6OV87D/h7gqx/HVwqzVucOLY/HhrCRhsHU59+wC76uG
c3YO5ASoVrB25tX6rVPWrLbGRnO/IrK5Z6wxXDAwd8yNpTGf0YnOUKNH9RsyY2fDjNTc0LXOp3hs
i/xjVFdnHS5lkpyi4b6tnLsvKLyNJ3tmkhYPc2wLvuO/M1cmxTcLJbs1M7/TarSNvML4pyaR3u1L
6KHcC9koqmOmzZtrcc49IqxQNDxpdaiTCO8yDBCEX6ZCIiZnxvdM6cDGSmH7Ial+dTd3ufqgguk8
f7YZHTerTVcaw2C2QlLcIUGLd0HHQ959nBpPKUpGhJ+3kUVGawiIxgbzr1zbpwxmESdhcF4zTuq/
K/AVy/NLLBvREMjcIzp4JJmK6piKU1mm6V+/OvHjUBApnAPTKp3Kjy+X158RcWk5/n6jfh5PXpDT
/t6dAnrJXVF3E/7SRJgbLS/NROuIed/9xu5yn+3lzEetuQaWo/Hdx4OTnQmq3wiPjefwGoFF8sOT
4j/DizcU+/9BVUWPA5dQkcdfkwUO8NHt9msUOy1WPkdxSga8ZXLSIOpnhfyxo+DbzIVCuECFzFS8
fyWA6ubv7uBk7ffl5O1po7b/ACiT4l9qAI6gFesTxhRtyXEn4JnGrPn54tYr71DHgPjm4RFgMNdt
2MJvWoChlqp2NNcEKD7QcsK0bkfpkZuhTYdJrGBejvcAhCVU/j5atGKxW6tW14sF71BCgqteQEgs
JecfGdAap7vGHMQDjtNls1EeCkVFXwo5aKC8biaePJC0lYEv+75+L4Y2LRvgOXpP0hQO5kz4m6tP
APIe1RIGgxrs7O73BUWsj7kKzJLfkMkvSw/Jla6rKBjFbcVBe44cal3U/5otgunEYlTt+R6eBA44
/+sPEuwrA6cXBQA5a77neweQ3T2Bv52hCcN7zWIU1Af6SE1jl2gZz927wE+BWrJEOG1pifDtG5Sh
6mT1RSLavhYjVjAAK8Yl3Nv+nj0VXvfXSSM05qEJZOj+nPsf1T/W1+C5y9pLFuCWopzt6VVG6tmc
rhIoZynmtfzy0rbelWrJqDx57GmDDX0bqh0j+3W8x7Y4dvJ2CYlL7IBfOTPZuSWN9LGKQzbh2Eli
qRW6e3iYH2EPuETAJpT5AuoM1Zbpw/dMC9yrMYD1qmmvl+/SkYF2ZVhT/UaVL3EDpFY6mOx/Jx9A
gjBb6Jn54IXNz4ZXM0PLpEQFcylciME3IeUOrv2UzdtfBAoHPeSklZw9KLs5nU/MXim+d32kc7L5
JJkS+gFSo5HoTCMPsLNByoAA8EHwlIyEH/OKt11AqUqkySTXNeXH1ggM/3NKVUrgjTg4OaJShG2B
eoE9NUiHT+GqJCM4HmQIeuCESZZyyuy8JyLcemhkYvvbShnO/MPsZxtLPdgljWpgdA50i5Bh7Sip
MLJN0RHoZnsaPvItHjRmjEcWJN2mDJRBLI+FaQ9B0HA5nXdMGim/rM6qX7G24zYICsHY2ToZj8uy
RGA41FoMOM2A2YsTPwhanZfxE/P336lMMkAlws9sZ+b8v8MbZk687/DDT1oCNSll8qtTuuMm2CqQ
Cw/biVzlqGfMKgLtScrBso55PHFPN01LbmL0gYlrdNtaQFgz7WeU74VwYivgCFCZChhYDkZQibNo
D/d0Sw0T8hoJZ4CVdMQvBKUWJADd2E7TWR5l6ptmnh7+zNcA55bFo94WWIjVprILSxi39eSep/7k
FLNPcp5Act54dFu2xjMMSKlOOVur06LNzjnOJT++kgPdro3eXHiqh+wYSvQlEm3aGVdLj5BwzHMq
fb3LgYsvX2wLnRrOBsOlEpjz8GSQlgCUQxsboIcy82DmEFPpbe+ge0x3eda5jV8iXMN2tqexmpvw
cl4weB5CiT5VFKl3PH2tlu6nzdIFX6hYig8K5znaLr8TCoBmdYVfnO5KBAhdrpUPCo5pPmAZovsy
2XGeGn6/gSRueEGqrjwAkF6eA1H0TPfhOgk8Z8VLuWuoSotnc0QXdZO7StCJmXi8qwPfmAiTuPQd
72UQGG0JZi2R90lRpyO7Ay1/fR5HuPdpwP61p4uWVGyPWIxn8G2uz9JHEDxoxF4Ln7vQJ8oomyCr
O2gPsH8LwKeo9wCGi3UKEoLQJC7PtMrACBV7e+C5klphSSEPSJkOi54oiiThuekJFJrJk2nf64Bd
o058rSxItGMqm46ytSWDhAwlKi2iZSrgMVEnGn5Yvx7NTNlhNbLbm4EW+G4+u6W0QiqaaeTRPKsY
38RVlL8vOthcRtIjSdIPQLo/qYIfPUeUqmYNhoWf9jRBqsEO2MyeUG7FsXAsa/sE06xoHyCjMb7X
i4AXs2OK4HX4G1ZpmmGQvsgWZW6z/3c/7Ew55+xWzjqQ8VrtW6RLpr0CYBxHFKAHk8UVn4ADrnWt
Lcl3VjehjSQYWv2Hky91SntqWdR9syLTJZ5NXS9mv2O+AyAHphPhBq5fbYe5NPyRV8PKB3lWcAlO
sc3pW990ikgAQIzI5/kiGSgQdZ3VvyIg4Swgwd0svnT2gfLmnxGzZeLNp8ZLWEBCWHLketQSDrw7
4y5O3/l9tRgW+ERPA/rhnkHeCEZSPmb1sED6wwg7NGXexJWLZlwsJVzX2hLnvnPuS+riOno87mDp
/VjCcJ8bUgRGT629UzvmKfzg1DVAt8VeTKrXVEVGzFGynoWbgHGr5J0F6Y0voJUxBSMoP1SonG2e
fCgyKtHkaQ7PFUvmgeZCAozsd0gGE7PoditgVdc5XyEK+1XM4vwEZfS6JjliUr+u2dscJil4yP36
/qAKaHL+fHQpX0VKAgZVicBIl0l8X309b6xt2A03jzKdnz6aN39lscOOaV1L24VvUuKmE3S4K/jv
kt5eG3gM5V+g+VLE+agOIbTetnHk9HvJ5LBx96bV9PqM2R4EfrJ/cMCCppjP7J3CPJ7/MUxJA3Hk
7oTxmBZE2ChMqoW8k5VP9muYPeDbjTtUQD4s8Ubm4Nyy2w7KHztmU/bHy0MN9bwD2VUhrD7n/HLe
fV9WzOumCDvgms8qCN5QWPrZwE6QvKyaXI7We2tzIrv/7FSRXbBOisRPepWnv71e3Ou9neuCVleq
EjoUQW7ljUiNTGCo2pToj7iM9aE+72/I2fuco1cvzvu8hHwTM3+0YcbcvG9nST9DNn+oK8i91xpf
tijW1gfAZf6UoMJqYYypI+WeA0etEhVNrTYLRZFLl7LmZySGpztUX7dD+wU82TlQBDVZO5bMsjew
7sxV+qg/DJiZ6tLve0GRg7jiCS2gLeZr5y8vIJZ4SY17ufahKD/SmrnMdUjuLTkxmWtdHfNnqgGb
mwDoMsdxXyDEunEaBfNFIH8ncJOds7sNgTlL05oyGVuLx4pa+e3z5T4YLLYlYUr2V9lIfA/jnILB
YcZrLRIxH5PsvAYeK6gUjIMLESZ+SiUKCNg4d/tEPld5J3h3nrmGWHtw5/v5MtyWoHBY6XrTxV0Q
Ar2bEFQ6jjvlfYzUdMcu/TIUMWGTwTC5jCWtL1bWfQn4DC8EUJRHB7QNVnPdobNykX1lCNY5usgn
5/iKGVZbk7Z0xMWievKCWMX3N6LA0hdVHuYw4x8tHD5vh0ZTdQtnbqp/ttFYuakLrXNgNbRbboPx
t98miBjyKA2hIisXdm/5+YesoYHGppxXz7w4zuF6G7VPaHnwiCiSF/u4bWvm4KnEeBUli+cXhthL
iWD2xJTZ/hanVEtBbUUTJEfBjmpoxuYwA9DxPc8YE3dJZOn/an9+JakwbE6WKFtn9qfi0aBtzf1b
H4sdx+hqc94Dam+t71yktbotDj1JQX/1jHTBt/VYrcHSiV4XXfodznkY5gkiDp7L8rp2MfI4wKJx
drtBm/QRn5jNkZ/+X2ETTCKmNePho4PoniJIokJXQki4VDolPbeW5Pz8INRX90ZvoLM8/5CBIrU1
HuFgattqaXSy7MtK3mmqL6a6I/je0B8b61pu0cNQ2a3gVqk0jK2Ep/IciBRgbjxAS7xfkFiYlt9C
eDWLUgwj5o8ArQDCuzipYNCk2/bpffS773LVPxb+7ypqz3StVWF4igee4hmmjDqt7/7NIZqopfxl
48HS2iLazKzYvEi04mR+KgrXyz1PEmVIqeIyLEVtc+WE7C2tAgJriNbNU2GtqOKnKSgBO0Zy7h44
EGrbHaBBiS5fX5mnUpEOaH/T284SWxqsgPsZ/gDKKom+5VCVU0yRVX4c7WO+Ty4NrWso3H6OTh6d
6/e/Y3gfwJuFzxmo8tPL6yu/ExFQffN/IEsCmbb4wbyhMsk9Np+4LWKMRaAmJm7jIvwcDMXvl8uS
QsmoOb7Dzfoo5KH7LKrtIIRbcRnIlWh+sQaZA7D9u/yCkZt1wbdCBRpyNKboBT3QeL+LQsRXXEP7
M06MNSCFv1lLyGWzDEKzLiKPWrQkOf2T2MKjNH2acV4LCO/DFNRJqIxdGnozDTAJPuHKiOjZ9pqw
Jt0jhMfc19S8Kn4xKVCA9ASws6MVsS4CqJCBsIGl8N3qb+Rgc0dzepxSvp8yqvejrA7ivyUQabuP
9l2ZeBrQQOnhvUfAXkjngQH0Vqps020bKUBJ0kF/rGHOtd7j+2bIQqkTSonfJPExvfrhGvdL248X
/zPMaIXP7uEedANsoT9gDL/ZOS8mrKBA4rNuCw0H0Icf7ceAbriwJ6tgzceZNYe1SCoXlzFaJyJq
6dNUX+DcZSes2oRXtJv2WImjbFxajaV1ZDtfg2MWLZKDTYA62N9ZR2lgjhiDI6cdPOEh79LrkJps
RTlZ8xtCAc/OiRaD2XHSgvqIcPi8vJuMtDGhuGC1yVPvNYVgsznmabqOUeOGG46dNzHr6mXMnzAL
75J6qYonMiHqxoODH+HfW2KLHRft90QDHXi1cqk9tstuk3kD7uttShFTAZbnN24WPda/7XySEJJB
CSCcDPXF6+EN1FlxXTphTaYpQXyAx07L1LktEO4Fglta8rGO8X7bXqT9bWzNW1cPyh8k6v3Ww+Z5
vyXafvzrYXnvkGIl+PDpX9p5g1PeVf04tQlLQ7mYnYM53wYcyhQLHtxehguAqNHLLKLbLEzKsgD8
3hACorN704CbpUb9S/g9HLToEYBTjvGCrRPioTNNaZQ/j1CggOgY/SuR5yBHyRwG0QN4xHtXBsdh
/98OQASVarSMqOQOP2cVhlyn11uTBq+Ld7uR4DRtRmzl6V2YUCAWGVXfGTboFyXTLk/ul2Z/p9EY
Xb18y8d21fWPX8lf+sBiBDNV50cutr5RdB7j0aSh69mNmzYNItkSkkdbHY3O0kCCX3wRNs0n1jlq
Kyp2TmZaeyPkK8WqWZnMWfCfvN9hov1i/Vd1QrKK7MIrMM7kjbqL241dv2Z7ZmcLQgWQD0oMs9xq
9nY35WJPMieCwcrNhsQBt+g7lAhZWMmwyl1z5X0BLFJ34lbVlFKTalbG1KRGg4GKasz/MR1Qdaaw
fhxa82W2/H3JeWuPVjx2dV6GSTGKvtArojgnF6w591BPxyhbgbZINfNKSMFDeJMgLS/2KZ9any+c
cYk1c9OEqm5MmI0zLaImCIE+aY8NApqOx7SsrfJJo8uAIHWal6Rf0v9hzWdXGfOdXYYyekX/D8nQ
HoGj7uEjhvnllmZs+Iv8YFzvIjkIF2Uw4yocCvdBacjAhpsrwEdtDuyTn99mOvJn6ptLUPha5bJZ
HPoFmVJuW/ds+44npTX3OqOHdSUmE0/sdB9UArG+UiIhHk5+kG44KZLGPc7XOTvtgTRAhopDcRfS
zRJibCXsn6FTY3YUf1fPN8Iy8jrf99yVUvDN2r6w9A6d8EjMUOUsTY0KW4MUf2YoGaD0UCjhlxdQ
uRwY8aaEjSJ7VpO14KgN2SFtt+lJeYNpXfBlrGAcfG9jvYwj8LZ43zWkWg7WyjTHEUP9gYiE3gg5
uZwfNN8wEbNyg5/p5X1RWI9jg71qRMB+S+YmiGij2xUIjOROLfqQNHAoxzfjQh5er3y+7+r0ovwE
Wsrq6SU65Wqqdl2Crz+qk75dczhzxEq3slgtR7V7sqvZTGW4+rOD/RGWpPO7d1jnPxSTobOcmPlH
mM8Jq3CvbHN8Wy3vRpmYeiSHMjqvQIxx4Zjvv392aarzMawHcMl5FJH1C39b6rw7/F0euIBVLEKY
btZ3L/r3z7sODtkZvOfCIn9pG8f+9PbeTXlSy/zUemGYXjKfoQTw86zRNw1R3muYPWZ6HpFTq1Yq
2GmSgA2S7ZdUoRGRxtVwIJkAR7UBvgSLS2GP0DV/5WaV32vrTIZ7RoR0fj4ETHfrL1zJoyrpYQds
M2I+z/1At3h18xZQc8tiFLIPHsaZOEdzzvnnn6TskdbFryAsUi1oYJ+dxcd9B0ItFXqX7J4xsb1m
48m71tbMssAY+sVXCOwpWGPWCMMtjJh8w1Tm/Tl701TWyol4ZP3hDXSuFxuTkZ3OgugwCzn4pftC
hLQnCPeX2u3VhMDCKESlRQZO9dJe/0D/pVdrjR8ADVXdJ1flsz8RMCyPkzXdrH2EZqYf0zW3/B90
H8JKDi3qH4g4qCs0hpeWxZH+ynzMThTxxeqUunoPVfR4wV2Hb/kBlMFX1xm2BwM6b64QIoqjFXOQ
v0W+fGlONZhyw4ko0zzT+JsDNTU3qkxMvbR2oiAfFiKD6/0RFqlMATg2SzQ6DkA3UZulC8gOSpcK
ZokuCyabF0ubXwAHlove02683+IUOyl9DYeGPbg7azuRnnmOHjkLM1wvVo7+LD/Kf4a8V0RYyYAJ
D0Ev2/REYMpaelSNhorAoLy/ZBHJyX9fFAPc1pF59gwPKvFZcObkdSawO8lkwkCAptyaqLHvR0fZ
kNvW4Y/OrQLN6hBHOd+Smj/10t+YHdegXXxsZ3teqD9soI7BDtX6kGw9hexXB3Pgq77XsmkK6Sj6
4VpHr3imz7Fb4FGS/3Lef6pO6ypT5jEjAty6gsm5V8aha3qIglNpHns/p2kYJ9YA7S1ItaNzo5cq
dlU72HJiQMC0y4IfLBLBQCoIX+lqitBdJhPBlzbhMzFsJGCoxE4uqRHiiCGB2YLx61i6E5JimBhc
Elfo1iypguK5y403hXYzaxBTGGRTINoG7yHu6OtY8VKlKQZbvWWOT/+nOtnTMaNhAmDV1wQL16CY
kH70/U92M93rGcaKnbJEZvfOQ6z/sDlom38/FnggHfZuIRre4eIYYnm03MHwsn9bpJfl72LZTd3r
tJmKcgsy3OJcYKwMfNe3eU9+Q7AImVlEdTXZAhJZo+jFv3+dLPsStr4jHDiVJSBaqLqt5pY+C91X
6Hu6j9Qq6kide0Qt6ydcMpXhtsQ8cE8XrRuI396ouThNxuHB7ZPPnoX6ONBqCxc71wm3LxoZubNP
urPTR3EHHm+UUjFZVZlNVZlVxSFzCULBffrQV4uxfysHisebK5YFy9hwDASCHAfaDwN0/qwPhYKh
AN/4gmG3VCezlfaOxFoyCIBdbnIBzn3bHjlfXdGcm3tNxP2r+Mhp8u1mxSdwYntVlQYO1A2Rd1QQ
XkxclHJOJYq5PCkAJtnJVGHBTIYlcvwYDS10oORje3QcnLtrMjnuPeS+4uM0QwA1KlFHMnvhHQfN
DPGBkpi8senLbTif/5zThuhRVJlWDjrnJ9VBDZitbrkr6hleOa4+GlpwX+qVKNvBB8SZXCc/7pez
GLCQiMXM0v+9JTKdKn4fJGICzA9BbLTxTFuhwDyTfk02Zyba3CvoPhN6Va5HNmTtVXMhdIKJRrRU
UUUxXUsqatv0an7Xc5YdJ1T/6hDYqJ4vAsXAqqKUAC/q80F3r6VKYEGwGKLZgsRWrqEweG67XVtj
HcqOXd2LrfPgovxgH28j1+bfdFvdOyq0gECoNafD2FiXfahGlUatM3InH7yyPG0Pdk0qBObwqF2r
dE2/LhhwMBGiDEpSzYxoE3ys129jsVk5UKueKxc07Lz5c1RTfYx17EqqCnHxWr/xyBSPMcxnZwvV
JUPlmGi0lsXZljqE8AkQ+5H9uDTKv0VIcsjiV5o4JFuuNmEF4WCr6rqHdxNZ5mwOa15hc2zEE0hV
K/V3LsZD5GMVUAmMQf0Ld4XZp0sHnDRnAgmRGryZr6tW2AgPQS2H2PlpKebZ3coRaH9RKoI8YfMl
bIY8mFSEUxNTi4XR5LaR7/tJU4fj7EiETEmTXTF9hNhWVvRtdHmrMLxJippZdcYepeA8FcZMxrFH
Em4z1zqCOGh5DfwFJ/VRTzl6349OTeIBXapQ33G8+Uny9w9bWipKep1mBWCXp+gQuFWinunu4NTF
Gme/SQca7nS91blIDcvAGtM8nkk90WQ/a+i1ugIob+1VikgcmOGrY/7FAYid1+5dgHoRidbDosey
e9AJAS+pOmqygHt7hlfQRl7BPS78DtcbMI+/xWr1ArvEtu1jrghRjZsYfSa6+zNW3aGGqcqG6V40
NM1z6SUB9HAKHfcR309ncQA5VJZPw7FAMYUpCR55dGWuvwOGFrbvEe7DbQ/j13KQt9eMoVH04z0s
mTU5qF969w9fu9wnVyjxLn2LNg/DrGJeD8bLiOrJaomN8byxDjtkn42JU39w+TnAXx4ynR4pJAz5
yrUjSx7Y5GlkPzCHTiJxZhGAg+w1Wke71CH2WQItFBzJV7WmljYsIBcds4RdhcE0Xsmz10l9Yxpq
Sp83GhiCWc7kSpBucZf8ILmI05Blr7iqvr4j2/qhXDcW7SnvUAr/NzjjZbfjFJFZrit4O3naoRaN
PoP3HxMDz+iGfi0HwHRV6uLCj1T7ymHMMyFFWbYos4Cli9nQl4VUSrvO2sTkwMzTo+Euf6dZv8lg
nNpBrcj3eNnu0PqNFq5pBcs8atL8AKLcowcl2EyhmFby3KdnKSV3jgaDbvknQbnzsBerubu3tgFp
annBpOWf4B5slZuGm6mSFTXkMNBcqsrwPQiZUOdUsAjyRM05Of4K7qEetimlWQMX71ID6SIhgTGf
g700DM1ovWBmkiqxfX+ayTzSIsM/AUfNR/mJnpwYA7kt41NpQou4CtIX5nCxP0Mz5GZVfTbgF4J7
AVSccN2WQYHZeTIHkL93wflyPXEyuNeyp5XPW+caK+Px5J0Q32JZEPKu+YZ3wrH/d+3hpZj+4rv0
XTMf4trPtY5P5TxVQJ3XVLLaSHYGXNY/prc5uIV6sfb8mFD1TLHGpu9c2XMV/W4m9gro+PC8qr9V
7XMoBabCTKMw9U8HHRuHCCeLNJgQ75clxTKDPjXfI7HGmZ36MS0xovYmK/wDtORZv77JogS43ikx
ZIZHWfIPQwdGC9CJSIeNbwdAXb7nzsB3cvtnu8STHWdzOCeE8B22XupeZ3zjiEegLVR+xFuR2j3F
gr70uaNHgqnhZMsZzEl7nxcAwnWBrs9QDcFB84dOtr0kW2XjqRDbRz9ZcFBS3GsabzQGT/4zrbVb
GnDG+zdpUqATTsiGJZhpa7eqFz4EGIWFKrtdhYdTrF30G8YDuM/AV7u7thkWovgwPOgSAQEV/PtR
+7T2+uKRB+S+OY4GTorxeoqkuV0thPJ9wnFSbe3r4FxFikkX/ztAg2F+viq9d+/cYOg6frmWL5QW
0yvz2DpPh35S3vkZID+suKHLdGgpQDbnCxo/RakuHiYEALxsvGj0De9ZuHgVTlbK4kT0R8ohpupu
JKmCtdjX0zbV0FBq2cmfsWh+QuvkYy+fHn48lVb3f2C03j60jWc8/jSU1250BBAao2Gx8KQwaeyL
cqlRPrC0CldtqCmEh5TUlBJzR7ZTmLLyk7p5/GJZ5PElupHG8OasdWzfFtdHSqXT2VfhRcBDKcLD
g5XOQtpe8dXk7nHBPQ2cyXqg+FvdAOOGLP6T2PRm4oui8pCj+ov2mSy42VIK7IwXOquV2jHzTYYo
cxnKb93luJdrHh437oVWblW4W/JUOZ0hxv98YD9whd9ZIIqChP5W8vfTBzzmZNbx9neVX9s8Qsjo
TX7uEyO/Up1U5SIhmwv4KWzgn7vws5ZIIMbLWcTquE+1xzyBcBikKF3L8j8XKHGAJZ+6wzHXsmzk
gBIohfBrguqJOqHFO8dzlnFjOsBlPhGxr9LJKIPQUwz/HK0Et9fO0NlgXIlQ0vpf+YrdfBWrnEXm
+LtU88gW/NxakO1+28C07hLeK/PUijvok9oIIiEKZYiWiomsVF92fZ/btx6EViA555TB+gzEvBZI
IXPAfz58xgUJwcsb7m15HgSNOZqi8bCE1+XWHOHmZlZq/enTpbvzhPjecYvRvG5cO/XwXn3I+kN9
8OoTHeBcPKrJew+JWZMUHffPFczVwWeUWD+jMWRHScvBj+tIQCgG5pLSFX+dpG2ys0l3LetD1A0L
EEZrcFBpmU41CX980se/V3ul6FBFR3cswFZv2vE3Ucj8mcwTaMhT5HH1r+Stl0BwdczRKbqE+yuJ
fP+G0pt27ak3mobej9eLmKMkGicjN9gUd2b1s/oyqyhvmutUf04d6eJI3UJshBP/13PZU0nuZZ/e
Ogc/D44+nuPEFtYGKWC0pFFg4qdF6Go7UHdBPlNh/yH4GqFcwPeouZsJYkSP0Cp/Sz7VtBfDyfqS
cUGo+Ituo/uOLeaF9Elm2vZKdqZ73Z6LFCLlPgGw7/+oV9de+FOzm7BwBznXmQYhexu/lTOgcCF7
JSZyPhbLIud9+7vPzsJqhW4uPxZJ9Kx6lbqTr5gxopP2VwdeLewvRQk1oUt1Jj2rTBvdfRWYqq4B
5hdABETMJ4NdOGjVOU3sAVOZLjPbDPAhnZgSABd2JZHCDHKfVi1b0SI6ikeaXMRkxNEVCYrrs8UZ
SWZq6yVgJYim+d4fJV/N48iwSs2v1NrLGH2Bof1dQp4+xzNFgOR1i6v607rol5bSBgNDkJFsMcI6
sOBdx+34R60PFmYeFh3lGjFiQMa/MgnJYpkXLzHq+Coo+20m+qSn+KzZ2ij7RuYIu8imYTQ0lnH2
dkuDXe3FmU7/1lHOQs+1TvgNzLtSC4eawq+LzbFd9MKex7OM2WKNMypEZyVLIriEcTnAy4etIh0I
75cY+wQWeCVCho/gNjad+M8p7TuLzvBcSRkHIIZKh5HzIEBiFBkHo8WyX9kKa/qZ3TTAiUAAcQ5W
XHHy0l1JfHvEcrfDZ/muAro/aJIDlErGEJwKUiy5sxIwoTUmPZP76D5vBt5fZJ8zcYjUwy26mNQu
J9crcA7bbXkPbq6kkdRd2maFmPdQ2yvj3MQVKZhZo0Z9lT/VkNZSsz8ul5NSzIUb1hKyCglUe+I7
PoGEvUaL5kjgfLADKpMSpoK2Wa4cGecvaDR7BMK1plyDe341MjkGSnY60+8D6RzSEeOoy9BaZAvd
mq2R7u8hxZTAmvwitvzg39vjnwvh80IpSeDLlDG7pmY08QdgKC7l6xWC+yRG5nXxsbhg7wEESAqp
XKOqoX9Am/A+mzO3yW6qcU/G31s8egK0JHZTCCz2ra5wy6ucMT3voLYdqghOdpB1/6GwyqlOE9tT
dfyreeWmbYCvdT7qQtFMu4rkfXA8bA+Rn+3mSejoqmiVCtBo7WN67FQ6UBmxvhVDwNmUC3twoPoH
o2EmWqHd92yS3y09PCaaHQnLaWLUDi3mPpvpg4DcVaGDtOYoSKqD7OeXSkKQY/HdfVCrTFnyZw2C
MUU5KjHVDtASWtWPFi/NszYxTDO7WHAVl0btD2lj6kIM8ypzzi2lfsIkv6XGgWE6F+dxibpCyAd5
bUxKaNhDCJwAQDrNlzj4v4HKZURZz7ZGFwm5kHdHyw027satAD5qEcQRov+ElV/Ax3qardinWcAk
hLVSEbkLQnqpufDcGlWr14V3xq1r+0hDOA3jD29viNlIkH+RRxRY9bcZ8Aci+CdglAZed2HCm1ER
hy4Kxjc+WNPgazejhVYvl66iYd9rJX+6gamLQgWk5Yo9k0GDrDDBxuzL/zoEgQXq3NqXi0bLHCEB
FD629LouEynI7Y9bAeACKQKc6XkjH4BdjXlhQD8Xubt9bRCfkpHAeGPedmGEWPbKKvK8YZFCjCIE
KV1v6k5Dls32sweonrIULXcauJs9SSfn360fTdkUrYchbgcPfYOUvrKq3dalsivmCLT3SrM7Qokp
HzIAl2S8PjcqUxAqSaEvnS5c8TbvMMfDe3ObZrPvB9FOYk15elFqiPiMuijXOntR5Uc7uBkaXG7C
k9CFxMDjTcJ5SNZoVTYVVFph9d4KQQWYlAqnGsOWONfb92vOOZ3d4HjM8CblV0+t23hGJIjb76Ie
Rl4xGpDo9LgxNAvn/2FVooaIWqTzp6qH1Fq5d9l7uEj0tgzo2cENYEqo8u5HRqK8d27mWCZ188eM
tN5Z8cm/gIdpdfPzCaI7WwTkzIx7JcDPv90OTpwIHFFHCR8F+rUPtU+LLaghRHAh/AXTNgTBL2Xm
1+eZQabzblcDgLeyYahlILdrl9hg1PWICkhER78ovMPMfjw6C2IUG5rn/A8fyr5VfNfkOiGoIT2U
IOmJK6HtLYAikEGzkET3N8L9iagcxidFD3IQwisw8Gj4pHdEWWUFKVWz5zJuQkZ6h4XJLceEoUPn
bYnHGt1IXVz3C2N1EPaG/sXySFBA/qwGWxMm9sZTJ8dJ4jrDo41pZXkfGrX4J1wMvZZgLWApT8ys
qfEN5fX9BLuspmqw0j057SWj1Le77uZ2RX3LAKW/JnjF6fglqzHkmKsoKpw0xUn6XoylcYyo3UFW
59b3Ner3DN+0wh6f2wuVO2MqyMBZWVuJsTsHX8ENQyxhT6dhqszMziJvc2x88h+i/hT4+IVgtooU
QEDz7fsrbKYlR69HH16phUWQ5bLrpwBX5ZE1nhxCkHC1sJxPg0LuyK/u0l2W5VtalsNqVso4fAhs
NCUc8BW1VGLnWD2npNqs7IdJcwq8EkTqf2KFFCZBKQkMA4BnsUVEGOtrkHzaViQwGtmmztCaRvHi
dJiIKjes8nykolRaYnevSdtFl6i2sT41AL8i7DeYrn4nPq7tvbXHVpo+I+JS9jwypnyoJrfM/fin
aotfDgjkmBscovFu6a4nHpA6tYYqIYnqjLsy/LjGLSG2u+ckB1+K7h9NqC0azD8yscUBZy7QWeG1
9e6NqlwAaMV2v/iGFLp0HfLnoIj54Lzmbbz/+myfYi9lXU6PRxlraLqOGi3Aa6FjJeRNKpDATRqR
04VAfXNgww3X6m8G8t9uQyoSc2Cu/0tnp7GjHe5tzmY3fSxYyO5TczyDFOo7cPwDGlfAHrXhfR8R
R6kQSA4uOSFX/6dabbiYAf8YUamIagZZbogeYGkUjV+PctN8+afmzWSvcYaL16FWgZMzQonhTH1M
3+237nLHYYtYiB6xq2tT5RNvNCUxHM35OKrMipW/Yy//dhZBc0iGnN/DiYjZ0d3VewgrJr2ZMjp1
hO1lnolESMXWGBW2+W7Ug3z9bzxXccqKkv7EADzJc/x0+T01j1foVXQCpKrF5QKiVlReLE+2N3Ie
esF0iVzpiBsoFQfeo0/RYE9mor8u3Cy25kPcYCiRxd2sPM6TxD2+fQG6c8kTpEFarbN47PuyHxdm
psp/3CnVVo5C7dljYbC9GeRVDLz3RPM+eXVndtwh2pZNIVFF2z5eBs6DgpSiSvFMwtBGtdpyqeNZ
IysHhOVarOsBQmUidw1/6q7OgKDngWODFpQcSw/OjKKxU0Xs8y4hiUEs+AgrjHa9Frus0zTwS2dN
7SsOQauG5SS5PgGHh0vUMfR0PDgzrLVrZxa5PUoxZu+ajz5HpqsS/wWbOyJrubV+keICUlCWxI2l
OaAb8z7r6Wy1IGjeSx/GhNpWUAAe9e4dDNv9htT1ACdTE7/4QUYtKQjZkNoEJX3RFWSEhBlkIPQf
gb7ieul2ZJBf7ren5dXI+H9/Bm80QdeBAKsa4DZINHhFVVA+5IrPeXmvf2PDKSHl6P5IuLLjiMS9
Ra3k9ar4urICCtc1u9ExBqzAXIMP3NDNjBBKkAU4WThvG+e3SonVlL7FmyA07Wz7rbSWSuXhXZef
zK7wzS5lW0WHPhg+KkPgR5qaqreEqVASMEL5naGZv0WBeH4g7mSyH2Z7qXUbX1w01JR5keMQmjuK
qEg5pqSRZYj0V1veTwLtrgeTzDWoTLnpb0Jl8yRlolbywkt04S+87QnrBfU7VsKhRbKZWsmxwjM6
SdSvqYjdxenreXAlpRo4kqFDdpdjpkS/gfMbHJvlino4r4FEIodpnwYF1h+FrQzjF0oGYMyRjbtv
yagZu080xOPQMs9SqcJNeSFoonO8yqWH4+00p3VX2/Ppcl6WfY+eVq3C55t9w2r2Sj2Ygff7HTcB
CPv+GPNGuKqhepM6eyWXGNv6iezsmL74sOTDjAGc1j2hGBEYc1J0txgdHjHnJpgAGJpSJRnijCFK
B3HBNinFoF73MGyPNLsFLqQDYHOB4HKEmbw3ARKKmME5g9CYOFQQ3s5APwnQiFKv+Dl5/KdddgI8
Mb7MknlC5AozXybqaRFBR92XDR4Pv2iItWuMALhBhAQtCcb9YAAKqwI0T+m9r+G1pG+9dCFpeS70
eQlGDz6NdUU4xr2fHiJR5AfsE1/0DCVSVfS7u0E0ZQU07QJHKsawsMPpaONf7M/yrPBGW3N91TEe
5TMr8p14nWm2ZKhHRIF/gAaRe6/s3BMY5lELXr2RFQySaYS7SiIGOf5xw59dp77vr/8vyE5JmBDg
RaJM2jeteeoF9DW6fFVEs35HHMbNS8o9E0BxzkT86hML4FNsLaufXgaSk/cUKq4HSTr9JEaUCy+y
8fXdgLPrcakx2ScIXFmmexv45V19u6P92IGQiiDKyq9iCxwIgexvZ4m2hPhdVBuI0gUj1qf68+0G
x6oKiyDHAeCwClyUxyq3sFzzh7wiUOHYaiwIiLyIvW098U9lO65DclaGgM4E5lcg2I2G2+bBx1fb
/XjOyyt/omjzuYhlCSUDPgpHF131BK0r/BHU5FHk3piReF3gqPd5wQ3LhUEuc0tjdYrEUrpSOkNJ
49ucIKxKen7igR5aI1tsokwvNUyPngJoeLAY4BIMPvwf5zhFrNvZBwpvQJ/4JZeJfRYSugR2JTr8
qWXvT4Apru5mSQQRZEut3xjXZ9nM/YBReKCzvWDkugcSLp03rOrejbqigKVejG9Vyfs1P8Y0qSnp
YWNOu/ce18Rl60dId/iei2d6flQ1snZXlKjgf9I9lnkPZUs7V9zkYCknkoJlnjgjNTFS1I8c5c3p
j+KxJu1Xxdcfj/HAQSluAFJoDVaJEB4nexxUxGzRguwAi4DbvGiQdkMEh5tHEIrwlHNcTWhpU+vT
TiyFQ9xxtEXYnUDjoJsdP/pTbCXBMpRef6wc9ZsPTFd1iTidN1WyPH8WftvON1fg24vdV8uzJVp9
AImRDWLkhzwquaP5aHqB0SPVkoZCTkw1mbv7BmJe4OZdjTGhFGUeLbcWMMjNh4UpOEVEPmmQUgOz
v8U6Rolo3KL60WXDiUrT36lVgGZ4+0O2RqD+ChHedX0EiUHkWD//hbN881ELwPkbfUKIKommeY7E
Igwuyr3y+gboe9DLRG6cxbFq1vGM3i8CHJ8tfZmy+r28+Bvcvtqdb8QXGHOX8CabekIGkus8MJtM
uCItDh26qdG/+0v0zbahmLeEeaQ5tbRzR0zewJT/FA2I5NphHj5IRlnT/R/Jkp34y106up8NhRah
0kZd3NiAdQQKGLjpztZQBvkTwRIvfLSwUxhj5eurEROYkScvSp5G+AFHIAVU0hzbszS0deq0libe
OcBfpUPAKIJcqJFHmPQx1lNhxsbdBrbzJQ6wNUqkuDscjIplLVsef2JT+MtJsrG3Hazs/ODjqOKd
Hf4P6LqSEz0fYG9dOFNtpOO8UB5+L2pJkPIrcHVbWAZEdvXI/2D6ywaZjCrkj2PNfUyO2QZVaule
6omgeAWIx4TMcIWON8YtFl88gHWOV7iEPIDkQc5n73JAE2dVZgUXpz9EMQ8hP5zWrFgHkiPGAMxc
DjSfVxpLl0Vvc31wuBJtcgvq9jLNzDvO5DUG35AGD/vp+g1wqVFrT7MYU8eTVJL5/cijC9DkUT8h
HZsiO226di5Cc4m32c5rC5PbdbRqAePEWJrlROP/gOtzq+S7trSUL6Q2rm6LbWtBha+0rpHAU2Ru
WJ8wRu9sijvp1+U/mdkQlXpnwr3hraD5WF8S+Gl+G6c8wgaaiUFjBLu9x/OWMVUhNpxvDNcXRgtY
MDrgWRjU92IAgbEbAWdDu6igH8GTm9MTWHik/3/ETqkZ55ti05ixCAeuRrg9xm68SO41X4IP5+Fl
d1TuIIuC6602DTy28WM0tLi88ZQiDNL6TT4/zlHUjDeU/bo8LeKnT+BI5RwPWOL/gvCgvmtjE9l/
O9OpzI8wbjPZjsT5JzT+pu6J7F7Arj7gmgRjYuSmLSxHW9Ccx3xRBLzyY7OTBa304zV2skwHzkzS
USraHZFBdUNr5MmH2hPC2pTOIHe8MTg8L8wa5su8h/d6IhE/51A467WQi56oqafSaHyeOXAzGZ5r
CYUN8eCyk/LVNA281BpY+arCeL1eEz+BXCrEEnpOWem6knl2f5iR7ezxg+VBeSb+h9YwaJRwwCug
FOB3PrcVTkuzn6IVZ3EPhNuFiYoheXpcBUFQ5IAhAAVxxRAPY1bVEPqF968wJwA2x74m1pELaI/0
d92zduDHY2rxog9w2dWkZjU+Qsv8RJXXsdsZUJZGtlIukWjQ5Ti+QI8nr4AP+1KuSCY5T8mv83Vo
4FnNMfYwdJW4IQc2V5PbB4DcBKTaL9GDeSRP5QrDHolsideTaooFgQYLO5wjdKsyopH1OjKxaYWe
9hGefHysA3TIOLdzzlegkyREZD7QZ1aiAx9NnPQ1EJVTwQrBHt9GdMoJG/zayXtJ/59B4+rQJVf2
VBN1WkurtE6HJL3DrPUu4wZo9N38kd8LttjwmNDsiVsd86IumpNUlSmq+UOr6hy8mVYRq8ChCP9V
7eFH0RPrLyP0myFJ0JmHm9M7BmMbHMg0AqDKtzroU2FJkn7RgC93o2+IoOU4lZiOz14m1XcMSK1O
7UwoUdlhMaKzn4/IRmCqpxOullK0gKV5+Er/Rhcy7239tSCdV9IZ1fEqPLivZgdCL4kUsp+hes08
Z1rvFO9tfBE4H4z1OlL7RrrQORPKEAMgsLhaj4FYIK/+ZNaGTHi3IX1L8rBM9oxflNN4yKxc7lYf
i+5lc05ILdA3DepatJnmb7EsXk0yiD5U7XPK2oiuMsEqs2QAvoCW1JgMuJ0WHD/8eGJ4jU0bGQNw
pka1WeOB+MxHKCU3lzQB1vC3CjVUiJbd47mBnqYONx6UmTfG66uPjSC1bx5g74p9RU48Kf/nPfhd
oYcEjYgfByPtJ9xejeZsnXCppl4JBMnKaP3esPfk/uvPTxGVI/gLPvTL/gbLRb51xSbPuIZsuOLt
Tlylv8XpsOE0yDSGMumIELRrH5vyrUYikC9BO8+lmwVdcjQFUHMi/Mes0zGUccBnuO0/uoczz2Sw
U3y89aGcV1h894Wjhio7reuUJeKPZ3fTn1rwFVP0+NgVagSN4RCcyqEj23oxwX46ZlicRiWQRjm9
0Z23nDok16uJGVtFEIytxQbSw0MIMp3Ykb00xxJrexQqiCXABZ4R7jGvVnBhUQmF9/mVLzHqr6pu
rKVOlnhVqIraNbWidyzBqc4vHoovY2W4msuHD6B1q6I/dlsewmx1HlFigMz3s9IvmtkzF0vOZCGB
bUO4m1bZ4HK4VOB7po18nm10TFcPksL4dvXixAh5H9/3NEGVxgsWDXtGC4GvXmkIxo5KFm/GNf+Y
w5gE3O3TKuERYcm7jX/JEmhXX36j1j8IArGQ3EcxyuAA499WpI0lzQIEGfvVwTao4mhpUfTu3RtW
OZEMTc/nv931F6MHWufcEo+2W8auXoaB5iknSPhM4r/ITjMXJBYOApJ+/6iuFHuVDJ59EeEiqk9I
Ru+a3392INZGflxVt+jEmXJywh8cQEi3Guig/CpBztXfRYw5LFRYbvWT2y1AMdoEFE+LMtVLVKZc
wF8tnJTmJ+Z5fRoXW1K5mISksdtXet0cUN0h/21qA2o52RtCKIqOetdkvAqMlRyGVdG98tbadbAx
RCt2fVrnGAoiUmR6H71phC+5CXx74UcrESpHT3eyf/709Smf0S1T75kBsiQsRNC2bAMmvP+QCAvI
8OaHft11XJCawwqp4uItWICjHSfIJZH1qVFvh0VCx5quhMSshfD/w/0W3zrofHrmxrHur83+Mc49
VpEE8o3CaG8mviJxvYMc7OvXi+eSUJbbaZaA5jLRldHOdfzhiYCvyMKJdcyzrRle5exrNTGKtdVZ
jy/NkEUtoceJ6tox7Orre2uSZRXj43lJTqGKe62wOrNDmp0wiyBhk97I/rUx5QfRjihWuNz+RLFV
R0AaB8sTrelGoPugqdwe4Jp/7HQF0yjaTtsTdTf0/ALaYol+km8p8wJTsBOHXujz+S66eSqpZunD
Zoik+M4IpSdMXOZcUi5L/aXvA3uBdnu8Z4bcabU23fegLF0nbwRCPd2AyDG/1IRoGNO/WrCLhQxP
2fsKVL61b0q6aQCR2w0rfE2NCypBWaYc2i+jWusB1/WjsLGzLutSKK+mkmf7EKFI3RXWIYI6GKtz
HgQA+nxYUWHHKsro8X+SKPvdjNcrFzSB3+3MWLYgmw5N0UezlM6ToxqJUdWc3OM5m9ctGhLndMcs
dLzY+6VU2LOiO/NunvwcIru6faDraPh5XhWOgvaT2AfN02ZYLWJEv4XWV9YF6QDJX1V8g5DU9SoN
M24GC2hKlVeWv8G193WIBse0lM43mLpHX4IIbnour8Z+9sg85xwljrb6ugaqZ886/bNd7b0J/xnu
ZOWi0bu2cVxDSEVpG3bCzJLUqXR2SVQ0l5NRMyFgovEjDVxaucB8dOi4CTtd0rgI4qe+Dyp2HkdR
eup9cXWDySNrdxtSwGKq9bWA0FtGvOL57pjnwr6KsVJB3Me4VxsMaNnR8cwSddjuGej0fvuImhuf
0rBXIoxK2AGanO/NbeSnpc6PHpNTB82VL8pNRinH+TZ21j8781nZyM/bvHywNJZxFMF/CQaj4Cav
U4PMW1zyZkzmB1IfV7P4VwqEZznarhBeafomDRNbeXjXKB52FpqXPhqaGKonWw9GdEKX2iiamM7d
tKlBMr3zY1cQapzR6HKLFc/6pyMR/lNoRWbJRrDCFX68ODOunXAKTIX97kr7Yz9lAB3JGBzN6DVo
FGeJWeI14keTj94F21BiRfsnEOTGOrHFAvK5UmK6/bCq/fWHvc/bmp/ZDIMMjU8GoklMMjXke8xb
0iRg4Gvf7C7WtiXVxLkzGRMYGI90tYHAoqqVj/n/CSMXsX337YamQXbdzZHq4RxVgUFgywIH2vIn
69lslZR6tYOqKUGOApL2vOzdh0fvva0N29PJf0fsR+maO1W4Ku2v/USX+adkzdjfL1BpKsKrU471
1AtcVqq8fyLX+gjXV6nM82jt/rkDpMpPnORTh1mpOurumigoSalTRSFfjrdte1DGKEVeHCziWRdP
gwwzAl73kcBckaQZs0D8qBw8gFAcl8ebj1MbxuB8MpKZONIatQLhMkNfy+mZ4308VFGt0ZVvf25d
VlxPVabqkFWBSRdlIovPpmhxbeoFuh5ePTPBpMYu1y1EaYJ8p25G3I9ERr0lHnh3gw443Oi34Ku9
xmklS4UZQSkomeLI39xzS9ziJQ1i2eSv05UOxacJ2TZgOMzp/kJqnRlIvmPiGI7JK4qGBmCvb2wL
o1r0yeF/FqB/7d+zGgUnY7FjoCHhX1aAplGx6iYRq4nHTwOQortcWORo91z0EYczRuGrhiBA1GzQ
L9FE3EAyi+1AWlKKPJs9VnIMihUAMwmsk2b4GUeyGmmWqaOYbj1+ygbRXtV/tf+htempMhhFP/Al
Ry25NWzWZulRR4aSeSkIbKWm9iV/5jSkzqaV54xGzXB0VXnIz2TcWlUqzn5s/706FyDU8GTuGFH4
AKtFrtUQWVuyD5/7lvRorFiB8wj6U5pUdEqZeo0X6rEsxA+UoK0f5KPpRJy7ANuJJVnQBxuBSNy9
6v5o5HkrBq1OLvB3+22BSmeRtHPwKRilcLNuC0N7j7N7O1WRrQ62E3IvIk0NdnK26xAnRkSNFgC/
Vd53sBCNyjIryeJlwLtDnhbdKipCQVEYbzlRg05Y0Jatij59ThjKylBrAbmnsqmUFykT9vB7bk0f
A519uqQxlnTxrPhZVCp2D9BI4p5GAgZ9mp10l8XQnD5GNdvIGl4L1dacRqa19EgzsaR2cikZ0Jnt
xY+m5ARjN76FF0XzLmx4Xqb6nQH5bHGp1WeuIlVIEU0xcppcE7TnxRQgFrx7lPEthySNwzFKHwDF
MmUrsvWDwEOD4cT/LxQQL5JB8DqCikg1R3pdE6Apm7L/z0uzc3RAmAo8xQUcfUrfIPlL9anHOvHS
X56q3c+FRv7rpI/Ek8zHXYJq+IQ5RthrcDflbcR0MfHhBwewniG+STFTMVMrTk5VZSyi7LfARoiB
ijXzXx6iHNuqmZhwwVX3YWAexKlS/8/SfJ1M20NOWrtkEiGLIAm+J7NjXxNwSFv3xpK6Cw6PRkMS
Mq0JWQ/z0hYN3EUXt5LOdO9leprxa+VyULL9Kienw3xhvuNRH0lWcpHVjKAvKOBbawQYMilllLIO
Jxz4bne7nMXcGir9++mybLTmM5/m6RLcEkKQpdu/SbPpHpERDI3xMZqcVZXynvfLxEWa50Oi3ndq
A6WNXo8kH1r2XEhoz4Zo5hHkXQ/cf9BWA7Rx9+ywSQVEg01IB7sFBqVCXfQFkL7WLrNpKVrs4EhH
CIANn9chu4wA8PiAX2BPls31D9H+OwMN7qZirJNZTSn42+Nn4/0nfyaDthI/PD94SGmxkm9G/y9F
mZ7lKB5pouKBI3g10vvnm3V3KEosfle6tNyDhL96GInJ5nLVj1ZlSqYibxrUFzogYkSKD/H+HVvk
t9mdaNE/HGPXib3/KRYbg20UQKCWN+4dXv/Id1ef7Q7CGNLw9v9yX7hBWRXPKOhxW1yiccJ3D3/k
92XJkV5brnMrgwW8RpOdCjjD/uU6dNSEJG31nz7DEwM/JkhInmWQTAoYuYmYDJ0Kj+XUkaUtIGwg
ObO6sKj7rTjrv6UKU/Y1tPEzdnwdjh0V/YFuyGmDzZcDR3km/CCoKtdkpuZyppF2pRfhPzxZqJqc
xDgwkKJU/fNxsEKkHzH5ez56B1F9SEqYy1cST5e1pQGmo3SCGIB5ajZp2PGcoydC43lRq9SNnGOF
lj56HUAXPhTU2iyTYUugBZtBM4J2cgVkiP6ZQUa6VtEgM0jvzyBw8FTBs/VNJpwoHgcRF07VG5wn
RTLKe+hhwi4HLShALLYtvAWFr9TVuZHKe5ZeJw08hxIeK/Cm6QUC67LS923lGNgQo34iS2+pn4d0
ngPGoBT2gbW6bkiv14ix3MxF80wQuk+3ztsGpfYIGCj+T1jxzBBss/6T9g6MEgY9/lSrB1O6FeGn
Phy9HgXpJY0byzLjg9h9KpfotC1qwN44sAbUlXZ64UBQ1kv6/YwxnjmNulupv0i2oOQWVLi0f+Pz
LBYEt+ENMSVKVP/7170JAbjwSHUBohR8eqGiGlxoJeTkOrk9EqGxVMgxS7p7B9XGXRIvuvYP+wek
eEmmMmhXwohMW8f4JqAKp8W16TM7mgaEu9R8EGNjkwPBx6G6Y/65uuhYkw9ceKCkfhEBaKGevE8I
zkVxLpQvMnGip9ll2bvk1CrNxhx5GGunLkgxFQEfjGx4ifm3kjVolFV7KPsad9Q1zJztcLmhi+k5
3ihct9iG2ZRi17fVFcxl74lyvovkDpi3kyHN3w71Imq314ArOJEghFJBG5gFpjsrpyy2HOIkgPXD
uC0+5sJHGPCQ2NOureQuWOuGtwORKG9bT/Pn6YMJMqjHrpq+p1XijUVT7Es4KxwNUy0grV4mC8ns
2xBTkLMUx0zQaPDfAxwkNYLm73SetCa+V3vMl6gfli04AtTXZvrTggmIjahajYRE98A0hagY7eBQ
1yLbfwTx9NVrubdmn6nAYs6QcPJy+a/+3a8gfxc2QxSPDFLq0JPB38cvkzBanVhUcha3kTYdvwBU
PfcBnaw6gbXzT/mSHm2PgYJYrZ2frR32DKGO1QhocIW2+zy77t8bGPZ9XVor+YC9cJdyw0+ewRMM
g1s/vcIvxfxEppEQjJG3sX1zcfCt8EamScf6rWXiKNrCU5D3GUIk7vwmG2vMf6CYC+1+vEN3qe3Y
gxd0T6wNvGCggy2ZML2MflkyhdwDgHWP3vifZBTRf+lmVJvbuwtzaRxfKfG5BLMBfAj9q709o4tz
jJU3kkhFKwtoNs71yqu46VYLVnAbvq/ZR52EpM5AfR8TOAWdMa0t8BnnL5GgcUGIkfn0Yey5DJiI
XeOUUNcmKrXat7dMWapGOAlF4AUJnLo/aKiVdSWYrHxfp5YVI5MYrtE/WftBT/ZNwsIA2pN8YQRa
JkvdBnnsRPoWeCm0wks34P0dVHP4kGnYvQ7HMqBhA7pbJr3SSmbZbf6xsNC2LwnOcE08FfAIF8DS
i8GwdHrBCnne66u+hsR/S0udA+XBiXXe883XiHPozldjUg6a48WeILcJFilMphuER3IqVXpwBTej
1f3IgYN7IbGOGyQFDalScb1tHYUhhIgj7VkpgYL4Ru1/ndnScXtJGU5vp0Z+sDTIo1W2AxOC1MH5
/9OAjYITXzVG+sYsaRZb16aDUkfuaO3w77myYBTCawqSNFmb+iA5PH24OSxNUNMEVl5FLKNa4Ayd
t7fiDxRZxVA/M+C7krSD3UxmdRcV0n698rqLfOMOBkeWhwWZ6d9lrGQBcjuAdWUU/hzXvdYeECqz
DCZrL+Tfis69mg35wI2k+dnxEywNfqNQb0ONekV/1lLxjV7sPz6zTqCtApQl8dsDR815x9k+BjDp
7XhKUfCG/2ij3jrDnzqH6uifKdus9AF9JicloJ5/2iJIff1YYRNdFJx/Yrz+gjKFvBkFqerw5SpO
SEqfRs3cSsiGrFpGHLH51LGzT6zFv498n+GfVHny19+waDpCTMFrl9CzbJ8HIX62Bh7SuH1zeeYV
4Kxk04Gh+fBPM+Af8XNSaTbRU7ZZDgPio6weBuVekkhp5rWP6UCbzcG63D9sfVBTmds6UeCZuxgL
Xz0Z26VP95Wd5URKQk+YDTIkXb+DEJ6VduRqyo+TZou5Xz027dwke7ODcXJjKzK8cDBhELEOq/VM
wt/PceEoitwamAp454tMvSJx/Dn9P8GnGVecmTDVMdZwTTbbPXXCIWfUNOzdhCfhwUIBC3Xow7sb
WRXhUyBZ+IYVwAAmoPusWe2Fy9+FI8gOlSIhJTKHc69D1yJm0YqkbOay5xis9EYQZ7tfy8d7X25C
j8ozfs8y0TYEQK4HBD+21vjPrMvLO5dWHRpjCcfbKaqkZuqWrTTQprgf4hwJimLFBIsZ26G3/VL1
nTDLnSID3cudzXfJYnUk++4P/tyvoXpckJ5Q3qIvGGPbMcPmTKCvM8DtAZO8Ny5aBVZ0XSdcrWPI
MkLdkWetaKvEyHm77J3SJQ6nOeWT/V1WP6Qz9/jtG3bUmGm8iPuJU0sVT1JRn6AaRJsKICs+l5JM
fp+AyfAljwlDfgHLJudJNqfHacfAsm5ekkqsRxINo0jir2BiQxgjPyKqim3S4/cQFatejf/443jS
rCVbxq4XAM5N1OeEcoMe52c3OJ//BhiRa47ufyyiOwvPcvbqSlKPzt+7L9dXZQi1fqSkfAo3LHXd
hds2dm87E+T1M7Ed9UZvRTlsjou/NqnPIgUegU5+z+2xfDcJGHHw7f8GOIUsnvt5kAGoCUPUbt8h
XpOYfVw1XHBcyEl3D6Kwzvp9nijpS4sNVUlJpTuHz/1T8hl8ofAl/bMnLV74QQJTkedG4+Mk9/Z1
sfgItpecDlczE//RrTavR2iC2aa0TCOsY7veFQTe7GiGSiAg4tGbIR0lFe7oQ4afTL0X60PvkR2Z
xPhKkacR9EpFIurzJjEuZey/XOw+0IoOhUS5iCSnZTc0IlALWP2Vqhgdlv22i3qHKz1nPAVs0uzS
dzi9wR878e5MPTFCZUhxw8f1jbWCpjxOJeDE8zweQwQeQqQ3e+peyxNdfN/owKLY+29u+OSlROET
XqU0dJZSZjMfu7PViznp9V8wOEWZaQYfjGSybiS/tD1usoIM3sC+AbvxT+P/bbr6EM6F7mbbzLye
KGbLyxscEtwgJvncgaSr0nIsEsEmx+jirkr+whBDoRhTwdLlvfZTGididJG1j+tzYGjKcVIrhmAs
iKrGapkPpBv6jTYn1QvjWbCi46vScbxzXGTekt7S5BkuYvjZsDLrppKgYdCbtoQiqvhAwb3dafjy
psdINo4nkplO4n3HTyEl1mO8P3ySFWd720LQEa32ZtJ50yeBRcpmDIPNTk6Nj+x0HKzFZ+Iy04Ui
qPOSw+IU5qrcH+Cs1LZUe4jRf2brsfgsQrdfkFS8QR54NREbvkMoXXgSm+CZEOeuMGpLHunaQBOe
SHQ1U5h2tJ5RIOTbMmdf808D/qhvlk4sXbz07ShAZ+9AgeLRGyIHxr1m9vORwSC0BsMxjCMXuken
SPMWWVDEdudKI7be+611sSdTEYXXgk2k78/AxvK6EcT7zv539QvSsVjdhqYh0iUU+fjhy8dM2qbr
K/TaXYxynCYM16xGt4lOTrR/Jv+Nxdcve+h66ZO5XpgFbNiPB9WYnvmDkTXKqBdCFhF83Jt2lG0a
3e8lBw9UhvBKcV14EFVjHHJWVylXbduLZEg7yp59+nkYVgaf6VC2U07p4K5eYaHKkv2hfA8BaEvU
JEItDmPXkvguyMcl/GxeqS5ZAHqQwI4b3QrNS94URi8/X6xK5z3O+qOZevYS1Mz4ZOQkJHTR1Ifu
G2J+YdGlgsurlb5pMVPAISNNpu5wMY0EVtWSEdIM2Cu8viBkNowm3aX/C5BG9RiQadePLUy+VaE5
+wN9vH6oFFM0SIrombNRAhISIAjPxbIoCD5X5DpdsO42ldcitXIiRKASK6qFhWXJD/qBLjHBS4lp
uVaDv9T8xlLAkpfnJj05XdLjg2G6YuWn36Lr1BP7FPZGVpxfOWIDW7gn7gdJ1KaIOOIZ8QHVSKfg
a6TcDS5Rizst4uibWLpM7a67DtWZB0oHcPRWakDYWMiAh6+HKks5kAIYLUJOL1c0mxtPkPKLKfYU
Fj4GVsuus39tfkwrMw1XYp43Y+pgv1nzJvc4WdREtZAA4PHdQvtB9tsP/1ZSTHz60UhSmgQirmOs
fVr/UCi1BUT0xEgmPa9z8jXDZl9bP4R+yJdIxbDPYqXjFDLGGX2VE7g71YTM8Y4a2E6ErBNbqLRf
Hutx06aJQ1wCkfZgJHhn12DMrud13nGCScRxK0teXXwzQUaiU3zSj4eCYf6zLUmCurzvbysoHdfe
EmliMf9v4BrHjzCr9fl62hoAaWwVQ6QksJm9AX2gUpVX16nOFvgi9gBW9VQmqmvlfpNYhN9etp6T
3P5q3ffZltPj+V97wc0hOkSMuXnSK2T7aMuIhb6q5fnNcinl0glJAHkO2ohyb8ulEtguOQyMbFFN
5mVpR3hDJRpeiYZdPe85TM6cdZ8rEcUIdj0U1kcjjC/OOXlqYeShReu6DiYy6lNW2wwwqQTwDlwl
a2/0H4EY6JXiBcGJ6HVyDzabzq+Zo6KdpI/fJNlAgSv9AyUFQf5OIjXIiAASeTXOzWdO7kaOcmMT
AlKdzcvKIb+NyD7ifUeujGpt5hPQqARpvNqur7NXt7MZMwoNmN6sGVnfSi0AcAvKlTPY1JYwjUj0
4MNhzce5hJ4QUnjyrLIKOPgfgHsKYs4kCZyaJVdwqKnM0stxrzS7H5eyYjS26EnhveP4OFPHwXu8
JQXB2/2Y1yBp6W4QYyiPk0taVRl4R9sHt/0Q9F3ACINZ61o86MbEqOQq/WsoStt9aFj6jj7wioJM
UCwanjuLDwqbfQtfaXkPkBG1jbcKs3Uc1PTbmEa4AeKBavhUjhVDr1HTuVrmaJXzGv34dTbXd+rO
HzO0qQ2eM0g0CFagjgtq9mUivOBPaadfp8kanK2u7Istni7V1nfl7SZ+OuEAzudKX56VN0UBPLK6
lgqHW7VkTZVsHPgDPC81hOjdJiZAzCPw85sOddwxDIbmDWcPN+prYTbPLkabTQ4/Vt47YlaE7kxZ
YpoxgdzzBS85J1LceGbiFVHSg3+wZ4kQJb14OujAxd7KIQ0Li5cOscVUr9OO0KDHfC40VvQ1fQfz
68bGL//pfL8Ztb7iIX35bWILpD8UKKaGqqVs2w1iw7V8X0NfK3psjLgHq721XORgHqiayYxPWnuD
8PAvSiHfvG1qy0+gHT6v6lWAG4Nia5U+P9KWLyJltG+zXUrkotCnhoZAhbFWr7q3mRsBjWWo8nd8
0j2c06yY5WiqoiVRzGooj071kNFeemICLalm2GZ+yae/fALhAJFaFjjmPFMmtJoVD2Yjq16Cf8TC
AH15LCbCrlMOfN8gxdrJOaJeg3sRnFFqLtllPXdkRpN+fX7Qh8JHH0/OTjAEHBDUXO4F65C/8or/
dRo0nxORN9xGod1ZMYJj1EC9PvJEzy0DgDPJoZr4OCgJAUX1VZbJsI1clMGjGOFkxucfiKpxcZZ9
fy5WIKQth1GW0a+dz6BkxdEdPCtCrFbYToa0g2UJ8hIpbBfk5Ni6wsvOoWot0cVZJ2EVSFSQQ+ES
19CTBrC1CajNVYDRPVeIgX6IE1+XyYaWnlrbPx+CHlPJG4BRyl5kDkc9v/et1lyI945/D5PzwJq1
7Qthf8/c0vB1aigV0LMF3f1U2LR1RGGDHbFo8PJofkjgIgPiHAZv7ZjqVRRXS/jvS6BygiUdsCAv
QERi/ZGWctF9xOD+Y01vRhEZOcyYWaEol7c0j91FpmtlZSt6SfOdd+BVI8WpFVgad8bFv0apYCvL
TmXIQg2LNeQLy1Z7kNEz7EDoa5omdKXRjzRuxFt5xUPEAh9V0ikrvcDbs9yNKmagpYl+oXvu17xj
9vN3DUjXHf6VJJTbe2IZJhKiz/aPUTBoK/3QxeWIlNoX72lgGWXOtFNob9Frj5CnCHnFM4j58DB3
62nYT8cHthKfmNsWG6vdfvumDOO5h/iWs0Yujz3e4eoF3WkKNabiE2QjS3kTuW/qvN6fjS75x52l
QwTY+irvedyWZLbhye+iJSzvtt7Mc9gHJ4S+Ps0II9FVQ178KHOTtHR+iAcYO4nd8WKm2R4F5wRN
93oc9SSp6mnb8ey/QADlSBUYCzSI4/pM3BpgVR1ffW3TGrs0SjDS824SFeXgx22e5K3lQmh2Neet
u3NBlvyBPGdXzKXK1QxkBdqC5vY2gyOaCynqgJqhALLmBOqpUgkviVABQ5oXRtGvmRuA9HOGMzY8
2xO6RHiT+exwpzX7YLT1WitinkG7jW5hbRz2xNGogO8U2NMeta+sDRyop48+LlcJxHLyeOllTZsv
dHJ9nlkwCj/sA/KDhITlP1I6+/SbXFUSrdBYUN8QcppHukaFV4Vyoj9IyFVUZCijl/y0Ij0C58si
eAOTSwL3gPz/8T/5UDvnw1slMrD2uBkcU2G+IOdT0LUWLcuAKLM15iN0cZLde5d/K1ooDFwRjIV9
55a4NKnluHUW4e02IozdBmPd+Lkdyb1XSa8y01+Hg3xi5Ivx1dN0i0ZpWBGCq9baljdOTuo2BtlG
kZ9HHpLcIAG+gUCi1/i1gxO20y/M4UN05fcJ0HxzRbEQsvbny2omrlr52RIAnA5FRI0Qmxm8KNqE
q3DPzH7sC8f0uM0gQ69jXJFB+QJKnVN9tctrXP67gUnoE7/XAx/lT1xUJQgTM7SxvHYoqbqORnqk
otV9R15X+VXINMl0uuGewrBRV3H6o2ySgQf4FBO2UOS8WRsF2SN8fqHUu5AAk2s26pIUxL9MXm4n
/3flDZDM8q6wC6N5nuifjFAZzJ7RUbZYZxc5aPkjzbnIbNB2OmvN/OAN/vGZSn+r52xM7m5Uzy1p
DmhxUN05cWvxos62sp8+jh6BG4xTx3egHDGbZtqjTodO8hz3uo2nTh2EZnoD2F5nsrOWXp9kuCVV
WuwUMHQEIJDk7jElbno2OoZW9Onu4khIf2fTcJNEGHvlCvuCNhtHbU20Gi46mJ1zxnNwBo7SS5LS
krJ3Bol9qvqx2WnR8EizujVjYZEbgi8C5rDNYr4vzu80xe0chxlwMwckBucx2t3JwwuYzHA80sLI
1e8tLrDKXh63qh241IPoTK4Wj0mTpLmjwdJgyYyyJZB9+Btgsjo1qsBrKUIKf9IwIbWopINJjyQ1
8G6joVO87abbSX9Jomjzu8P8pZ0HubmlA1LkdlVkgLJ5m6EhbsetaU5Edt85SYBrZ1bV/YnY7DCL
Koa3bHxMmnwRXzOU+tsLhDWbx/o3UWf0L78s5Ds8T2p4YMH2wx2TOsAU5a/7Zv0Q4HfIDBzKRaqv
Yz7BRFTZSRA+5lFeMLXHS2A62UsdHvprstEn84Mq2vmx2FVmMKpEnWht54X56X+LV9Ys1bnfA9Iz
gQDKaDbTzXbxMCeQLBKcQlldVdTsFOs8YweoeeXC78/d9T+ku80Bdbm3FA98uduIW47F1drYmbbq
iZE76UL35H0ZyCG4MPk1YzfHe26LJY0Fwf1KQHCSVC28i7xPupW5fAajc+pKDWUjZDtK+poWsW9b
6DCW1mqRXyEnRBc1zt3Wxd6nTabU5sIy3090zoLfP43Tk3Ayx39GIxFmClI9U3XJSOZ/A4eAUjli
rYuOae6IEh+onTQPesTmlnMu5yABtGdVREnJz5fVFhAIHPHf4mfaEZlluvCvenpHTLqQARB6UKgv
SErovX0FNmMcfLyMHKT6leAjqHKX/43VeP7J3EBQ+SVy8bzHJf/5BOcxQhtaeWrjHKjXY8CH8Nry
LkoH+Igoik2hCnV2o3DpHlzFAkvro4aIZR950GHJUNYfIZTf/99NgR9xkSl9FX/+GlhXPxNCX2ii
QaKWbndrhCp1XfYv8I+DL2XPbobyrZr1GkESP+omdl1mDgUjxFJbjU3hxlyBBm6vuZde/sC5yz5v
yP1Af24fxnmhhNz3SBzl0RvXnRKmW4vNOFCyQQveZOmaDs7HrO/s/5A3nvZ8DZO1IItA4WHOgmLM
GnALPgRQjpOeQXYTyytR74qx/wXaF7tUqlKDOSWVRAtpcBFkSaZ75B84JSubIhi5cRUux+Q0BrdS
ER8kf9AXFyUmK1KudORdWHjtfMxdVLC6mZLGHOppKgXWRFdcGJbs1gtL4uy2nwIyx0cd6AFR3Dzt
WRl/dB318aYSEvKkIiRJH1qC2H1dVbHyHSY7cu+wgOTwH5Per4towKhkDPMmKRRKhJGd2g5tRntC
cQFE79w3b7Akf6989joJ0NyKH0LUHVBVhC19s8xqWJ0SUiVwZFDByudRBdyP4PB6Mcwm7ym7B4JG
8HlIxyu1FvQ920iOfKifcu75OFIIJtAsVXLQUwjWgraIFsdQRizJwWsHzj/GZIuN3gk3QZAdVqaA
eTKYpvESoHogFkxRTHc4Qf/dWZklmaQRC69rKLtEoDXceKIH2vFoSxSMfwq8oQy7cFHC2VvlUliu
EdqbaupJ4vAOViJne8L2AcfJvxNLmxhgrW5U+CB20kC0TVojUAYvSDSRU/yrjnA7Yb4t9cERtWM1
QqFIpcyqnoGVhKPS9GNnx85G2YuqqP0hW3w2W0EWgP7J3y972A4QuDWKWVs7T+XrJbKD5ajd0bJW
n/HP90yA8y3JqfP4CBuNq6bX42IGtUM3WP7qOD3HapCNi8bode0GW2LQVKZi6sty/nwkhK7/8sDB
MjOXi0R9himboxggxowIrt6c1LH2dHvTLMP/LfMNmnpxcxHjVK+6zBh8SAl4nwY8BtaLifZsVFnW
g60BwDQVunvYGf2xd3v23AgdW7BT9jpDSW/CMqy5/QMycyC0xjvGiiO14tbVd6XQnSC7H/aMahj/
yNumr9JUn0JTR2+E5d2RmcfRLCaCLJoqF8O4Tu8OFc8vCsV5LGvMZ+dWtBmiSYzss3QK1X49x2YT
B8JXf4XTiYig/k4r7Ox8ajnFhI6zqByMi6deSrRBYj0AlJOQjbnwEqPSzWmaqrDrRWf48QYviXOd
EJi5jffVRx6K+869Eaz65DoxkCsn98MygZ6gORVA3zM9Z5gEPE+hp1O60s+43qe9pffeQoQ1HL6o
C7I9PMta4iLcKJ0aEH8xsT8jWIJ5eT9kFHWCbE935gvVv+FHWnqvdh3SocoAdDcjNzFwvR+JDDFW
k9rARBIzn0b/H/YDm9siaMvKPrmYu7LEZm966UVki7gsj/N6/7aHCZWFwylE4yQpS+VpBDIWNJ/n
U82+K2R7R84uS7ufOHrFvMOGDnABm3NXASvSBV9p5i4Gk7WgrTLAaLHNlVk7No95+gx3DkvXJeJR
fLlHnjsxwxBmduLhtvxBYX+tsTZRW4zo7GjilFY4kqXI3vQHLu6nF4DwjAwFO0uSoNXCdMW89fLV
fZ1HcVIq13RWXjM3Be0tZVazEGtxSldcVDi9FUAGKAPxSshTDqt9UVmTBXMuvLD9Aol/7n35j/Dh
2HnUXp3Af3RRVQ4uVRtTKu6TGWVLghBrSPi8TQUBsmQVs3ho+fKfTEwLABPW2xrdeA7/Dfphnc1P
QUcou636q/c49LzjP+cvyRl/AwylGMA9ne0w+Q9LWK5ZlMqIL/6e4IlUekd2dNZob7c3FlLwo202
JF1b9SjDD84KmpZCwcJt23Ro3/Ni1W7UGu7Kx81ReFmB63hr/edkHgzDN4UpfkLLFTsmtxw1ZLaE
jmgmq+oN+/vjg8HFyKAkO8L1/joP6YXfvhecyVDqEyO2MRhlWhkzXrRcFVzlvS68l5bJN5L9hYbl
sEE01ZnjwhMZuhs2x0o0KI09yon6N0IThtHInYz3dUi3XIPeE2Xp++HU3iIRCJm1M55353ZdeRTH
5lGJIO+rMNZtL8uyFZrtygeD929mODAZoT/4dFohkGC51vWI4+SHpF8lMI1Y1r/xeRL8qmNHX72b
LnBwKmb0HeklMPeg5PDZXDQRbmmrCdHcaymx0oX3cxXMk5KCRwBS+RHnZCUh3St1kUAPaw6PorMl
slWhtns1v8fKfnmNCu4VETh5BAz5XbiMNt4Sg3Meyu04caA5jUPC12E0eshEryZYwMPsHdFga9FQ
zuPsL5MgYuc35RGemubiS7Z+A8Swhp0majF8wc2bvV9NUNeRq5vdtkkYJyJS2D3pnIbb/5q5aPkR
4MDy+MKzugU2HSLBStT8fubgmQ3wtkVs4o6IG/s7zik9WaqZPXTCYkOTxYNMdv/n/Ww9JOUsA2o/
Sg9Mm0Fc8iZgpvnvZWmkrieWRQfl15iyt/j9ewJXziOvoPBydbPimiPvBHvPfOzwlxAC8OcQ+ORw
gN2C8g7PMHRJn+Ikn3ZX+kiIfSDyRwRjHHUaCl9RPpd1tKmupQlukqBJxBi8zFs4en/Apvl3LLm0
g5pujnnILgeaCJB+v0qGC0hwgLc0VGVjjKgjqC3aTj3sPxoL3oIsDV6e7gSgRYTQRkCGQKkQ+pQo
F12Oyb5P3+KjgLrHCVKXBlqb7n5U7+j/udRYZ0d9OsWFTX+qTkTraUlSyxhkJ9iafheYWd1M3yUv
nNT/kpawpcoKVB6lsz+BaLMXb1VUmX7c0eQ4H9WjU2P5iRnhmHqi+ep7ZTA25SkiWV4PINgPJgDY
p9xsIS3QB2JmnvS+IROSPgHsgMTvQASQsA4AXp/X3NtbHyJD+3kTaA0SWwF+CB630AZZeWrHxanY
kYMIFoIBC+S+gDnedkhPO9p/jToyz4ZxJBiRw5Znc5MVoLB5uV9ypeXPKqYW2v8+cXCycUYGGEP0
cNNgrPZVfVk3gkVkvhXH4Bk+LggFQdqUApM5vaerI8fT+NqBUZwgmi2c4BhktIQbhDDntHm8a1Wo
E8Z42OuhGGi5aaIr/IkIXJtiwT5myg7sJRSkZuMdCCh3NPtQphMRlxohR41BQ0jT/y5MM6n/dY6C
KoYd1k1hxJHCzMjinremWxMxNzTOv/MTQ0vWHKI2tgGSr4NdcbKxxJ8UyxRpLspQmB88tO6nIai2
3q8/ihaUPANVP5UT1kqWWqx6ZmvXT9OxmXjQgq7vjZyTmkDnhtqf3pgCUj0bV4cBksm2w9aNDKFu
LvJn0/7LaR18kBtLKNfGkIl+S6LhIOSCAGZmvPwajXXq6930azENrQrHzgcOpTn/R399JLp63Hk8
1kbt8Bf2fFxz2GCIRtUmwW6978kc8zIJSeX6/Zsu3oFzimcFBr5evANg3UaQYYMyR85hLLbGV2nk
uHA6p135I5261ceP3tXCa1Eo0FUgIHsCJkSvQmZdlYx6HGYoamZXg0WU5p7ufHWTo6fvPyqv0fVB
BZMSKXxB6nXCkfRkZq2c/o0tFHHYeGdtj1LadKlAs+kPhR+c1acEoUgS2216dxsgXY6IiJBO9aVR
uhtqRilW6y7Hik1xsuz0Lb+bm5K2zKpv4nGgfO7bMlHLvdgp/pNY43c+YjO6chNYNNGpgramAcbO
uMFjLHkGc7v6aiiV5Gtt83XPqCxnV056z4fFciqgmzWu0nZlYZKgLGV4VysbQyOK4MuYBQJkr1e4
qgZjEKLc6GZLxHNEQVeY2j3jTQelrVFpgfxjNVsMkd0U1Dx5k8ZbbxBh9q/OGBsj4lFUeDBDg+do
8VtBHNym4xpVH0Vtq5MMqZMY4eBERejJmkBdb1dIETAu21AgFQ5rtwZMzRSEWbY+W4OeFZjWuycy
bgnGt6CUcyTeydIf1dMFRiM/5e0uYdDGJNbOkP6C0LSK5vkN7JEYjHqofmvLIROYURzwARCMzp1z
+iI4C5r6acJxMMfwuV9n3B4auradMsL4hdCopumnelk/AK0HmCQJUCihpf34MPOBeEWvBrhN8cWi
cw6+cDYvXZiysTHvJzNsCq6iWirBX0WB41YBFxhzFq4QJKu7DHv/UVcTmAIVsk0Cc6YWZHeTMC2v
sCKhtufyjkL2nlKU6JbuYVotS5CPq36of5oLyeHlw5SauN4suwqEOUkJXdTi2Q9uMpPYOaXGpHzS
1n6fvjse/GfJ8aEgrU/NAfprlD9knWGOq6IBRdHtnhTmjtYqPf2qBqLpZWvszql/XIPwxjuIbLNA
J2sRLAanje3nNyoLv09nz09ClrD6bBNBHLosG6W8OKXxw5HR6enRipBriW/+HztPezUgKzCyzRRl
iBRiQB4DkMl/KoigqwxGOrOD6Wz9WSQAWUx5U6wj4M68mOBcYpFu9pK3onaxG3w5e1rR/ByQRrsg
5FFJVEfvuJqpGBo9waf5s/tgq/eV5GSDdG3NRFtzSaigCoVGK6D7RiN9qD8MiAoxCEwCeB7EuvlA
XDMr3shoRfOIi/r+Fj19QtrY83ZDF5Inl6jlOxBtG6OfgjSYPehcAM7BwyGmz569gJ4n7f94mXQ0
W+nZNvLVIQN7urCiCzHPDUN+XwUdlqzQL/Ex2d6v5ROhy29hsD8+I34NxsOhENI3PJ8HYJ3jOf6j
X5oadnmd6ut0nDLc+3cNxL7Ets6JzIgTUuw1KbDk4jQIiDPeFwjdw/n9NpnA8Hy0Z6PsZPaSPl8z
4htLTjMiNom9n/QL9RN3d94fs8NGBQQOp+dHe9arlbLnJCvUJ1B8qEmWwXU9RpegATOI+8bgAYLl
IdDKqjuAcfQfrKdtDRcvQ99EbkdFcwVQWtGRtlA8Y5Gi/kFBiMa6ofTu1kYCVZEM9zaJaM1OVxKy
gWiJcEEKzXgrYVKCXDjgstxBBl5g5D8pvyvBqEncLgneGsVQGMkAf3feosnJzwm1eYos6wiC7WbP
nGDCScduBEjYOIF3veaHXSrgr2D6Ehy+AyDXpb/TyIYZeHdY8LYiv3sMuu1mQrIdgRZsaiHElixp
/DQiNdeakU1STOzz8Pz4ZABAafVuQmE7ZoxRAgbQD8TL3/gDD9siDchwTR1+QadUFx/a1kc4A+tM
DUhWFMMDupqqBXuqsrAStp0OtAZFsQDVkVDeUZcj2LXtuuju6kUCTp+ZZqgW2Y6d7+45oU0VLrPf
FA7CyANyrJeIY9aWXfadrFWdTNf6wTNGa2c91aHAT/rEdnGQxaWAPuLn9mrPTDpl/6wb/JI3dVx+
MctHYbIx1hSZpjg17uWYx2CBm8KH34czz54Nti5lYU3oJVqQJCpSQoXpcu4K9AOwRypFAdaIcVee
JYaE8Ijob/ycFzXanfiRUbEqidIyNK5mpq1mUHqWx1k/yQxbBgXuTNmrwg1wXEJoI3ZcMZc8y0yS
7xNbG1D3F8Pd990zNguivRr57eRl731HaPJaOAsfmZbDHm1HLAmosUsZnymh27UmEEZkzwCD8gWG
Ni3FcuIeZ5YDZYYnfaAiAMm64ekrPtHurokXkMCpJFlJtk2ol06afwAY70Flhef9fHd/OeYdipsC
DrqYDIf/lQOc85P32v4yAvbdJfkn/lJykZJ9dEgvSNxH5R54NsrZQ6wDbEwKMqaQFYJRoxHYmHmS
rSu1RPgkRC0ul8vdkyz8MRJlBxpmNBVbhDm8WVnK+CU9iLyQYYNh8jA8C9CzhHDoVhjf+ouiKr5s
Ef7YCtSFVktFETCJRA2uim06zzaXgnanLHWiW8hGav5xk8dMDaNKtPeoeL9j50rr+GZkXyqTYtrT
K7xlo2rYIqTmkpSMNAQqKkMpTjBZsTm+qI9aR2E7xt//VFs8qtfFCJOBXNOwzm/tPyg0+Qthgi+b
JYUCW05AhibKPy/hYCKLk72DBCw+nyKSeTm9c4AVvEcM2qUR9u7vx0mRdnrQ/STw2yp69lJZXoga
KWkbT52bkUpL+o8SNCqTDNKv+dD+qKc6q2nFrl9Cx3jUTmzxsQUWBMC3GJ4EJFSqsdhJNBZj2vEy
b5cZO0Y3Tu+U7/JvYJCRBmEqFGrURwKERtgxWdUCowcNnB8Z7s8BiXF13ejH9PY2IC0uKngEhn8v
kRXND00SMdztGvmXQYQKJTqVNeEvDSsNGBcdZ0WSEsFOczhTLZhb61fR/QH+hHoaurRB8xMcDXuX
lYSxKAuow77Di8Go7MZHmHap123lLgHwez0RHpjsFj+2Sf6sKUQIZZCymGgxWHTxM24p2EKcCDl9
A571yzhYijauMfxGxG3/LQqi2X23T4NVWMchD7jcFDDaCDuI4Qux8tbzKKBHszI/gVlwaL8qpCE/
hV5K7Bbvz9uFASPXwFszG08ZcxTczdTjgDA7e3asMqagoCnYF9SwrytzTcN88Sur+KsBdIZleGTr
u2Tp8a6eHb4uv1JlijS/pDK/y8x4urk7Rf/UUS5n2RAAVulSgnlOC5qpqurNCwguXS4Pe4NQdmhp
Efgq3UGwTNDfVUaiR5sdUthevjT6cDnkwPBpBZnh1AAiw+w6uFy8F2AIH52waclItI0u8WkPBhlR
4iXXhdcdloWDTAXlxq6uXdnppKAV06u5pAseB5SKlWL5M2Z6SjMpUks7y2c+uGbbwyQaaWFpV/JW
P9L8/22cgdtcT5nSDr4SAc/fRL8t5uyz2dqegl2XrXLPHO0cb3wnwI/4MYFuDGlMtlTNNZXbHekH
Z3FsMT7o90vjuMmNjNL66QhHyCMKXpSQXlex2nrp7c7bT70xsd5dv7AX1mYaTC1YTKj9elQtKNlT
WRuPTCMO3kuSEmye93LqM5UdvCksJap1oE+cKbQ9Y1qeuU9zlvAB0TAdVZIr+8PfZ6o6RY7Bw172
C42+7pjaqQ+PFoqvmFYoz8pMTvecCWRvt9Y5i5R7EVRSC1xkuZE2wPHGYIO4AAPpdBujOi8QVIjv
y2+1uJUvJu7nFzjdZOZpoJTkUEGUgbC7PL2WlMhrH38314TbfmGdA0zkXC2hB3HW5hfI6G9ca68L
ETC6KkKS6gLkavV28yTda4d9Bjr0HjuFlkb402JoCzfIPmcqgROzvuTw8lSkdtQVrD1Z6xKSs4sy
FIdk7XKtraGgiQA8bYMx5wHATQF03EKtioo4wd7u9HRe+Hlj9SgzbQsyQV4NmBC1iEdiuLX4oRhi
iH8eOUsg014vU6SY0+IrQDZ2chf3koLptjExbo9vXMkp674jTE+R4D+s1LKslhz3rXQQyjVN65tr
aK0au2e+UsTyvlj47pBMKz05ic+7yAl/31Csjj1x5+97M3dnvUhk/FftREgD4RHyNCw3OtNIn0Su
Nq30qrfn7vg+sN46UQge0/3K66Y3P4Ls0t4+GEi878hJ8TQ9teYvigCu0/HterJkAmzShJSMMLvl
aS2cOXksnuQ+1CL+vVJBZ+Kh1sGtbwJEKz9uS/OJzD+zc5v7ssXBWlkar3Mn04RoDYX9ckkBWrYT
iu9iude7WNlgM1Hp6BA69GU7sojR2I2gI6TGPh9SJD4WAxuAWnX2VrEHI7E8985V25lzaPfHxAIy
gjhH5X5i4ac2tJsWAZQD4u6TjlqC51HyfnadZ0J2ZCgbrTNZ6vestLck+Aw1k4mUSZGTyCya8pu4
Im4KpyT0bpLd5kTdqi2Ur8ee+a4wly0OrxUjAHoPbGxgM3Z3JM5RPZqvYUey2zhO/2H+77MrHiEV
ndtnnu/I+xp1lTyp8Xd3MACXgPVCZ8ZT6ynLZ3ZH2s468rBBpMYrK4GCpEF3tOZhtX7AdN22GCsp
+pG9esbKNcnztI9QE1Y9Qn97+8e6HoESn8rJ38Rt07symHDJ6VsvG5oh1zjwVDRxpzlJtK8ihjsW
QqoBymMkkVTMKCTf06VzBEPdHv/63VohUxB0btggYxsX/+R9AvHH02mOBtT/XeWEomWxbXPDO/na
S9CTQlK6C9MXnFEVcXpRYxZezYLIsgF+Iycj6UbQ9jfIERtfESsKZlrtEcFSmVeEFMrRhRLmubQk
T4fTfU66yxJURhMpbQ8jsPszjtObgV6uO4Arf+fTN/GqI/iVoxErJgGB1v0PWyQcUAVMMhX0Cp46
zRBiRSfWDdag4AcrIDt5c8WSQui+AMoQEJak1B+ZhDLAu+8G1BufguEpMghcUTywjf9mRotkL8eo
cOaCWS4bjqG9H7eg9V0rgux3soXZlivFtIZzG/5rSL0irgXaB9C6eY8aeIwN8J43VSmhkuXi5qn0
HFVkeeMsUlP9rw59g2y8z67BShQpRm183i9xwZUQMuEeEWIu1IO9e9vBQYUCZCQamqaFErllNL3g
dakjH+S6rLYxW5vqSiu4t0rjBx740k1uf3dM3+/rcYYtGYKC/ag5On8H9bFUXuudBijFBlVSzEOW
SaDgiWLUKM62lId8ZUKd5Yi7MlaoFyOHJmN1/boZm5raIidPvxrktVP2dofsL0k+au3G8ghdiK6W
NNjscl3JHB0qA0hWnWIxdtFfuGp9GkMnaTInXAxj1w3Rswxz6TJ8n9MpZR7/T6pAlYw9sxH14Rga
5fGWxg+B0LAwmGzRneMGSdWAC68p+yD9mFAOdcHXt1DBWTRpce8ouLtC/lO7IS6/z9LfL1nbgIiS
8gSnvcPhmEuR50tR1JxwxO45Wjye7DyRlWaIie3FjUwOUx7+SHz62s1JKTSBmhNQQQk6F8pYDPKc
i2yvlUc8xnMy3ahbxCDeXEZmypYB9OSVEDCiXK/8QeHBB+NMYQui/DABL2qz1gIuJC9ogEGvJHBt
2d6mrgKCU/vvgSRG5AYFIvOQG9KYO/bgW0yoD+Mj12oHBPIGhVGGwYpiIxPEZxQgELG/ceOmIEz3
i4M84SD4NfkfbBcz55VmWrCHVFeMgi2BB6xExvkd3sJk5Iox4SB67AJmlsnfWvLhmBcKUzKCQ2Kt
f9mu7bOIbpEa+Yjzikq3FMW1BxNQeVE9lIWWdv4wHdxSfs5i/mdrW7zSywbO5OoLKDvMH5NALZXI
P658FRVr6/5Y8FGgkG8Q+VgzpohL5E5za8oUZ7N2Ibby4oD4Fe5sFPuje4dQEGVmtD5wtCPgpX81
WttKRJgT8EjOFh2cIdFE3pCsHtNZuNOENQTapiwKv6W4J6MV00wd70aJcodaE0IOjsMBWxxJsFTS
cnHOv2oRgg5YkXVrdooR3SIDdZa/1yjHH6gJaoKP/FisHJ0QDSyhGeuFHL0D4P/TWy5HAnx+RbKC
lZdcEZ3J0W2YKA+MPfll5Blw4TovL1QMdZ123WmgBtk6OlhDPnutjR3MCWnnwkAWU0lr7VS7uE1g
j3fCb2UugEtfYuLXSYwlzuL/EkwDtzP9UB4QyAAXkbPJ/8fdotxVsZjraQLiaYv9Zqi81N9luaHp
sN9qPK0ymwjI1wDwFzmSD2z74jiLifDaFbMiVDGW96KyTP2k+m4jYAO60xXRuo28bzTzr7fKABqW
pQZzNIUFJ7+/g2W1z23V+PkNW2zcLdEB9yilsdAYM+KTvDJELD48+KsR29moH+eJ95HvA3K/oXUR
ttp49CPamC0Y+8AmTUXW/u9+5zLX32EqD01g3eMKEz9ju/I6RfYrz38YCcGM0uLGB1tV90KhpM6K
Q658FRsyJ0QzjEiNbARCnWhhUqAe03PJW80nfYnv4eRWRVSTGAwkMiAHuYNVMaJjf47R5elGFCFQ
iWQ6NjFZhcOXAcItpxeSACxJGMOWy3YLlmtBAyfvZxzhA3LCaPMn0dvX99OIU9MnoTTgm226TSaG
P7+eJzDg+Iuliq+qCpI/ia7B81lOyClMncwEiw/J/b0/oc2A2byYIhbdeNxEF11XOSxRger2792X
vqTn3v1jY6N6JmVsWMuPyzxN409G/HMk4q6h+D29B8Wsh1vAQ2eiBa1+O+KLCGZakFG7QyjD+tW+
rPbMd5WKsQK7uQXUkW1YTSxlRoWfowrOc3T/QU1PtZJ2XBpe90Fpk4Mw2Up5RWEVg9Gm5Ec2SXra
fTJ6CZx1Y9grradO1bjCfEOM6VomIfXYs3LfURqp5B1wOS9CG7X+BtZU0vXPLxuVORVcoNe8FSTp
Xn73qwI3JIo95scOBPxr/nMZhuGzsthlnwhDfNlwYCHMuFlWvLRtIlhcnUB+ILuEsdrnP9NuTVyA
gHphCvOyu8tgFbFA1oAX8xcmVlOOK6pKHNg7o02Op4kgqa3OYAfqonlrTRdEeHv+7wfy4YzZQ/7m
CiWmN+ELM7Sa8K69Ce3AdAauxa2AZ8z9EHolWhOnNyO4wj1fe+hR34q81GG/L/N4s+zRCHC9zjMX
mOhbg6NuMf+LgyJQkfUgQY0F6109EWQbOkLOSEPpvfg8V2bYIDRAfxiVMOk11qDFnFazivBAoZRg
NqA79sKw6m8NMSOmjrgu4pqjEElW2Yeci0Nh5hzfhrNq7Z2EfS6Wv//oUIjTGEno1M3yCz4xIdf9
kNVc1i+gpmOr0DOiYC1vxmNOmJnX1rGALiRRjRVMWHIATv4AgnV/gL331mAcS+1pVA1tSDvdHecc
tVgNfxCmmTIXP6LCeMH6O3f2KhAsW91099iWKEaQkiPvFzEg2LWhfvDN5jf34FXjmdQPFmI9as+n
g+eJ33/oCsnK+rHb7vGeJVI7EwejzdxxUqkkJw3mTw5sb1el2Z3zhHyTKSuSMSTj/Tj/iJjAsfl+
P3HDrQU7rKOJ4yOc2sRllx5cfNYjrbIzHZS/YNDNquyumrnGvJW1X5GgqFSAOBJKkOXiOfkxkrQw
/jgbSV5gIXjaqEPJ5uMQeIE0YY5J0wYVS7oncmy7tR4ke1KaQ3hIYAKNZlI5FLpwybKLbOvjJiuG
zd0baaIIOWHOCPyKy6ER8Zztu0ieo+QfueA3SMGKk08BXKwU1SD5BVmnVH0c26pYZCnOsW8ISpW/
6KO2Mmr9txHhE/wM1S9v3MRAYpzS+PQPxBBHKZF3rHJwpW/lD3n0lcmpM73Yq6kx39sO+Oms6agw
UoiwO1CHK5EZe/V4h3PbKhxFTyb+tq9Q1HRe8j5Hw1ZUF0X0RXb2JSh1c3nN5eilTW7h/ghgQgGl
r3Br6uJVP166KGvjG3m5U9C/TmY1vSmkUU/+H6AL/9N75OvrgRmdkd3d8c1jUMjPat2E3DK6Hp7T
k8b2biQDC6ChbBvDIKtJ7IhzkGZStBsnxxC9Xwm75165zXCUUtyMoc0ScaGde7zLEOaCeQRZ9ZRO
l3Vv4BJ94evkeqVrZeXo+Zuc/Ew2x3yn6WUbvjdsYqQOF/oHMiHq0fjWxxh+OIJfAbpDnwdUMKDi
DfM6xBdNO8ZUHIcTuZRH+dEYpSErZeyu1Wuh7GtGyJ8+m8BWbQWUZYPi0vz65TC6C7yQ9fi/SlDa
QeIxlLMY1N8vUU7vjNGP3yFC5uqM+Mn08XhawEFJ6yEFOMJ86w/limbfE8NP2wfA47+wDa4hn4nu
la3PNyLhHP4yxYUH/qxmPUL8TsGXfpVk46FV2dAffoOBIVhI8sLSBLhJVaodlwjkFGfrfwqCQKKi
C3KRWk2K9IB9ofWAxoDhy+zHRLu207HT+YNxvI22jLSklc7Z0R1wFu2afwTmWYm6ewmnTY9PdsEF
86RfQAS15CaJFFmGBA5CMrNO4qQOidu2IkTX/cm+op8EM2t/aL3kOgmAtcN556LvtqI/kToxwETH
fhZ0OhTW5A9OwMW+4QxlePCHeFSYz4y8qDa01Ox7ds/M0WqXDqmkIZFxGqsq2XBIZzK5U0OD9UV/
Er2O3YH7K60Hzggt4XnSg2L3PYJSxbyVz9pRlIqODPK7SSYbHi91tAD0NWD1wEdHQidOEvHLG36G
KUpnuHFdbbDopq940WncTBIg1WWuOtI+6hUcZUQExeSPlSdRX9wvv5PyRHveTFrafJNKaJATT0xU
dDexzNCGqGUO45DXGah3rBs2nGqSh7JZsJmcCAN1OHUcxqoDBcd+r3f1IVr1GOovUUWIUH/hRYS/
Q+PgwinFTeN+aOqV2VoeP7zefTUKugIMdXEQNco8aDI/yKLJ9CN5s4Ri2vSwdO5n6JzoBRlud26J
T/AAmESW1VHbjxLKWNs5D6dh0wd2CDn8Yi9xDpzcr35ToxTi+5waIPH76oOSILaRvPnyhkJZkYnX
WpH4L2q/ev8ZAQ8eypqhPQClL/PdjLRuBcahHb27ujemYSlICLvCq2gHhJquM9k3zcV9T8ln/gwI
8eeTo2LqqcC0ciXfNzXb/CVXFksB47yuBa76oszj4LIaGXcX4wniSxuSmV2TXeijEOyDzBUJ247u
T5iHrVArh9NaqlPMWM2M7vfq47pu982pXOFq84hHwkG5vAbz30DX/YtsKLXMkwV4j0ipl+tVz76y
5vJe/pSS9E8dVKfQGRMAiX5be9XGcY0g5eU0f3vW9obE5NpAEh4vftcJCJyqtVFGXymyMNR+kZlE
EIUEDyDLdoAbFsbOfFl4GA/jjhASF55lv9/nIfzwxRO8yUeNAxNdzlhztu8fXvO+1/w8JYPj7xWS
2R5JSyn61R6DPxuj4xYsrIRThfvQKm0KZ4UnXBtqC20KvBxeOQpXUnH5Z/WC9kilzYaDo157WBFu
/livFuQuaydB1gWlAwelARH3+a1pLUXH11AwTtXU5k3Lecsszf33qgodIDf2MS05wqRphSr6U4yk
/M/9OcdTtqf93mMc1Aka2IbKAfQ0YZ0hJnSrJVs/MohdORzQmern8VY4vYktiDHD7RmUQPJMhn8W
BxUajHozbgMWad5LhkrnDmxYgtdUxbFmz3QbjoQ/bYrloEfj1VViTueFYG5LpyclLLwOIl3Es5nu
RzqrXPHIhoLhviHj8TblGdoDobHQYnmgPL4Df0ZMsxzz+X03i1DTpL56aZ2LpMkfCCs1gNA9JiQ6
PnFYq4iPgnQhxQoDG3nDNM2Aa/0QC3DhUYQpdmsde4hFz2R4op5T6a42/naze1U9KzK3E1H9xhh5
xedZnZUUhbT63QFEW8lpvO5caaLoV8Pr/flqlc/tKhSznDUuIngHj8o/I5I1r2+4ZBBZpYwksvF2
VPAUWHqFbrcwdEcqGMS3/2GxUjSJxQV72XAtzMMXl3miv1lvbKgWKDMk7bDDqOxjqpVu1sZzyzIZ
8COT6mrHiCXLxnpVZ/cSn2vwnSJPxuKHVOIjx7hsY1xbPUds1SqOyXYDGi7x4Df6hDd8kJxm4rp7
Tv5TgzsI9idBMmt1w5Ls3AqcPZ/ETcy36yhdQSkx9a4oCI+j8CAoxBeDiewAYGg034O6PYAp3r7g
AbzT5b039IvMrh6pBfSoY/eTbA4AqFYlPK+0YnBDXp9QpJRxji8OTi4ucFU8+g8GPIaxaz9d7HqU
plUoqldCqq+ZZPvqgmeDYo03mG3PX2kiUfXvm+rU3anogSJK0bHvmmiJg/EfHjOpxEWtMmQ6yi8E
HA+opcRykSbkXtPk4bDibcjfv0/rCPeCnwmx3Xoq+/zS6iQRPbnfxS8RbH3lFKI+Wr4mU+7bq/du
ra8NXDDKr1Gx5TSgP+5ECrIyqd13D2q2eeEENXW5/1Mq7awrR7Gv2YKClZKCELeEBiqTg8NszQpt
Auzl46tgwlLhv4s5g0YPPq5T/u/V2Q44MS76f0JacA1z2Mv3mKIK6IeoA0H0vtH2YvrjwVGYijj/
ZqI48Rs7l1XKgt/iLRvZJ2/OyXtlJlVSeTYEoznRDMumbvHWmf36bBNA4waqRWBKDD5P2t3tVI/J
DzAXZa3HkUS7rlrmpXe3ZoX05oZUaAY9kH6zz8LHXQYmGEQv0WcWW2mNDSNHdMOTps7mA+efIthj
bkqhamBFBGayyU4Qjl2KCXPa9ylifAz2qfBW87pc6l2+lwyARaOYuZXfN4fsJlWecVsA+ylGbFhr
6lPlyaNv3fIN1iLfhll7NrOX10x64JxZuE0EBikUPqBCnwiRlXJIsPVv1uTBloOmC8jgRcGB7ul3
+WJQoaOaeVPEHvdaaspCaXhP5pnUlZM4vU3KCp3QAuO6VprlcCl6X6sxDAqgvL55mhlxUxal3ESm
6b4ggaNBFq0krruuOxJf/kxudE1DqJ8i56zisUL+pXJCyRtkEYMVPLR12YBn3DGFN2s8Qk02clxL
/yEwzr/DYvVRSBQ9uqT0Pfss//KORL2FoVP8sF8OIr+uWvlBQuXUufJCwDy4yCWOIrJ2QHA0DOvF
Sc+mdIH+L2zsuI/cGrMVO1jgfUVqB0Go2eBv0oXFsyaywEe8bHVXBSmUWH0UifbtwxhfRbyo9yvp
TqOLJvp/OcvuhqIpxfMuzhosBZQSkklUyoW9YICQ2SpxgtmSRgzmQ6I2196J2MceLS6q25VX0lEH
J96lEWmsVebI82B+2usHd4THENzcDdSNkSeSKI+w4DTo0h/J9JkRg0L+JEzN8eUcg4nW7A14K8H7
XmT5XCnsg4yA95MyXlKVdiFLGBH4V/DpgAr4E7ElZ5oVOzpVdtQsInQf4VLJOsjvcuMz64c18TkA
dowmVH2PBj9VC/QyD1FssssX9Y21awEplGTN7gD2bGO3h0XHZfRLIHsi6wOKlxE+EeoJBFUr3jej
+dGxEFQnZFmcHOm6Lm53kivH9qEpG4UONDR6LyxyB1sJ8IjVhCxs9UnWLusO9gGwP66MkTMQtesB
T3eHRrmVbWUERJBgrMo/Zq0aG5H8Kf8hR0QUGlGBWcYp2jXJngjtMWyRgLsi0e65wStMQ71Fb0tG
MWIkmvRkLAhRb/mRjv5F+dUaFTMiE6KzsYnVWEu8Z5vqiS6igTlLCqJZhvTjKqukMtP4taYUxViU
pS/wgQuBqa0f1Ra8z7OcthDoRCIt7fr2X2idmzcEOBv5wR3tlcU+F6SVeJ5SN1R2RiWq1RHaA0Ie
Zq2qGnGTpY5ahBXlIyfproZ8EPDDR7TOEPnOkp+NynliKaOKhL0XCJ3LgWwxFXFSWK1ruB1MT3Z/
DUiI8cabdtibWnteeFcYnQmIFw2hJQnefVIT93JIowRLHSLZ7PBFGV45MQc3ej1pzIhdirA99OI4
Ps0TXMsqtmClqXUhJI3Sgcl4sYZc0cCpfAW4sku9XCWfuKgC5g6rafgviZPk6doWAWP4PXaTfo7Y
69rCyzt0Eep9kMHyL+Yl4MQapiIlxqzfjm0ZVOMgIIqfMmny5ZLX0KIYSjj96Bq2oimC5xWc7Lpd
FIaSzoQLT4W9ELEqWVvzoggAVTELeYD9Kbt4iTfoBPs5uQXKGhxUrWCiJekc10ELS5ZCU2mNlGWM
VL0xRNCosrOl4c1/p0oS7uyzmh5GPbw1pVmdgrtm9eSMeF6XLRfI29qGfwvCIaa93FPmoLTLcbgM
3BcU7v+qIhQi0nq3AARYThVU0lgOO410fBIIfZqdGZnk6N54xCli0PgPq9n7ezQch+zIUT72hOHG
1cm7k2WcfB53qDaQ5MPJ1ZLDnbyDswiPEqpaZTPZowOs7gn4KsdwITgJPuyGlKpdSYBmmzLftecs
svcrFsn9ZUverkBUS0ciJ6x9FTecJPzXEA3W7NXSpW9BpuKM8FLkWyzoG00+7QmqSneGLw/AYUVq
OLZTAJxCbwcYNlThEopxqgY1tBD1dTPuddCSbMU6u1Mx+X1ExJKTXK1PqA6wXQ2fscIjas0sN3pr
fvSA4zSAuTRiasFRWrP3UVwe5M0aiOZLla2NQVJwOHZNHHbL3JI7e3qDIb5Kaqtjdx7kw5V5/aDh
0eiLNWqF35iVAQLF7Cm4ZnGMphpqb1L2mIA78fIHZFppYJca6UppMWHkidMi1jPAzTQ1sXTkqGKk
d1/jfWZQnFPrgLsmcYj5JUBllJBVTbg+M82QVxQY/ULRB6maE+KiYalGN01exiewRM4wmVPaqjZS
b1JAHejaZufNpiToaMq9Mea61Y4apfOj7kEwqua3PYsDCBVhahxBSFX7i2CTANjXcBuwiBw6yx6w
oEJ/5/rn3Kc0yUZyUsmmag8inyiS8mEfPtx/Q/1GMsqdFEcvxhZk2Fzl010PQurJ4iDCU9U4x3LJ
PHWQPPRHffAlbzlc5XzLd6sQnUlgv3OjSzclvrIcXz3EVu18zsxyfb35ZHgLI0J89Gd9iuHxuj/6
HCjlxBzHoQXdtTYLoFwRavLmp56aY4ngl0HXVHZyGK7K/XjbqJjUPurpS5pRUK1hyLPudUEMeL9S
CDZ9t24ppo+5oFo8Ot2bPYD05+tSROTPECq/A6CeXn6SIAZ/JmVibEHA/Wd0D5HCT6a116PVDLKo
IYAdj6DG03HBT1Y1fAcKtkQ+zVYzT8lTEzkR857gfEPefSKO0SPN8eQYEK6fAIS0j7scbcQzjOEk
5xstM1z8+AQNZ85v4Tml/Z1uLHPVtLcMcpFF9a1gPoJnlXLuUv1HiZMcvaiS4nKFB9QtYZvrHRu3
yE0dM4fOfgVqUcRlepFC/36hMZ2vRvBdrgByo45EhB03CgrnDKD1nvAR8LPvjxbmUSgGeIdPpME1
0MEHWieQwkduk+t+4Um9pTsqra0yxeMfsV1tf4lRiAhCBxjh1aOD9TmBUyZmeLtv1oiWTB/uYZky
+OQJUF9Lzk43Tid0wfNru5yT71nvLeSwHT/0p4w1x48X1wjOQScclsXc/K0Jc1X28p8xQCkpBP3i
LhWePVolLw99a5V6ZYRLNufgVCsRoHTxWlyWvMquuCTZS0GH1ThkC49yXXMrDXlXUuy4K2+RbZ5f
4LNrIMYxVeXSE7t9nd5PptN6zogvePDijAy45NjVTaQ05KdUC8JU3bj0st7X0MIOivGRc7cSRLnp
W78tLm+jWMfoHOhBYR1bfXCvAA2MJge8uRbJMlCEZjCLm31B9c9OCakDJLbkgXJ08b/AJVq3LaWN
rnr/QxH2h4tvJ5TnGQjAaf2qx3BJEQ+XtTAu2G5Mi3LBu9uZmj++EZAB+PBF5+3WXQgjqipwo0UY
Rx51tP1CSIzBMp7hubaTTN5tn76HVKd4wSiCfbHENIC2AT0Qe2EAzEbYGjxJN8yiM460OtJr3o1t
J3vjtaTzJxRBroqx94BLrZ7Q/aVNzwqYUJIHD6qGOF3P5/Qh5xESVSS/vbWBHwTs0sCAXCUtjfJa
HvJT2Gn5gHYJQGwsKt/9LldGpshchccQxaXoJK6OA908x6NukAUwzBo4wV7IyHX7GkD/fB075rhl
frx00I+ACTmF56uq1RX0vlwX6RfXpOFqdTdKmSPCZBVqnlpwkfm5c/0b7o59G68633OpeiTN3cBD
yV6KsByx3SnR9HnEXPU4VBYJ0jrpL4CuEfL/whDczOBU5qZZlbYF+p7BCLIc5sdTyemsE6m7wzQk
qw3f/lNbsKsLIsZAnHddrMakydA6se+pDkyYE/Xn9joCm1eqsK1oQItgVbQKzUOvzwA+3Png0meZ
sgOskwTiJrteUE88bF+GnzT25rpa+9bsaNfs1nVkdMUUZuMVH6uyGYth22W+JpYo4iABomgIg1gL
t4gaXin01G8znnJXRT9RROPoxtkE4zKgkz9fr3JDwpf1zkE84GwRVASCDCUxJtcPto03LkdS/9xa
8BWxNyuuDTvJdN44EG8VRhslsQDN4nbh+uEVAoQb/sfw1Zpisx1eXnOc9DJ15un4aP9xYjnX/KKW
GCT6aTa/63SOiNrAUfVGjoVZB1XGzf/oGZhvGq/e6h4PmaLu8hKF/lEtWEt3jhrrV/jOR0MIiiAk
+ZM9ktK2RsNCanle5I5iVlSJtNfOV4pLv6BxnWMfh0OgkqDOkh6xXqNZ36L0lMuCl+n1Q1UmMZoI
qkfQuksjD6UT5yIIpVrCbPE78r5Q/1XuWTwDc212tSE5FUpxPeuW/TsnuwRvefvBosZ+eUW2A6m3
oQ6uuYCEz1msV0DCAiTfDkT7LehCK588Tud+VVq1JBW1weSvlkZa+XKi4lh8T4pyOmVdPKuPgrWa
NywOMI2aNHj4eg7p3zxRLUQyXE4czDuy3i7hqzGvaH6WztFOU6pQf5OEzkpHGwozF13d+3PdwQ62
w/KX3XWeLs7QHLlLfvXOT4ks+ChN9Y3H35GMpChxR6A558Ot4o28E8f8V5qRwgHORzlnUigATdSC
chPhKa+cj4uYk4UWxVglXd2OqpEZzQeMQF8Wq+jsh9Vrkhs0fNlZn+ULdKgffBrktdV4Rnt3DlT0
bvaRzOstUIbRLZfMjG/3zVGTHLgmVQ5KmGg/VlE/IjPpxdt9MlogzEToy9/gA2fGloODPCF8IsFJ
OFzXAPvfWYzn1Y/8qr6tecUmrorHvyu1NAx7lqEDaMsG9aWJnkKTmN8ypUibVU6nKmMQUlIbCgdP
BAy/VYiYpFHBvJzzKbVakD4C/zbCnnY0eajp/jIgDSsTzk9c7EZ9c+/gM/G6I6LKcIHjCx9/QaZO
5ytDx22Z7bJ61Wuo1JfrCG61qzH8Spxr3FHRGASmAOqafyiOGgnUUvfexZbUVRARl8sAMEeCS6z1
2iFcy1w441Ij1KGUfcxZMy6mo9s442S8sM+aMH3mKITqthXNrAzXPYh1lsogzz+4mGwGCZKGC/YP
bNHT+JfgLzsDLkX5mCefmwu45X5PhBa/VIb+dCoHrdmlSey9b7VG0J1gidik1iODxAJq/Cpe4CWK
eS4vmNGNbuv/mqdvhmzKa6rYgPXgHeSys4LguHRcqlmLczjzqATaSYkNbY4lb8POvIpkPx9bvLei
RZAr9IHUAhDaRYNZq1t2ko1XU8nog2d+gmAD1wg65gsrj75MgXm/D2gLYq/+z40G+kx7yiQyn3Ee
IOvaDeNgLEeQMjdkMsI7UqGQuyH3lJwliT4JT27DJhkgBr5e/K/iVKfNxqTHdpLUnYJIKqgtjB4Z
vFPK2X6NXW0KKbXBm86HrLL206jREIo8nTVxgHz4IFVZP01DB/I4cua6oRc0ry09lLqugaJBcbp1
SCVFFAOs/t0CGcS6vUopaClohaLiJIIhcWu/6VH6sJ6oRi5WWcyFwysUNbkcnyyN0TkFKZsol24z
3BGHUHuimKCNtl5TlX8jxlUh0T31L+OVL1p6yuUvlJSEcv3wOMWf0a76g9qUmO92FiSFXX4bVLAT
bPHdZFxUsYGCykU0JPvXm1AA1vkza/BoBQbsbJDZRiAsxE7hE0ehXHsyDoDCNXz3vZDd97t9sPZB
wuXlMMqi0Q4wTL6ctFuAddytv8iiodwaAIa9jhr9O74PnybtULLnuAsSLUp6+BF0KTyKumFmt08l
RqxKHuGWs1QVg2PaioApPZ8ePLGn3hGgYh4s+3/b9xllpD6CZRepgS8oV9f7C+QoRhrV7qdWGzlD
aauWv3JfnSDKaB0sOZ0YGolxmJXT/U7KrysbsHlSVXBHculSVxxYUBJy9p2UaRrU/TJKesPkz89T
MKu8ZU2FV4ySD/nx/iXonwTHS2o5PEZ8N1C9V9JwPWUpxhPegv+83nNfPavFvtO9/5Lj4klOe1jC
nXyoMGywd7tZFJvbkkBTR/c9Db2xiVGvz11SR0trCi13jxYCe5qUrSvTYKCSiN9OOrOecBlH2oE1
iDwLnrfkUYC20SfHyjJVAyx7AYjlET6dQReENURyrtFfaLD58C+feOfZbexgNC3qPBMN24mmYLrV
M7DTMVhq+x82Q1hgEJ5LsxEmixlnQwdmWMw5u5aCsCLRyBi14hPrAKnZZsRQWt3Gv3Jzt4XFWlAt
YXdtFEmx3dOOvY16/y6h1bQE29x32PTvaNvwHa3PxhlCOmGplieo0MYRYCdt4n5EyZkB4uXMXVPe
qUfDJ0X0gj6kWVHhXbVYaR7Ud2FxsqqlXCuFT1nbCeINL39l/3natGrDFyW/GYRDGrxWJ1NcTTDJ
FSFLYacYAtS4JZGt7c6hekSDdzmZdGHy3ONey6ldj/04cQG+VxTjOiqZDdo5fisAyNJcMeqtfbQO
At0v2Ym4t08g8/fbjZ7KQHKB9LUM8fKWmIO3Z734+I0AfkWArfl6VfySFzRGrwnVloO301J97IfU
BN6ITtKEBC/GLskKswOcou17HkVyuUfQJb9yq0q2XTgfzj9asc31+07FfF7tvNkR6d5FDj8WugXT
LJZfO5giMIbGVq22/Yrp5MsZ/lAJK6m6TDJ9i8CrbWylt9CaXSx7uIkJuOYDNdBoA7CgLyCrU/xz
wB8L60hqR7v7G7QDMBoyatvOxiBlkKL5nwRo1CzPBu39ekFV6ozBMO/OB1Fu4jEDnlew6SL7xhqn
IcOvBuT2EPAYY75WszpJqgfNKTpwlfo7kR/E/+JC9VtIs8MwYPCW/GBclPgtndn3jxuR0M+ZRYc8
cxF4RjfgWb0yev2zRLstuwKp9mlRWiUsFZuQOSjOED5IwGN7PXVqW9b825qKrYQdaY5GmBLo8BP6
bsmrlnqfL1h1f5hT5hLfJ7PeZT1K8+9bxZ+Z0AB1vp5w7Ez+dp3RgPdQi4iP10KB0Kyf/M/46gSP
SpesH9X2KPxYqfjtxwX3kjqIitT7uaU8nSl0w23G+nufLGDhyJhheNqRACSevUfUyNJioA+jDv/R
pSFRik58cvdd7AgQE+nNAJCX0rJXFxocJXHOVrnZY2HVX3xgMJ4iOaGjM6Ucu0VAqSh5t5MIzSco
MPjRTvcymS0v3imjBhyC9On8ZH0zzRL8vB9YnSuiNTlGpYWOMfBzG014H/1oSdgbigUIiwz8NtJK
BL6wJUToqMGKrYb1OOE1/K4LkFjxb0fggkQFuMtp/nnVOfCCbrjINg0QJkBWC7HZVybOzw3Wyrrf
KDEn5fjO5Uq0F+2kXcvi+DEfqVP/FLmRg4OVXTUxKfm6NTJxcV4S0/Aoe9PUzpukD7K+KzasQNRP
hWhetmMXUsYxAVJ7/4W9NNsf6Uvr7YPaBprDMZvRHo9p8sZmBIGK2heyfuf7SImSJo1rKrE44QIu
ytxJqUiSN1ZX4s8ao/WLT+5gRU1G4YJSfsil0bnxW7378c/hkPjWlZRY/28QhJee0UZf4nlXVUiW
HK6kjNGSYfvqB1wdqc1fpfT1H+ZxMiFoul9YN5KwdZsDvnfYNVTpYcAzQJbA2oz1R0M5sc6/GK+u
XktxqnltWoM93VaieCs8GSDZAcxdD+zbaFueoDm8tg5IRV7dzGPMpDNcLUhmgNNz0NFw1RaWyFR2
tq9pEHMRFqf100hVIpZILE3kcVSpDsLi4pRw6oDnzFEKbHq4WmuWVJ8J2GXiktrR2DteX/4I7x4D
fPUkoYWfB4XaMwdzYnf0E0YHxacxPDuyPpH2OAOp/JvzPh1k48lAUZM7WSXkfH+KkUb+vF48ohI7
ckNxbzVD87zARj2cTFH5YnoPe910/ygYO2BrXeJI8OPmjIH0FmrMV5U1RhEBteBQ0Gv/8H0KUx56
fE5sZRnfMWWgFCrgKGeB3Mpg/4xCggMJb9YBPAod0eno3F+vGMbU55+1g8YCW8MwfBVT+QMmMfr2
upl+g/Uj3/vTCjA4jVbwQEcbhHFAb2bs8Ewv7xDDaJjFaOd933H9qvADJfTa7MU+Wea3xuJvxGjL
wJqc5IZ6F7W+F/ywx2tEUyrw9AqS0C6Xt7MtDQTOKrE2doDBPHtcUmno7hrTnrEG/yxtDN/L9QHc
FarMVO6uUwM2M2ssQP35neIVtvlaZIKabu6M+c9cPCTjuGm3vB61RkCKh7O4D4kK8tjJEuewF4wc
2AX5Sy88J6nD6p3xcDUQLYGBmAeJTiMU/Prb2CtBam7K3/IJRAwZMIctokSYE0GNEa9CWADX5IWT
jzfNSP/uc4HvQxTrQXJCpR5wAy90dtk7alTiQjzrZaN4DEwmWpAT7u5OKet7R5cMDO/wVMtsDHPg
MiEMlB7X4LvK4nYrBq0dmw9qRJQlssNisYetLcYUKdfFw0tSoVrOMwSqEu+Dyl4KMkCrU5fijP27
7nfBd6/TAGrftdAIlOqvPXtks0J0xwqZ1Wv8ot+9dqYxPxqvjC96NoYo3RD14Ti+7mIqTZrxT8ih
u1T/zAfbvWl4cr86tlRPHEPfMWUJMf9V4Gf0tRUvbbJx18sdVrK6KdtAQGUQ03RT183earaKMdNQ
dyd4/E+MK0cIwKKJkN2wxEpuIovijLgjDmSel/7PyVGGh3xQz0IQt4hFxkM1efYOHQDnCGpXnNbi
tE8VlCepmqoL7K9u37DaYI9Xaa5i1CiCui29M9KBLW3TOg4/2hJKEmZGdQ3RlfHnrPNWPIHxNlDO
vJg0bsCnLEBTpUxFNhu+cyWQg2Ci37n0/SEJZ1eZGCD933AcvEGdtLRbJZfPBTLQE8wcyNqTClCs
uif9Gkbrj18JlDYr2xzvaHtMGaDF9wiAYl53PhXujb6FkVLb+k+oEDAvP5KeK0LaYiwogXZc70fL
rc/1CUptqX8mF6yMxstxIAPr9fDbRqiEdy6yXalQ1e9IJ0Iv2iM6HAhr4XGcRgnsAWkonilsqPBp
J3xZCogmgXF7nthH2fzDmwrB5PN7zU5n0BYXp7bA38QKVYOe/oboYrdUZf0aRvhvvQymmy1maai1
APIuGcbXwOov6GJWwvo47POSfldJgsOzR++GaNVSdk6OOp0N8YY2wU5FVVCxJFL5ah8MYn4PM6zr
2MHW/Dj2LFM56mFq5A5uXaIALDo5b6UK7sF36LnYFOn7X8XCt4B0yTamW8xaLhZApNpaeyliVXUP
27t44KxV13DU2eyBsJYHT2z7hhp6B2YbBHwC5bk/hG4undrJqdVXGLa5q1TyoWyf3I/8hFst2dxY
Fozqn/RIhPfJRhzUI0UEEoNYDE+fCxlhEvyQ9hUUmXQxRO0uYYGB3kasFwKEioDXwx3DBRjbpYs9
dOZcVuehKaNMreZfeezoMPhsTv2CcLwAh9teYOMyAQZFcPGarxz7z391ePhOZXNzudLdNLbHip6g
Dvh1MKh40MbKijHXtwtcJV0s4P32Dlb6aMQG0j1YbEl9bapzruX2M1IwVSmLZr+MZsOWC5u1VSPS
8xOe9TlgcoRgeb44v95QfzVvSeaJUI2Fig4mZbFs90Sap2Z+JsDf6T1mJGJM9C0S53XCaAKUx2SJ
A/4xSbwpBZVJr8Kk4gFfE2IIn7Pn/HBlqt8IVxnlvCgdMu2zDqIxsP+CGBsJk+btqpwY7b64FA2P
b3ltntf/2whpn1xGRRzGe4jFKGU46j5byN7Q6zVzrif6TL2KsrlusuGXNYOIgh9CmiNRdga9tFuZ
BNAUFZiHPiXDy1epuLmOHOPB2hrwrtdhIiBhSxlI9MD57kI51fhKQzbendVfN/mZbmBf79cedFsc
OJ7UqCE8Dq3QSyN/mztixC5zwOXVCe6kAkXvNOqlOcW9RAW1ZKfO68xiLmP/VQUHuUIT4dWV68NI
oIBjosV/NhwGdDs6bmvCkpLnzcQFI+V3G+S25+n8QPmFPhZlt8TrbCZXUePCy0Y0cYWVdsaVNLub
prRhoOAag+gTFH0vt+9pul3iYGEfOtjBnpfKtxqBW1Eok8MS60IK7NeFX9HTUXqWR66bqIMbWpzL
KOsHUG6vbfA3FKZKAKtbHIKJutHH0Wu3wT48+4FngcRZkMF4kPrtYxwb2sextS20LXo9R+kiiiJp
AhW77FHR3RMz3XEzuyCBZflJ0Jqu/18J+oHP9A5rmVxIUDq4HL3AVQs5JHrgKcCfFoTqsLewZ+pA
X6gR/NTLJGeappc+PgPEyCOa1N2fHulH4ZSga1sg68YN8SqM78M44Y2O9VdKmq/Tb7vgrms+Ufzx
uR+5hrWuESfhaFCNAWiHjRGPU7yt1KYUBJ8GVKLlyB6yfYoPUIATpxbeXWKEIkaROBYUihrE+D+6
B/yXwiwU+nV6EBrS+U40tNnAuJ3eGe5LEq5qPEeDOdRzdeXtq5iipqTkACLSsJpu7SHpp9lud82m
/qnLsP5QjTwm6a6NzrzdxdZ1eJJQQ4T0ZVwyXK2DQCMj9BmRVBA5MuMWEu+JZfAS/HsfSExF9iQc
y98uSLPXFneXJbc/geI0pdppDptOjqK6FKqyw8zwJ0KCXJ8Q1375tZ25mXU8s3FN9mrw1pMKixrO
sGxano8l+TzAs5eN7eyyiCpywk2oIM0q+Bzb4vL0i0LxtZbjbJ3b3fGp7oJ0GHUE7L/Rtt/sHS3V
q1dPOCBM/Eg1X82fUBGo5dDr0JK8vgbhrUpEb0DYLrfTkYZ3/k8Hh8L91gMU3gqv/sQL+5a4fD0Y
CMsxdVrvvXWdNBOVUGBi04JvBlzZHGczqkNDIS0ewIRD7cxGKjpYC0hMvCN6cN94UDGIhGX8eFiS
wQgv/Bqb3UQ09l+KjviLbKE4zimPwObFbfQsq17F896VT44oYUCnUK5Lp9t+fwpXATYzh7zWTCON
SInPLn2gEW7FVhotIg0aPMz2ekfys99sc/EdUMCM7KvwMO8yWS4blPIN5o+4vqjZJ9BFXpiBRfx+
pEKXlbK0fA6ro3fGECKqTKeTJr9ebgj/RGjCwkwFDSvPW8vzuT4dQLG3/DNcxs0WH1WM94tNCxob
rWnTaU7KB4y634/Mk4qSmxIuTqN61zAKkeKz/V57nf7Jle9T7Cs9RUGdd/8wLoDH7n7HjfYXMUch
RZZgJKLaKuEsoHNE2iPhLTBWXoXRM3WiDDshYNJZ+IJN2fc/APsG/id7ZaqPDSHjvPi1AObtjKiI
iq/BNYXnZ+jba9iJIHD0vSMcuJ4AajOuw+sQOkpswUHZcUNZ3uPqxEchiACzdhQuswYsnd9Bl8Au
Dn9TDWIkq6gXIxvTwTHBAsgrHWRXkkFQk3F0WOtVHcAtmjO7v2VyR61tS1p/hWnsl0KnhsjkjdCV
KQD9KBdAUKeOtuYKHs7VtTWO27+1fdOdo8HQwnFmCs5hrQ8L0lRHROh4qZe5IRuyWJjoZe+m/2Tg
9ZbDh0gUuyEubBi0VdJGQEY2Kcctav5yl+hNstwGJhZYMVEALT1mLIXsq5pr95KiF0qU3ebB7JoD
Ymai2gWvKChiZ6/DIj6jBjggOw25mZ+ct2HHulYO3rhkL1mtSjOgfkZElM8b96Pya+kVbFzKik/Q
5XxdaSD9sToxuy8m+D5r+N0eAPw7JxgTxd3UmMkps1kAKfJPdMmj1e1ecr0Yj/OIenya0VPK0mn1
NjfLUbcPQxfTDL7Yh21+9HquVo61QOgXikY3VjIiqnOcotLgp3PS3/M3DPZ48XUBOjeImPW99gsB
eFv/5ZLCBweuvlYYy9ukAm9NHKPhchGl19wTtaTsKVq3Gc2ShYx+YIGcV+9gMvu5BBA44NUJfYHx
Om72cs0WHLb0P/CheuZzQBI+Wm0ThhJaRjZAG7MeTJ1T2geplepz4EZJOvAuLZuwdfDsvPQDR3nk
wS74sSeNmHf6juMpo2re46OHU/SPP1FwmUWihhiT4lq1Uq+nSuou/d0VXdxyWeCvgSDyAIw9/98E
5t9e58VQvyOUJQmutriXWYpWp6JyhSaXbcRgJmFImQW9jjaqctUZ3m5x4nQGq50epT0CrYZoUqp1
Eid//JKzBwGaurS3neLkd34XjnHjWob89oZ4qB5N9scgYZC3RT1OOtN+tYEbIC/E56d6elIQYjPq
qe/xyN5IoUfRzP/KXCOIyvtfc4kc32JqB33HWbMpGAdH7dOeb73JbosGruLRG3ea3nychL6OVO1f
6k7/wf/1OXcyz7Ra5f/dOvPTClI4ordqNRNfDQZwmWMGBTOcbYgN84vW2sL2e7Erk+5e+iTxlSdH
fubX4ZCXC9oV3zR4EIxidNJTcRa5Y9/+Ijz/7dwlxSLiqD+Ntdww4ZyZW8aQqN6leS5egWWrflR8
4iNBVP1Puj8rulkq5Uec85aKhsV2LdQW+Ig7QBG33aKjOpTANPOykWqvFToEqQlMIR9SMrbMkysG
TvcdnMEquBIZAwYMTi7UopgEbJBZIWXOEhLAdSURp/rZ3TdxoEmpF8ybdVoD5QdGoLVai7yzI8Hk
sGEqPKe88v91Ue5t3RFa5hHUHNZ3SdGalra4L++UJmmcG0F11YqUL/6Fwgm5fKNKAWGpZ8Vx9Vb2
8SdxVQztarIbpvaqqeAnb3dEXZM5MLKJI1FyiK+tKiTp2l3hR/ikX/TP8W0ROwvB24n3EigGp7hP
oC4bkUeuCYYzhfU0cLUoOtvvDKXNjCBj9JQac0EnJQjRauiBtut0QfpIIBP4x1bs+wtXjIpzXdux
YS1sxp+4Zn/hpPvjpBZW7ZBqgEp2YwhllK27ah17fN1c5nNTaFR5srLsBMioN96s2DKb3kI/nmjj
wqUKV4UC5NEmvbjhsMx8MPnEHzW4L4GYOfqDF9crnHSSBEtolLc9+qq8lmVBUR1QQeXwGMbWc2MG
g6A//VY9tOVklV4KwC6vOLM1FP2FLtndHw5Vez4UkBR+JHIoU0OoKfaxhVdDKWCAkjy7u+4cXFjQ
JaEoHfuFRfImJj7fCRrYIms5jezw0HQt2lBrZXNhH2mLJoPHbAFJscdKTUa6Vc627aPHMATPACR2
EwWsXJtbyzNuqPcr8ypKpNPCXXUwCgp3ktkVWy5D6dw8Fxk3mVdXsmV7wRkDZuDN6j853FIlSKHi
/VIkOo2kG8CRyd3x8bZYbalq/WSBgMdbjEDtTHN0rrsMil+YZKjK+U9ObGof8zMj/Nf84ud2V8Z1
Hccosr/qTmnLq59MBbCR4RgUbRso8bGa1rT3dFzE2/qBnU0wmIQyFq674cUY/GZWa6goRfXrW+OJ
pQDxVjfyiMmtDHOvYyp+Fmx5Vw2IOVSeERL8HMkt7vRbdD5yEIkbbUO8Iore+EcLp8msRV+8JCxH
oXq3u0URiKP+qmUwLr3ABYix9qchImvWzCrOarUbofxRRIeX5ENSk0LQYZlXhsHOV2c/6N9KazQM
3p9FFJjag1vJ/epIENd7ltCAiGInxlcn81n1GR6Pg8wc5X/q3icPlN94FLKfmyq/CVTM18LLtg3D
9vKSBqTumVRjCTgvQOmzwg00nK6UnMYr+tg2o7E3uzg1z3TnB90JB+C27OhoQUBLr8zKJbjQoMGY
i96HOVjhbs1LAaTyYf1J40nT1fuqsFGyER12OC+65ArZvmatT0BCboitU22h9uPl/4hpkS+uK/ej
FYp5ZD7apZ7/JAqsKrsHZ3JW9fDr0JaIi13wlJwM9vesrrUsIWmO5xDEQovjdAEbWV9uhv2wmL7J
OtN67dTaBC9h0uO53UMC01L86mYWxhIp2jIdVawy7x48h8M66m8OorBoMjJs6LjiAdrJJYpAmL5c
6krEKnCCasR/tN2dEW3tQgBXwex7vNodADjemu7Wq73XkCpxWlM8yf/PAV0EcpRaIhBBtc4v8g1N
MmNIt4H4cBj/QDAI1cmNNJEnGEQdcUIWGcM31xh9GwPZfZgYBsFeuHhH6M3Qxvt5K2NfneIFRkBE
SmhyYOwB4hBYUe++aWvvG0LB0gh5O/LM3kFhnz4dn4EtIqSwAKb4J+NexDhr9JrPjg0yEuLYYZt/
v5seOGn2CUf0K9V/BenxvkTuyAisG7nk8ol8CuqebEHz7TrWm57glHb7xDZccM23SwWkjJ0utjQ5
P/a4KNRbj9JpIDNfmtdDKJlXR9l+ZqeObXPj0+usNR/5yElxzMRpUeXY7GtfkzS01hAs1XaZoLCm
mmq/mPUez/WBqdbWrAfTEvfGr4I6wepLuWfCx+O7QKue4fxrvLvzL72hHiqPz5EESPACzOMx56FK
D0EVspHKvbBYt+9v/F6r0vR4F06YOlPe2DhcIESHmagBHumXqGT55GI5DuLY8wvjveb5aB1XmTEC
i4wPPQqI5AgM+25xy6A8oHTWLb9dNw+NUWFFlfSjI5KYOesYAoGcEyiLHounugWJUMPMbRJcZJxV
+Y4qOnCJ/XHyRQ5a7OBuZ33mVj7sLa18AoEBNvLNiLcLksWbF8WHiTrPTjx4VKmlcWB4CV8eJ3Fe
aaUWaFxbdLOu/ZdpyL7z8aq7hkzut/oNGBy8n0gs2+P9QF7SrkDTbuSUc40NVgbogVKLwY6rOsa/
qfXgXdt01yg4ptU3AtqyUz/3dJYrEGvY5d6g76pBFDXKh8Fc19wHD30KTP1BN0hwhj0F/mqpgBVs
FsUg6NEt9bYKi9JQP+L1Mfyv9cM/N4LK0BMkLzUCvCs00dCTv6sTSgys3ePyE1/dVRv3E06jt3QD
YdjS/r5jHArreQzmDXcKqbCbDDT9HdENI7qCnTnnm6LbXJAsH/9/4KEz54aYMcK8EqCWW0a+Qhdz
6mH6qOAeYPWnmKv1GHbaWLAyIy/vM9uwPnn0dBCFIAl/gCzMkwJVRmwB/XuI4v16eaVX++PF4asZ
iLnOKgTcyfjYm8fgHHh1B6gW8a825/C/Es1JIyq4P0X7S8Y+YTDUH9PWGZfRrtM8mYJ3zlIbgzis
ZewZYRACM9GqFoTeIVY/a21fS6Q+okDhLeFmGRxOWXLastkV81vzjdziZTL2V2vr7jaZX0rpUvlW
WFUv0VpF6y1l5LBusF489bss+xa2EgfqDLqleStbTKg3Ld6Opz8iM19yxwckyeQgnbSP36e1oNOl
9WwosPcbQKUYpWj94v4lQEKesnZFEi9xSMH0hQKnZKxd7DIYL42+BvRjGiu6y9K2Trx4LswpL64x
uvbVS/ZOu0opRdahefEUjXwpcYNZYVOXvIzqkjbfL6IwGzGj8Vl7y3z/eBgAeTS2EUmVjC8sBM2f
/Tj3XZa8AmPrn/ZrRD83cn66D56DQvQ0SdO+gFKhgawiGYsot8efH1YGul/e3/vcQv5e84pUvyxe
CmQT71StaqutTCkrMUNKuT/NdpmP5kfDUEMkPpmX0+U6OfdeIt2rDFHXoN0AVkvzMGF+3+4Jzacu
F9ZEs2rX2OJq3HPLHcU8zabYvycMeHcaltykx03NvL+f1BP4on+8lNyVJ5o7cVagaq/w5ibrO2Oh
/1zWXIAXtErsURiuYm+Gid8TbePhu796ppzBZSoQdOZGLAQFMux0gxcwSRW9cRSIwA99r6GOb1FD
e7Dbey9oSunVXNJJL8VyQ86HuPcSgvHIMHHBxPgxpE8hXWKBPqeGd2SNxX3C8tYjh+jOfIEkWWIf
gtNk5EWORmSlLH80R8UwY0do7HviJsXoAdjQMpZtLi27d7pCsJLsEVLsv6q2fw/bePcRo4wFPuRh
G/u67xV7RKX2+ezSt4+Fs549KCyK8O0ZZdn5MsWzK7tyjUfUodss17JrPSLNbd4ErVYz8rWJG6dA
m2owqm5B1+gwhcoiog63lxrndQvbAcdewUUcluxZGzrPeSS9Xwn6UpwBDtGGr2EDvF9y4HZeZVQj
dsHX+FyJ1WYcl2FnuHerUsNGrcOe7PRrBf23cpq63dM5JLChfN5j2GrcFjXMtp8shtbx77A1HLIO
suE4czsrLEqCSvIjYlTUO4vYvOXzhEv0v+Eu7xYUfRuec809ovjvkXp5RYb2Clddcj8yZy1IUpra
/TsEhzEzZ5Y48eMLxZ5dtQJI38hToHOn0XGd8F6keF/hEuil96M+AnuPIJBTSBSqg8s5pR1ivvld
BoqSyOTqn+sQMll6AQ7VOYSCpx8ocr4gdMbRebso0pje+hcPY1g+sUykXhGILMMeTHl2cddJ2MPr
ALgxpPYLWRE307NueenxXZLJo7/tn4XBDch3Uz65QyGeSgtXZpEP+uFV3dpXI0qIHK8omOSd247n
YRbgaaQX4zVCw5yoSnBBASi9AvFAmRVRrrWW0PQopMqbSEIckq1MrKKTWNy+TwZ4SNzJ1pjB6Psp
9V2qXPnKijSHwnJCdpsYi4VcVciwBPd3r3m3CIJ75IUiuIYt/1leO1yW44oh4ykFO23+XXZmNGCM
Pl+utHlo9P/OPH9+IKnEv8Ps4Yhz4A5WnbaPu5R99ykmTDlx1G+LufuV7dbRSOHpYxUNqgK4qP8d
3ZHcCZnGaGra8mYWylFVu9A2ovsqp1jfe4I4mnhEilvBsfhwK+ESPcnbFZPmHcl8rdSNDl4r7Yrz
xsKGZQO5KezTOvvZzXebl5R50b0Jwm7UAnqjLdyon8u6CFDM0IcAbvKVYUV1QF534kwNujcxUFhW
fVTYCMzV4J5TmYbKqIFwk8/WYdlbV79cqvl2kIswmm6Qalfb/FvQ4l6CqxQzITkXBLZJc9rEvXaB
ku2WrXsS838VkAR+97K/HZ5mhm3arluAmkR331PE3+h6aGzLQAQimJGDk++D0Jr6pkQEe4AumetR
Ah/YmUlchwgIeINvcEsZWjqWf7RWa+KJdY0F2XLKqPtmKOIGPFwA4hQaUHKPUoraSjRgXUAe3Stv
BywE8JFAHfJgNxKiULnUM1JKbZkh6Pora/V97TvG/O7xpFRXptdmp24oF8MUdxMnibEf1xQmRWa7
NPdNBJPxduuyKjcDzd5d8liUFz6HseyCzCYOUEN+iezyE5t7RMGm+5Wm6zuN+bEUvH4woD7ztxjI
7b+9tvpJgSGtU4NAfhc5SfSZelYv4b1RlNsJCLLdxM4nTWMe8lDhgxqP3LthFp70ExML6QYlgu51
py7tsdt40NfwWGwnrk4bu4o3/DMjHfP7vDgTSBqwRKo7xXj9+g89pGVmo+cjOS+naRKxVlnS2Jfj
ei940yKS6GRtm9R3906qDTSvYEdmJBjX7GmUuoWPrL3u4WOOEiLE56Bv8YLHANEjFmCYg/QWmv0j
Gmx4EIZclk0J4FuJH4kgdyrtSPihyu5/CJC3iAY4jdASFSoZL9uoL6i6Xu9AkA2ckUPhwFtBAIeb
EU9B01NCTK+L5Ci36flngVYUcjbOyLBgsBd1vH8V6ySMC+bAscIJT7sVMMlqPUq/PjHd1ciLcasq
mCiNO1CDnPeaHA3vUhNWMWDK3tFSh4gbH4f/msaH05d5bqSpRBcYtE/+bbv56bkDSzjrhjkaLtAu
1oUXBMp/S+To/LNctWwMK+kG52TdYEjHhIUjOTYjldqkWReCwHsd5fzde4xn/hOTvUhs/oH0vRIh
S6GLWzRYCN+LuJvSW0XFBXBkeXoCMejQxbOBN+vy6dr0fYcYpAxb6jvDlaWTuVaeIHPn+1S/tTVJ
5BMRmQa9osn2r6qkATQRSGQ9glWl1bd/tR/yTlnDXUif5RL1JsY6vMtaLeplp4y/wEzYmHVLRChf
m+kPPqF+Ot6VEwjWucTZlwXgTHvbaZKW8ifxnQ0tn+IOn84mZUrkdstIcdyG067ZXMuT/Z9/cM7Q
3bKHlJ16q/R275rKQkGO+gEQqeg+FoDlGxVKD4zL5D6+Nlkxgj38rbGurBDtYlhMV8a94x8okDns
UvDorRwBSmOryL7YgJCMLjhtlZm9aFbabVY0mKsfWWaSz1pcn//FsdJ3oI9VQo1y7gVK39OlZ9QX
uTMOcrTrTsMP7Cws/Uc+T72hI13YFEVXyS1j/0J4sfw1RgMlrk+Yj2el795GFkJd6ziuBXZOfq6t
Czr6vN0o9N2FIuBfhzUpeERKEWOj3FyijBE+QZQ4HVs27uhNn0Z/DEa2PGY4MCIYRXMSqrxNJe52
ZtEy89Ube4rOvYig5xoOgwt4BBDaiIaCWEdGcY367Rx2dFjXPmcB7wDH538a3ze1q4TpqWHpIeRc
DfYiDjlA7EO2WuPORYlE7rYY3tCZgnfXHTiaoi2tlX9ixBnohJu6VfgJm604YHEfq2Fv81K+3T4j
6B5/VU4gYY+qdPaUJAebs8NvEV6mOInrsKv0HthQ3oZqgkTv2ucQDjKLG2WVP2rAHWeTuUdF5tbU
N2AdRAm/I5JtXuBj514xXuD7zYc/ZlEGSt1VnXjHrtAMuBCgPi58gTWFNwvIaUO5L8o84/MsSMMm
aN0mlKF1dtW9fCWnUPwYSMLKMgSIZY1LFkRDB3oBfLoDWCKvWoI72FAU1H2ytGdlIvG0JbU8k41j
q4mG2K8B03xJK9tiG6d3R8YYHdnj290+xXJZt1+iTS/ij3VyPM0kN069trA15s+ewddHtMOhbBVc
W/vTeW++EaiCa9ACjzRKLfGx/lmvs5KM/KcBfV419s7691yFHw5TbEpyaWrrIJ5LcRDJyUpFKbtU
TqBqrBva/7up6B/Hm5eb2B3Td9LubKMq6eneykBK7SnOf6HJgqVXitjQsM2hYpjf69dS01i4Gpww
jJFP2QpLe5yA0wosi3REnU5west1f51F4IcOiv671ShJjii+tKVx2va0m+YJD3zeXrpmDGZLqa5B
P7km6frRX/iyi+5+9M2O+nz3AphSp3iAzTBp/Fp6/KykYKSid+i6qEpTQPLcefA5qA4vJlfpgnh/
/beMu9BalpHkkSb+B1MlZ0Fvue+B46WmqbnuOKJReyXh1lvlWYAAA7CWGEDfGQmLa1PFoLg7wu1R
eykWyHVTOiyDiwNlh2BhU1JIC8ws4fkWYBlSLwWcRS72ynPdA28gyOQiHXLINirINmw5iQRwztck
uEDL6V8pba4aQOEUq2GpBOUo88s5YOs92KLDMzAd+NEg5NONVDwjGcotEAU3jpsUnzJ7xzIoRgFs
yyFbjq0pcqzlaLzIq51rJt7khAva0EV02FzqQdJDtGbAk1EFjeDjeXRB28moxzXWE2ls4PNK8K4F
Lp6bcU0o904LmbmDcHUbkepIap6sqOCl2YC2Ai7Au6NEEVfCTJR5JiyJx6LqSqzh+9DS0q8XqCH8
BoKniZnDkXk8iQ22SEggfsRDZqfywDFDi5bAwQkolfqevBa9fFW6stcK3SuI6wCw71/3gJhtGaZS
VMIjTyWNnDQk0pGVGDFzY0uxdSRALlkNOFHSsonEaLelk1IG40CnOyhc9BoDmP6LgXFYDgtKg+NI
j4DhOWxCBqcDydnOX5ByrCaLrSUgek9eVUZO9o6w20wR7QqjhwCn8WTRCiPViZCuA6MwwCLvRx4z
VZcjHRadC61BX4Ib9k5OzAe5IOTNIrMunqBeqN+SRJ/z3CII6Ja0bYq2EGQSakjfOG6CVe20Nng6
agQVh2VzEfKNqdMXi4EVqkmEjk2DxuHkMhYIyQU04zbC8jLDcsT+LzhwJqO3oBY/XrEpm0jWzq8R
uF6yGu8eRutD64DJ3PPrBsUwKWDEll0CXRNkJEtwd1cLwKhor5XD0IadN78wWJOgFertPpwiQYDD
dOfLrIvDIf20hkUHrzSgRoJqxpURpZWRi5HJSyjp6E7gpgJr226U95bKUzIunYRdoqv12gG+jBmw
lW+s9ssm1eL7ct+gIzTkyhp0ltsXnbb+A+3I1/MKP3oUV+MsJsJEMtMA5nUFY/4KpHTgWXnoVQkd
ihbYCaGEl3qB0i/Li614DLtbWGd8xgzRhvjNKgO/3YF8ldrlVDDSpH86GDZ6kvqLDo6ylsjX/EXU
yFGK9zfOsNGGGat04XaAfahhB+0qnq8Q9eHpzXxwbb4zaRwM11XyL7DTWa0aCGIoHs34pghVBBNa
5xVRHEN4gL6xqnRHiSySCo2GNbW4dp3M7VeCXjsAPsNI8Co7e5nxuJLtrI/pZRlDXASHptD5QBS/
jKXSKVVSySDN5BiLF+2Xa3r4A56ABhol9Zhin2wfzcol64Hr9fUlrZNhWvy2nPDYVTbIg4sKnfEb
BqNyb5AlWY2Azx5cJL9YaaUmW4Gmx8OPfy9g0+SYBeSs6H4vPDxme7jKZoDLWxIiO0O0/i6hBdD0
hdj+CkBi5uL9s2Gi5oSxcROkjjm1BbDrX8CtvMyIxMgUVjvJsYoMCCo+67iPaR/4kFh40pZNru1G
eo/eGRUTv1nnOBZpX4BtNf9sm0XyBeEIu68IfMXd20vzvRSz3D1UroaA78UjPN2bnmKZQF5AB08A
3cpL3AYhRtkNy38VdCnd+/0FEuLo+w0djY8ZSAnhBHsboQav5BU4EKzcw+3sYEOA8xqKJTTyf16z
sHMdx7RYUhkO6XUOKyI741ICIFOZvEWfY/5tT1znswkfr2/hhS4rwgIQ2vkwHpp08/+zfuL230fw
ktyqxVpjq9BOPcbBGKb7MHJIYGqXBIG1DyHmHLHUZwCTqsIWbuRkmBEYB92oTNzOvaJzDGCv5qxD
OIhSh1EFyMBRbGd7GLK64B67zbYlpLQ7OhCa2UAyrDdGnFIV/zuquq6CKTd9ixLct+JGF61Rh4jJ
eW/sLOC4RGhS0hIFo2MDb2coPP1UcEnxx50U5x+nItbBKxRQz5TaDVv7TU6TRl7ZgTsDJTdkXecE
MAEpPXw6xURfm9M+iw2tRhTrgnlSMtuUh/NwOFjEnHURlnigkGZJsQsa5S8gYOqG2IsyBVp9HKyD
p0vFCfPQ0hKwfs7hoYtQ985t9EyzmnOPv7/K7zDGORsK7VXjGZVyLk8/FT/cqo4ShSlwGQfPA3aq
EuKBuRXoE08XFZ4EkhCBuTZ8EXTR3VuCkhmXI6G0Qn8nbMHKqzVUr9KFMfOk1pwgHDVDPT6chp+I
sGM/ibUn8NfShUGn/NUlZliSNbhlO47VlPFqHJDU37A/2cvyjG8dpHXW22ZRFpBbNXe/SB09vQcH
EQMAI2SwA562OHHIZwtq4ZUf6y21cp0w94IR1afPAJubn/uAEFYFuX/hGv8t4mCOSzvLpicUwwja
eX5oMrsKhi8c1G8GchKXixkm7iUgQJabcuwihRIAX8SqQt0AGCL6n3kcQ1c84i6t8pJE6WsVqScF
L1tQQgvvd1vBq6wFODs1PQtS6utE6xaO0nrXb0IKzkeYXp3sLTnKOCiGR4P0nvs55c8oWOLHLD33
fpqN3Jel+UG6hw3ilhQnZwZoQauyOuD3j63Pafr8FmJATzDLzdD9XbRsmwMzLSTUa3TyaE6sXHBB
5EymIvRl67H4PHwhkGmYRpXl0DpxovJQ8wnUCWqrSCjn48YUDwezHEGPYIPvv12cTEJx32FuYUDg
4CIEd+GH/1uPHMFlH1YIbGISrQkXfSchlhP8SKkGy0Vs/9KKZq+bFB/ROboB2MhYTP04Z9jZTu/y
KeBPbZvtqZzXlGwjqYfjUl03se5RO3QpJ+fDKtIVMzdhoZ0IOuNq5z6Q+LtReu+kW5TKQgJw5TSn
nheQe+6PRZLX0C4teO/mxoeYVYoMzVP6YzJ3WBQjufLZ7z4Ru6zPg28B7S1s2wL33lgCxZlaKBTF
1nsHT7rs5+nfbQuBp6JtVPwd6wcxA+LNcL8TsHgxpms6ZucfHelNMRzTi7IGOLLQn6eKAfNTTBCZ
DrvPjjjt7Vtk+mlrTRP8Odk8yw8UmtlAk970/RXN5Qxd9FLtRvY6iZ1ckWb1KMRwYtzKWNOqkxBi
aAGBigmUTgDSKUz7lTeDfB65MGbUwvsGEPlO2r9H6OWxeu/ks9fPnFsuWwCHcnhK6etjxpNBb0vX
lqMtzGeIe46qfUw7iOsdtRUjsIEB9DHGQAF1sqmElBJixLmNSmM2jkoM4MPFncyR7/z8skJFp3aj
882ZzfElOOga+hD8EwHUGa469HzY51qRzyXgFB/72CJe8rvmDa3aS9nzOVx90O5wNPT6yvx2r31i
k/6m8QWCpzuFiEzsGRXzEgxE1WJWdipWvCD9NFJP60HFRXQ/d97P7Ddz+DMMZtSs9sxuOMUPANxT
wB8ZkGVE+aB1uhcCXWy8YXgn5czViQ3agEVCaJd0XEDTUeap+dAM77xJ+DKhQrm0j82JvAKl1p74
tfEVKUespVhWiFIZ+a/MO1q8cOUFH8Ogb64fQpC8izL+ttDFtIHk5VkQsabfTuj6f57WkVioYrYJ
iGVCIACaIGmn7e4ynrDiuM9shCqO/iapgplIO86zG2JRacftaB4jgSWT79jJXBo5crjiEcpzgfzT
0fNMIk1+QTqF2HZObuysCLlJb4/fbGM25B78EZKhkrKc34pZ6+ep7VXvkcgIGeI4GSksCbk8E9bI
1I2hpYuS3R9KCE99l7whCXl9g2JkGYBre8M0+65mjlbJqkoGGTMsUcw05lo6N9m/Cd382tR81twJ
eXkTcphQ1OgmAQ2AyPnSAZrDI6+7hC4jOB/sMsqRJaOUfNmaoizxWcgGa1QodtkedzRC4Cx9zqz9
Swb+S5ZYZzdlP1AKtxEqi9czW2DR3v3TQE4/Uc4bVvPmsDrOVdbPTtgVwQDe7VaTh8XbO0TxyAFz
Gv5K3JeZu15b6rzJSsVPvowwv71oZGkk6vnA3PpcJ9nKN7woActGRsGekZiXQbMn0i6+X1N/RJlX
54IBZmxqYktW3Mmka0138dZCMmyVZdqdmIk4lDB5sg88iDKK+Gcn0/Po0OpiRpVBZI2JyCXx9ZTy
xSs8aDE2+1PAsrYUYT2oYF9bPtgLbicdvqj48M68o0hE/5xpxUYHHzy49fbUrLnmkJy9srXI1u2z
q+xl13Qiqq5RqlgdZmehwiGVLkYH34MK9Lbu2lHNrOURRnPYbnyCyYczUNAwSGJEJimFJW4mCmL6
77q20mfr3lfdDK6/RebiIcjeDQGx5pcZFDUt0bt+QBbPDo5bEe6+m2LlXAN06yt6sZX5dElu4uuJ
AZWBo5FabGNXzGbosjFPN1U+223ihxfe2K9am3saqtY40zCn1YxQt+e2Bhbh7BzRUulC0ppvmCx5
PeWsbyBvjQZL71scLlrQ8GMtVNbZzeAnLlf+RyubEuvUgNKSAJRBMUkIyGxbL9WahTcOUGvmesa8
jFLmZgHY7iA2gqqJ8f4DtATXv3rmXjavJdKblgr0EhK7ScwpoVpmTR7jEkbus6Uw+roFDfe0q+6M
A7eSVENiBZO31PLIqlYj+oxSEcSrQowk9n/GvWNtvq1TGJPiePeqCZBqm3VerAync/88kwcNYqmn
OHhEzi6BssNNE73Iu4sgFU1tx3FsNPz76RMYT7YZd2JZmBXxq38oWCwjizRCv3USP7HvT25ZGwxL
lxYi80yBcgpHk8Zjt7wOv0AWX8uotTIhe9dKcEWGVqp1bKq/Ullbj0UqWiaeib13QC6l5msgU0uX
cqet7tmGFutDMZtHD5greqxw/IpdS1QC35oWHghLPjX4kAR8dLm6Fz805BQmcvw3SC45Eakpf6I0
/OMP6uOZ4hehMTkRpYKlR1xwYyX0JWGhfpOSsmhVBejXrpwiMapip1UZeCnwQW0PdJqQDO9A+rEP
ULZSkTEUSbUOUpbkImZ13MxnjkI0y4BabRAorxa3yYczwuEIixHxmZ1TtiUfP7QEeOI3ucfO+bCK
OIyW47RD4F97RBxR2qMBUvWoWOTeo+8HZlhJ4tL8gL50s7v2WraD2P8f54CfBhK6DPAqy3ykJimm
Wg+HtwqWu8jntunuWa6P/JXP6+LYKkBn/sCwHoTzIk+A6hwZihgGMfdLAYaGG1TaYuNUd0PoDYJl
/kU9PVoh0iHip6DsBuOnPxCLLH57Xh7CAVeYrzjUgK+IhOG3c5j8GvzmVUWOvwnKCa06+r3eU6DM
ah1Na5wlLbSAQQytlhmLPr2x2MAsHjoZ/2JX9Kodj60PAEACNk+aC5Q1oVdWVVvnUN2RD/DSUHNt
Zi2+3ge3BnNMahdGezqxAvr58EbAbntiGhMB787+iLd84hQTNiHK0Xm2l1UqdTn0SajR7jcaAOim
Vh216f6AMF71pcH0n5pFN0KSlJ8hz7pnbYNnSqISCNcoi6ko4qbvVF5nyLmM+skh8OY2rYiIaSlH
OvKUnzT7+Wlpb3W9w207Ylr5QxwryScx95PabWwOwA8QVu8eyBdsZhtpYDsoPNBEduH+JtdFWEev
trsOGln6iMP8qrDBC6YgDYQHo4xAEMKsaWEePDpT8BVqd3C/X9hTHO3ASwTuLc7hb90tLHqttFLH
66G6sH+l2onQYaILWPXclr3bXGMWgpEAVq507dJBR3wLi0uEjWxDdr656Hvsb88MajUnOF9h77io
YtgzLxCWSttHwdYKlxPC+nxeXurzz/jDKcanjo4bMgMxTQAD571IRWspAhSLlsUo8ieUxinS5Axa
45Z3j/RjCcnbVR3df87/k+HQcpBbfxiY31AdBw3rofggZqMf31psrqTXQxC3vBKiGKc5tNirjQ7P
lb1FMpsV9Y1qCBJXrDEPJzrKljefYN2XPK14VF5cmN5IWYDimLa3Bo9Vrp7ZqfuVWyyv9GWwNQdB
7grkkFLlVYOX0sOsGEIa4dF/kK4Z2cxjMbK5RoaRSm6FQUe1LMZSebLk/45WzCgGAJWCl11fcGeT
P/9u0ZXrNp6DMPDqkpitVk0B1hxMN04ZQWWSi2U4ljNFYcbtFp9ABaDpcB2ROOY6wk1IdMn84Xkl
ZA7ho8WZ/the5LcKdD2wUkcbtgJnBONcHiBwsANpfuRRljaPQ3O4/65gM9DOSSMmCbA2cMA2WNLG
/+CuQzOraXaCEZxCnTDAbe3Vv+PWAa5k7KhdU0LBHOBmvF0wDVek835KKA21yhjOBKKBLX6ic7T6
JqwWo/KJn6kHMZm+WC1DEQvfQtbFsOH70GfdZ4/fSNHpDajRDpLDqmhDySDF464ppQo1WuLSmRUQ
c8Ry/3v/hmjBo1oQDGqc7o5uweuMWDXap6EqIRp0X3eUKIZ0u0IXLkS32m2BfMormG/uM522JQ1b
6JgDhTjmK/cG8P1ZjYa4GeNQ1ca7d0H4rcmVIlfuUicAMvZNGIrWONNqS9FTooLlOCuSI3N6iW3O
Ppak8BZZ37DD7nLNUNn1RvQ4LOZlBZWNfihzG2RBNx1bAAWNnWqnuTEAfXOy2o0PchWDXtXkFB8J
VCTIoQKXZmd2Noy8y61bzc9wk6iQS70g7n2kyY0eCGpq7JOiEqLiwI3FNkE5ruvU0AOeuTfmAsak
X9zep0hFLtl1qhAFMfjCAZQXN0USrMGuk2fOxiU3ANtmL/b6o7To9flwWJ7b3NR6D8qFhmIhcoqF
6moKhI/Ycw3ygZCFb5MCGQ3MU0CfKSIjmnpJCZbRzO+yH+DN77tz69kFzXX9WAjH1UVmGtRtMqkI
7lVt/uNeR+i2sXo255DCzglbWJQDXki7l/TOD9DFLl2R3nHLGe3z8x3Fo9alQbeu/22U1ypnTMdT
39JCtHuQB0dBn3y/C4mHe4mR8y6xNUV2/XH4lDJUlwsUuWrMMen1F0Ubx1755KvdVBIkQDiucGv8
8R1QqYs7KoGgLKP7FBWZFjdbvsGsxPbxDD+HJPkx9yqlZQZGH4f+XX7qcfZrFepyES5Ys+2BfJ8z
SyUKKQymK8Wneko/+4JkcIb88X0Se8t93hLLwqU8c+NYhMpEXx6e/E81TDF7PaGfG7sAFN2Dfs4/
QLR0mrQRsHqZc+LpBH2QtOx4b9e4xIKzyoFybUop20oXMyGxqEfyFNbLDHbv9ckDJRTT+Ygj9LXn
MsSrNsSpCWJ6d0EkExTJ5NNZLpRAb4vnGGxhq8p+Yj/1cruwSgXv3hpj7NNIImrdCQARnu24jHBR
G44hnLwMo3Kx5D7JhbgktrwICbqoLnWOH6cp1CLg+oemR7n0NtXsl+gg7a8/sT67KZDmfPl6jlPH
QpUGHsRLlKCliuFAtXUajqhTW60rN33kY3NxL+ez++4orKgIwdL+4Gaqlj1wLUL9X8HKcQb3KOgU
FzfhtrNzWqxDsRLN9sU4MfwH2opJc0/kkWndPDjvHrGoL35KOLro2FtD1O5vpFdisMCm9G654nw6
SmabpW83TGDbP4Y7fXgPerHi3dBfpKtRGghfYenPvOfU8KCkbY5/Rs88FfF3KVrXXhv044BWAozw
lK6bAw5sXQvxNn+aQ+hNCrWsjW6KdB4xoimanzi8+OrAhSWOZBNinuLOWR47t0PvXpL0Uemna3GD
Dx9VxwsO7uC/5/ZTzi0oQy+eK5lEdzm4seCTV3AcOJG8F5gudhTS8mrApYFsZiYEfAGZrGgpT4VD
oa3JbJExRWUzkAty8q+95AP/mo9sE+bnaTlk+xX7mBnOWRkHjSG4cG82lygIak94wIvfqtsl0PyQ
+biRL4c6MY/aE3v8cLcQft4/l0eOukK/cAjFAzPwcJUgtMNc+8TCUTtHlr2eWOB99beOLMz/qH3J
1iU6UE/llti9Wsg4Xl09NvqJtep3sD7gF/7qLjYp2iPOCmxd4J4Bmwr5LNp5VqT4yb1uKIGCs7vc
52dzKNJKKbrMgWZtUk/pH4JfxtiILpbpaDn74+z6CC7woQYlyAx7YBcu40LQl30QB9UcXu/U0Nvc
ob3kvQcBRdkSetRtDKh/du5gEwg1sJ7SL1CpqWnszWVxElqAnrLfqO5wQ8QhnqaAbbDqQq4AtcdN
1wlYg0WyEUL80u1Du/1r3hD1geRKuy2ki/BL/lgnCAlkYMHuz5rNBnGkJtaRn9cENxf/OabAKC2O
hooHx6BtVHM+JdlBaTySn85tbmhddq/YELIPZISRxWrrQ2jCr4Wn/qbZKMSX3lIoRn9h6kO3a95y
wJAxzZpyXppJNH7aCST4oI6PeBGVBcpV4202eLHQ9DdH7v6xV0ynD1mEVpE6SpP21kuJnH3s0fec
VfMXOT7h2PbcMfp1q3Fec2Ql42x7YTRKweFA0Vo/AUpZD9pfSH0Zpz2XWphkW4xPyWP/I6R+sty5
+1D/GqVSBPRBN5LOEeOHpj7oeaZ1SmbjNFn8ELhm5hqtosjD5sFwOXlXW2tmtTlvePWN/JGzWpOf
IgyYLCwM+knPBWfqCyM2sjKNbSkHeI4W/1ALXmoE1fQCjO5PvHd6quZN9H+VDCEGLXGuemQODSJo
pN3cyZHLL3coG0ZX90ZmnQ5RHtUJN9pO2FN974xTiqOM4zDBPHLPpt9BhFOKyCNFXu3dsVOrcCKT
4Vf7wwgrRlbnQbTuvK+EAeb+8WUd3g6hU9jwTmIgxo8JT1RQQcLpWnCpzhZRuOTgwuON0IHwHHQv
OfllxlaIQgQbHvXiLEEyPIMqBwz115qDZwRacD9nVFctlsQfQAkUz7p0/Zh7UyrSVHyE5p/JFwpU
F8ihQ+p7wrzMQUdYDx8PFk4KCxV1wGRo5ZLjCVqMnc5rfwAS+GvfZVtEZtRr0naAisuvUNmbkN5W
4sXuo//xh0K+c6ORPcFK//G6XGjq8U53DDL/uNpvy0kIXZR3XAbKdpdcs3zPBxpShP0+xBdnr1Cr
YvDFFuil5yo556FlJ1x04GEquh2jlzIS481txIvF+y3un7Kw30hW70rH6WqBeeNUwcXo0qXBInx9
bfkfOo3fChJR6CloJmDXki4XbRP42sby1+22P2kdeQos1K0g+7GMeQ53AQkJr2no0y9YAV+BOvk6
scfdqexZGTrVtJCLIv+WUxRA17QVqvmTyrgYZ111zLAJaWINulJV/BhvuJOzQoO6cFNYq34srCvk
JxaHn0zw0vxkNMYgJTmhXr2/xmHM9V/9Il4AK/izmsE57JvwRfCtpUTSMtYX5vmOgqHTqJlL+o5e
t035px65+2WIS4ipfPQ0Tt/Ke9w3m4oNJnhEiOOzyWoz01uiQiLkoq/L5hdzuXbprRz69OOOzZuN
bkjAvtl3fgaC0fp82ZjxjoskYhDLAEgS4hqtTjC3xFkmPDnbqVWpXLhLzgFfKuhOJHHv6z1ht4zW
KupLK1sJTkyvBmRLirJCVdVIbvX4yXYVUgifj+8ihpfTiX3iKWInJzhkxN10P+SMEPkQ88FeYAe1
d0lVjsdkkdNRkE5G5li4kK4Wox09OaN3FDYeSVi1SdvrlqJnlaXA/7svS4+ARiwHwm4g9H/mrppk
MHCtILZmyjx85fjT75dHd1UkI0h5OUXYpA2+KBc6LGULpzn3Mz288EWs4w0BPPdhWsp1wMQ+qOta
0blLIVlY0GJXSyn4C6h+3UBhG2HVDgOW0jdRK5fTqq4sC4RK9SgdrUHDpCBxwmMxiy5RwT+/F09O
RiDYC6vNZWqvmC/OFjYu1G6uo05su1El8pJkJRSLkR+LGRmonQydhNKOlKFq40WmJliiVOXv29Vo
qGfKfYgpc9eZu0cVs4biZQX+0crguTuyJ/dpG1O0SKGlnt288jmOuw7/ZDDemqOsaAB+auf7v+At
6CzOj+MuGxGRX3P9NIj3/Y2bw9ufBIl8x7TZny7Rxltoy1RUTo0fdrevLHSmzoGcIKi8tnwrg8l4
m5kd4/F9xsem6iFwavKZ0ao23Goen492xKzrmNJQI6dU9uO/rQ3jgorqO0a1c6lsAQX65zAFijOT
WCbCQnpZSaViFHOcxMF8FpY8obXtC6xz+iX9QAr18U28WDOZSk381nrlqWrj3GGSKir/oBfc5TBa
vF3T3FyMKR4AZUwrEUD9lZ0FHnlezOrRmlp1SBCgTscisLPK38ee79ScYNueZqMQKxD4ohhDxpaz
1rQRcBhVjeWp5pA2pyEX5VU67XnIYxGg3nkH/kViSX2rS6fxGlo9UKBk7ChObS4Cqf5rixEU4nna
bSdMuAphUIpEmTOrxkZIzuNBMiMgeuU3p3i4JLq27YCCTtouPcjbj0JDCK99fbEPFpxTSvnfQlIr
NSSNFSr56h/kyghJK9guLuNt3hS8BWL1PUotAULJQx9ntNyjO3E56cJuJ1t7FjightG6HR9pq4g6
4LZaK5glHWmfFycrVI+sFzUfSwqR38JIsNHYmK9c9UZw+PpJy2oPRFcC/inQ0EVJKsPV5monfvbh
0hq3TBwOJUC8t9jC09qlf9F6gRr3oPaTDuvQB6FJpeu/jgjIzmotP5dxRjBmqOArIRgzHa2gtFj1
0lioDTvuy/DHPrr5sed7Q3Ni8zgzU2rECTObpTcWfGtx21OyJswi3Bd/BwgjiSZhsYpEb10yI6fE
IjjIQQiOClZP5PXVrjzCv7rtjgXd2xnqUhz5YjJRJaIAilJNpt/Z/E4cZPLWdl+Cjo5pJesdJWi+
TX8C7n9Yg8C+h5pgfj1qtp1Ihja1RylxCCf++4ShGNCbPkIDPiuqBYfSTFrRg0YT8reua6hOyNQj
4BVm537Xoxr5jMUk/tBzKgT7516JM2DZuGApmBx5D6UsMlXrSQpkr241ZzPJ1LuHePHuTNHgb3LH
nrI0j4AndPa84biVHDo89zdV+t0vvYRozZaUBrLPAZ807ZdFNwo3O10KhDXEZ8RrTWyBGb22efEq
Hu+ob16h/gSuMXg/x9RttJJ9LoLhteGQ+Hr/OwP+xbeviC/qpaw9GhZc2nkNVu/EcjrurGfzTU/F
FuNaeg2uEYo/CaWRBUMOiT9v0SBlbH76nVV1YIYVn7ccNkMcAy2RSth9qCfC0Bjd/V3e6m05l4oj
Ig9/5s1MjGQDdat52hBls366Yq4H5+iCqz9js+6Un9ifUkyIa5oXy31XnsH4zXF2b7C5srlMUWkZ
zFwlHFPhqsUT2VC75Tzaust8SB+PobtHF1WD5FiZTbeOBZWXpqQ4qBMhY/Sn5FDBAEWhfP0uApyu
IK8puSVtrdWlxUmWzBev3h7NG/zP3bZ+Ldy5xbTTlksCUCENZFuCck+XACRwOzj88u6371WmWsvn
nKuD7tFm4NG/PhZRf44YzmMkwyrY4N0GvjHaMB7eKzLaeaDVXcYuEhI5T7K2XBk/SGGIc3F7nAWa
OOhN05hpRpRwp1iCCHbWpUHGXz590yHnZCx4CkRL93pPBQt/+xV1Xn/nq4sH3ten/jEJbLvkrXRy
ddQxxLZsp0ZYgvYaRHq1PlrrjV/cngfkXnv/xt6RdWAP438TC0e5UVGSrQa5Mg/OXhlAxdwWJw81
6MY53Z1ke0Wpy/8Eqv1ocD4ETDOS07YURCl8Mat1+gmnwqyNcQofMtFjZIeituILKwjNU6fyhhP2
iwHGotIUdNSBS+U59f057wUyKtwB6y14xDKK6lJq1Uh+HUqTKpoJ0I9SradXaxkkCgsmupWWSaT8
GzK7FFhQCRdN07XFK4sz7RF9oUoYYuMPRX+i1sA9lEUp/mvG8NJftbpa7ixGkWcsB5wFOoEBuIdZ
2xe/EJNJWkiKx00+CIg1r8+5awkiikSKnpkDw/H873SeoBHqrgh1cv193fh9uwKv4yuIHUuNSNwU
fEL51eiN7rKDhhonYJbXM7cyGRJOmiLwP7EaXWbVDR9Hp64qsAkxm0wcVSIm5Kt7rMwVV0zTxnM9
FrCWoeOdwU/pisYSmQnbqYPwpdmgE/DsggMDVPilRaFuMUSwdCAxR5/jpx7v/NUNAAw3+JySeSu9
idzh85VC1QbL03v8onrXMAaK51WZoMpuIoA9zuink0J+7sC38M/Lz3bANHXSf0HFFkOtg7i6f8h1
AzcJQ4RhzlwRoXgoZURH/1OYqs0StGdHeTOUyiVgMst/BCRz67zRDSB9GDAnx2/0+quNrSvc9pI5
g+OyCZ9KHK09y4bu6OTl9TshSnk3jlTjoyGJfKqU3v3Ok+ITpcPDptSzcScZJq2svdnUXL/nMzFk
mVr8pG0NE4KpZ3LraEz6eytniFGw6HBjrVB6tbxzcJvMy49PIX/hhi3Y/p1Og34PIGyoczd9p7VV
EV4OYDVI2y9Uv6slI4oMbWULzfsxDwZYfSEydfCZTyG914eSFEzg7B8uiVhSI0gUNxdXgBLzmcTN
YbbmPulfFc3FRpa+oAAsUP9tNc1EKWaIzTLcUfb081KfJkaXZFuP0gK/SV9nel5BRAtazZ0rfn51
WDJtimMl14kf+DEG7wJ5uiCNiANRFACAyjmpSoyxdQV6AQOFlViue0DZkToe6/KjV1ZuRBRcDP8C
sX+eAO7D4W5unaTST4RdW/KOfPsquCO3EJHv1/mlG16z0XA5yGdT9IAZSqJ5SFG295hrxGlS4pU/
sWxDPG4LgzHS4TldG1PnPI494t8wl/bGbSRFrGerVHfUsW0xBArfyptbi0yvHwiizE5FqLOlWubW
XhTW7Hde0++u6Sgucb7rUZVrvVSyYC3WqBF565eIRBfCGNVoiuxb11aPnSs0DRHWpP3h5ts2tPgB
Y4kQ1bRVldQ6srVLC+JPFaj9Si7SNOTPsXCTz7UyqwQqmbz1chQVLO+NBGR5we+gKUzaAW9e+Evr
LcbGA1L6wmumnDpqcXhSZO4iC5eMyQhTz5mqN7VOyJGe1jSemeMKLcQYqqyWkWJVBoI/LbKAgG3A
kHtX8cdL3w5oewZrz7kc+kkX2nzJf5LsAX0ejvoSmzBdPgoVDEq25+wrtQ6ndVdiIfwmBQektHOj
FFGKA+UW/kX8uJwfIycR9TQBNpBomrTrDK5Mf5pOZRPByneih9Xl62MEZv2MQaZgjXGqKp8Rdiv0
4zUpgnAE+irKXR7VEhg3/xP1b+Vmf/q/gOMJ2PbZ7PO67IJRnW2n6otj9kzeMwuUr/yg5NMYN4Jd
IGzeGnnPkUMIr3/dLIPWh/z2Q9c3H2N+EIUl/5naKvUyToZX5pj6dcYICycdgrU3p3TWvkToaP/b
6OnxHp0yDXebRbaXVh2YoqED2T9NTp6WDcO54JgNCciHQq7aFqrRDw4TeAABU6zR305LwNqFSCk5
dWjTysGy0JEt8SXsLwivIvIcNSO6+Stb8rJpTRg4tYddBh1ikY/OXiBi2zchFXpkTTOneTNYrWx/
NQr0v6VFv07hSu+E+LVwwcjmhlqf80pcobz94Hc5/kmUwV9MpedgQg2dSd6CNKF/YCvA/cUzaHWW
xKqkzZCLcaBnR1clXn57HwiUw5V+O8fWX+hm4MhwH7gqffAgBJbNeyh9ngvdyYVQgPDntdY5BrKX
fEyb7ctPJMnvCNTHjTpOr8ULjxlKOgJi0qDOptpg1VIXPs1Lbr1JRXNRT2UBf60d/f2QsXGmzS2a
angOEKxj2ca+GCtUIwZeFebWVMFLecmkRD8PdN7E9sLG1G6J9cvc9mL9ayxQZoCTwNgS5WK3/mQE
cCLAtq85JcvAqsCZteorUhUSJA4hEwAlALepbRIPf2x2EKkyfMHh7jrTqaLITG3qOlmIvg3oQxku
kPJ9f2O4zTQSAO6QKD1lTOEB0OKHoX+H8+8HxhRwqBqfLccfGCbsoQVMeuULYXh+qGfKDkyo7Oos
1r6nHiaXmxNaIYChJONaCVuMZTxgQQgPtP44j9+l0pJZNMc0Io9QW2NN46ER4/r9lIRXaMwy0VRi
Tq2DDvnulJ/fvyHW0pxgOjzRjrTDkHjGSGsA4vOGwNb+A4xenIomNMDc9qzsCa8K9Q+l1vVwIOSc
sdpVG5C5D69rS8/qWyGy/8MyoJnGrF9P6hjon9znIe8/v88KjSS/t/H/KAI7k3Neubps0zYyVC6c
+HkxWwMmDeHrHQwW6yfDgKfO/4J+tdZWyosksY/gfCLM5eKdWp7cjoh5J7QtbD5ZnT+xbVOs969u
QXNiGOloU1VZvwsQ2+IapgTlmE5UDgAq6COaOY2mQXUQtlWte3N7/xmoilN8IJV1wW/BLM9PZPUI
ayesRiLZilwlztx97aslgsnQbZ+J3UlJIig5XyJ4kLiPljOWsdrN0ZWLc0SUGek5eh3Buy9tikJS
wQYNdQojagmNPex4kuv21R4/Wk2vMaRiWOuRSezUm48JoydhPWy82aW18Vm5y5Jg/5Pry3V4E/Sy
n4xO4hwcrsPxPTUjifXJmKAewu52v7C17sZ4eKIv/sXf4LQb+vkYuP6EL/y454pBHupqeteK7OPA
f6gV0WH7fOzUT5nYMWI+TbDsmM1vzs9B4yz6hNe/bYvc/1hur0v47m5ws9IuHqzk9yr769h7RO3t
w5iP8iNAqJQlnhFkpCwVIbxO0jIAucwW4NW6hWhj9imhi5URfdAAMfAKreYEysGweOH1mM9n9HRk
PTddzimmEjcdpKcDmACEHlXDr20SoOfkPwaQ9kr1n6I07o0eVuWzn9xlkUtfu193egZrOvHlRf9Z
RtyhPHoK04Jo3XqKqsdrbPoqmyBLJXcOvzSlS6nv8vjgZIlTE83XN1AWcSLaLxlKA7acuW1GtIO/
LTIgjEcwmSwyCneLVIBXergSmTgGkVX8BCLsrTB3ta5Kn7euulr2GX3DNql6H2dAlDj9pa5Lt7TJ
ReS3yvZz5SIgP2HvCLgPtiFlTW8hgGMCOkpmjj/Cb9faHuDflq35xExvIDFtYtABZBu4GjX8cC5+
ox6/4PUX4ts+Qap9MSfnwXaY+t/fXZOR7x+wZU1wdAo6M+GR2cJdxtZ+iAsxgtm7/jYTQcu/Ksg6
zosQQ17XDf7c/KIHl+mkuRWWS12hikAdDrCUNgkwxGAkurfWtt3UNbNyd+VPLRUMGXBvuf5C7aZY
zRpYYCdFMkm/iLz8IYlN+KAX9MhVxmmufKizPVQ+5M0MBrraMqPDjoQ5j7vlG+GDcs0a6FQkJ6sf
UBs8H//hUCO5bLP3XT/9vlqg3JUuYQzHk6xcbaLPHZfKzq8Z6m0CsHzKGzgmcEuouFba9f2oyvMh
Evg+PeGNRckwsDAwc0uma4gN8bfiLe0XC/CVN6Zg0ARusRHgciiiqQpgp383BkVmEqwFQhZVCOPV
JYyf/5hcieSMPZNFoCSTkgSiYbrXfglBOPV2KQJx6ApyLCD7YiJHT+k0IS6wHc1yLPTVpZ+CsSWC
suY6GRdr/zBwzcTQCGO9JRWQGvp/GDY5Z3g1QqSYNuMsiPToBC/OSigrqCi+qngDUdSWH+3jepfY
yIZat3BXiAdJw4KXwSgqWubS4mt5yog1zaKXw26CPrkF2gUsQNtU0l8ldY4ao1U5QN8uumE3T4g1
azXEaS+7GTSzqCMgA2unb7gPqxVo7tJ93iTYHLlFBFDRj51ZE2dbUqcTVYHBgDgUT900JrNHcQAx
bMZKM8RiqD99tg/7GtmhQPFQ+tLuFdRzhYIpFWqXHD/71UIU95KPSajNl0lGIc9VdDbllB7PGLoY
7VuGFTgadNVXkvuBp+VDIt+egF1vYqR7PIiTwcaKIvVDcoLy8iOLVVXpuW1H8a4zIt9lu8emQ75U
j7xAkx3sDsGM55Ib8zEjPOxDtifVUE28hHpzRa9PeOOOiLrovRjpHtms3rmLXJcxplyJLHwC16JF
lH5pAnmZbSqCEwCJOhdbujeLKQIK/eKKPue3JD8JA83aYnZ2C9vgY1QwejPge/jOWsHWrGLZG6ch
SSthfPylJDpVxWPYTsYCzHZ2fELVtuC3FDfEF08PlKWaQ8xOdwlQ6jM+K+vFBZLkb/+4mbfl5Mto
/ah709Up1eMw5rKAqVD9+Ns3D6kaFT3TUFjJ+afwdkci0Hk2LdoEmoILjN1AULKpcesRPSXj6WAs
ARKAzPq9lurkBOQuOWzpG3nPLU0WLO0XtpYyiDNYpGJU/Auo8QUPhiYs9RWclwPU1/QUFOmiMhsj
ufvYOHeE5JikgbA7+g85whu1RXgqHvWCWklGNrWluNImM6zgPVCSUa6WX00sO3TCpJsFxMgZyTAi
CFCT4qj6WYSYHHLq/tLMUEVa+Tk3h5OPGuoJJnbEDHVtQFdqqmjrXqN1rizk0/wgJAkOFEe0voM7
BzihNiZ7BhSDcXRAc5IcSAh3g1YVE8RRKMjjP7VHHghJUZDiQVduT+iip3nf8Wc8K+SQ5x+4CRqw
nPvcXazR7Gb2Ae69m+RYsSuA8J7mF8YPhHMzj1g/205xRmFMdqIq15AwZzbFZNtP7fxQC6ZtLGwB
UA4Y8TJ43pwmFBvDyGCkLxkoacGMRzoQmdr/5grl2I4sNonViD+zNLoglKiGKoFYE7IC8hi4N8/R
MByzK2LQomMZAQrYD6aqW8iQ6ApjainorunghkkqXoFGbMrm93mHaUbv5wvuN6NiuPNJadARCxsi
y5grrTO+OHMm0hIICsv4Fawt0OO2xVGDkGcJgJ7tJGYQg8XarpUXo2mUDfxL5W8/xUzOy4TyidJ6
cpcJqWiPXuutYJS15gUhMuyHxFTANvyStGPXA4DY5jnqyDnsMA4OLXv5sMQvb2ZcvTKbHjpGX0PA
cINe477nLmv9L6AVb0x5b2QuBSOcc431n7oPP9x2cvHFKsrKe2m6fnVKnuvDJ+8InnBa5iaNDupY
8vxGL+o5Btj4Ul9bAIdNaXbATdoPt+df9D+NLHJlZeFxg4BJGzjUmeE0QXfgte3dC2KOR/MVj7oL
WDJyflSIBdtQL9DUq9Ey1gCIdj6GN2koqz6S5Hpa9k2YpdcxoNfF+fniKtaI+6t+lbOzPdzH/gR7
T5xPtPvjCEVS5MtLlICQQWb7xQmoIep2oOsTWkQEx/rMHMCumzzG96+3LtE12Rdmioomrlb9ZQbD
KBnAkH3u669ewENgjXYK4pf0/eVANbTzpSL4GNcNrxv0ASQl+Gj8HRRaBHZBa3P7GrENLrsRoiuZ
biAd5DL7fCtqDui8UF6+yeLQj1x+z/L7F+qoSD5e7VC7qej8+YAKoVv42kEOHPzVK7ChD6xZqSJi
G4apV40urickF61/OKj05QozgC0+myuazP7kbkIlp6tjM8TSjkaKHsbuSkt9zuuNSUA36d0KJi/l
m8o8bi9VFopmrenwpaPo6dP2XgEbH6Y5Mi/hoqNrB0aJZXby5lVv79Y0JnkjWax2b8GALnQdCW0F
G4G36EbHMAhvGB06eBtwhzK5VrZ86IYk76CrvoApCxJwxzZuWmxcSATCXuhPnGEethiZ77pKdsuj
qPqa4dVZA0+kSsgIot/AwEdEn1YRPXHrYr2hcODF593Bm2ivDTQHcqT9lnbaKt/vFFWxkFSYnUMM
k/g4CXrPaSlMF2d+k2CUzvBWsYehytk4dYn1WLVic92Ylpr68DsyPSHFFkRpLrm0E7VdYGZ31KAM
lAkhI84rOv+dSGNkfOvhIN4XZXKJYyXGl1devjEVh3FtceRhtzH+8Wt70z93dQLbgusy7TBW7p6D
C3rD56WcNigpiwKq3aDZ2Ff7Zwjoe+G2ja/m9a2lnKF90ZuUGrXNj7o7Tyx6LwJZkXjld1z2J7mo
IB8X8AwTTUcbPPpZXCYiQSpTdtq1Pw+9fdBiYXc20Ry2k66W3N1VUpKA3vIcMrpTUnjH9GvJ/Fdy
WWZE5SKcJ+WSiiDxJ8B37+0EHVk1YLAUGhIxM/iH6O4SCG+s8UMqwnuJOJ0+pZyXHFWIjHsTZ+Lz
ADysuyiDmRMbNExcA/aKrlh/KBZV2TGdzgXCBUvr3hBNOCRIOUw780C1SQMHNT2tUb2/eiYwt71V
Xf9mhs47bioKmQGn7Z/gpyXdMFtv03EZOGHzvoWKbIgm9cWNLC6B6vDHwnaWHEu6ZHwN//BhM7hU
liqZBHcq/n0bK2KSXrFr6slRfnFhLT3BbrPV7XkmtrS5AMV1+csTVpHuNxhfKU5LVdtUG/TexD51
x6nnWVPm5ap7Qicka9e9o4Q8gkCWkBDSKOTRXoPu1K1Cb0XUnsx9hDscJn3c8pm2V8uA048JEeY9
IoGhJGoyWx2PDRuxFbnN6w15oK1eLPAX3AcoF++4SxFgBaLGDBX53d4a8IS73TzjvMUc8K26vfw4
97ce9ZM2VDWhzDtnE2QjAvegXcuZpc1v/T3aXuoEkPhV2Z7ZJq1ATbc12kWzakJkoa/IrL8nckE8
zjMOgPSGKtjSSOqFSuPOh3unxHfJGuP33GQcx6ZNMnhmTpHNbq5Ycw/hFwQ4GPAGSecpuhJatedG
kqCb53laohkJ+x5UK4K0ozjq//5oWjbJLIDEdYTbBzLMUy394D0pqviRCyYiJzWNzsnmRVd2JmPp
ttEY1tZ30MydDpada2W42VATJY3OE1jLzeRWegmOtUPtzpJd0ZCmQMXI5RQKkx7Elp8mrxqmcGvs
aVMxE+NuV9SP9xwD2It7qeoq2LpVm+7kb9Ob9wVqkTQKaXMhPwrYM1sBNuDLff38M9OWFj0bnFFH
sBQn/miPBMHRajtuLv31tRM5t0Ya7WDYvGvPYbLZM9Toa2/hCSJ1lf0vk2l9c4L1UTsedy3ou4cg
vBCUjM8Lu3RLt1AiSMpR4efzOAFORZWTZQ/jaFcoht9NO3r1DoPAO1JU0ilL4C6wKOce1uzIkhTz
yon1LbA0PZeSgdZ42f3FHV8QUPJRDTGk5CmFtvUk16HAoIfMDRxocPp+o3QXBwUcQTPnI5YVqy0q
tI6HzzwDjHR3XYbZ0gu6TwFjUTisx1eRmr7cUP1NLEcGRM41vr03GEj+6tY1WK9A646xHUct0Xtt
DE9KrEriMzPCoA1Ukhm0YXpGByLwBTHjRphMLTo/Jb0Jw1nKUxhk5YQqaOjW7jSCabv5hTNCO7jn
Kl/q2d3B5QLY6mGcUmTwqmGafhp2vtC23UoQHMPG0NdnZZ068IyoSCGRZTG52yeunFMrB3TsQEKU
zJM7H37QmpnqVGhS0Y90jjKDXoyVBn9M47X+NTRqTYUcEoPu9nVc65yWHhuIIhV9wXVYB+gIWybS
/ainZe9VRw+vOA4SpRa3zbowQ6G22x9lvUb8x5tdFkZMi3JIXR0eX5RgeJVGFyZYdfvS/zCeoHtG
DhMP7W639IUPNZ7bnyITKaYsuQyoU9ZB+8CKRB1Bt5DHrr2rUkN2CYLrBCOIXANHT8T2iihVsXHO
x8Dl8r4h9qqa2KLIjbQsca8YSXZ1A+zy6rcaAwfZ0rZMZVvd0nOE7dNqjEWt4Uw73r4ag6M5bSih
owgc8f1njkb48zmRRd09NjHZGzoEftCR+kkslLIS6hwegMlWILH/eyrRCTGi830Qztzv79v8rGUx
La0Zs+XT4rdrxFpJUtb9CKFUjIcI+Zwv5DZlgg/lIIZ+/n2+nBGfgzGLnNb6fKplQ+rWIgLm7u3B
k4jVyc2WsQhsvuIiSHDUmKXYZvvCfu0nSOBEQRa646KUcdZbpaMcatUgA6Td6iFbCuBns70n8sOT
hh0prI3TNR2n3QPRWFib0ies9y70sloNJkhhHhjP/VfCSonVXfC/OgJztr/fcTUMiVFjDnOQXMDv
a11xWy9PzoAjBXRsj2NGesxY/aUdLU3cbOzROaQG+FnviPARgsvNqN4Xa2zLJRlp0KOi6Oz7ihR8
l22G5ejQLi8RzM388Ox/AsIWdkhRMXNul9Pru/3mpzSQL/jM7OlTLBsqnw6i5q5opg5w1Zx9KmBe
/RDFgbqh1nKctHKt4SQb1YsjtlXCWeBfpIBO9xpkZVr8o6oVz6Gbc0vhVRXk08e++UG37Iur5buh
b/suSVtLtvDvdxWD8rk8XX9AjkDkVPNLPjJABOhG3Rdi4m+EUzBVA7nWK0LgpX3p+e/9VnSXQ71n
qpJwkjsWyO28WLR8aODulN+cyOPsCd+ywyEK6lh7z58qcK6m+jkG0kwgGgjk7Csu8UTyOt6bVRYN
0G3amS0uEAfqknvqAUahor4wgz9xAVq0Y+zkSwGA8XZrY6XhIgDF8atR9GI7RO8pG1e+w7Yj/52t
prfHGCmWlsCu7TuMVbv78YVfEYnodRdFFbKWUal3ao/T8+QHvijXzdZhoK5je/Hxhx4gsahwBJQK
kCGnKUS31n5dZCAFRLkddPdkJ3ibDOYVwvRpJbbQwAP+S33GDhm1F6CWr9MlLjDxBddhRuNZuRcB
WTmubNtrr03whOrwTrZC1tSdB899evnfQZf9nClA5sIIF/JnFXhkpazV9ptp8MNs0eUS/o/w4JoU
i/QqTv5L2vE5uidj6kadeK7PoY/Ta+PHjV9Gte0fxcPacgMzQL7tY8sgGETbXCBcWegzmadQxb2R
OoObylIZSPz/gLDSCullBmZ1JIbaV417GI9FP4UtgcAvGDWLGuJaN2wUQg2VX/KjBbVwTI5oxmDD
O62oe9B0FGpfwVlEDHqgpdUwsj4wz3n5IZ2jxzTLCiMbaNY1WEzrEdf0Re3CHbGe1Sa2yP0+xb2m
533te5cQ17ueHH/liDTJr0wjhdiqj0yMVf/INFgf5CAXKnFbgZ3HCze7xulkr8HVCGAcHEXQyKLL
mZwYTp1BfmwzVF/klcVQ2eWW2SJDT/gL0DtzKJ1EqGBevsz6BRy5soZg7/wPf2Nc51pqyfXxRcg3
yyBI+jSZ7Qu306KYN/nGWSZKKwLZ7L1h5isKAXBdezrbnpXaR/ixWbAWEeDM4n1hYbmqkRFUOmWC
Qjz6kQr7EpWNwpctePT3sB+QqorZcR44F3ObgtwmuPCid3kh7OTmfe7dqDKFpW+5d/GfzZeb9GXi
Oug75y4yB09Hv1bfG8t0y/WC5luV63KMUiYtxj1mN/Wr+Kdd2iS7xPCj//IfiXjfPUTFCVdODoo5
30cNe7SA8rM+r7NWNhJUII6ePDu2OCMJF2MhIBH52S6Ahrv2zo6Y58BmAJsDzzyRsOVnhkao+1f3
LzohecqcCI9PpHYUWrSsqBmKgvQ6lCW+QPwWrHfVvkxsEtj5jpgsi1R3oGE9j3ikoq26wJdDpLgM
klgp35vjsBawB9dABBzITRU6Z1kMlOLEfqt8zFC80rpV8V59WjYTS2pSMhDlw3LIdZ6RjqJb64B4
IXYhTFTMRt2NKhQ+2cOTr0U99JDuAqM0JjH4Y33qEJLN/nCwcDTG64X5CKHUptPTeLnKFDT6903J
4oC5+5wPI3WbfO53OUt9mxB5QTGDHvEbNEFyHMH5++sz7jPbb3JOtbojuvfzJlyOLVt5hnuBJrhY
+jBTNYkw+Egt32AiaZHyFhCH7PWK9IweQwC9DA/KdAhXMTSMlYkR5Wr0+Ozf5U27sOEsNKPTJYpH
zqsTYvL4tGIgH6wcR3Od1a736FQRwvkqvondoDA6oRnWEuNEc7XFgl7gN4d+OEF6gHDT123jdcwv
ruXsjKqAxGCXqMUXP1bX21+VTEqXCyPdatz2VEvV+SO+tvYtjUlykyQnuBxIa0+JY17iu8apzPRE
dIw/agTg/7GGuIpSzn15EwWHH042y+qYCAqvRVjl3f82g6bVTXv1CL2tymzREN50H6Sx+OhGsa0d
6KznPlbJrypXRTmP40vll0jm6RpuQIN9ZtA+Ht4oyyGl7UCtdNZg0SBoNskzhwaBkURGers8CDl2
Irx6IAiwK6+vJ5XYDdPlahiVg81BoTVXVlSFAmswtSP4vjILJE8cR5Bm2lFfcSnSgejBeOZ2xQcy
TSGyC/+FLop2mbPx5dKJYiPrgqEuX36epjF9gfXEEj6jjvvAf7PntnfBasBOlVqgUMZ3Vvz+RlwU
YPXRsgVDUHqMNEEiLkB2lVXINKkQoYe/IpFU5SrGgKmMoMIb/Xs8Pv2OhIKVsrxkv6WrNpt1K7Ya
F68WePzfNl6h3c31gsNTK17I2w9BJtD/7vuwXaOwkyDke8YfrBRXi4LtjfJpq0ROM+jkbPytQyv8
s1aldKEyGY6EpMT9YnJ6qzdFY5LR+UVeu81nAjWBFuw6snwqklG9zN+NUWTEtPIFj6jb8zG3BCex
GSLQFwx6ScUOlZaOUTwccNGs3hGytPAXICjyCsYjQ+qGpKexBQ4RUPUXvtH0iaR9if0n8lpqbfCr
K6YZeCexljU9ddpb2H1KKvNOjUJeNWsBh+ITpwPr6lM4LbB9IGTjDiL0dWpLh8OOpYprkjB3ZUMn
sA4x72bqpxB02vfFG53tY6Ur8x9O458RGtkiVdCJc9+WHzLibOaQsrgypOqk/BLtmU6kJ4Gc8N14
MWRIX38vJHmATvTDLNqDMXzuUuLvawhi6im055eoLwq/aQEHQarjVFYKs3cHNutj/cCTKFDqopGF
IWIX2SAgsy2ys+jZ0kafsP7IkWp8GKMy9tlY3SPohUlZ5pPbbH/o/yE1aVby5g7gPT2dsf2nmKre
zjri0EO4MAPWIKe2PTI1Mm0PmHyhlrx8oCjKSm06uEbEUcP/O4vv72SzgDlIYzhjz0YWeDjemegA
d/etXWpy7EeAvLNYgddCO33cMvMVUMTJPhw92S8bd+UtOW9voHt0/uxB6pet9pfQxciqR2JL+/P0
VTATJzdJLeX6tVO1IDOLZ+jyj2bXIftHofjZZoTjSImiFBcI051MdFDBTMlU9ez9tuyixbTBt7OF
F8wT6w348mCzpCOpVenV1H4W0dxPFn1EKnBGEX7KyzE0owYSkUHkepMxIrGALl3ttvdmjplAIPM4
i9eupinnCnIbbHzJtN/hS9RXK7f+EteVZA1ikJE9TAWHBCo8ehDJzkSZpf4Nf+5cwPilLCCSEodE
qPc0xbP+Y1wAGRf3XBlxwZhmrjyob94zibn9e30MCSfn2qoVhWNPKuoThcZhsGFJiKnAdNWSVjb7
xj4ry/a4BbEnl+McTZ8aj6E07LqealYrSTk1M/jvIVGRLIyGc1xNNKlF5AZwUD3VlPDJmL3qg7Tf
DOtqULlrVcPd0lKGP/GlWToS+ofFSxOrg/0LLT4gCl6IO1WTUh3Rw5wiveTzWyE1qra1q7oRZGVw
PQ6VIVERhUkD35wyLwnwNUKAuAEYIIvF/LdSbor18NcXOb1lPlS2qnRDqyjm9/MawSeFv2GJGuzf
GoxQbMFL8avlH0VC9KBT+Z13ZM8y6/dSH5Mfk8R1ku1Qpd7ZFlbIjifX0CAki3lHXbEM7iRJG0t2
pXKjMHLWzE+61g56oe/gn3i/UDnjDFVrr6wRuvZQwo4xVZ0D+qWsJqPEV8F5jDnJDgdgrh1zmChJ
Ufcs5KQ8jQNvjcOu2hF/RaUTXMM7gdzqWDED2TgVF6KPxTQyWUJ4SV+yq6WwSWnHibYEqVvyh4jK
+wIFn2TBZca41M/S4ztHf3Z1x5/m7DKy35xmz6+jI0JWZ8HEPzgNuPesgehZ6sOrRhcaqd4RirJg
ZsQVyjNXdBRlrFrCA20aFYfYkBAtPmiSCRYhc3wC5Hb+kZvNxA1yShxcFn3lVtNAqtswZo4PjHKG
l6GZ6kmFxC3bl0jFVxlyzWX1+E6uR11Xq36bMUHxxSw+V24TzJbu52pEEocahf6DoYr8BrqQVOMm
MTYPTcVoXApaYBZbEGJ46YcYTiUCuNeciS7G1oMSLbL2iu2MC6yOdAkc54w/OJDLTMBvBPdPxgoh
HXrNCQGuU8/shT8f+VPj9nZswIGdpxsoD6s8hikk/rlAtk/WoU+XnIu6yYJ5WxbRpKFf+uy55nxn
yYkqLRAPNt68HP5evpQosUrjDBdXM5OFAGF2ugXOrASL/FfkyPnmWcaEtqi1v6EVQgM01tY1E0/h
7F6b/91q+6JgDDgHvsBnt8YgJ6wxk3k/O/DoawINoteribEMPa+Nm+KmecWCPRp76Gaed2TI5ejC
4fbTm8u027wCEBPPoOuUetGDuQqqPCjOx1JHqgmMhldwRsTqhFafdGszLCG7ICDqlKjSsm0HzEnV
R9ueaYSwe7zx6sUXsKeBJ7Ougjvhv+91iEfCkFbZoTA24+NEWKEtEQ9v6+ZX8heXlr+fW0ZDB7xj
Iwr4b7Mp8Jl2W2vJPG5ai9kIuvrtA3SXq2E7FetOBA1n75Iv76yq56jfwX9HYBuiiydppnKiwQaX
bVHv1cJs9A9QRm8iEtFdvFlP9Cxd9w1hpcbE4CrXDdE+WBBw0KQnlWQQxxw5lwoxldsDrpvhdbmi
JZDwkVeotR+WMPZCLG25jLo5XoxQHiDbMsjYi9OiBfM0M+xp0FjRUG6CILMDO8OidqX986ttUevO
00/ydpSg91MXYEtHcM9QNDovxZH/tkaYWRMdtppGMNjCoOzuUMN9w4llX85+5ONRAZKQi36DxmhZ
Irrr+D7PywdrgyaAPycbch+jHe/+mGwtcd2odOd5ruW5jF7g6O8fb9ffnHmCgEkorNwdiv1nlzaG
QxIDPR6d5g76n6fJni0bSfqZG1jQ0rgEckO23KQHKjphoVX4y88EqJGc1XFJSM8+LsS17aJ8bMBI
yROx1hDdRRDA3x7k2KRTwfV58mkMLXTjUVTGT3yoWI6RVqBpKK539bqV+53EwU+F0INf/1IvNiLj
XbldINX0xHl8DbgLY4105yIOlMNP3h4I2UwhGwOAtZXA4QsAI/AHakgyOkPDnqRNjkWD/FN9Yf2j
2ZOyDbKUygrETweiOMMuxEJaplPOHbRVqLrbywFwLnCkqPSWP2Sx6jzX/dEOhgI8RJEfVQwprKrC
tRZ0zTS3iKDNMNnQt0K6o+fqKVrZuy7V3k8lTHpUPrRMU67+lesgMnXuTXzXRD4zPNaFcQzmoFx3
JTgefTV/q40RQ9a+zytEl8fXNNapo6XUzNh22MSRQcuwG3K7dLjCdvxh/GPATiu2jvg5rdUjU6EL
kR0eQrVStVkyNarj7Bd0kM/mPCgUJQNVpF6omjBrBGVLNptkck0zhfW6ITuxSU6z+jmvgqAH+M8x
gyxQIE+LRFlMdaQYEPmMmC1ND4FvvXp4CE6DUilhuHrgFumOppFwgnwID9vHsF5aTHCkaF4CwZcg
XAnCQVlivdJpu2aAHJKwaEVeilE4aoOgg7+zJyk1X8zLWVEBE3FaDepOBlNYPtzI9PsA7WfiovQu
G27a5jJ212WaT9IFNAeRL5x5Qo03CS50fG4tpW4EYv0RB51HUVlCtWr3LHcZXx4frfgyO/naZbUd
VU/rdbqQYD6DriXC2rAne76I/3ZEj8zegIljQGCyoYhkR7Wv1zSxx5XHyqqPfItJIkWdMQEFp131
hUrMCR0/75lv4sYkaotzGWT01jywzM7y66T9vSZK9vWBm+A5H284VBwklCjArNCaDXhUPno16Ahq
LpUx/Cqh+P+oHIU2tMUPJWUaDdOMHn+f9rBdhc6eSkFOrHSHozMbBY/jbpW7zh7EQ6FhUvcdq8Jy
OK1kXYhgZAeKOqXx0ObtG2VyTIRxv6ihbyKwhiLWh46R8pHnYcHVcOa5kLKPFUeU+joz0v4ol0eO
df5bmgyW3SD7cTHZ15BaY3CbNKAHTGtaLhblxJfIyasaNgpH+lvX09rNRdYo/t0X6QaxyhO0pYBd
Zxm03TkYhG2uzFoTuyMyHtUAr0CRw/X5+LKTyQKAKX/5t46oYJ8St+9q5X4zQ+/k6sK7qSGie1mJ
keiQWowwkhFadJE4Pv9t8NECHd2iPDgQPs8y3syQplXf+9x8BNJW2bbyNkkUKlmylkYBzItUPtzi
rZr6MwJ/xUTfOwwmIJv0hCFThbPBZnW+NobxZf2IRSsMBX2QGgxcraVCOsz3l31QVnEqdTm5b5CH
+mknGZV7bHXsFAqtukfODL+nYjhlRiQq88zVvBuRAnUdkaB759bPpM6UNR49EcLJa0dqHtNPMmxs
tnRWvahpTp9fDmLbVdCZXvp+gZuviJMM6RCMLXYKV8enUAsvCaswY+8O1LZEc8TSS7iLMiSl6ewJ
z8ziUBnIqvQaZvQriLEcPj7FlKGp418w7Gy1dpu/lLDuYkbvwJGOHp/Eu9yLmXNroQ9RafWDICjj
SJl70cTfkpXKkrSg5hCHBz8pD3YfY9oqykM+MVpYDgBT0QD8scclimEFRYyB0iJyjBlIOAsLoH2f
IL7ltONgCLJm/ON1c/LQMd5NAI3sNwCL769LbjOtchIOe6a31UD2PLyQbZ93AJo/XV1SVhqlIaa6
CzrImtExTVk9lWukxwxrM0q4MLamJzhYiZGo5qS5UDNthonjP9AftyxVllJkNiir+jXgchBzT7FB
SCHo3s/W0bvL0T1sCzcwtXNQPym2OtnxhRM1wpxsWprV+LpOJJX2n/WSfhTJd+Lt9Mg2xCiU0rwd
z4uZJlywVcHwNBLY3eb66gzP29vDGr1Egiw+4+1R9QVn6herhDyipUn6+Wi+Fff4KIL5fcBRQe7M
PEvmtQAC+HD+wRNc+KxWTrlwV1Hlw4Qik9SEw4AGp0L9rqhTxuuK/0i5WwqT6AKeRL5FfCoCI7lS
FjZLpzJziP38ONTbGtGc2e7vwMZfrpP0bwf7FUsqBNIaHGPXCOiqndqgiP0xKJD8bGUcm2N/P4Yx
e2SEg42G3it3VkawmJ4PzrFOnGDSmQOIe62hYoqSgmlh7FQb6PuNKwzsYO9q3BmQPF/x1gatFPb6
af1qtOf1mGXuHUvAa0W2lbOXGmvPnm3N/YsO+hbfj17EJo0FD+BsaHqXJhAgG+0CIQATzjRr4PCd
2oXTUXDQTO7P4C1O8kXLEAmB9Pb/E2iomRejL/hGk9N83A3KH4cA4D2XNCfZ5quKKo0wyOotkhH6
6AV55UEkdzQE8uy8+pqgwvdnp6oDXYPYU44dTeUq+PEVlV/xC8GqIUuj7Ae+2RpcwNFaQieZfZyl
M/xjKJcdoLnnQk5vRLCgC2KM6T7qAIwC7/bIm7dB4rlRdf/2YSu7Ldh8JH3mqegTid1KzhRcY9vF
A9Ln3AzPHld7TUkw+uL44MKWaUZXZM8W8p2jKxk3WWPSy17SfDFn9mTHmkAnYo2ZfcEnf58RarYz
j7kYu3jkmUq+1rRUYk6EFSV5DKhsLF0bbomWaL9IVdQ4WhQW4BbUACyZ0irncgnC/0uWtJsHWN4I
rS//ZWu+Ylvb4OI29Pr0m/peXD7sGrM1Swv5yBX+aSpYw39YkMIXg9hridMyaLKfKQG4wkxZeOhg
not2Bvxl0kBwPniz3Z5WByosLHMK8UYtwcbqRDfB6s6pAacO1uXhnp2r7xtKMaorKlen+2RGEjhh
yaHbESGeDIG4Wk17VjgtHbSQRQ7rXuayMg/xS3FBGHe5BT5cpslOyGN69eEqZcyc9vuZGQOfMK/L
6rHP6CXsK1rIXydLN2r40lIwhPU3DXoSOLQXzfE1XgqekiLDo9046JWc5jz3KmN8QKb0NDxDpxtL
nMKR0bjI4lPDjp0Ta3mSIv+E/jKzkeCB+BCOI/pMqqNFTReCIYSioQCB7Qy+Sg6bKJthUZBzHJ0C
8hQBnRlO4Ca6RjTORwyFuR4sDCg06As58V4UswXIO2q8MHMcQa7HTqcit0xZSkZE+liWXwWLSkTx
3d0vitoatt/KWKAynmj+JD7iV1uDyxUJUTWv+UXdpFGGHUWoNE0ids/CrGw+dSQU+TpRerg3gpPi
6LVIFJz73rr8jTZUoBfpN2Tzxghhh29YQo/lYkLRY0efdLnwjkZr5YvS2WKl0ddDPhClohtu3Ra5
ThGVj6Cejwq46tqE2jvrvZCDuCD2Q5wubzMM12X4ZwN/bpkBrsOCK4UQ4qY/KjArXEcPRXxPj4zZ
ydj3/GPBjsdxvGFZbE6h5FXu4pYNrXOSpg8yT1heIbEr+ih7NrTRfRC0K/ThJ9uYh3nATrpTAyAd
YGBLchy5eaBy1b6LXIDQz5rKjiBm/JdduqoLvSf0sLgXq+A/nHdAGPx8VSpTglzMocfi4JawTw1Y
5YQRA0hFjeg8MgdEAlbPaSATyqEHpbICPAlyOgueikOrioNaQAzpCIJNie0YbfiyurrLRRO4Oj5A
uh5Xptj3O9483sFVS8hAHmBL/MRXG0VvBXwuC4CfcYRcDEZGiJHrPWVYwPq9LP4i/uuJF7HRoZMQ
Jj+LE4RBYjT9BRsutlLgkaFM/ql8laS0+TSaTyLQnW4DsbfqO7qoE6h7YUKGxgLuYZCCFmjxfyVa
AkZO3wCisAebM86QHj67jbPma86lGh8PWqOxA+RtnAd3eXeyT2Q0ewSNXcXiMRpdB3Wiux5Cddes
wS5AyZoE65CchUQfJQUNdm3r7OdA7FnElLfPixfYeD7OPs7LnZf1J6yxwmW3uKwTPjfHqujt3e74
9r6IzrcCBTLBgLCEiar/JRh2VXll7HoRwDcOppF07kkYvWfDcJ84ghHLeK7epUyvk7LsaXfXOdi/
Qu4sNJiGuyiD1erCZ9pUr2BCAzsZAiA8f+PF1vH2Y698pgyn+NZwQd0rBor1Sa3T+GWzw46R8HTa
KXViRUDP3eiph03WNefjr8ZEKa8Z6kPrM5gv74gdJDaebWFlaVoqMprxz/MvDb/8uTz7jHOpb8mi
AAVnjpWuMJXsfs0O6wa7PoWXtIYXIZ/A5AkMA0kGXvNa752hT+mQfQvY270nkxzPNJDuKDUhG9pT
BBUYUF8L3XMF8HBfsuj522MxQbxfnW5cp/If751cDMxSfCnUO+nCJTE0uP8wT/g8T2yUrZ1YMYV8
Z4NZID04o4cmYvfJT3UBRB/SqMUubE1Ddg1VFtzHIoDpS36U6a6NdYgO9vuqRFkYR1oXH4VB8cPi
ZdwdsJ3Hx2EZhbJceVfg2c1mIxvF+OOqJ4rwb6r/3O0aJAwZwkEfa3iAsfWQ1LZd3LrNfjujdxjL
o2v2eSictZfIO8YTPzKzdv3+eOsyeIBv8NmtSjA1te8maC1Cf+Cab2SwDGqXMhGHS+eeg9vBAQ5w
HrJdCaDKa54C8IGWnhXfnUg1FK6Co/mgxF6pxdEUj3hEXvYusFpOCpg3/V5Nuav3yVhIM+cuOVdd
Lz05/5W59BH34Mb/4ZwR9UlhRcIvwGqDni2oI6ENxc7xWL+NmOQ8y1wrzGwvuQi7he/fulyCMZIL
0QVv1pgIw0KkSsDJ0Ho13HZAOC3w88mErbZMbApnZd4p13M9wyy8Zi4aTMDn20d+NopHWJHeezAo
SWHqh3CjQYg/CIAxMOQ0NRe1cMG7xGaKy2+ZU27UTPrXF5ZAKCxUdrxx1D/RjgB58fkhRdyBUGNa
h2+1vRgUFe1M44agAC+uiAk+h6lbIfQ3scYBXCc960/yTf0kSYz/uoQDY/nw4Y058+fejtGC0Gb8
dqLUz1wOM+ffYBde4jFpwebr3EaQRpKPpkJ8MULBJ9JU66/2st67qtJ/JcMlcMjakDUXdX0+E52a
yii2u/2esEnt02+8CALx0GWD4mdYTPxAPEENckUWaKvO5w7kRcOT30z1E+aXDVCgdKGEy2vglfNS
LoQb3swBm7lbBaHCMLHFsPY4md0XjJCVq/0+GU9l2kMMGge3QziR+Aukiv0sxtE2Hzo2AfXV1Lbx
OvT95N29L8z6UL7yWk+kkyNAwqpPmB8tBNA25PiRjB6RARq7wVOvY0kwsa7HktfSh6t3JfUStHHC
9pMDUEB6gF6TM+AdbWu8cdt8G+fiiUPF+4aV0U61wHfgLldGYpbeZ2BGGcQPsf5OpY34rifhlJeK
MseG6GRHXXzf8kHfLhnVZtyzg0opaUMB5ql7e/KD1NdvM+87JePOZuW6WyR6GdN3DnZeJ6eyE/ma
+MqJrn5Smw8nzb1m+5t5svhRie8wKrfB98sRExaKtUZ9AZ58lFA5mIi7Fge4JhZQ/H56S8AMXgr7
+KBoykud1bsfjG2KahsRZtep+3B3hfYnb/5ABdUxjL2l7mmNvOyJAE8+wSp2mCSHt+jQaUN2SMN2
ewSkTc+UBJ5EhcD+3ZwMjpFEZM3lDPavRO/3NtGmzlU65SAcSC0iMS3YKSEGth9PsoF1wAk2WToR
Dt2gN3K5IPfXc0Brr7N0ehIldW+aDBjOFOQ/1A3Gn8tmJLb9RJGfXCVV9yky4dpR/0B79PCiE4mk
BZDP5B5URQL8FZs5wNo6t8eRcBIEgN0W6sFCvHpIn7y4Z5Rz3rbl7Fz4Y3CUWtYlBcclZ3UiggDN
l66WgVJJ4sakKjfKCC5/nA19g2+g7eF6Ux77nUbUxeU+P6OnpCSCXDqlFfJsaGBM3dUINYzyeGup
UntSWcYbegVujUcgp+wut+3s2jGotVCtnvrX7l5on7T2cWJbTTyhEocZTusNccot7qpm0clPMaQR
pNPI2D+QRbRJYV4ryDC271OFzQR64LxVGRqFj1TJPnDguHaT0ThXTchbDbTbRhamPF4X1qtdfpAm
D+WikSeVMGN8ttFfXbYHn8Ag7WNA7tzZSsdkYZUxtYjAX5sG3Zm1Jl2KX+IxQr98sgwhuGgsZkEF
EnpAo2+7C2zu1DOMihtJf7I61Psxc4gf7Db0HcwpaIXAxbLt1FN1GV4SA4ZC8n+bEsm/cYAN11qC
omXW1C/f9djqh866HkIdS6hNdkSFZQbHtx65gue27uaXtw8FEdGiiERrt5X4vpOBxEUneAUwNQ9e
fx1RFpOG1UyHc7gdUMi9q7mT8ClImNdvHOfOMiytdkaNC0pPelkwRHthK2ilGqz/St3M9EB6X8bc
4spZXu4Ag7SMATeyvPneEXN/qDbMtGi/9WWrwv+SSjyhm1DIiXzaPOEdz/efs7Ziw2TYmKGQDdz4
7uME4Yq3k4Ohv/psB7ItLMteO+AKCdQ+uWyTsFJhLoJCViEC1rlTDaceUbYLSoAKa4a8LBy3Cblq
6hGGuGV6DiBfjVcEN3rL/ItkuHOhUsEbKNh5Udw78WzIABCQPEM1ka9vyCzs4C+56FyHB2mTwMb+
Z/bBo2ho+XF5jwVUCoFJRo0u1/4cwNm9xj1wPvMgZoRpnTcNB8hP3Hw/KKp/jN135qnchhYtNgru
TqX70dYH9uS0utXikPBDdxmEYvcIFsE8NcqqJx9eIk/UacZcleRfkHBIDtWqcodtzw7eQ9lMb6a5
hZJiyRpDhCU1NQFzwzUpabhjk3NxnczNNjqMP7LoLbLHzgfc5nEkH7oeiBo57YBiR5r32/SKpdjv
Ior5nIxWUmGsNC1tp7ByFpDLm35YhB5x/MttStg93EP395IediHQSDnoO64mUpATyId+v7g/SJZ/
pFxlYeBhak1g3oopVTu65G/X076HQGNT86d8VihaDmuLtX5Ti9QU8HTT0+pVeadhLFeev+/f+xsI
I5DV3YvuMzLp1Sqgr/6Sx/2Pp6jM2gwg+RQz9DUeNTdP9UV7hY1we3n0Rljk+rxIDV6XiHFYKS5a
t+nvBBjaAhgBPkTjTFh5WBDzNmTH2ksIphFO9ymM2FrUbIF2N/wCMmcUelWm5EySoDETs7v2ek7j
r0WC94gnxVFuMJUcnxxl/nQy2s+jVWU4iR2LYrUBECMg8MqrxL/lUvQLX/fExX7UcZQ8EVCY0ZTh
vE/knkqy7qMx+Pz/kMSn8qcZU9wOL4fmHjt0KXL1kQ9jNWrzzsGxlUzOAS/NyJ1o5umZz2JqU0Jc
n6D9mAg5BfLeUDA2A6DYhIUl49H3l8+1ZHJtuq3XoffRdraCwP6rkxXTilWqENKzFHo5dVlqbEy7
io6bqyXhjYOTTHy7vUfiZSk8vVlUspSrfDkN9vx6MeXhRqf7SN0NBShDz2FNdJ5Sc2zQ/nsVyLDF
/nbmxmG4pNtwuDKXLs3qL0nXkhXjT9KlCe13avrUMuQp8BQY+PHI4IWmxd5I5JxXdMhzCoNpr/Tt
n213KL+N5RjZhiaoJI1xObF7w2jqBZ6y3dUV5HfswVK/5kp3LatMrrm2OHHthGETzlVmVUa2ebFa
4Q7M0Nvthk0fIpJSbmAUuyiJLD/a2ggx4G/d1b1rm0nAonEgmpQliBMnjcAkXBZhbx5uxQz3BOtp
Dvq9M4mBMkpDZ0hgf8NWP/Wk7S80ZtqnE4Q7n0Xj9Np9hXq0CjUCy2h/AhlskrkGk+GqRryi7uWy
XCSwUJNJHhROMIjlIFOVhZu64hYDA6uCwcp3eXYG544nCHunsWGV7vGEFAp2SOgbc4N7R/fev99j
VkRbxK+6x29lvnDl4tu0RhDkX4TkpHJDdlsCDcXjUm+ubr9gFGgbul8vKGatIzvw+mt8cIWdGEBa
uihGYoXIDGun1FWYHwj5XJLibENxKg2cd+KMSLGpvhUhGCToF2QlPhT2sXrIMh//uNlT0dc/r/aq
Z3F4yTWaFrg2Bujsim/0rn4MnAoSAjitJ5APMdshYt0VkLcqcIstAif/Xcoq+VSonq5kAwojzkAS
Oafj2a0gQFlvHFxi1FgtHhMwVxFEhjL1V7aUdqcI2RUTa1gsun8EL5u1s+PpEOR2FrKqzaswWDM1
7v5gn8SF5wSe+/R8cUfPSjL15O98SfrWYRIHbs53rP9PuMgeq9+QhL3HHNfK6HUA1FtLryGQxDJp
QPqxZ7qy/h/zWp1ocS9M0gWMa4yViuE0m1VcxZp0VzKSjw4+ejODI1LlLDXHzp1STvuL+hYVCQmO
l1bdGkzq1fgcmHeMZcxLtSJ8+b4Pkix8pFzX7jFGald272LT5CkQmBQWhE17z+NF0sEXGcMj1MzO
LaXIq3DbPUmbE0A1beqwO4+HVou74WmQwOK5LE1ibDgaesaGe+qP1uuqdrwneSd9IEwnknbg3J+v
iYG+ICFsLmgZZrw0CF5kcNVU57RUqwPd7KZGE6o8daBRrlmP7ExxavPUI52UCGWxyegtU2EkZT5k
M8tGUEUjH6euaxrMD9XhrQlKn+pV+RTxKMD7MBZjnsuFTGdcR/eEpU9HphHOsVTwhghgQO8j+BE7
bB1CyPHoHbezFhRUZf22OZqNMTS718corxC5F1XQWEuHDz6n6HMd86/0cSrSeXf102BnDeaa8W9R
6/AvyqQ+bP6YhkUxLWiqc0wg8egrp37/3VPI0/bBFvDM9LzEV2ntxCX9N0PpNH9sOqacufXH1tYr
pyj5mqLU2zhZWzM2w0PfoZjUJkhfZxWRxiVjuN+yHkiDk5lShHhOj7LYgsRkRISqTRAVq/xt1Hdg
IPwJSkeGtxUdMbd0Gdg3TJLj7Uye31OJ0oJ6fZKvXV60DGdIIoYiAsTI3totLFHNU+n0HVLYqtvB
Hv2RM81VrI9oxjVQtCVd1QFEySAR0gOlom/V6b5H1QGpwmFPTVGHH21ES6LPSoR3LSIj1GaOH/KS
9k+Mz5VvywaOCrc2oc4LwyYBRN6pUMsIlV05K80bo0jyMnssIPSqQQ1KniuKVE8Fc4pMaE7euDeY
FITVDyIasKUgh4mcr1S2R6PTB6Sy+OVVPS2qfURhGbKhlxmRFYcCoIaz2hdXeqvtbCXbOTLCNLuX
WEh//4/wqomJj3nACjwe1UXEBZKEDQ8CKsk/7DvEg72lGrc69l+xOVxOtj73JOXxPShrOLZ5RUrN
MIi5ak3ciZYLki0Um6E0zShcMHben7l0qdHDrzIA1klwkExS29V/9CnEzqtKiOhOXs0DpI9KqBLz
EuOpR9ydDzcOBExy1id0lTBbBzIXX7zB791F776fUjYm5DEuHmhzt6f5M/VzZntVfIynpTqBljIA
eMxtmbNj+O7IEPQM7n9hc18qrLgnoCENMMSE0+dlYqxrOA7VZxkNLTxl1EFu3Poqxouz51sI4HUf
vF8GtnckDvu7VnraPifWVrBoiNo6TrJXEVb4xgpcuO65Gy5qdpNtMOWXf8ouhkL+VN1cTAeLr7i5
CaD77JXSqQIVs8aHblDBORwxp4Ctgfj2EwN+IhhofRhVqoDgMFZ3yA7LvOfERMGhs7nJrzLGyGGu
+y7UtpwJ60KwHIRDCj4mf5xBpvaDGzv6z/jTG8FrV0+/rvNqwRWv3XEtxgwT8NQpkk60ViMfD3xl
eSVJbrlFDWsJD87dLOHVIwq+eBu2LkXAm9/0aRXWJsRqAE2HxHg/tlgUad3I6GLK4/p0jjjxlEnH
KZZRl3V03YNS977QEtMJ+C34FcKRci6MkllS5YRe1F2ABNdRdm1j29qz6vcb2xG+w4OamCZL/iiN
VsM6q4KGzeQoRELnLjbovF8mylCLgsth/sS6tP+8HCbqm05PvUABv6OgLMR+AoSmUrfUo74G5t0F
vhkLAI6lQal37x2veNxPmjTYeObjpnIQ5l/EdE/tBd50sP3DqKEJtcXZukw/il87Zd84BMo6412E
owzSW6tpkqIXnT7A1c8Z08rdawWaH4+z9j9+Twv6JYA1rb6lvb8HBAByIygMo72GzNo0Xx5enXjM
TVVWDvnD2X79kFTSxp6vi7duNSu555v1AooD3KQsV9lHC7tTBS1DIBeGZiAdGRI34eqBW3665TUJ
9S1anwr6lpcIgjspKBi8HElHp9Kbsz1y4pVEPGigvFsbO/ePLlktPO2AgLKvc1HoRmGQ3uMP9lP9
vHnVfiiSjeTmNtC7dEEwLrMOB40ZblkqP2v8Q/zvO0hAh933BKwO93pswGMK6QbL/HyXHN0wJ90g
Gb3N9+dEDXgEaW2QyPE/Yzo9druXRbw3mRqlJgL8xm4zWs4lY7CVKPb+hAerb3g0o7Fl2LPjk4iz
/Vl+8iMUwEGdWOysVE6oWGhynkK0nX2jE+WI13C9H8SRJKvho0K39XTdKElf2MsIcg2QpTiUpnMM
XV7+iinW8JFdPmnUlHNyQUKYc45yxp9UuqNGRr3BaU38dnWfK9hq7EFYID4vListY+Q+7KBU7V0H
6D68Q02taDF+0h6FNPxgUa6hhcGzfvQSrfS6vNZL/eAKd3rG2DUhFWDgElqtx0LA4t/0pYej6khz
ihYur99wQ2ZauImXagtks9E8Oap8Dk3KxC0yx8lTqhyR5DTBmg3zNZWbfYoqc7Nt80keZ7f/dyOr
JZCRZJLAF+OFAdr59HcxJv/gackC7F+5kY8HDEaza8COn9Z6i8JMvM/LViY9v1CquVNziyww3wNq
m6+YrK9szZB+eGreR9qwE30qw8TOBITnOHLZJHW3jxJL+nXXQPEClUow4Z0yJmMxFeLHZUf2QFiE
gAmCRrb33UlhQv+o5U/xiL2cOAvuYDoS5F8a3nL07v4VYb7AHqFqD8Uez/93E3I8jkVz9FlJIrFP
rUxeagVBuX1xYBFo3YzOaP1K+gqfkDwIXFR1F2wz1u678psNS5iH7kgAbqDShE7kK0mbhucypz7O
Z6cefK9RxXHUpTcOBYChsojZ+HaEd2/2Uuub0fDkBJv7vPYzjx7NHl+Iv1des9fH749xbQBy1rll
CHIZG1lcmLkib1DgMxFmUNIqZmpzoC4dODr77yH6BKSlyH7gyOr8LkITHipps2cuA5w4tJrwhB4q
nHQC0yX3Xnrnmw0d/ZSXO0ljKQ+KsiVWXqiBGRJ1tLDaHL4g8+FKVb3yk0F5yZI1zQbgXOS6ZJcM
CtyVjUlILbEVRant952cUKG8CHiflWwq8L3+mOAV/1V8UlUvlwA539dLNtcgf8TIBYaHCEc1H8oC
4swASinQCw4RFvmfE9ciI92G+KiVTqbTLmXFl7e/q3ERY03aM0tWTWlHZcXK0jPf00V7kUMPMxsJ
CF4e+M+zsxs0m1qJzazsq2TaGr3+RYi4CwUqnlXoBK8OP3o4BU+1lN344Gr0XHnelvU8Nq0pYA1Q
YiScxwL9UHiiQOaJrmUmjEg80l0TJA6zsHIu4wzopIpbOoksWsF6+XFodEiLVbJBd6sjUwUZB5/D
BxMZ+9NnKhlUMCqSm2+HvhJeNUUojyav0SIH9M4UnbMJCwF5j9AB9zhqSBRJjP57RW3um2xpw7zq
rfoR41mWDFy+3N9G9uHIdZdRIdK9QEJwNBXb1qH9sOS8lJMdNym5iVphhI28DCnIjylTN6gDOEzn
hRAK4SFXKuZa8JwXssyWOZwK/dzLAqv4mztwGLaJMshyB2CG+OcuhEqr8380vXYyp5H6s6FUqv/f
b/HprZntm0+Jub8LWcJ3ONcrCZ8fRHTv6A4C39tmh4dqf211FmGN2qK/8/4XkYXlmgk39slbk70i
pQSLJV5MA0ho9o+drUKFNDgz8YFg94SLAYGnrcauCgfATAtAFuUUp3s1CpeJnOhRRKx6LW9lDU/m
UInTFAyAs17D3830aCUgprjqiU2i3B2MIG8w/j97f77KwjXlNGRP9uMPFW5GLwqMBnoPhwbufKKJ
ba4J8CcU4uCLqAje/0aj4U+vurweWPvS7fnL56pvR48hnc/nTGzbgE+KZSveFirwote8MKOeXp64
WLKZRejZWZX1xb0AmvJZqvAfeTfn+sIKbZkTJiV1z39YyOpF66PPH/4aXctUxwuoLJTxDiIOmlwR
rqezkOH8HFmMqISnfuxRYXVnniRmgu1Dtk7mA990obtwrkKyGo/RHQDtmUg905NOC3asde8RqDkt
D/UowD1OG/F0rZ4gBw9LFFU27LX9MlMyI71PowQLDGTW1RQMFBaTozuM/irbv8FSVh3m81hTMqHJ
DcsyY0qSyqkzt+EquS7QktBOxMkR9NBEGNVS2OBRD3PuoszFYGMnP0q761W+ImYbCmrLGqZT4FM5
VCvn9InWLzfXFOYBpvxOKqSIU6GMenlMS2sZA9VsmAm1UIGot7RZV9uCizwUaW9VMkNmc79QBdtB
RZli6Vz8qWp4rvN/hJt1dd39YObff7LRqVjaYJVlSVRvlkDqr8yXD9/9I1cjFVDGiV5IdLcDhw1V
Cd+anW8HDjxcY5+BInYtMfwSB32HBs72Z6/ioqHZWjkGbi/ouEjOq/Y8a7/NMIjdQ5myBin2gxA7
n7wEeM8KeUoBgEgrgNBwIs6mG8XeukO1NQ4gqkBsTgYgdCDzNv3ZDjFkDyeJtl8ajpATtxXvIwMb
6IRGdfkh7lsigZnkxrAk5Ktbg1OatScoh2Yz2RvYlSOR4krJza914Up8b5v2Vr/VUkkQclzhuR8i
W5y5LGVP1sVUZEYinw3YifIPQ53OWTZZSEppAARpPtLStAvLNt6gCA5WtS+0zhwYkbu821kiYRX1
pylZsrEKilawvMXpLUzAHPVrm3a0tylcagDBKg8xFoj0ktptCIGYIuZ+nY7Fxyzl/2KBFI9vhSYc
5kdZho4o6de58O+hCki0loMonfzDzhtDFCUviTb4AkUJqHfnRFqxDkV1x/sdPR/GYrvYe9PgrWRP
g2pFQFE3HzP9q0FPhSclrqbNfoQYF1TjCQDCUmzVl1wIw1FpFYobyR5zu8Q2XnLyqGwnFYtYJKDf
momL//4paSNtHQi/X7tzZ7UY3kgIj9v65xMEZXd+CweGwtbSrMJ3KoDWDqEb9hcwZlipDHFJ78P3
qQNyDgYp85dO0QmbtkjO+W66+TmyPszh7Ohv/QxIX3o1UQXH1Vc1vig35vX8+8nGutYyejErsjEs
EP/MUOFXbs7p+n7EKPAqTqlx4Bye+XGeEuA33KiA8vjrWsJ9bRt+XGBglpON1yO7KjI6lfVea6cY
QPsIavY0F+5i0YQgjMfT0IPDPWMUsMGaj1tAIjX/xptZjZ2Kl/UurUUQC/lyk5eW3cLQlISJv4bj
kc4gDkt1UCPUeG9vHhK8TvOjfqwFjCasq9PILH3H6QmNE/rVZVABlV7IjuIC/dZtxqaDP0kBv+5T
OuaOxP1MpKN/ZpaaIk4/xHo3F60cU3l+p/Hh+im7lwt+6lXY+BYvaXxUH5w1hqQenLWMBjvaHuiQ
1CZy478riIhl3mbGGmT6x6zD0EhxJTn2VyvB5loKHRuIDBVQd0XOoVTntMDeig9WbrUbZk61aEzM
YJXcXXP/Z+SQ203ni95C5ckC38C1lASNMCnFqVQMQSPFMLW+/JZXc1P/CwRVgpl1tv6pkzvHUkRc
Qb3g7dwjz6mfkcWLogY0cT6jhvsv7WNi/Ih6s9X7Ti0jzMYwkh9t45ibi9k7JetAVvpK/Zbb6O6M
uN06IXD3U4hfXXas0u9ikC34dBJK5Pvbf05xvbFVBRsJVlMvPgFZzfcC+CbSY5OE0aCM2Xm2ACnj
NPZyaKxTCT4iQFjDsc4abS/a5AGKwngVvqMOjtgmaYJdWrebSWaaXb2yE4XxP8ZZ9k55dwwjYaSq
+2vSLV8Hqbsj1fEj51e3Gj4CjQilq4OX+L8Y5OGxma7y1Fcvxq1ipJwHQzI1iusyQ7hjL4MMQQBS
MC447nZRgcsHzlwkMq2Fvxjxlpuu9LCVfHl91vUKX3WQmJIvcMa5oEW8KTBhjZXD3ageUYgbgKxG
6m4TjeXD+aY5QTGGi8sNluStT+AEZwFp3yC2wDU3ZVrVqMySn9aAOQnacroUQarXyNcsaLkBnnxX
ta811GQXUFUBdyT+G9/YS9DhVShzAjrBNyCPWB+96r6ydYHUTarLau5U165yr1O2PTgYzx7UDoIc
OgM+iKwe946DmpF/ATI4y5/iMjlaqKOVyI5wBe2/y88CbBh37i3HS2ttPlV3lo0/SYH4YfFrwHjE
Xz7Kp7Fk3kNqoB9im0lhpguaN4RMT5FwxaKa3QRhaWLCGQie5cQP3yx48EAjBeqFJf3i9G1bPHHe
scGzSJuQ0MPMqVCmcxudncRQBB4Bn6HDd85AgmtZIYHVc0sUYzy84W+u4Td0VxckRx28d92Z4Npr
k4WgN3LJIiueGfowUQqrrDNFEk01i1ie54mnvPFVMLntnno6FH/JLkRQFHIJBfmA6t37dvUPS6Yq
ncXtcL8jJ8yGa+RztrBnODOuBbj005Vl1DpU+J26Vybb5DHcXi59VEcltvZ9EcIMJltG72SEeeXb
URwR2GfvtBCeZq+16/TdaX0b8+1IeCz8mJoNQFbKl9O1gCq5r6Xrp6yxzxn102ndNUR/NdVLWCh0
EUHHZQJ9rLw7RroZi1EWY/0irSXpV45XPnf5tTZ859V14rvMGGhnVqcKynlMQtPlTNX0AxGmT2Ru
3EndpHolSwj4OUtZ6NJRaz3lUpTkPiPEcnb6uwwFCidap6UtkVvtZWQLVhU92873zzRSSsFHX5Z3
0glxunFbwdbNBvA6coJL1zyXPhU2cH0i54M8hIW9ItcxM+yGHf0w0fgmf5USGiV//C7ztthvt+hq
qWeUPCGnRWh3crAYzVunt9xEoHRTkeK0IyqYhVbTNN2ZIDGa3NtrJjKL0nQrGIYYZHGyob7Txw9n
zqhKmfFIm3wUFIFAGSDYG3Ig6GhSlHZeBI5EFRhtFgbGpghJnWxo76AzxagYPK5rzMtBpYitlEd0
AucaL66L7iQtDg9svDc0OwZA2mQ6oJ9yXd3rwbK1lhOlqP7VqVWKLVmwr9OjREpvcklnmXON62bw
aVo6tkU12Q1s0B0beOTIkStImhNhzHJMN9cVkNQo2AZF0bj86ZcKwtfXYWelfCrheUFg/eBFZ37C
+tEKfnSKAXy7pKBobGy7lg9yJWr/lfYe3eCXisfUrm4OwZ46XWnStqf/2wU/DRNSb4kg4sEP8mYM
wCFYwrzE8R8P4KEDZARYXVFQbgufHF5ubym66Iiu+4R1UuJTS46hcWrEPkcIafmQZI7NTEWO18RH
/uUcdHnXN4lHHnK2WtNDjfkcW7X7BTDtwcK/vSuwqlDtWl9Vs0OUfbirI/Kn0qq8Ly3I4D8IWwwR
qMdvh5rN6xDTKaQQXqBfsuuo/Fiv5GmFhGS0zV3KsWbDRAXXBPChBJizB7MZZPGkrHg6WA+ag5wL
xLIaoWg9SBOe9j98aplVBA1eblE37xoRsEf68XEs/mbIRtXooRFtRAEYYHXgPwwvh7Mc2uVkHRPE
3P/UtKNC7vhw9YPCUNXyuRNNvCwul9+cQdIzKYx42jJHQ0rnkmvQSNIRUG/RjcAXnkxVu3e+kjKC
3ghrqhNMyXTlkm9hIHDSgmZPZdNCEJOjY1hmAq41ZBCxmPhQ19g8aXHgNjRljMRzRkDh8OBJ0D3i
zoo40UNnRaQhz3jJ4O7RrynBrCLNf3Ur3SMx5kw7vySnIXwxX4aJSQXkyzDlayPuV0YNd+6Gqsn9
+hRdJsB88iMR0uov1qs7dNOdqKLjSdkeQMfO1YEW+79SqoQK/KKkx+u2jJQw/350QPQDx3fGNJMj
feqS80mB0KkQRnxcSjPdAWN1VjoqcOdTSYzzuYxNXrli36lITx+PFnfQX+Ei3FCEGzBxeINPQGGf
CTGDY9WITWZfTo7KX7uykvzcvuavi2rXm8bo9wWmOHoyJDq9FWfw/twiXx+Fs+HtpDHmB6ZZau0Z
6tO6P/rhe7FNyq6JxZ68xOIK+6IOBAboToQK4Z9RelZNpCaJpf4tvLiS3RoZAlpfrFdbyKvFJ9DM
M63mnwgOe49NNYF9+sm6jp/gYvkDIcfj5+lA5/WP2A8qO8xhJAV2rEzDtda9s/7qbe4wMYUtbHb3
TbwYP/6j8n0PaZ2Dpe0G3kxC1xntRxK0QNL8akMFiQ0pKwpASzYAjT5V0tFlxcVkAWRTQKZHKAwg
C7XdSmut8iyuwCoW7Z9nYYNQri6y4k3tDZsJX288/X3xJKXZVQ8VWVrgonkEcYEDIM4wmj2Ex6Xr
n0MnK1R+gswIqOHi4kSMZSzpqQhmv4flhTXwZM2lmrmZqnwrdMwY/sflTWn7xCeNKiHaqcZYL4dH
hyoxFWLvEO2woxsWN3x8Pl+DoGJ3tH8M4R9wVv26jl8kk2DJbrVZNzt6ua2+3K71p8k0Hjv5ztKE
Kixy13DVbVopTvgq8q5HV+0Alk+lzQZf550VjFQic5JpAnw+5c6lBBJR/jZDwkR8S5IWeZBQpO/E
BPgV+fC9hP4P5LDciAGsnYVreVV38vAGKgb8nHLUx5GZTC5zF7FH1af5cMMKpwAXbr4fJ7uL+QOm
itxmacmKhiS2EfZoikFS/aUycUZW6U7XkzpMiNMZ/vMl/BrQqRX8Y2RUyoZFYzwV/f4mETt77wgO
7VFOM6+rXL+071DCgFDlt9nnj9uEU3dFbS3yIeCTdBolpZBLAb+QeSy+31gDzC09LjNa5vqvJeM3
R6XfN/ENJVUKTZoCxcVldT65X1BxD+hCUVOj6/SXYcZm8wmfbhEe3uDgaRs65Z0n3EHEdKNFT+gP
o4wVzVbMkjt4kU2RZ6Re7UOhaKg1CKgPn1VH31eh0g4peZKIBU36Bd1fd2oaFdEaaJGN4eZaOU9u
lfUSUKd48toXlunDYvJvCjVAFns1VsdARn63xcXK5lUTTzJuJZ9mM3MpZcevFIAeF9XwGx2+M1IP
q5ZoG/2wLGtW58RoH7mToaD31P6HPZD4Tc+uwZWXQZc6lFWhn/qKuGIk4S/j0+Nv10I8+ECaUd86
DMedzM2qKIdXXCYTOZJtkgi8pqGiip2156hdldD1X+iJ8PKuIRxVOwPGQDhK2yFDllCv+swMuJLK
+prYatuA59NgEacPs0cAJgld4ruigivLo3HiZZ6sIWspg9F6XRPGHz+ThOx1MPajZCadBj4vaaK+
BIRHT89aLOrwnrXRjy9W6euM5cK80ateRpXAT6/TV9vHqoawp5o0g40UjIfpQ0nYLYLP6ktr7q13
Pj4qV7aiR66jKsm9vZajqwj/4EJoYNJxc3tYH5BbgQ7BDfx3zmV6LuFveO670fvQ+yCni+6cRP7g
1xhoMblvy6xMMd4eZIe0TjdG95BgdslEjHnCyspPrLOHEvFlRr7TnBshueXYhqq+2i4Tvd0C5m7s
VDPZKdAev6T8KFRmo1Ibcw5KfGooD2SMShnDIgdaZPLO93+9gQy8c2D3Dkq/aokhf6rOBgYoihHv
xBzPxXMsHNMJS3b7RuCIVdhOsipT3NLIM4LWFkBZ64eOhSU2/NHjtewB/RrkDyVC5sewOeSSTaWp
REquKtuUUm9nZTSU07NEPI6imJ765NqbztBgrl03pqDaaEA8FRXvac4V3XR5rNKgNpLLB/IfAIGW
oW2njj5yaasJhwDriX5w9liIcHntbtqEmZTXyLpEXgONX2T1T73n6pTWrCAdiWviGdrkPUZK3O2t
/Olri616Q+y0pK0+EMNegQeuZuoUPgqm0XiLIEC7SL1YR9sBYtjoOMkAD6NYrUqIC4ucfa0hOtYf
EIDb0+qBiLoRCdek8PEX83sYAzS0eR1hk+8e3kVNAZc3rfVIS1HmJqzpXvpp7yxpFwZA9K7Fojrs
09YvnN7tXuPBl6IZGiQVwbSzBo0ZVJS6Hy3krrmwLDORJb+wcE7yHUxQnNKZixolnH+lmp/oedMM
aVi2NiadYAdwQhpp/6fa2/3sp1lP2R+9kWUjwn1RdLpfZJgwFchaSF/oO+zWgqyMF4d4yzOHnZkN
46Z7Pr4r7wwdVH0JBS1sY4us1qkeJkq7PzgW/ASeXFPZeUbX9xZdp319SWmRDoaTX4yMr4iMp/2Y
8/gw0eillzDSqaeYC9Z187q1ZdN5vbuNlkfi+wmqgQ2UnfLUVjuMFPBSwbUAdMUwH3hscZSELW3j
GOQg5WGEjQQJNTM1Ij8inDC/jGg/AOtAvBVpgGdd4F5zrOWpdviIlMbUAf7tUK1iqHX+k68Czv+6
gtjPDBNyX13cwj1dLOXBw/DKL9fmfJK9sdKBSBpizFInQExFR4eNz04KzO0Dsyf+/u1CdVKYP0H2
saK5CQDHeL+a+HEQ0wDZICzqUkY1s246dbA0F/ujMI8xHhL+KIo/RguDuCWt1zuvxlj4TdfBdgQJ
LVzruD120E3ke/9KGMwZAc9tiuGnbU/lC+KykdW76/Ujuk/f1AzkruknQZJwrFTjKdwftqh6REop
g7z1fSQ7vllFGe+rZDJuAE4S2n4JmmV3TMcqDK/Z9Cyi0qm3Jl4QluJNaggeiCSkypwDSNC/4WU/
k6Dy9zIpEGQzHp/cDRpToO77tlolBLcQp6/ORgEhnTLCvsZXK3sy1PyFkHFC+aDX3+ONe7IDXQCF
3d3E5Di2oFc2hLLP1bQ7tHUOirES/Lj50TU1iXYRiKryhlLD+U/ssj73Fi0X9bPiasVYFhaj2fAX
P/+lR2UeBYxMLF1IwthHqjrb7ZobIowz1E9fdjPPBQHqkkYNp7BfPbUbwmpCjfNCdImgE0Ru6iDX
8DSLaRpTSDsB9LHgBtA8/tUqtC9fMYAbXwbxzUbU7gn8GjFdI7nY34GNj+w8D9WWl9xk1ZOgmUEq
qMfZZE/OxgRK4IGlT/OuAGz4HDg+o+CrK8uIDJ0UZTEtACKAMF59Z6HlMODkmM/JbsOlOK9VCm35
K9dbp7YGs6maVDIeIri8PDNgef0u/mjK22HP+xzwPMh07C34fnRJMVyRQdCZc6b2IUi/Pw+UVGf2
Qs0uoLzUk137qIWLS9S0F5e1oUe2QW8psU+KQZxUvh/LBsYv3nEKCPyFENdw7j1N5Jzq5ZdWihcY
27Ez939xSxcw7p15RBZECmrQ5qZFehDQqL/jwCcxNR5tAheMfSpJpcL4loPOsmkikgRyix4mMVDf
v/+VUm1wRLN39gJBZKTKRAnZU7my6DjYpmAx7U/3DXQuG3qH9i6sJvFnTvy70a+XUcqO0RL5Fhrj
aJ6/AEfTPqn98uzQ30HWpIvjGtHN7wDplqAPStOu+ZdzgZ9KP571M4GKWntJN9bwGb1QNT7GRHLr
37Xb4aUtgLEMOxpEPsExDNQojVBI1JkGlaV0/pILLWR0vRFRVSijrKvHlADelyU7yLxFibpGi75G
77QVdb0fFNJ/hJlAQCfNzE9pUWPvzJMM5w1Np5C7shU9CPrX0Kgjpwlpko6S0zHaK3+qZIyAFz+f
HLNa3qsfdiFZO0hDDyqUHSRxoI+oTHYa+JsvAkgOtg5xhVTf5P0tg2QKAGhx6c8O4+T7fBzjRWgx
maIeYlqKxdnMwRSctfmd6N1cK7EcmW+AnrW26s702mXCKVl5RZ1Mxx6MeyQuZGIjSWWZkTNdQS6u
bXj3YX6bsmr9LEtW7EtzCbibq81SzwgaHXhwYAg8grp16DJyXVtvscpLCQfu2jQlyEmOU4hF2oDd
y8+D5XkkOO+wXnpnftcokDqcPHte9SpAH6UK8uk/OplQEJNJ3iEKbJCfezma4GrqmDNeL/WL5rAV
NH52PICF6uLRC8s1tNNAGSOYjD/8/DDTLpK4+yuL+typqu8bxVVY2gUj7jedemkekpU94KN6WKEm
riRw4inOPv7g9THo6MjLS4E1EMsKoh7TUSVywv+rPtQvP4eks61PiQS2vElIvb4Wlm6aKeEVOGOL
HFDN65WdjiMU4zdHyqhdVFKeTQ3tCXKyLc1d+8B5NE/4IJW1RK3ByzZalfI7mOxomPfdm7UDq83r
nvr7adadwWVDfqnilXgTKyLcH6T3a9cohjCJf7DRIuS3t+4F2EM0/bj4Yj17ojCMqCH58yB9kPg1
VIX66iKfkvOmdb82xyCTqvodsQMjwsHGOwTNiOuY6eXS7Be31BVpqtkKOVQrBRPRiPTnMVxaFsoq
a2rrc4P7K0vbT72Ja88RfGPNDxepYUsqJoS/I5voKoZ6oz9cMrunqqt9UrzzrWreHH2tA3KHnG8b
zUrBWSmA9WRtzxnlmx9LTtSk7OiHN1Vm8OSe0minfTOdW+fE4SIwyhv91epn/LgN7FAvkj209BDE
NcjOt1LjVuaZITT4ZWQxbc9bwtRIXCWUkvZpOSVuWL8OA7Y3dqpUxU+bEdXj6RDa67xpK7+l8nLS
s99aSXgah25gMIu2F5ZPu2AJqD8v4QCzlnzWA0dOM/ZV9L292WoTh1w/H4PeoRhWXV2UgrgdyIvo
aC9T7eMbGry7RkNDBdNhcwEf99K0DX29iCft0ok/W513VGPho2o2q00yToa7dTWczO/05Li2zlI7
i2yvy+1AhPROGxz51JyBz5rNf28tzZLZNwKn94K5GwgvEwncjoGmoDemzMSGvO0kDoUDc6CoUC4z
+EeSFCqCqRbrSkpUkxcPaSudyO1a7gSzlnhyQthoX89VprcK3sK8QtKAhcvI6hPkVqZhHblUVzX9
XyzS/d6CvFoFBIFLgFRqeSxsLHf24xixeK+PheXITeh1DC64AYXfK9yjl3Q7lVAGCQ5cqphLPkmO
TIgf4JNeW2Qyim2hrdQ/H423sSc4UMwUnlBGCLWO+FPxst+EutFzIURz7biSR7WgPzOr8qHh9rHq
zZq+66UjzckFIfIM9k0x3LtsId6z9/0uxeYue+by6pWUyaG79XHXy+hpkmjXLrbcvxNfl9Hjt/yf
94EpLIZmSBovE6vky+uWLE0guhVe7Y8yoNhjFmenHmkdUMtxQIWektOSJWgNpDXnzrDvGyPjlvMF
0FMLkTtCTXrcYwoFQHbm2lF+SAkTzrP1DIEsK49PFNyzOiM56UUMNYXKKfEq8/m/W92ucAC3+CyW
Oez5ShAYJRdrGMCfcWTq4FKVWrCSljyprY1T+NpLO7qa4z0ZEC2sEDh+U1I8WT6llRfA1T0IZrxq
za3X3/RFdwhQMF3rq5bmrVorriCivgfW+lIJuoZoUmDzG5ZIKgT9quCtKrgA6LpAjOJDj+UEp0Hk
HQghA4QYyEhMfvKsi6EPt2PcGqrqUPZNKvkWTNnxPSR00Ilr2O7WfaoCxgWMR5EB4Ic9ncEzUCqX
FTLVE0PNvQTUGDZDu3oH87vaeepb2JAQ2boVc9vLPMIp+ioPZWmrljhXUjjDkz+Hco0yKFD/zgGw
l2qxWvpi4ZJ1ddc8xHq1apEBc6N7Y+uuxfTOxkg4hdpUEyz5CCnMgDl1BpJ41xks916A4lZMUHs0
VMet+xm9pRpIUvlFecWHHU/6w/qsjiO7v1Vo+5omU+Jv8rxejkBZvjib/biLYAummCa4ygQ+w66j
UFlWA7rMNTogQVHYdjPxfwQ3nZYpmbWAel/c9mnlVq2aWcweLAL8PlRgP7Zi2swPuFsWVLHrSMhG
/Rt5Mp5/gcJZchz+PLRb0ueDrU8d6k63WspFJ5aG0lrhTu+Kc+E7WBuN+e/yNabAtM+KApem54g1
QDmpgkBOg9zq3SaDCbgsaqlk4dqYmmRZH6FkwYpmbumaYa2vAmcLiHgdR4rjCHmKDk4nNC46GUVN
HuCoW3nKjpxLuuRZzqxjBSsA4iYzBArkiQ3bNPKW+RGFtOdPts/kpoDpkesQdtwbXC5lM4Ov1kQv
7SuIGmpYYYddPg78hvL07iLTmggWUtotFXnEKjYsr9qgHI7oHOSR3Pnt28T3hB7p+vDjs+mcOpSl
D2bFga3xFiDCiE/43JaQwJyWIZT0sXfBxDu0ETEPw5emHTHl5JQn6OdhGQ8Jj6JM5ugpERsoq3ge
Dg8gCEKadSw9e9nBs+KEbHHsofft7LlOtOAYngVpu5umcI3eijK7KMPB+JE7UMuMO0jVxhbmMpBv
ZFDhI/hJQtpPVsjmyX9LRvmWnWC2lfiReqDdihSpGa5RqVBydIm6UHbMCWNlJSzgju4tuqKhme2G
Q29T2tq//u6jr4/7XUXq2BHoEiu2qEKpDnZIVF4pzYM6RI85spJ68FIgg5xnjkyWJWZfds7PMRJT
RePa/mXPAaD4W1xZEbcajlqailzi12z1yT3wlj2LZ9EAC/uM1H9UIbfMbercjR59NM0IbvJrvt/I
BMGnmXEujK+ljuNmPXwPVwc0NTdqeExgbfxkoImlbhYZGhOBf+ME2i1e9rE+zGfD05KheyS/KFDc
NdURAt9GY6R/nRnDdq4ZzKPpG1NMCetqALwSt92BSmVMj9AP4fDSfToAy7HG4bNVCCxmWoilXym1
Fv9pbYC8NB51EGUhpkqcd5eR5GdSktnRTL23lW83RczUfaCPpMGah3C66Co5L64prA0rWZlGM09z
vG7bqB15A/3FB43Yxhr1kdYKUSQkylPgBmRh/a/PsWNsVErMJGCpaMVBOXalrhZg2PHkqVLfPK8p
z7NQsOIwCaZ+VcBO+PHPU9k0jAmfspdQfMPq3wYLkvygdge+gCvNwJz3lzoXm6XdNlAoKFsrMub0
fJJ+hMbtbMpuIC0+ER35EqiGYArbuVPo0yaWfMooP9IxwvKqJUBORWlqUfR808TJVQMuNFL/vuNQ
YVbi4uyIXw4AWlg2skEFbE633j+ngD5SYG83KyfeoYLhUF1czX+D0m26C+LSCFVLNFb7qYuvmKLS
ehHrB3QKJbmoyOAbRPKEUTikAHrc36lfgRCXAW7AXT+LCN8Lrwf+NFT0NvvbPM7c+nyYrGx8yw1N
B1IqOkLIzjwcLuzrzMbm+yFnOsaL0jIEZNpmPjbu3X21KO7MWLvbQkkiUpLRkIgzamDGnS8J2RLY
LHTQMouY7jA8ePX7qKhryy/1GfAOaDVjlxh8zXYW8jqQIWEwppLxv5sLeJqGA6OccNE3/7SUEEYf
W/itfY5JKR5ZtLuDYirKttCPk1wltG6bYtkuAjNFJgB9yYzx43JWjjKFel0HOU3iiR6Sa8mEwypn
bTTtezhiefSYU/55lTg655vvmUNkR4UfdcOaI8tg9q0oYziYUDisJixGMXPBdivjPnho34FiF1Xi
UxgkYom0x7zQ5r2CyRNx68EhAKxcyrBibZqFZQEwO1kvcjkVDkbXD1nf27jrkwi99juSA+z/wqZB
hD7ZDUugnd4as6vgRqL7Fr4U4wUc/05WdvF2tEI9VGBWhpZRlz1hdM+m2HlKBxt/7wUq/Ssr8+qZ
Spa4tIMbhJvIkjdGtj+sphm+hmyLTeuoSnbs/fuyERzFmYqMVdrjuv8/I3gCFCSnw8Hxu0+AIASO
H82TgG1x3W35zD3KKtpIKilkFo8T4N9BzxywFVK9hB/JeCy9VJUygqfgT64g7MfvP5mI4d7N19+h
QPTwcO35MvIYIwPjVK8uJNRp/pS7dVuKZYp1FbYJovlA3rhjExu3bnHWM8PsFstaQwjTDRmx5h4O
tDaolkszJH6peQ32oPSg9wwuLhNEat57/ShxvOKkx9GaHzk9GULjU/2aHUcsLj4me3z80ZJDoZfe
iMJ/nAMt/cQxNvHUduZpsoZ4UUmC4VoXuYlr1rAq5vr3kCMqDGc23Opl9EGr50YgZAy9LlO6EB7U
fGiBJQXy+zXUeS/I+jLXF3tcVUZDWsQW6m0BKtvmu28/QcI8aZ6/ium4OZDCtFdFXBCOZyyifLP8
Bjeic5jUsPh9s1dRopZPftzXgM3zA34lw3EgO05uQZDJkO4gQY6vUiJUnAhzETFFaG6mliYwUASS
/cnTQZRKjxuoUCQpevnlt3N9sjM+rEcF44NkG2rP814yWs53I3i0vU0HGG2AKcHlanK6W6JnlRkT
wSouijY3gV2LByNn4zroyPC8HopdGOjM2PkXnfvF89xDBed95naKQgiudG4C1p6ITfyaXJnNX2wo
M411YocbGNzNNLadiaitLzOGcXe0wjhZogbGjfv4I2a0/EMqOfvNnMNLKN1cpXiVjmqyIcFlq4H0
/lWMuCjdhjnb8mcWOUbxFYI7M6Tldjdg4I+EjeMxC1EyvqcQh4bfdnHp5jScPYL+MT6b7024FVSV
+8xnZy01z4VYNm7dqWKog6U0xNoDjuy+r17hsxIEJhfsG5J65jRDxVzJEJTygXKRx855hi5lAmny
56GWEtnMtIv/xMgXp9Y6s+jTjFeKfbOCdGfRw2knmI5NodylzEXMrYViVprNbxpnAmQ3izIT0PUE
rniJ4vfXeiBTSpcjF8MUKc3Mv54o4eqX7fK4DVLSGE7/COFkuJ9+ly7hp8cu+pEAu2OCMlJMGrpP
8+ywWORS8Gspe1kkjRC/6XWzlJNb+UHBkvU9/axiuN3af14/BpJeH8K0NseGlMdS0bTZekFZf4Dt
eG+VcqzoUq1T0Hf2y6fvTDBq4+iBxzE8tU/mGxtK09iBmT1nka9YpC3IehRzXbznYmMn9UKKqt2i
67kgxsSh5JbyJ2gcZvKbASnLdWxtPXU0+mE+4t3UFEgtDrHiIotJ3X7czNOhfLzWCi4fa3N/ocCZ
i7rYjvNQ1CP6m/1GWG4f0uxg9A98ndTMQDXtGsU2fqk9JFlM9IWc+GXWXJLnjnIbxuYP7+n9NqVt
cO6FBuK0uQhQT3leylY6YuRITkG7/dCl+V1C22vnJaGGtIWShsllcBJLUl40NLk4KkRzeqqL11aF
UBRRF6GFMUWP+qqotVUBQul6jW/HhJSjWm8wmiGxcixl9PskbAD0lU9bLg9ww+7S48s9CWJUKoDY
VobgCSwBcheS/84gt3sz3+8VwaLs62lVnYBTlFOL5ohyaAq2f130DvCm6cRD2+OXNeTVuNdJ0XyU
DgiWQrBWbF/dmci1TIILLjXzLQLBGouijsvpf0Uvohuy5g/lJRI2eCW4h5WH1aB/PXXrhZZFDrgs
jzMcPdjiL2+JQOuUNJ37+HlgiFSEoly398NJbgyg+GGrx7pTLjILWJIP0bmAC3xz/O+opUHE3DCl
rm5FzIDFFDGPCZw8NgagblRzC/9SgcQO7rCpkC7ow7oXXEHTtaKmFWNjUk9+cgMLbgdLPEIGO/am
bmtszfvIJudZgPxP908FDzPSnM78QAqRaLk8Ye/V1CYX3VRjbFEI4v4FVwziHAsjGU5bi8wDkBoY
xK4U7LMIdKKobdMEd+phLjwR9eZ/TJEppl1MdLwYKV4jEf4+EzWadvpE32dV4zLssSC5mZ2L1i2X
4ZQEj07IU+CwdneNmmpP8abusK+agmu01au6VeSZyMG1ES9LhnVqVwHFnShf0q2wm81hNl4v45rY
UqgmvP/bHRyychNZTYi67/j4l2NuF87fIiBGeyt0dGwpY9HEIkWGIK1hoQ4Z61zzd8MQKcraXtep
72na/c+qJS93XlgvRx7Oy0MBgeeCb3xeNq+xOdWecHCVE9xVZeWhKI8qFNhVuxP9Uywug1GalN+v
BZ2eO3T3XkVxo7Lag1kciOGV9tRQpGwuSzjLvLUIo19o3tGMgnxjaaANPD415h3fLbCIiBrPV2OQ
bhhJCA485mcq56x364VOUfYEflB//fGJ66NgczVkNGN8nLmvBQGAutBvl/wiZ3psXoHNVKttafsK
X7EZThKqerWOfaOumQXxFarieuz8CpdwQVesUh9lVJYtNs0+lAsCioOUnI7/jd9adiPqEamMPZfY
NDC+PohD81a9pHE0cVoas7KIlL2gvC1XRMSIqFlCUjiGvfIwcdfy4obfGfyYgjhiAEu7GN3IiHYY
KZ4x7Gz/iWSUP3OgS34XyoE8lmugQnE6FqygKmdn0At4BkFa1VTk+XlGotF9GVf9X4mxN05S5Zoz
wcUn7eiyuq/qLR4rhD8XgYXVNQdCvy+Uzs+sP1ibXjF8iQVA2fi0h0EcWkDKyYwZGALqv6LOkH2l
qIlT2FOilkgkRzX1RAWSfljPlaCszoPpFJfpobl92OYNQ/JOXZsZG20mBylQCH4waPNpoMJSIIDL
b1MlQEXyi5ND1ftIOW8RTwktYexQ5CahLFi79292Bydbv+fgcQo00ACRzFVBdJp17AqBYXxajL/i
LEnGGGBY2LJTFQemXL0bITu64k0MCbgmgV+4AvjIyEc5ToF9m5iGRjFoT3MgWDRce8Dl+1iYpO7x
V9yRE+u6sLtcv+HPWw8mL5NTix92TECc9brZAWbVOm+wCse3PFezXYpCDPbyE2aM3d1QeoscWD+u
PL2HQlsWsXkNxiWPqNRnoki8iuKVHALMkIO7ELh3MJ7K7Vyti5ASxr5jTqyW7jk8d1HPq427vgKk
fVI82uvvKAMXi1OOI7OcLMH2Z3K2SZLqbVlZhkdrIbCvP3nhc6DWDqDVe+zBwR5e+Izd4CMNqbWi
RKvApbYksuC5lrMCILuKqBN+4o249ols2ZONtiL9tVf/OMoKSSJsTFr02+CDT3VbRcLB31QoyCx6
uE0YzyA00LGGyi+DRIUBuyo0oDu7GK/vsCuyMss3BLnHayX2o3tVVgENfhh/lRFxEGeLu2U4g/GT
lTBLAzKcXhNOOj4t61C4gFh54BBbWd8L5QSPGyn1lPv8BNkm9bdEh4liaAYE2RiJ6zCw5RiDZnjI
L/5LwCUlHSkUHylAAeCU9G8mNyKr8clAGgBnXiAsr99zrwxg8SP5fPFU9N/ytDukxjjWjdRrXNas
Dn7flNHiH0xhYAKTbTOHFidTEoa4BmRmkdQDhh9PF9/WWIjBvcJRoIHLOXzlMksFOZTLiDNV85E1
pHRGP6vR5/ryJJgZqKhcWu1Jib+mprBNajwuLsfLM8jmWIIDQW9ykxljY7ZZ77zXe6Yxh1zxtJRu
YqxuN9Wb8yiBl4uD6uLFUNDn0Ozy03yF5b3lv6gPXOOhG0Nv20C+oxQi/Gw/ljKwH55fgRz3VR7M
JNOJcSuz7AAxkGppkbKB9xuQTyXHI4/+o9KyHcn1f7nFKdwks4hh4DJHBOmmv4MZuL+jeeFTH7TP
iS/UI5swkzOAjnk4wd8F6lGXGtxDdwXmXOLgq9jr7s2hyxFyeiQo4SLxyH1pYXQ2iYZTn/rmysn4
oSUcxe7A9gI6hAuWuL/rSlbOUj924gocoqjQ4ET5ZvduE9MQ9aacC2RHG5n+as2VXQWW2nEAG6zZ
oZrvTPvF3C5APjBUXKdYTs8/dlzWhKWjGnFF22Fw4uS2C1F7uBVfUM+GNKyTbkrDOWY+E7d60J4F
9eJbf/7OLbPB165ODp1m1073E1j+8m65edr0cvFyPQjbkxlEmPVBby9Bvj2Yj+vhuuRJMQswUzg3
TRxq2PRnGmB6qnEaMnOygOwGpJS0hAkaF0svwkFmQSM/BXpiOcx5TapiIVZP5hpbAoQzDAwog8IJ
G9cAcN70kPW4Dw9RDmwAqs257c1Gnt3+8o0Zj6NpDBNmGfqWWUtrXJRvTTAnk0mfrMLBJqgiKoDT
95IR5534ciV4AV7zNsY0YgQ2hFwyfQrZ11UYclFHxuX+jYLwawtERRIADIt/5IeEFLSnjrr5m4Ar
QczpJBKJ3LYKJkyz0a85JiDamLyf/6ViUTXIOrBGdHuKQeNZ8pKxbArW8kkgP/zEQ/OVqVOe1mUk
RlkMaqibS39PsifkuvLyEpWn47squtBj4cCocfA71zw3bD+9J3dN+4ljPOqcc9v9yftobHV5TPZE
CRcfPDrAVxMOce+vndqdmErj07Cz0nCJxDYcttIoVC3nDrQ9/c6Cah6eBVQPpS6SdrLxfeEbQ5OQ
KurBGI34PZjwZrG7oKN6fklBBJVvJTgSjQsvXNizNz1Bjh8YB5aqBl8jRjcPCLHk/Wh/e+UVZN2z
wqBqx5ej2R3pZwedR6HpqVLuJ+zHMUvY/5SWPjioL41uVeO3CALcBvi4Xm2oGXvar7rbeJhkL3Cs
K5MavRyYfyrrFf7Vr92sLhJaZ7m4Z9r+P8sj9xbQcVZBWlE4DQNlbUyHnqJrO6GSAeMbmurEKbC+
Z4I6nPUgc6yiH5CZmc8N7NgDWDDVxNMK5ISOncjYg2UTvmqxvn5c08VAVLWe4wCO+pcf2rPkMI/P
LX94Xkt6hAnpMhf+AXH3lo9hyqkCtInh4kz423p4uBujzRvXcp6ACKxX68c93Z9+2uR3EopwFAml
Nvf8kt1r6VxqLFzQ/HIr4fBFORzfP5MdUJnzfFuSWf4sr7x2ZVdigZ/zrKJ008QOrLaKlgh7HelE
0Tf1U5/MGkZVZlCkesW+jEoBW+6lVkNOxJf97PH/1EDKOr4jjUanUrL80U9c0ddZrn3H2p+cxiHy
415tdKZ16maAaEWccFJiL10Y1XChLh+yWdDmze9g2aIx980qLdBtZoIw0wIXRrIuOlTt4D8kfp3P
nGcQFQ1wjsEZXQB1BgRNO4sJfxmUsm6zCYkxh7ewbg0QoK3NcrDl74/YeNmUw4PA8JpLSeJ8nML7
gE6OM1n+tNQIDTuip0ZxDtj2nM1fLf4lKMJpDU06CKNpW1s+1rIFk9u6ZLXFDtDZlInqg3xWmhRz
bIvLn5Xw0J4JCXNlKjCtprlyO8NuXWAzfY5ymHS4bPKLhGvvPDV2g8HBmSfmbBUgAAJcpkkf3gBs
7+4PFeL4jER59CCJEdOs9LZeebDcFDvGG6KI7+t2UGAA6GYjA+C/mrWa2MAT2bZazAmlX3NL7bZM
ZOefBU/8QtWtV6xJqZo95yYDfB48BH7PLdRSalpwJ41EsbvxLE6tiPTDyBGbnwAkuqCUlVSbKXUL
dLltEL09oh9vi0k5mQ9NusZX7adKOz8hSeEpQH2qP4adagRqcGX6HWuX7sDSwGqM2Kjz4FET7ry9
ATRwkWSAUdnsBSepZzv4k5tB/YGZlSVLJ1gV/B16kKgqt6lGw+bSsp8SCaPhmlxTDz4qQI8EASK5
osxN4HhVXM9P+iUhe/wkwZ7UrEVFbQbVsXoIAgu/oRyc8z7fdIFqKWgdedh4U0f2FNMXe/FUj3WU
q+lJNqLLLHEkWW/yieTGp4GHSBjpRubdDq4woqu7qIrpwUQE3e1+bpeqHQt2sDRGN8FfDtMKAVG0
fvO7p4DsHfSwuNNfxHbloMyzl3q0WhDBLoEzqo/1gWCfX1XePF3/64vzJPMayh14lQ3/FXgRbWEC
G6+fh1PmNchTKMNmnJTcGOq2AC881Txx93ATuEr/TN1I3aoAzDayqC9IkeE1StMNhORvUXoKdAtE
4lMugcqgrpUF3kLlQi1z6jKAa/mDKBte0elbrkdnZGtcGqGTozrrEi82zn2mqaXRAfLL8LR3/HnJ
5oL0ICDnPtruNBuIJFXzi+JPS5QQ6JWqiSRRPCUumEOYq2d48GMFZUpaYXqyKJL9qjKluvnXjhko
AHvJ4KjvoirIT11PTzvgkRENrXiP8zfbS7oTCviNdQebSlXz98UqHT9PgwitESxDl/6a70EcMTLj
fz79TYz2JI5WNq8lm+1li/5tNR1utImX/glVht3Fs2+FeokZCiYkA97XfKEOHQYWHg+lDUo84bKr
rU6yaS35wqWJ3YdtdM8jkTkOb3veEsEUyiqCNMymAcuzJV6QtURWLRlVtULJmj2NkQU1C+IiCJar
5xtfwbRgFMwcOK1W5WsBbL0ARK4HEhsYDny173wI0m0+GWTDEhrLSmZmfLod4Ob0uTmFftSuDC4w
jdk33nSg++PEqc+xFdCXpXRbttiHz8hWsX6XS9AqrVHa8vTUamUJ22OyCeGn/BAnyg49iqKswA3I
rb5WLkgLgV0g9qX6nfRtWqMzlFou/vr9MulZMRzRFdv0+46h68ne9JVl+0ZLVreRG4ON1NB9IBDe
74vaMBdEBiY7EAINq7ja2BonHRe7RZ7dMq/ngFqBep1f9Pribj2KR2avDJfnpHKNzTyxzPEhD8h4
TCUQGpeZoJ8/QSJsI/DZ5d118E6jjtNe9EdmBraQ+4PmJQo6iKOKJZ4+EFhIfhWg3s73LhEMAI/6
vSu/qpCzI88uWWYeFl2GNRB7K0oe/oDyCVlE4rYRE9RG3kRX91oD9+fsr/ZS4W4rUuz/82h+Dibc
qNAauebIZUYS1zmdWsr1nVy2ofN3QMQOlOShWoealPfePDjSY4puUeA+pV2/oCNJ9AF2cXbdToGW
GltkN0CqoTzsZ4WPaKhWSsYxTLM6y4Nks4tMKTpAzSYHN5JKKcwy9uVAwdITu9S9Xap0Ye3yOgLm
wQK4b6nNEOZEt50KHRGBqOZjCToHKY11532ipaEjiwfVgJBSyY6oIqBAuoeC/HXekcdCaJl6lFqq
+xsZaoa04nEHZGJhrKwwW6x+geiAcs++VngoF2rfYe0cwQnOg4EhS7jqMI9Uy2xpgn/4p0DtraS+
VpqW1f38tLBC4XLOOLuvx63ct/oU2D3lPf9Kiv6/fn+KTq/5jsIxJLh5p1PascJL0nLzKNKuT54y
aZWGvpuvTQrSztMf5B5VYPRZZWX8EVRO943Ga/EAG0v9vSPnVjtQYZwKNP3Ejud7Wcxy0fhSfBdZ
E/sZAKvzeGkWLEC5JcItZ5h8ov4uUlDOuowncz3wkxLMtgE2CV3O3RovdG+IOb6PORejyFHk6REF
4Gg1gsulNBj2Hw0Hdfuyftp8lqlwibyE5b/gT+CDCxCsm2eCH8ZPRE4rsKvbLBn2coQTjcADA0Th
wFBoRBLhNRgm9pNSLbdN149Ia9HXTRQM5HCBcGHIGvl5zWvi7MkRchcB84UiTv3KSCP/kWIGCI5v
psBjE5/OM80ADPUHFnyolrHJ2Xw6HzDHMgfreV+pC9iH36cY63jjEslYgJiXZFd406pN0+yWNN+F
Fp0WNC6xlCRYcc4S9qpfXYurGvaqq8pzCLAqNS/b5rNJvtCA/T/1frcS3mfum7HToXbkB3miTdFl
8vsf9v73OOGfCKz4BFHVjZiHzIz56FR/TCGEWnqh8pda96iPxcM6dZKqbUy0BzZ0SlGHYb1ipykr
MZMhGqClGf0ctXZwzP+cwhIphQT5j+j6Pg6XlmBc/7Nx9KOS4ciIK7hdJarEyc0bf7ClHayj+FRk
B/xzDb6NwGXWIVyPPt6ZqUo/QOqM0JKVfJgikIaoW8i3nVdYUiTZyv89S7b7bJeEUUnFkQd4G0JS
ITCakvBZ/S803SHjj1Or/pqa+H5FrY+w3kkraPlpF8d1L9KA+4iuQmCTHR0U+rvg/dTpbhuximBM
ZMoIq0/9Rtreu4RXZ5ZCvqZvPWebAPpGRVEU/qCR1hbeZvnRq5bg7XZm4Y/+OTOoaLJ76D+t5obi
uq/NXusBVtb3A6Doe8kEHiwcARmpUUWI8ujti1IP7kGg0VEluDbMKwKjC0EhX7m05ltXM2v5Nas4
Q1zWsjSehi5DD23QM7TINV4dkJhg1nU2lXp77M3d7UnfPmuu1FfzA0PAXQizbrywYrgnzk30njgi
vS2N8Gl98Iqqtt0+D/StR9N/nlBNJvfwK1jvIJtPWGw6zsVTrMEfI0C3w9R7uZGURjIAaq6p1Wdw
h0/YzKq2tzG7I/aXJqrpnb1ONqOpIqUca9jTPm0T49iEVORltN70sy1uNb4GVeHmdAHXCpAS8vTa
AiKOX+XrtupNlgBKr46V4g2QQMWJbqqIUMsN9FRPbKBG+b3Tiq3FT91UiVUpB3zjAaAE3pAPzabO
katg0grytEDZ891o1g5f0oKY1IcPsTyTvY0Dc9bmvfHCsx9fcU7z6rybWcvClSq449h4Q7GuPeca
pENhuNEKKq+/eu3P8AWoDSdI/KVCujDqUv4YXTOjGnfq2TSTsyuKp7m+6qabdfPpTVPd7HYZzQ+3
yJb7NjddRILsO0qLyJVaHkseBEbO836kTsCr75oIKwQMTwtNwhL6Jiy5Mx0++HlSqLaPVQn/kLTJ
j+8NuUr6uiSLrcQ6iRiwBUNV3392tI9aTqdtXB0Jfrswv5aoOKAAso7SZa8MCULuDB8D++/36Z/B
Qz6IPESYc4xM+ULRHzXhWTHOQYx5Mvx+YGU3cDGGkWMCN3rLRil5iTj8sPOTXk2CNKRbcRQOxrsF
g92ooc2f6PUUB8AvuTBNs3vEu1vqODG6p3xjgW2l+IfbQrYXD0UdSE78Qvj0VcYzrlI4Tg5CpByj
8DoZByKeeoQk5wcDIMRsl2v8bmRjSAK5I0PO7+Brgg+jJoNtlBOaqNVxCTr8o7vFPl5comZ0zTaP
4XUWEhhRPZXGbfhz2717T95bwepAyGbaSP7wJeOKawlYSKTCFwkyHcYqaCz93eAGKIrnv0VK8QBM
FNm1Qa/+cFhLDklvIpBLZJTDD52wOPmoxmQLiyo6s+UC1JMxXuYUvY8M/Gr/5LFo3LTE2tDSDEuc
XkOQsrZg6u/nWuwN/waLOdvMk3t+39W72BwHtnBQzF7/wnFWQsshHH/EFlhfy/fzxzXnhdzYRGww
PG/v+tjsS12m/QG+s5eS2a7m9SPqa4/gwDUOim6AhPiFv0AK0qD1iY8Xk3LQhQJm2GXNVC6JxcuT
o6CxJKyRR1ubpLNnjRtCDkK6FRfSYoJO7kDoHjb+JSa29o2S2mJwd9tIAR9P+1r9+GcxlTRlZc5q
/xChZa8z2oZpdP1tGgdPCoJgVcb9GolEFSWFGTsNdiAFslfPg5IVNvQCFcWhFIgafCv5/tLTjxdC
w66T6+EJOB3sMD/J/rBOZIFvPRF1fI+rRyQBS6S4npcYROifIMWoAj1BTncWCxbZl0FUXGoUK/Nq
+wczBtxneVRjCFpu2Xppxhi6JWZY4Frb7efbKS44cSCt446K2w2zPlJTo2Zh6bj5lPM3Zhu6NltJ
F+QNfdUgCBG6tcYMhFVnxwBBuB0ejiBmgjaszVgHbaVE56zI6Ophd3CTe0EqE5QPTJiZ8Vp0yUck
61NHCLhmUd7t2kJtQkF66e0WxuEr3HAmz9owCQHG1dXEENrlBGT2bT3tjmdeTIdXmvKLbNZVuheL
v2IC4eHyqrudLX6LLWPNp/KPwSG4i0MkR9wF9+1tB/fuSAcDNEpr3mXypmISUdR9Q+1qNy1D9N+/
cDxR5ipfpxaPEElGhrwRpm8Z0j1kp3bQA9JDGYL8ELn0QuOBhCLIh4SF9j7tmNB8kC8OLlBTIUHh
zNf2gZ0q56g6Pmi7ckWW76Xdm85cTqVFsZAb+HfkP383YaHNR3qrXr/nR/QaFzL6lwIoisVTMpum
QKWl8fJX0rxxy8BhSS6wfITY/oLwbv/DRxXC3ZnANg8DkJkJykCJhyRpUDDEPsQNh2fRwrVTTkC6
YeVGnV6A5lHTG0y7gzbpxxhtiZl4PB9J+3yPXnQKkH52rLVxngrinegxuBewC1zblGY4XCHvYubK
dpdlSKYoBpyLP0ZzZ3mAimrkhCT3tm1uEyzDXB/nYMtwYZ7amTgypVUucg16FlQsP0AZX1uifHeB
4c2shOY6ANBHCwVREuAf5gLbZ4oL9NXW1cbo7792VZcfgGEBwAT/zzRr8NriOt9c70OKDGmar0Y9
BUHeD/0yggW7Dr20Q+rfAehBC1+8q9L1Ggy2+gu9QPBVmgJxgezaCKt/FzulYIwTFIhr3CxtBFfu
MV6mpDjyOmFhbN5eHSGAp8J+3uz6UKSXBNzm0FrapFW2xSpCmPyPqzlzi10+C/1XHw3GBNEkpDdb
UjuBUSotFeXx7YCs+p5WtipFjVotWNT2pGZzJzsfZpibnUFU63uJlFKwLZSUpe22szFWtUKmry+K
Itvauk6EtLoqIYojHeNIa+NC2IngSvzJYhJXqZe3p95V+9TFj5BnF+Y08C7zhbvXTn/b/UNXel+z
gA5Zzif9Ca1Ju+MdnZBTUPfFQWGtWbAcgnx3XVEAJ+1BU89eNZ45W2zC1a0/svxjNYySO0RsRAUD
NiWtJnL4buKJVI5PEP23gszxWKIk2HLWfSx93qAYipYSuuDzKfrKH34IzEFeMvjhOu4TKeN2D6my
jFP4KgDUJm4K9o14ilpPueL7Qux8wNbohApT+K/mAhV/PMDDYJ1VWNsZgngain6pspYLkvbgQPLM
3FC/wYj1oJuNnJEyWfsNLAONu+PDXBVndaRvtfupU4svvUYmLdq/keDXlk4cWgMxfAg8YXpPHEg8
aq0ddX/W7fewY6/l8qVdb+MaRUb0KHW/krLHYQkMFY0XG3V3GAR7MbgcZGugIsVOXTVdWCyUEduq
AuXsBSaTUZRFathviNn90ha+pPITYgDtNolXH1/5ZIjRzBSBhfnlqHyS78JjcSRiPl0/OK6veGkT
JJrRp1yRZX7+9kb1ZEenyQvMFQnPLWB4L0Ruttcf7HC2XQV59xSTj1hfeBGGMu5imRVxwWSYaSxD
kKC2a2ldqXrnjS0z0E9vh+zRB1hxKlyK9MA/LWFItdIBEu2E+gw/xNh7nPv8qISCWVME1VXnB/4n
Z64NN8RXw4hxV8LCLPxioj3vVL3om7tFsgqQcptifUKrbUZJMnEIeyDzV3XuSxAbKlK4xr8MogXE
C9Dilr1M9h+dNvSb7BCzcj4enH6DlJ8v3GeZxSTi1vHaC4wzNnXfEzSKexxhiVVOZhzMFlclac8G
vlzSlgyW0IzlRiQDIypdtKDyQrm0kF6d3P1Xu1p8qAhLyDnANEmjizgt6bGNx1S/j+h42FCC70v7
qvVX78T9Kv1qeVRGMQpDq6WmMnozphji68ZgOOnX/n9b7NWXtxva/uwrblyJnqnh+takTjDC6fo7
FDZKFjLswdd9v/7PYxoFeyeae6yeEHBw/FRV1pnLYxu8xpCnokz00Z0J8f/bifmPbqpHSxcPTk3m
ozOgP4qXN4yDuYeJLTRuUl1MnsCxUK19/y+m2kswwvS8VKrT5ODX5r8LkiuIv0R+/oee+fRJD1Wg
NyuJHX0Maxd/Kf8T9JKVXyWYUhEhcm3peBcwZ1lFCBiLaaxKJlquane0kGTXEawVYlkENIk5EuAw
thSswnB21jrxVF5GLjxxhlsH/C+ikCTmAVoj6Yo2gUqYbTL3jvrrPZ9bhzrs/XaEy2gag9Q/Sk7q
Zu0Vn0Q1+1VxyVT115K2KsOK+2RP7XVNXxODDrZYXvfhXDasur8WoeVs64swvIp7ROVH5LPCYYTU
638FoiUCUyslgLuyDauH3itPV1bjHZDG6c0/ZnNYa3WM6wBnCLCqiXwMNXM+ojGlDsdyTVCxt0uO
K/fFTo3VDgnmm0UB7/xN5I/WuyRb0zvaKHbDSgi7yr1n5a5b0TtAYc/9X/vsZ2TX3bFB5jGFKb6Z
b4utusI77/ze2XzUi2+CMtVaoP1ufJF5Zd1GhDEfop5QYX6RtJoUM5SRZydM5d8sL0qmtpHg3+a5
QVV7MicjD7bb0WffWbCLw2WiKDBueLsGU1+dCuB219kTjPeId32BjhL9r732SzDDeDJ2ddqJUaxk
INjeLPPxcnUBfqsDC03jYIuTZHEuO3OIjX+jT4VeN7D58Qc/Ew5m5MTpHuuozSblWtPKlyOjUEoK
/cRqf9LVInIg/gN6HlXzD3q4RSFwB+XYrjn1RiOGea1ZCmEKiVnx7oazUZnBGVp/j+wZoMRch49/
pRpnY8ErGyYbxwtZLOo5hy0t9O9CswjzKCpx16iIldJ6I92RCYGn4zZ5T4DR6jkYrWcuHWA9A3v4
xnqTtA999bTI5hgHoOxbjaj+ppILC59Z/eP5PJHvYfQvE79guow+V8/Ey8pnAmoC/rpTVFLjOYnY
RNeNJkyzerP6muVDs35p9yzUekEt2u3+M/27PNcju1vSRddIx7OdcEuMSgtNRTzQkLDTp9yDMuy/
6NlN6QDqbHYV4a8C5NmmH3RV84RV3QJpycucivgZM6ihDAyS1VN49DW4BnWcBZIvX+7672n2llqi
3l0emnwqQ8b+xyKEpRHfHErGyayMGtj4EpvCxJLvWYEHc8OUnDUZFeIp7geE7k7SfZtiz7hFQHxn
jknIt8XIUFQJToXiMOACs30TiEeqA4rXl+n9kb5RTU9hi/veb3XW7oS+jAQwPacFmOQUq8vOByAe
57s4PWjYaO63VPQSRaqLj1ab4ogBjvurP0JNlL2Mf2QWVDSSds0XmgDJNzGSmYd0zG1YH58iKK4r
xDI5cjiagrLTWwsGBLJMgaM9o6ZFdSeae/Al6lM9pqSsqqRUD507799iY+JDSML71BIgE3NBP5Yd
QxPJGwcS58/HAQunktKMxJCpo0ZhvX6BGQbCGWEro3UClhLfhqD+7bV0iIWEz5J/ziHQ9rh2XjX7
nu821DR7qsw5PFyH4oDk++Os3p/L0+p2A3gSK+JoJQK6MOnRYCYnMIVtvhMC3bsMW2GiHciyPBBU
Fc89OmzBfdgBuvQOidRS8zQP5DgIcO0+b4f1hKcwJ1Y2LlJti9Ap4WPeLmbEzZt8OkHFqy74CR8s
8+X13iON5ch35lagYttZ+r0LwSsDNjTHHGBKkwEWtQJmyign/j9T61lzARDzwcDhXnZHz7IsHvS3
MClcuRaDI/KQjpxzmFlmpXXQR9mxbhyym7y62ikfy9GkL2naFLpg4aRbn0GWXslL3k7R2ALhNsVa
ahKS9Ku1PoT5ePvDNrdz//yGc2SRosFW9STlP0yhcEwiUVQ4FqEvEKAW3qP6IFRp+Sz7yawEx3sh
JbKa147MA8JhODoM/OBNtWWsKvizOridpTJQBqNoqRMtCeleR/bx4UnB7mZ4jctPGx4rjfP+5CJW
FpbfJ/hQToMuxz6iHwk0lldYHww+A7jPYXCzrEWn2o9H4+vOOpdw38NTuMneEv0M3xeDoG3C/QWd
l8sRvzSv10fKk+1v5kOYFMNxEwj+aDFKOUvUkLYTU1k45xMvvmohY/spVUWf0gEHTyWBfet4+NvX
awDyX4bZNBjA3NOh5KeTvxWqnALFNqLC8ChOo0lVQKea864kSK5oIbSxQsdlNGXrHEMQVp5l06Dh
v4v1QiIVno8XfFXsmCEN77/hJdRv2bkaNHUBqSPM9ncuY+xezO86SS/20Cc+VqPWQxNb0GKRLQi2
d4xl6WxUI4Ie08P8WQ5qqXgYk0nJIWElpyftvVn0eHcV6Wk/0VcZ6mLMDTggC1JuEmAr0xCTauZ4
gOIOFoGhJ5JHujtCL2IAOqf3vvbSObe/ZUt55TF02docXqpJZNwByUl2cii03QVDPAiefMXRFctq
1ge2g2FnLLAYpZhNmFnaEsidiCqTmBdhghyL9ZPtFrxpmtZ/b3tRjML9OwJVagz6knUpgKd2q0Mr
yusuUZvwbb73XFmtmDyXQMxO2OuPB9oLdvxANju1wnwN6XNmfRdLUsVzGKof9OzEROhbEdiTcLPn
LVaBmkrPvVauU0/WL5BXUsYQr+cecXPe5hQLi2KBIG/bJG/QJfyI+W9e80LIUjPJb6Lv9CYX35FX
Tg+1gxpnnyOO1TWub6zEXT9gw4ph9R1WS2gSpSpVEpP93BrTDwxzjOyYisFwtXdV23SoVnRBb5Se
HFgfUyC4c5PVdCpsw/oGjU325b2FpfLb5xRe+yVvc/CZQADzaP1UfYvBRoz6S/0qUCZbbSzUgiNi
ijhzYvCKcVLWMyFTy68E6VdEdgZqB+UuAIafD/O8yovAChF2XRBKpkzsCR71+fmridaPrna3CVXo
ftXADXQwbVmiP5aKWZXpFA5w90bQxQTjoRh438YfU7bQXt6DcBE0UDkOdkq1Amju0MQDSI6FbPFy
i9Ja9944QY4mdJOWO1pHTeA9C/W/5Mg7UjeOQy9Arl2ya67zjlpC4PhS1KFIlQLKYbINjQDfSCc3
Lh5KnX9h6EoZA3H8MmLr2MkIef0LlTWRB9GhsUgdhkyCdRVkAmv1l4a/TOV8CPDHgjuK+Vnh1AV7
AkRshUfM7NN01n77LDvakg8zPTzm0wrEx2AMPTZB2PlXvF9I6jMsCe28PP2DpC5iA9/Qokg5ZGK+
NsSs+6y3mwCXsbEpjKC7emuW7XhEcNita+A615s1xDbhm6CxT+CIu1ge7lv55PdPkqs+mDMsUo3C
8Z2lAJjbeA2q/Hdt3nNifvP78dDp10rBu1I0vrhuvsPTa3nmz3M7BeRHtsr2lDg9qzpZyIOw88hb
sgeTwm26baHrQOwHBZf0E0QTxpZLLnfkt/ZuDzGyiZRvczqGyVaBRXjELt+Q0A6XxgSvIzW9DAZ4
MjOS4J7Tx8tXYG6o2SWFXS7u1E0HKwzyQkYEYDl+DK9zdJj1hqE+hlb/2oaTDj85Wq0dWRjmzrB6
VJXmZ9sqO+V8nLR3g3zDDB8PRbf24aoNsQ6886dCskHxMRBjCmlfujmFrWKfX3SIg4hv04AsRRD9
RwdpHQiBkerWcL/uUkGIYP84JW3YmCdqt0UCrC+988SZo0i/CRueOGxE0c31ohUepah6D60vJUX3
1r+I2uebY7JtJTaIZHpzXj0iVUhn1TqBrzacagwwyXknPhZYm6tTfK52NKsM9vYzytVkdzGIN+0w
hG7gd9yM3jrofIrh8XV9DH/tqrH9wx5Eii0zW1MyXshDxvFCVeD6R7gZNByn5frWNrd4IjJHackj
DcKEqQY5A+x/vJu8JFQOOAtxUeFFxJPQQQ/o76i71wY/NIZC6FMQZutuNzpTyRju7s+2oCxKL4ZW
FBUvIDkpdFUAgulxpFcPoRuRb4Pb2z8LvLDMKZttKWHTMuS4OqkK1jXVFBq53kidKrSxURHFgNn3
elw6Zh/DR3/kIBQJoT3AV+mYt4VdKElUbFFWF583REuycYJwKU10hMbc836MKNd22dwhDdH/9P2Y
tmhPvKmmFI1T43tyv1wTkxnnu2q4GCsc5CLvfH6G0eKDnHbkkDn365vAGI9Pho3HvWIhSHwW9rSG
K2w2fmoPjQ1T4QKaJcGuoJdvGRows3ic5j3wisIdV+QM0ECyb43X6carlLQoWs5Y762LxgO9V6II
TauNBGt0XpO/Y89QnlagCpvPbc7MAmixHuM7yveDsT3AVN/VGNFHyHGWZEZNaA1HNjMx0PK+bElM
K4KLqmpqvL0f1cDQuEIxZ8drNkpNYVt1sCg+loMLOVT4B0m9xwqkWPABgq1r/F6qVbuoIJiOis/3
Jxl+O8IXJeQU3v+ZThWWGaHLsQ/FK2m028+jaeJDz7U24YmunP3QtzbsG73mT1ZZQMELRD+qcr6p
Y+GYshkIu1FL4MHWKSekX2ULprjDIKLdf295Ou4esIdJI+a2+i1mfNvzXa7Bn7Nkky+bFmL8Q+6z
/nPcf8/j4Sv/JQX39fHxd4sb0Syv+hFGEYHHHKkzIw50IGyRF+htZKXUarG+VNLRi2K9DWfUXerz
OKuSllYvgp798lBY+1rRqH0AKGM0tT/nGy9npmd1Him/aNZGbytZ1l+d0FloZ3euFusnysh4gqlA
RJ6XCcQwgRZyY9RLogLjK6skpUGz56BXZWm6xP/k82le9OOtmuWjUW6D7zvWkqCGn54z8g6rJQ3K
dOI8/q2Yu0t8CMK1Nf1LheeJCcFOVfyhIohwjldCs31YW0NE5j1GqqR4ERLIDp9rpmi/bOQLiyk3
YYyRkyKiVuB1vuCcWkGXLMkfrHlJtOo0lRyCvsqCru3Sxjgg4rxEgf27lAkdDAq1uW693H70WIQC
i4vsZRj0vj9pao355/4pZdtT+in8qIdK+EnGa7vsYYAmuWj18MUUJV55fMovf11NCTzJGnKkRz3G
G2jESIIWIcWjTB593nyXJIp9Jb5deEsi180QJbZMSUNztqLwuYTgvZYSOtRKi0h2nY/nkmXiBPwb
2ECtzOUVDINjidtJbh6zE16mVTQU607bz19vxpB/D6BZ08HCCXQlHWBm75hezwhLLdTu4pfWqOw3
6Gwz6aL+xIG5DuxCkv38DfosB7Bn7H92TwVsAaqwvzGIf2UbBSbFQ8euz4U408wN7RPRlJvT3JJY
Z1D4cZz8+HCTmpidOlu9M9BxSbfYD2L/QXacTmdh6Hy0KBCbWobbqzhcq6XeySIawjLYsrYdt3ei
ZoMXQ7tXBPplL9Hh+bSv3x2GIOb3gEvxBW8VwJ/AOtEhCDXgMPMqBF5UUMOjBY2d/ajdIQV66JbI
m5A7CYUCAeX/7N4izmQjkkaf/xuIMpv2Z/4qSjG8lP9tuJ5W+gsKL84516+5fOUQhZbkUsEnr8ol
iNPmH+cXSxac4+4EAV4nTgTCj/wUWd6a4sZpyFLXNIBOwTc87ETLLPgEttvZvPFPG/2Z7oi//j8l
AfijuXCN3rYbib1aPkpjoG1aEvwXO5qh/PHZzV1dKigGg6b1Uxy1bzN5+1P/Il2IFj1zt3RGNFRv
irULRfyWvKSUiUQGpWWBZ3NJpL+s7uCuKsxUGzAGy/B2asrHIej+Fjv58sK/7p8vbCd1MgJ4sn+0
yE+sIrxo0YPsdlNBwcrJJ+AxcAoP3MbvXSDMYjJOjMF+ylGEiTxCb3Fc8pNdccZSqOdW5zIRddrb
V6OF3uwP6Hc44XXBFlPP8pU7zSTeXJOeXADebdeCzt3715Y19UXGVxhz2Uju7TmIWcedYEIa1ymH
P5XYEY2fFyFayHmojzKvoZTUXEI2RgDfaE2efR9/D6oaADkdbpo8kc4epLsvJSRm46n5DqxNbcWH
spGb+vzIoR33d+3NnFtOF6mav0elTiKt/N5m85I4CJ0wHTYn8aIJ6BZipcbmdBfxp69m3rlj+pkd
6pqxg/DOYDf6Y09ItXmiKfZa9H93CMBmein/jWBiL0EMsoFQtGq/oMpXkt2MzVvcLZZcBanMvEui
KxvHZsI1xGUSxXZKgqKh0W+N4olVZPINx7tWKi8diQ5N6l96kdMdgRTeH5T7FwuxzdnxNrXxM/W1
mDkBvPPa6clurYbEHIcWJC8p1jBih0+jkrL4OJV4pfm+kN1NINSv80qT60L1Hy0Jh4EJeyAqOVxM
TFHQGcv3efWS5e/kZ6JrzLVwknArSDZyzpwJqjD7F4VNz2+0LoIAMFcZdnlbDvR+iSwt4YAlqLUT
MUG7K4yG9NTH2GgEfXD2gZctmf2+Fbqx9lODyelSZRgYrAd7EuBXlYNjr48FAoJse8N2/rU0AzV4
eDn0Xkcv0aDrZKoTnOjuvzsWpLggLUQmW7j2GvgZ1Xapp+rRxqjz0P2P8LJRiIu10XDy9aALeG0J
oRMTe3zrbAMq5M/uw/tKokFez2q3DLHeGoQE/x6/HQSn/bU+CvQlbdSoo+w/g01PvUh84P1s/qkB
8ai/gb3PiW7C/1V3bXt96MyNy060lIqqq1ek2ByPF1caFEXOVnFzMdgwSXUT+6ci1kXV2MhProYr
0Ap75Q9WCJtJwBdxv3hITIbq2FTdo3yOy/+jR54P6HVJa45lYJvXRKCR8ISZXsniKSaCvyCJ6nHf
wJiGdUUK5d9IaSKgGr6Yq1Bo+gxkl1LMTOjP/JR5bjoR20nBvv0+OqMxSDJOfAgRLOFW9uZe0hFs
qSRERzCpCHCLlqVgXWg7sbSwaIa/gS3dJZNWEvYSaHRDvJwNs/0abpWNXudljcpVTvG5bW4l7voE
c50j/oa1/ydAi5LKjtn82kz5DlMZ0ABGJc3HfvivpfaPcmYWpu8j+NBrALFuOKAwKFsTdLm5GSxW
Jw9qBO6jMreEM3uBusMWnXYy6KYfOZEn4ZgodTWnO0lPlF8N+gs3HIx+CuzAkPGT3/7NlNiDPBBL
AE0cex9dnOFwdhCxXvmRAOcNq1LEIvzYjLN6COozHSlZo+ePgcr8iJajmmc41A8+cAU1Q25jgK/3
fFWS2+t4qqQbH4FB5BkkMvRrOH68/PNxCAa3uhbS/XmrNt6iGqV9AMB37LKXLrmByzU0yGP7VqeX
jvVO40ThS0dy5VkBOl6mFweSxuVrGGbGk7DiOuYHCX+Jm7F6qpj2ZTFS2JJLuc1uEI08j2zIY6Ed
L5WWQuZXX//13UEImbCSWO05uJY2/G1uJDU0evtmUW8YXTo9qcEjZOJheTtRdvw5LqrtWcA6i4mJ
e3jJfjZYy1uwKMupcbd7xBLvW/2F5LGYoJXRT2gCfKj3UNZnYG5oh1tcKQXFeOHrgSScAKfL7LHF
jdALZTwmNyhGp0dyLn3T6e1K8X0P0O56LbNbb+FbxyAPR9Y8dLIORKk8ro9lcmy6z3Dbj5MciOIy
JnJsNpXuQ7C/VmHIgjMAI4vqjJVd6TY8VQ8W8R0dGRkFh+gIsUmKoByJprZI4UPyKYY9Vx95fP6S
Q5g65Zp+qE9uKlfw/UM1VjePlbJzguxBoMunGyNtwOgwkCtcUFMO+Jafi8NyKmCqTovngmCFMZ+O
vmWtw1vzDUiMsMknCpZoXCPJC15ZAwoDQYavWG3mhdYREDminaFsXhyRMNqajQ6ZyP129j7BimGT
dMpn2HDCJ1unu/tWXLIWAX1aIEGrlQ+PNN8DxeFG3vcJq8ucUlf7zRq37FOnaDUQO8ibXfXdPu7L
EXmLsHHJUui9XlW2Id9YCbZRnKKRBRZKakVAZkApPXR9WSg0raoTX6hbJ6HRXz+7o/fWt7G6mPKL
yfGv/vCoX1RiFeJ1oeHJzqbIr8JA5AYFCkDd2wzoIctCWdmq/wrBhfpNtrCFsTxF7ZtrZ2DavZ8T
fChWXmNrbRVwx+4h3mwB9wac1irRTEtB4KDH6XlwL4v0bVVvOwO6dqdXFPHTLfQAJjCPHT7xcZaS
aII1y2GdKnr9gVfln6dhuf+6BdtD2pxKQPlk5xCaVdHoikrjd2OWzduHQaVpbTOidI0v/HGZo/p/
aQNbhzZq3dFZSOjcugv+ePzXvJUA74N2QfbVZE6CxEjAE3ipuA59f5gErR40GdC2TX+V3wHEF/6n
ylOJHJB5oPYnE9GGmpFjdF8rDhU8Y9pVgSiWzIXBREM4ED3WxAqtWrEs/eXPNzmrA3agoE/Bvqip
dOTtHbiWsvAb/9W+nYjSgP9tPrUthmat7TDTcdGT3HpkjWxRkEjO7JAkqEgkjKuwSf5ckUWA9ovF
duc7XXvevX0a1Sl6cNjwW3XQtpgFBo2Sczh85fjpI6vRgkBNM/CLcHyDViJuZQo1nTP9vDqQeaQa
Jv/nM8yUwRgcnKuAf+BXrU48ZMyfXfS2gwfaDWvICqRFWwvkFFhvhnFpIrm0CPg5ogud97tUBNeJ
ykvpsuttTY84pkctGm21rokoGOsnOS2A8DB86Vy1VVC0bG1pJOzgWnt6CivHv1IA2P3tJWXv+RTu
wy66jcb4Ki0kSoIu/u0pTYizWLyjoNUKRvzD0VZ9llEx8dAPxTz2eE5IsEZ4/31XGZ0hKSTG83sB
pryy8suWqEJ/Ld8XEeGdQyoCmSWxlLGcpf+1E1D3LLjkuXkWkfBNIztFBzgmxaH2TiR9slmj1UrE
HM5Zt3jKaLbMQcLYdYcHpGfbUyuY+Wao5oAZtdJS7OcjF5I8pWO/hGFomk8yCeY302FnBPO4GTKA
SpuNvmJmmboV5RmTUbd+OXB0tEaQY7wCxmAdD/aqgEnu6lfMraqiP+CD7RA7fKMsIMPAEQMIvCfF
1OFHinEyxPK9VLcQnzdTDc6iGvhxC2d1QzbUk59O+HLeeVmG34eOuPahHGMIfsvFPLjPrXqG2EBX
hzK7uqrv3KswRCELs5/H3lKMH8LbCpfTfECBdi3A89tZ65KQVT5/n9vSklTW4JXOEFEqEcB/c/RS
r2tz6GnLMf41OaWeWciT3HsMFPuer1BzCspdNYW4+x4/yHrKZBfseYDHZGvXwDQxOWlDKXg03PnN
kISxF3awXA7P1cBjVeHu5CKx97bVsNImtaplDEMYtQQLnVmDzbYdmb0LUkMFqXfQMKPP6KnY6jmS
JlEwTrsTNtFPtBvMXmMxjr+Myj7P6L/Y1Z+dRjcAWwNWpuf16/LiR7/0w3nDzUiccms5OWHpfFca
UU7T33vXB8nglz1HznEvygyQMqsNuCLkEWUWptt+WvKpHeNxXRWB4slt27icpCuYo4MbUJ9dsfKb
FVOEMJwcVCYjtBp6+njxqmNV8C0/bC3xJMBrj2nnxwXj8ajqZ7JQHcOIlhZUn7RihC3q1fjPFgPC
XcDlpSMtHEhHr4/Els6X68yOzx5cpoBaNFsLZsCoZn/b0l6WYcWPIjeOdVJHJBauVUhafrTeVZR8
YJOTKy/EwdThDWDxhQfnJi3kmokne62HSDD//O0yHbUn1FN5517CPNWcBLoZRfDJdzeIrMZA/Vrl
Ra+irWfD3PvNlKgwOBsmAO6X83HfwOuTObk4phNSg914buZMpMSTPiqEQtACW+QA73jCWGlpAVR2
Dm3V8DQcwACzB68i9wn4qtDjEJuTPM7lk908sd8JqmzBkfIgX1JkQwRTeSYeZCeoWt6eeQKh9p44
q+/WC0G7CuEaW/0NgXpK53Pk+Fbr+2jQfaiaz++pgzwcVDeQLC7ANWZswEl3bkL2RvFB6dseV0Ib
pzUh70Yjq5T4Y7R/1w76A8gP5PDy4Xkrk3ifLYocnxn8m02lgUSRUU5BCuNRxBdiMUuyYaxLk+/d
9ktaJc8GOKMHUExm0JG7jpBaYSyPGKNROrpnvZmTac4sFFpTdkLXgNrls9oQGioOTg1o/FLx9IRq
d8twxy1mfW2aHdRDyTmAMtWqPbhOJB/zIV65AN/kHOrTxLxOSHsQu9QLjxRcfh/2NKw49GsvLNyT
hMj/WHZXOl/YxRQpbf1ob/EOjHqIgx6kjHD083s5XkJNll++UEVUX6Oxo0YJdYi1oHWzwgXSPMcR
5P6P8c+C5uk+W4dWgtmSP0jvMUyjKNazkHVc3WnWHRlhmWqzCA7qB4Obz2sLq/D6yOzGGiw2amGx
r6S9OWBuX2ncm3VoZaaMFauG4LeDs3jE+uN+WSbkhiRo/0HH2GHftYlub/4m2aWMIgpJPBVocoLW
JBu3rJKTjE2z5ZifXpkMtrBLTqXbUQMR2HkK9XDQKfzjERi5o38vM8JbCE1HwOc5+pKdBDMZ4SNM
/slrno0/Nv4mSRdCTYJxmyJ7PK8UrG5+o1qv/3jUw6tM1d/HRH7uIWgNCUp/y9UVEQ5fEV1kPxi5
Sx4HxmIV78PzPEL34L4Nxm7lmlYeN6pqucRsWl8EIdMxU79nRiiWtwM9VyderfA3sINDhVYsA8JE
28RmZdmytImFQwQV7npTyR+00+yHxPmTHISN6XolocI70SaZwyzTdoVyGjVsvAyrfWcFYAfnxohK
AgUaHuYk39+pu9AcUAsy3jpVm12TethTb28WVwSwypfjuQYrhyzCDbpBKsTg5yf5I7fMfMQC/aT/
XULUdT1nOs+BcuttPkI1whrhfb/wYlp8n6Ll8PyYDt0nmS6gmV2exKQFSBOAaAMkLTZz2Rdvg06/
pee+vnv3ClUXEPZ/cCan/YFF08W1hzxJ/paW6bhgYoPDV1Wz+WleNtZEQG291v3YDXgAziBKFPPb
OZH/1Y28lgCNciylwl2N88XNTRgmtGhVrMkZPZ5od37SSs906Jq4NrYqqETu+ewZK08emRRVjwAv
XD5teuKZD7sUG0xa7B00JSnLBRFfx+8c20kIuaU6Dmkysyr7ixy6M9Soo3xOurpzyx8KVIN3wXJf
6QkKtJoPi5GJLSJt32BXV6akGkuNeKb6ohh1OU4H3dfwBnhQmQ3J+scIpGvlCXOIz6Ky4VKLiIi4
2EQndQoS50lV51Y3o4MxS0fIrHm7Ip5928lEVgRsABPRXlChpHQH836PsJc7/9g1WI8eXih5EYdf
3XU8o9UBCsKI7M4AnkfMBJLBmb6pvn40vB2E8NRVfE3oBP3QMOZvaFhIbPQ3jrGftKIb+J9G9pCz
o4DfUl+YiaWzb78+kemu7fCJEudwW2P081zuE2IhmCbw+HMN/Sl36QkXR550tYMqU5tDf2oPcqQi
S3EcRVsSBiTjwr7uFWNYyQsP36WN3gqde/F5zdteKPjBPJTO5677TZg70aJRH3Y1PMscBQBAC33u
StK1Tja6/J+o6J/PZTOTJqCVU/jlzbfdoJxY1O47Z7Gp2n6vIdUFeqQLoOLpo0qLZS8DlZrXyk09
43XtCAHqz6hz3WiGbJeE9/6k8ssC+GuIRKedTAal9vRmOj0nFDFQSklvViQ33Vyxp3x5JDU1YqP2
rA2qhM/KhF+9IJ7vEpK9J3dRhN8/sVyvBpdFtV6gh7w61h3YoNocezzpif7pEOhJcxW/Ib3cEi0N
o0H8EvCx4cjYaTAIzCGGmBvfSv+rqmHDFKJ7gjNkrQXLYcFVwlLyphTN82fPnP5kdtI+OTqyULER
nsmu5TZWaI1oJHm+KXSp8yxnYEOgYZaivsGrADozefjEGQlCVGxrUhzpMldty5EUawB7pGb4hV6h
Hl75mLW7Z4L8YM6+uTQg6XWz/q6v8R4Px4B/61XalkHDdf8nhGKXiaD53RiUfKJaVCq5IOX6TEAY
1dELXXE1sly98NHVL3kfLEhKsL7VJZ+6AE/nfCH68Ou7k+ildRkOlOF7Tz7qv96By11W5OkZVVeG
oEa3/fGliFoqOjiSx5VDDs/N9W0i/2KyZOV/3lwjyk7JdGM9kj7nbPH9qg8UtKD9mOPZiZ0q7ues
MyzFdAye4dcxdWWUg5rNwMc2QwFDMLtjBGNUkBNyK42NVXlJ609wyKGhaCpKkBo7xMasDWlx8mzh
NOSL8yt6MMw6WrjErp7V4rTvSxAaK6Q9Ge7P1J9j5wXUBHoaYgo4pLSgATBClvTyG6LD/cw0YNeX
L6igyTMMYSUY6wcqJOT2sZrSsWfjL1DB7CiutD2z48wN0AZIW1ogyHkiZvR+hIm15ZohhWvUsxdi
S4v5iNO8XdCKrCs0rXclz9pUDjXW/UV9nyIOiFj8Ka+fgmFhomMt0w9HgUVsZxueDBqOGkkH7Cnm
O0GLi432id2o3IY3rlbyFYyn5aOdPGrEQv0kHnRajUSga4PP8OfkUFjY0rhKrMAsGKKe7m4EzBKM
JmoZq7wh39S7ePn1SNpnFIfQ7TbVS2wzhAsNfveCFaubctrvTkfHcH+yVoVP4oarh1v3Bgf6olnN
u698D9epmAfqOuDAxLCwDikncR7Mz0QZgvzzsAJmeLL2gSxT7/JP6AOvDt9yLWTWnGOXQ+qjzx0v
X/QQYCZCbWD3OiZJaxFusu7bdY5n/CeHm04wo3ddHPuEvQyZ2BxyTMQdDUKQE+9IeeXRAnh03swD
aBa1X607N8oXnBjOb27v2OIjq5XqzO+CdzT/gQoMejaeoRKv4eVBtrvaJoFNstn+Hgfawcvn/N97
SbwGAZQ8vBJiIGFEBJplUg7SVPCglYLBxge63aiM8K87EknIU6BfxdOyWS3OGYfszs/o5w0jNSPy
IayoqMSDJVSmOcTW69BzVwbmmnqHv8j2R5cNfdWA0i3HpaXVvyRhV3vWWSosSL0I31utFsjvNfN5
+rsWvkDjRcxsApHvtVSlElSimgNvwpTF24zoDrx4SJPo43TViVd84Frf7RPUc/UBbM/KyqD1lbhQ
4X0kh5RsV6qUvqxPm93iVywfAjshX0QOpyNciZbhs1jWrYfp1AYu0B7qxtJZ/z6i6Oj+r/IJxxj6
ywG2bfuYvPaIslRBPRJehjo9fmlY9q2XrKi6VLQ+1sn9fe1f9uUJvTUDy4yF2tXpaxxXtyjI6r58
5YffRxe6NrFVNJ1F0GfBC45aZMHYSAuk/H574RZS/ALUqPUY7edg5GJtZ7gdbUHoH5i/FM8/0mVB
isNNxM2GWkkxJg5uaHVqXrhGfeUG/lXFw0C2aTWDtE91Ia69dXn0Hg3sJM+7Lngkmqq03cE+RavN
5ZbFp6fr9WqD4rvYoH1gN1mwbAgJvXcWmgJ9sqwcTfeknUqnIMPfIjIj1thvqmRVlY72ZkQGqpKi
OktG+qz5iowrJeXGdiPL6rKiWoFBlvoZ4E5uC9dxvV984aM2pwjLWLmjGDGzuoAC5mVmKhbHoG/d
rgX6jDqAkNl1ZnGsYi83BicsYHA8vqg2DvHLhDK8FRyLoHVnFbPHcUiVHiWmULRk70fUiCNX5/Oo
NLu7I95hZjC7mDVJK1TnP4VgCzJalKUcL3xUtE85ZypRg3/eyl3MuhswdzlPMQVoBD6ROJ3zWycW
GBLjlrZ7gduc3VoqRE1SLhYKxUOb+4AZmnMLe4ZsTVX+VZPo19Wk7ppjVYCbgx0xZOKimVYPAoOP
KVlcjB2jHZXRGPY/VscJWH6a+ngVX+s/5j7x7RlqRb4q2FiRAG8tbk6tYCJdoEfNZUy8suLPD3Xd
5BlZFTPpIy0moc36TkHXCnkjRvqtKf7wYTE+73/Brdc+/pK8sXgKbo7OvRKjDLCTq75CGzb9QdiV
BTW8NbGWRQbDkpB+CP54mjbXJC3YOWRhrTsPVDOIYnjQbSim9Op96Lbj8Gp0h7rCSWgCgDivq7A+
FYJiOH4Pv+N7Wxma/f9n2bJ7broITs0I4kgoUUxn7VHb9hwH6Bl5pUC8+hENg0ODbzJvd3+dEZ8t
86/6ZNib5tY81Jmt9P4blmv/ek7u2skzEwIW3dpAZGTv0PHyIldpPZtjgJJSbyNY1yNBtFrsQHOa
VKthJpKaZyY8qQHXEROrSTdIOY1GTVwD7tTGhiUb4FMPgvDwd+6Gv8EpLn45AzxqyZ5G4BV4peQg
p1ChHBmgmxlsyX0uEbZvaIuX0HLisF55R9aRnU0mZDQZ+3keuo9JC1bcSdzyekHBvno0PynRYIp7
9j/smOXRXgTIujORGHb3OnByd/wuuP7aN6QxQlbCxZKs4y7CCC5gDmhZTUqdaMCBv64TtilE6ODd
Fte5p1sF/Pc6PtxMODDkgz3+uHDL3l2VNOrH8wazJ0dbWd/jMgnYjE3qpoUFJgVx5Iz7BOGiwvAN
eT11fhZ2yBb9/gpFuWaIhJ0SS0WdID6ieugnnEyKi+RA0ICIg7thXOHjWYkKksli3+PJNEXvrKAo
fIM+cqU+EdmfLb1lNw4q6XcGredPFZhZasVz6yHuDTK3P57dxqtBnDpRm4ieFbx3HthagKS5YtlT
Owt6UPqPwL/nptXLUhecFyZqgGhAkBnstQNuugqGPw7LfTCwuA+1CNwK7OV35btWzT3lwvo5axZf
X2+57DhMWS3FnIPRceFXuAg/T7z4zctr60GmxfvzYXm716LsDur6VwKQ9GSHELNQwAW0gIz6YgCP
n82FU3lCGLxwidG1l3vBN7J/EupfUoT/uJpTd9bpMeAoqr+EiHubs70lc8+70PnYYFr2fQrdfkeG
wHAK8S3tQZa/YxFRGLa8VjcSY5okUIhoNrwtzZZxFgyK1ohSQRSf8EgIuGoia5MoE1UJVAkQRg7J
MwVPRrYjz48/Cq19tewARKzZqMarXIp/wgG4GuzqL11UttRBR/wjVWxgfJn/45oDILn8U1xLf7CR
ogeqe7al2gSfTa9TeVSMucja7H0gopNhofAjI0at0//vI6Wz5mHVQ1ek/tx3q7CWX4FSeY6niV3Q
3Fzj08RFHZ1PFHhRk7Vj6J5zMQPy4P0eldLq2dV02v4+8EBewaGYHzRnkKO6+jJGAarxf7lN0mQC
5QD5+JSdvCkzC4GjYLt5R138WDX7VH/XrKlu6L4ZqF/3yT4hQ5rM5oq6wTn7133MsAco/GqgQD1y
uy7HW5mAqZ1N1xtum0Mt8b3ZHznUPXP1FBUYjq3QOBeyk/8qWcPpX9vS3XSOe6YUYx85Jnv12m+j
blJ56+LdPKV+CwJZRMlI2kAATI1YosUob0wWpD4MSkOfx42sGTkRYShJ6coHsXQrclJNA7MBOm3l
vSK2JMehOyNVWULaGVxR5aHsYiR5gvPA/Q/ELCXdbqQ7hBT5bHdhkP3SIFoE4lYfHJuAr4aNrYpM
PCGMFGn8WfKsU2TMhZ3MLro60CmaQ5oRfzo182DTtW7xdGjwWD+WzoV6H22TbCAT8v5e+zTOXBzh
+UgjKyuvJFKy7JiLmesC+ViomGs01TL1Sdq4nViE/Hvth8XZqBReymbBo4IIYZOJ8SL6vyxBj8Rx
FgcQyTYvU7wLcE3IeB7PapWB2I/xMByCw8P5J5UiadDt9qYzDwRhzpY2AIUn0mFbqjiLFRHlPHIe
Y0lyRZEy7H4U+/QlHPe14/kFtCYcJ/RiyQEmLIEKDaXihVdVjEPV7Gf3ku/V93q+FWWqidQlyUSv
bCaAQe2e1xMlIyZWxVitKyEIHo8lRAMJExwKfF19UKfU9dDvdQiMR7MZwEjnXG4rZx/vkqp/vAsf
kht8+XUHT5fuC4uAMdtPFpQ99MEzBw2dYBuQ4OtQzIVGK/RQNKi7SHD/mTJyPJOZHx9T2RJaGONO
ErdmDeFs2GjgwdcfcCC21MRj2HU0HnBcm8di6R8HFztXOxsYOz7/IWgVXvMdZyFFlMnDCS/B6ocW
j5tj2hnXx5QJg+g2PC3dgIf9+Kpf8Yb+OCiRTtCJUVJQrWeHCO1H4H+W9bn1YG5f0iqUo2KDGN0/
uJVK1q7jcm8k0meCrIXN8G9qoHFgLyGDYxoxaYa2KJAC+nnMeDkGZMA5MOZdTo4NGMD+dtozfo5/
yx2qmAvvGzZ3dvovtLBKOSy+9GA07LWr/h2thE/vbR7sjnv5oJ7BW1xEmPiddfHeZ5cn3Q3wtPkY
TDAx5DELoQdOuUOcMbFSXh6H4VWp+P++TjIkWcQeul4qAvxqPn3LwjxVQ6Uo0J/DiHeuS72YRjAY
FiGWsmvdXjHx1fgNwbOcYAHGUbV94DSprzCr3jzn1soXPwxVx/ouzET5K5waiW7SeNbffCFjAUt2
QHhdtGqsyxXGtK5uag9sxarQKAV8Vwk9GqzqsEyhJKn0WRKBNOzbq+BHPUyiurZvjEwCaPv6w6sS
4r6gIWiuFPc4wamdsM07FdCf+r17tiZMAFEwWGAzcgetQcLz0PcqYVikrx9NcRKQUgr6AaoZzY1l
FhsK/YkbenPbImmOtzhXUMH4OwprSmFNEPAxqteoVgTQZ9ZIY4Am45br9Pd8MZx904JYPEwyKePv
eTiOyoSbgvL+D/kyPWoYniO6Ut+jfiLTkjiu5puST3pe0hkvCbdGI6rguLOLH3QzyT9N92EIqCOl
F/iOX0rNKVz6Z9uEP8twYmPPMrTfbOWjFCLzsEvQ/1nPE3SfI12LbbNwI6wCCdRkix1Vr+AGVHmD
4UFo1qze42o1I70S/dFqxvvGOxsR1/XWuVwKncoxGv3D9OAn+WXzKzw4UhLvXRnCVE5J/jHD8fhg
6ijYqubeJeDwDBUq3jo/LOqp42ch1laysokKu9SVH6M1VSO0+nR0eQ0c9farEn9skOZm+Zd84/mL
QeyncKBUoO1tz19xi16f/q8hsDuEJOsuND5F4urEjCVh+mG0XT4w7DyGfLLvXmfeZzMKZm7JONtk
zOBhIW1v8NBv62wDEGGonPn4dpx/3RGSyB1m8rBNUlJD9inzoQ1mf1Y8mLkdSwpMLG7yizykHmNp
4fr0bq04IHqYFz0JXlgZ/4qDYw3gnnakFF0szmyhwmwyumxxG86V8iSk9wCei19pnQ9iIQ4w+SI7
SRWJJjFxMX6q14qjBVsZF9DE/gF94JG9p8v8QTFEewOdLgERBjcRgk4JHVHSV2uBXhdf6wJp5fAK
DdMPOP1x1BDUO3W7xvrXbLtd3HQ6S6rgGIZ2CHPe+C2m7PT9KPOWetSHdo//syEiQV1RtO7ZWv+a
w+RvQXb4tN6/PHUg1RvmoZYW+tqG8vwb5OEQj/xnLkJDhTmz9yo9YhPbb8Q4pPYu+XTCfLeSlvOI
lYDOd1OAU6gte1dmgVOi9VnNTP4M5el+WnMbmIcnTwQYPevYcEfnd59x2Pgk7nw0UMdsR7prKXf1
2kG5LFGASX2J/xzMfDMV/nnwIY73WOwPN6lyusKX0KLzxeldpnAtUbuc0LPKy1fGfB6uHbJdhkxO
G7yHM2tHbOrQCziiL+m2TCU4GdHhed9d8YmHPiV/sKQeOyGaxadUB1Rs3HksGCJgAA6gSzT2N6+R
FbQK1ZbRqOLAYa7KpkMSNWuBmQ80dATITAXLWUhlQIvzDqnaLCtoRZBVz1STkYWke3sOhig9SnmV
UD7C7737eOk6bUZVMxm7fA+MD0bcKS2xQvyoIhJ6af+BH8+hDWzLwfBa2Ri9FKnfGsVbP/avC6O4
2thgIyzkXjROA19j88jq8oS4uDkkryQUqNK7JV4unhMVBOu/mNYbqzFxqLFlS4Fx0Xbib1qvtnU6
wzYI9Vi5sNKwPEe3Mlq/QIHkIvfssM6iRqg4xm205p0si30Oi7OBRCHndQR+NcviyA1q7GxgWTiK
GChdxamL1W1O1RuFGDlTYh823G/4DkTnNIc+kwAhnO2FglxFdcUWNy5C/nUPtsDmiS1XbbwD1rmT
FcDxBcpFC7lJkKKLxucPLFuML9Og6G7rnV0gn72fmhdM52Uc6BJrV6tRSJLCRBTsXamx1Z0tLcf5
9ETGFiKhxbcrqFJ99mUIw6lAVozCKexJGavr50BhaFozS0da86VZzH4NEnTyYuUwNVIBSvEEZwJc
pKZLY3S4BHDGCdy9V7EgeF5whAo+ODmCIKI0Y74nnePnGEZCmM9iUWBKIdORdllBhL1sOCLkx8S9
zTJHyAFIEhCHPrg6G1vL4Xvzc2svytjPzy+7SXm7+LUvXe+7tjZHaXcOMbae8eO7GMrBRDDDy9mo
fmFQyZST+DK2Eb9k6DBLBZGLy7SYOCgWEktX1khZl0voPduGd0SKjZhGXWe7Ti6rt3reclOrKynq
bypvOOMOsYjgm3W+T94nlGAXB9DkMfWTGzM6UEiZ+MdFTzozYV/+Ek1Mk45IGQgxHqacFhf8TVDr
61QOdbF/GFkzL5uxkBQrECWOCfhwOygFIYQ8OF4Urpbu89cSNloqFwwlZ5huQh2ObqXJ97N1gDyJ
B7EtkrjhVwy6pcs0R/X9dgCYznr9NuchrvdWv25/OYZVnqdmyTUOQx0wmVqD93s1OsDSojrbWTT1
y02WH7KYvtnyrU/OleMYe8dXagHt9JzDCTkKAFYxloYsqpk8DDcnF4PhqShEO26zn3Y9sv/9vj8F
BN/0RHvfQtfmR9aSnCj5Z7BeU5gLVo9H9/350YTEwLjve9PgJCSA27MI5ohXzoFZbpoAHvOVAWNV
8CjCi4bCoHIj4gS6fcsDZIvu5mIhx8uuT9v2Z/zHvxqsc3F8B+cnMZ+wG83vJcY/rzA9ZLSobVYb
yx0F5OrUYczmOLCd6/HJPUmW/8JMrk3tXRodOg0ssJYPTcN9o49AVO+1xUnFhY938AskN/2E4IzT
gCCThmBaXqjiBeAr6PqPEYazYHR/F5zoiFVnxXDPfy4tonVyZXvt0+R7u/7jQ3cRkC1KYVr0k6Do
XSveYKc7D3ASoRZFMjcZaKkuMeGRup52ykO99tuXi8uABtUEqnKbW/ai2DYSQLxVK2W5zL7B1EpG
ZtfwkpRSTpX0DSSkeBzL4cLhTQup720HpTeyHc4AygKr1a84S1wzQ3gyTD6YI2NOS6koJsfP/uYB
+W0rQiZJCfR1BO2fTMtEUFsLomA6DKV+0uLsiRTKi7IKNxVdwPNo4BN+P+/r+EZ0jU1vokHdla7o
mym3GXm5ApxE99r7NyHLuhJoBFBMRRTBeyqd9d69YksUgp0x1A7n9p1mVP7pH1m0BBaUxzWC7kWa
Oi6E7FHmw1/YRulKRnwGHR77WuhUA1IK0zGMQtJmDAjeo/TavZaFCji9+PeFYsDatVyt5vy7sI3V
9N1UvV5LKjawerFQ8iy1opQDJ4qsNGTf5xy85H2NfJPK65PWVqm4IhgGF9p5sMi6ThSMHEb2wXMT
TPYy0g9uDGpGWC8OwhGvsVY6CaD5L9aeoOZoYKnUdV8VIfK6NwSb5l68vRR1Z25bBOEJhRhDlkew
C4gQkpJuDa8HvSa9xAHEC3DesJi42f75PtA8P5NifiROdMSxHxodqiyvCza/6QgKgZZ00kPcxTlf
yGT64gh7OU7RYtiGp2Y3488G7KaKnSlBlr5s+XpNE1tv1YsPBf8w+Sd1H0cKLaEABMQd2XUBKCPb
MeE3IOHvKV9IlsraMTpc/rChDoJHcrnMDITTRkZ+USHIfD4CrazLdtqmXIR4Xa3NSbNWX6MykVan
8QepqMugiBJTuiPkiKnL2wsC9HfkW/KYEXosjj5dO4vfWZN/sbtmymGCqPYO7nMlam2L8b8ducGD
mpqDeiAz4GcWaMjahRgvH5TJF9y7/SFI2iyRDbtJm0ErDdIOsZ2N9G6J/+QY6cxqVtblVZDOxWSr
t1egGkFc9kTMwxRpzBLD6nOrDfzTMJhd+AM7aBH9fTFW8COqfsjoZL31Qs99+UfU+ZwCgMcpZEzu
by74BlrkHSPBB7ar4pvjbzXoszNpbO3QtaqgfBrVFGmTi1qLYf+V3uHQMbkzf3q76BWsObhdiHmP
3Ooe541jmUgvRURtIYO+O3u+kAmvpkDdZVK8D1pr6J9ekH1YwInrgr9FmGnmlZ8qCkBhFp6ngwIn
KXHUfReOgB9CtRDKJIooE1g8nKF3NB9dH2KZdbBlihbum5NAWGPawPPeL5GFDFkzfuU/5J3HdNn1
B20DmJSbqO1S35TS8HWh8IAyZ/w5/DI9jpYDxyi7hM3J3Wjm2XiRmb72pVNohEF1t6zdfcExeO2a
7W/ZenGcCm/NdEvaS0A8y6vMzzXhkQmPuFUGFXG/IxYNz0hnPXgalstG+acQ1lLNnVDkrDZnWd7A
mnpBHgnBN0gWFKfErYlMmvG44bhwMloBtu4oG+kJdUJfI2tRx6cjGDu3FsyWXNS5QjwTHdgyM61V
iHiyGd635vOC1ugZdKmGgL7/KLWP2R6hNn9lVuWr/2BLWAg4MBsTjqz5RLhpL5V5/eK6daQ5Loxo
ttETUKmAitvJqoH3khWCZd/8FBexEbdV6VKMFWB4F4wFNTmAbl2IVfdYl9A/Q/e6H//QQ4sS/Q0/
awpaIFtYIEjyVAfVrsE23m+qmdYzTA2Y7JMLowOlpUvtUYSaUTRUkrx/eYVr4UzueYOB2yWePOO7
I7QCZaytbiq03+9ISkA7QdbCsc6zDOuTBojL9QgCHOWAZ7pJb7gKag3fjE2uZy1RCig6oVUZW+JY
0k806WOoLC1l4Wo4CVOGPSGmjGo/7bzxlngWcis8WiSKDW4wL2mUIwppiTJQzWY+dMW92Q4PFDk4
tqYb7RhmYb5Cb+Dqd/ABw8AyNQgnDO8hiJxsUPf33RZ1EAn4I/svVpUyNV6YcP73kBha1VkspG5q
l2pBMlUbOK+uIMgQP3fieq5P6FV9JhSLDJ7IfXOxUrkO4Nw5m5KbbeGS9lfQjngFHViqJafL5CbZ
zrgNigHp60zpYm9+I6dPJqxa8UViW7HIFyURqq98xCClEJqlwtwxc/9O2yiQb2eczv1xCXrzggdg
SvrrPtjFbKnPdDrxCwpywKrVlPif7Foztv42gLE/5G9t3DeZfBVeed0THBUQjyWZtH3agFWGqBtk
JPUspZUp4mvKQnog6/WsPZdS5r2ZioiDWkSzTqOGoy70ALFZCqr11ynUOyiGOfoPv0fQSUVFxp/R
Uh837FCpzFH9mu3MDFsU9kl62+eEeUQMjzUeWhNVKAtgBbXns2ggU3VUthE3bCKx4Uvcrru6BVk0
nB8Twxof5Cw+U+oJD75tzL0H0tlu2MFT0cAcEaEJjezUemQ2er+oGdPu8EaeJ31pz9P/S0vzlPZL
gpiwZB/JkzSiBHRh90Pu7uBkVVGG0ai02FS1bgmzgsK+VNYLCW3yUCSQ5CL9uFBvBoIx6Mzwweo1
KuQDVxOxpiivP0wJGb9NTVdFDB1iXR4HBrjpLNq2SG1Sh+HRCGZxAvW2CfxoaKzR6WnQInkds/Qg
JDlU7nv6Z3lg4CpAPVkkNxJYWERNCrwRRjlc1b8nxJhH63LFQnBZn9cLW2XIkjUjPR4oD5meFLSM
6y1Zb6dYRv815OgmgV7XR6v5EyoVJnhKaLVEdlT3bVzd4YG2KJ4ipI0SaZLzwfRsfdsGlCsjY77V
v4j+7OmLBO9vkh77F2mD5/s0iU+2mFdK7ecVzGeqvCN4Jgtk7wVbwP+0vzqM2Hb0U1Nl1G/Nvb90
c6Ut2bE8/aaCJosOoJxhQLSQrM4krqxEmOJB7k9jy0mNvn9GA79WKCvVdHutlqVBvbpEO1Jf+Cde
gus0UWMdjkE3+7z/m4l0smLoZ3Q5eD+6tXlU0orTRAvruiRl5ax+kbo8by/fmqCA3PcRMvb6JLT2
jhl/jjxDHtPCOnNh4aSira+tORWE+TNy9PzeF8JOi7KqD5+ldszewKfm4mpCOotHP0ls/d8foSsn
rGwXMpBZFUgqukSpPPpurR8dh0GDOddWE+u5DZQP33Rs0kzLubVoWnczqAV8v2h9N5scCop9u/RR
esSI7JevvRCRkCU/MjbkMrAVUsg+yY7RJl/klVBYLPU7o7ILf/AZ/HurUbEXeOvlJjLZejTVfKC3
kphg7TUHXc5WLFITsAG+uJ+syefMHohVfF9zPZxxE6VKHGT+3nEjgdA+RgfApY6l5DIYgUgtSpK1
0GYJCPKbQBibAJC6HSmo9w3zJf6cEykwCZqkv9U66jtZmmebeD7ivHVmbIJDJIZjFbGkmrhPbOzt
VO9m2vK0KeUQruryjAYKieFgqRwe14ZprIhvNJOH69RbruLRJQFkhweLXX4rT8ZGMQgqf7a5ogt5
aROCxVG8PGALox7+hf/mUnVKNg0CeOdC9tgjr/SwlDC/7NcchmEyxHYZEUXo5rFPSDa05QDWlC66
sjw7SUpo9p/cdFHOu/FY196M8n+Z14uvNwtfNi8W62ZIbiX8V5fkRDlZ5gou3XZYXWM/gZSEdpiB
3Ulada15+OIIPkY//XUuANpsRXMbEBEAQ+eLz7O18tkLi6Fl2nnrFADgxw+OjXGYOO2dK0+l24Jh
0lRzO+BKDx4j6qsxp73QJfcmDkSZsH6sA4hC6drFp/KrcY4inra5t510ev5YBmPHcShA14HL+CZy
WsVf8/N9/g9vweg+fu5jjoFpFtozHUZYRzCWHc96IiqDO9ow6aDu2Z9dk9ZeWfNzgzR3Yxzd+ZV0
t2caSEQA6xrCORAvUgEF1MZG3qxnuiXrtpa/Jn054PtYzRkIvmJiAkDzNgbK7Niuq8Lv1AA3d7XN
hhPrTeOcxg2sAygK8meJCYLpzDWznzbpF+sa06iLxTYmiUl0WV3ovgZwjNXd7nXqIi888mIuOZXr
gS9fQPGZdmWX2HZdAsssu3tU1nFolL99Lob3qZDkr6okmd8RtNBkN0zsDlCgLpUcFfwRUA8lKAx5
/w210wG/awRNNA0Q4M6Yja2AaTs+1zgS70LXw/9Rm5ryRVklVETqBVcsZNJPRfDQaxBT4g5VDHaI
N+A1uyVxX39wP+KKJ2onmR/OkwyMHQQfelOBaTZgsT57zoA92gJP2SgcNDe71rJQzGakfcVFourz
CYOF99zLHSb5CaSC2hM5L1jhlpUBREWt+vyiEbwrGvEY0Z8WLY3TEWwaJbFyoD4sTT03J7RA2zT7
m8qGkfjjpXvGw4u1sy88sIOYumhFuZhow2hoFFg/WP175CplEYl4waFPt3X+ECf3nfEQ/Oz0Gozo
uRnkpyqa8dI9FEXYUt0O87JOgRc5m0CcheKoB+a9RjQ7OxiMchmwEaIvL1q43EKdlHjijlmPdlMM
JM2Vedpk6EZwsl0LYbbMRP2LvzJMT8hO6PUZ5Ekk5dhqEThGUWsqNF/yo+gEV55EXUIbtLKMw+iT
TpmNgQCZG5BGa4YGcMdhUSFA1xPT4uf/N/msvfYC8Y/VY4RzoLI/WB4PTAvr9yMN23cSHuQZNYuP
Nfcl74GZ//lGWcwJYTp/zuzzmWUNQyydHw4BalnhFIySaEokcJ6uND/G6jwgBgkzozgtgirAN90j
yJsHcMgzkzwPuGfdciikEJ1qWVu/iXf36vFG/6H1LeTh5StRY3FLvKUVl46gwaK0EMpF7cO8TcUK
47+BPLx99Km2R5Gl+xZaWv921CUr47UWzqpC1F8pla2BgFYMs9k69QK1ZenciJd2RVIQXjOvWz7q
PPbxvu51jmE0i5UBgL1bNojLSko7bTtCWY7Z7q2fN8KRcUXF4QI4gIXr1vqAfG4MxhkD9Khb1D9u
FoVfB4ysFbXoO+9+MRdPf1TZTca96w+0vCaOX0BvCk6UvVeam2neG7FamuAYW/qeA/gFCCpGeSh5
PIkmNwzTqdTy8FpNFqu2+oN9kB3tU9WjqsDeNsWBzvGSgOFZ+bxtQhc5TDzg1S3lmG6MAaQlO8gY
mfK0LT0Uu5DZB6lfEW/HcUkh1VjdlGr2SVe2lhZOG7bl5cKO1YaOJUk98Gi1VVQpFHBcvjYA+yhl
V+1ugVFIHJOcY9jG2oVI28C8Q2xvT/PW/eolknEwdDeFajeDS3hMu5iVArMTq4J+1azfPBHTVe/z
i+UFduzoD0vpt8N+6Xj8rckFYsmX3Pi7KRQ99mSiACcJaoxxnpzNhuqAz6w4iCJeKkaNCU04dRxh
5jD1OiR80Yc0RLYu9DBENfp8Mam+Rh6nSgDNTeJqptPbtA8LtcMb0m/b6laDe5ES8BKpwMT0989i
+LnnuV+5goHhgG47efgpvThN6eVs0dmaawHGWqFmdLDCfoWI6mrloSxCm0kDn5ZLpdN02D4iL86D
3ukCev5gsZe8A7g0haRdf4ZN0zH3N8yPRXExB5Ui2kDd/ur5UuLkWSvxsjSAdYBsMm5KejWk0KKD
fbB/qpuM9WPJ16SUoAEGlKsrdBNs9pQRD7uYUMVFHZTjNKsuAbpXP7AYI4JVcN6DuJUmnwyO/TGx
VK3Ajm0uvb9zuwrIoNP6h/LPut6xOUGkoYa/2cF4k1h4Bot3i1rofcTILwn17cdtijsk1RiA3GT2
0X3N6uXu32EZ/zPRG6KCMBM89eR6ZJ61Bcp3Vyqishj6cwd7A9vYAjE/UiCtVPkdZ6qFsOq/it9g
tHEn6Dni96E4Kv/vsBoQWatdb9wPltjPQtnvDnp7ZXYjoEsuW7yyUuwoaxq1ZY1PkeQMVxKWCnE+
35+Z0oIB2pj2cDnX+WoO6w/Nf0tn4ibyfQgW1gowVUNFUbjewK1BsRZxmrslsHJ0XpqiyjJwE2vM
DBT7CvRuOb1/luE4rQgIiH5GrKAEbaPyqMhXf+R4zUNaIAcW0hpSiOSW+GWWKDE65oSlgylVDvT6
gmxljYJcXXCQfd/8EslfuAeDHQaYdIuNOmkBvxx1pQI1Ivy3QIuUw4vKsI3/6pwazLjfFJqviQZW
d7soagYDVrdwer1x988f+LDDn84LVIfAISkLShN+U5NmB2kIrmnmTwmtIwTupEnkf/xTw6321SfZ
TsJIAGqRH0yM6mzH6l+pGG1NHxkRBlXErkQnwQnT6OqZJeyKt4XEU6QUkeunDX7S6lG3+RRflyKd
/lOZpJrfvWVFjd1WJWWZItLq2kfLTyDV/zug1a8YC2W88ZDB3vovrgfhFOhlkYfT7PuYecy+XWMI
b44kjn9zFWj5sTne+wrxaiN8L/FpWCAK8dxvRdj7g8N4D8Di2m2vNdN+58P+8KcMx+15dcvNmFPI
uH/5+QzazM1k5qb0USkbamfwoNF0kwd6nklhYqNK6RAy4ks2Vzb2A4ezue3FP7k0dmsC+Sd/wy4k
wVQ1yzeLiK017QOJrs16W0f+EabRT2/2zF4RvACIhmfg/eclky/2neauGM/l3COmWJt2GEDqVi8d
uOJvZgIF9gtARi5MRfM/kMHqXCsV1kWpvel+lblSSEa2daYCPXJEI8gCbSq4BrhbnLOFHwbnW/nc
DFPoF5c3NGYW20MPVYoytEdw2+u0ggcVqtKgyJ2H0Menx1qz0SjaI40RZhlwGpRnK7M6ChTIGAot
vph00FwfkyXvZWyse6JwLbrYykfANo7EaD81i38hqosJKKZzwI/V8kASrJjaYsqLjfzz5qrXu7jq
JtxM5/gt54YBJ5lNpkhPWLE3dHtqgO+EnUYbod2nT4caDd0ZykABA89Tlq51tVDflmem+rKMlsHV
w6bAs3pTbgh0k/bBxk2GD4uPyNyevDw6hAkGtLL3+l/tarOLWgTMttz/0Lo1LlVSgJXThyBRhKsd
Z6na8BONZNUHuemUfaRrEc+45zBQTmahviN3WYdOmC8uJlYgj1+Aqyj1CkHCe+4OjeQKP0Xp8Nmz
NC71xioKvWxxYI39fUGPAhdNV9Q9fIwJAleuikkByownQtd9SOfvt6LZ6OK2KWmu7xpSVKOPoT9J
QpztC12cbYScHiAi0xosGMqqR5hfmY0mVUfntampoB4BeMjKDG/86+ks4sG7UEUIBh+JZet1KS2X
6KE1ydG0d9lh0eZvIr+XJR32afoeCOdOFttoD50zh0/dC4JsZQL/MGmUD/UL+uLUG3mHkNuoNxfi
q1Y+zo8k9iYbAFeIDhFO0yoylf/xo1OdIKv5RRtLfKQKK2ie01q7rK2xrkUq2moT3Bh7p5+x4pH1
PPeIGuQC2T7BzyDEBrJ72VyikAhiU4qjm+pLbczAaOojSou3rlamXeolWasA5tMsDu2gCLqCXgNi
dPaE9Ll6IUiWrUhK+eqIV7j+je3l7i7jyX8VRWqZdIFGAU4Dx0skU1RHV87zyJMPMxZS8scM/Zeg
FXexYCNpuHraJbmXQkyWjJHZU2QSTvWbizaXHslGE94aoqWMqQIXOi2o7wQv1fesUV78Oy0RTUnt
ULL4S7t3K+pmMXYpXvoM2BNisMvfSUWeC81L+JnHZSYJiT83dC8MKNfh+tihFkUktup28HR2RdGJ
uN1P8YqVYQeUsmXZ0RmYzwWAzzWXtiWhILB1K2wUZC8EdgMt0gjim4Phyo4fCnSJlNdQqtTeHUDk
Rie2pm7J0yRmDEXqtAESf8XlSbkYCAu5Es6gibVicHopg/ctXrUW4IixbRrmaqhk775f2mtqgBfq
dOeJDQLuQ4oxTZ8e1u0yizTyrvo8asTKQgbE28C0E2Rpx76b4MPGvL6D71jyU2UI4qU1Z15o3eWX
sPtHF3U2PDmqIBByko5Cl+W4/y2dy/rugewu9M7IKxTJ3eTraJb2lpBrI2eLYciqP111kSaD50sd
CNEoV+GGj7F8Lj6XY91Ya+WWtVQy9HyFwX9clh+n+f9FEvpH1c1dps5O/xHP8p1x/AX/8FXslL6s
iU1Ecbd36CjvIPbcvOR+HdFjuqNZVINpxB+BGG4f0EDE9nURfVmLYP3XS7OzR692J/Q1yFRbI0tf
D3RBjvgw4n/B0LEfB6EHDs+ynSuoLns4T8bqR6AMd4WG7wifVb4bz1UB6MoxuIdOzZxWogb1WR7B
KO1jLdCc5mGfgAK9/FJcDLcIHYt6lKIn15267AwaY5fh5l01BS8VYHlhp6tDQBaVtO6h/T7usMeF
gO2IA7uNVMXT2mXK4M5Ppb6q/0W/V45pTI58wg0rBxQ3dYlMBfkfcfChDh6NOXAPRYOa1NIbII8I
co613G2ZbKFi7NaAZbLdNwC/ROJ26LyEN24QV69IMdkSRKvYK5W7Olj8k9K9NsZOPw5N2IMhJTmx
vZ9n/OkvT3jCvayW/T6O+Y0NWNVNYkx/vneHDroHjE78XkY1/GFHE7Fudj3lj3naA7A3JEx1u0r6
G2YMpwgpVYNzboq58QAlFvvM+ZFY6sh6WMSwEdNm3FIh1AeFvKnTQAyICFchFrBvY8Rz5mnhtrci
wszJjU7QZarsg7Ybs6AhkB2Lp2wCYz6w4UKuGiAMJrG2VMPOoPIznfv0YYeLgLRSRkHMOBS4/P1J
fSL6iOy88q/Qi7rR2RKAacfYq95y86eWVyOTQM8yUaoghHRs/mxRLjSqxD4mKXair1Hq03aPIiYU
EGj8iou6kzKaxzAq1TAP7GypMLXTZ74rO9aJeOhyGQbUDYNg7mq9k4jVl9OoKQE4ZKpB3BmKe/wb
7g8iwjUnd2r2/BIJqnV/2p+G311+6Vba6SaKBivfgjHXUtMD/rExoC7p7JZ4XInCNhTZgNBG5w2P
OgiDe70JDdhn1F7c6NOj4LxpU7K3ej4cLrkSHiyZ7OorWpuz+Cs5gOu9KbZmffhd2ciWadCuECj5
jMIwEKgx4UoPQauikn2UaPJzHNp39hcJ5PgCWnhNOjNGReecaEoDzfuoAZjkWMsT2UqwWVg8AabS
tx75Coh95faVTbEo5iCksfz4V0+Tsiw/8dBfdqdsHoId7l4tC+BYDaneblvH7VrrRuQJe3tzwQkl
B+xEKF33L0TNziOsl1RxQMbtG6RUn3hfYDNmTw1kO5JMlxXHNo46FMdv9VhFp7DuibMV5EY34q5S
h20QoVyMcCTL+WptxKvLqFhcqEeQVF3L1glLXs9LOMze2Yukiu+CFC3dHitQxTXHTjsV4XNtAAO5
Q+4d4glzDfeZ12fNMTubQIXYOC6yTNrZnA8+vI++utH3udV1TQ9VMB3egQLGDvAYd2gVTOrdyLwu
gcK8tn+8LpfPpHXCSS5i3KVYOkXFG3Os6eUP31Az1mnHvikMHVat4292yXYnT2zMAXdMjEXDEOQj
83GducxaXeiQKwn9TED1wlkM4iwNnAqAhxc8/hqxiQqmxdqriGN+rTju2jea74w5hH6aerqLDSWb
9ZJotkU59N0dqpui2Gl8JoQivW8G8msgGP0ZeVTudCYcTF+sQeL5ek//hAkAapNccKVp5g0323ex
3jxVuzYfNBjzslaRnYs+BsMfRaeMCrQlkjlhsOcJT1DQmquujJAICrwxlOwqVGTF4ldlnCH0TKZ5
FppN7lE8cFlZcyzLdBCipHRjKv5HN2ZF1lBgDWevaemcya1Rkqbq7ehfMUyZoJge+e/92LAk2WBX
cUGnfCKqQWHxfvcQwddRVdzlmYn2KnFSGNVeANg2+xMUMzAAQyswQwZvTdX69hKTzZ0BwChq/eh8
RZU3sB1lTB+w821GQkBB/nXfykMFS3KUrHBe7Je3c+WhFIoPL84G/6Dvss6Y5cp0rniVr4jjvr0t
IaTXqDWnwmy0VC2r6CTZMkSsXscx+hYRKpmkPwNuPbKSNtO9s/WxScc31khCu9j1kC0XAPO4DMah
2GjOInMY8QNt2v6ycqPWe45PvBQWw14R/ulvBxKE9g97pFsJZTCklO7vA9VHqIyEncZwdnIz4rKx
MVDXWqCg8QljLIhmEFyZwISfNo/WNqTT+jUHxk57Jy8d3ikbnDVRZSclDw525gz/8Rl40c2iNNtF
BemOoXFGEEgWFzA7LB5QUrhetCffJ6gPPnYPS7BUOdvk5ypg90XpedCGvlKdcD9mm5RSi6SWiEUa
u5oWj+uUTm6vbYoDftQzwS7kZ1748DPWH7oWOgdM49aQgUfG+E4bAO4D42f+gFimnxW1OeOhk9cL
9lso4Vaf4HxRPdvbEDcgcLhOj4y+s1KG37NEB/54NiC4ztHuHTfGc4emKOIhGI+li+LJTDr8v253
vzt6KdJidrWbrTmdipmC1YYpeX6S7PZ1vXmmwNZpbrBVVc8srEihg6lm+EVGm2oZwY4/wuRbEEl7
RiVJcsv5GJBT4j9vQmjjhwj2skEe1jIIOVaxPW0fzJE8Ibdoof/5p4sGGXHDvh5SBY7UuW8mGc0l
5h7Q2b7PUoVk7hQ96NISzYyLEzAtbA+NY+rAOmMCPWJQc/NLBs2lH9S7L03A/9laGlVTZOKNUe1C
U3she3tFL1GXgUiHyHBmy1Tb6NW4EhN4iNTq9lXS12PFRv8W/Uxq/7gfNVhHhIIHT3mZdpnDD+B1
Yn14Sn5MmknedQzDsEiHiq10t0qXgf70octl9r8ig1p06kojIAVwdInVtQi6wmPMsVr35oXxEQYu
jAJbsRbt/inYmSueyAu+eCLDjEIJwQdlKVrVyQU0mLhT7f8UPtUvf++HaS2DBoiBw41eyGBrBE/3
+lNkVm/y4sU8w6FO26F3VOyJX/HD/6L/HTDVtYP1/1Pg3EtwbGJozmRcFRwSpjgsfxQdp5EkZO5/
SEx/zsNvYVB1uDPE8TX1uLKSwZO6JpmTYXaFB5dT/6FwJ7U9EmgyOtlf1rqg2f6JKDb+cWovmI8z
JOW5x8iWkXoMF///nqVFmUDBRGfFEgGuwa6/fGTs2Z/P0rlucaCdaj7g0wZnqhGZw8Fpo3zChbV9
wAFWJtdlGKZRxQ6dM+w/KhHOzeMo7PgIwik0oXTLOF3+LKGOIPVOCbu6eCt2nSva/klTRxx/c3LR
uvSRAr6cyIGnjxu2QxFpxEe9vsdfvBYS15aL1aQVktJytq/uawKRKt9RudaUmc0aSEnxirqsRtg+
wENVRP+iGqtiLm07cmv1nUAtbDYH+dnmjP314maROisihp1xZ/Obpp13H3Lt/FhwBSgJoHp1mLAb
9SgWw82KGlnBOW7JE9ei0NzKkfpHQ/o/ioq7NSbr64KERWfE0zMTUDxYrA+3wfe3Q3G3RXi1WiWI
zohhAjjHMXLgZkgzyvB6CE659Qu8sQ31mDU4Xj4l2IIIkWWuBZmsyZKzVVddtLfReD1RCHA/vQvq
chClPJm1Xx1HTiR02QJXiNoRKQTVZ6wtVU+urgV2tVZogdPKnt/+aKWU4lNOr5H0k6uEWlgGSjMu
trNI3fHJeQNhxfFI/PUlnGnMkcKDGNwjYjBt2cl4v+C2Q9o61smbJzcgW1UKHcl7Grwwx6XhHF7r
G4WfOytLho8eO/kTaFr2brYxsRD/rKEfE2XXMbbhB+DgR0pN85GVQeqTVc2K4DrXBrmHZsO0e6Q7
/QUtBd5pIeFH5xc3JOyLapEInsrKQHa4gYIuFxAXVVCe2c2HNK1LWGNLaauEtSXtekyJqhbqWQZQ
7v1i5VjaX+4JO6BrSEGyCiUSPSB3tWXaXcqDw4iJLesaWIxLhs5sfR5gXyHOCqRJBVsvysTScXdP
UBGg7EARJhScBnU21xk6geOUpcDi9+lQwlduF+rV2caZl3cbadlNHNdO4cXT/JwBqDRM0Q3kEzEw
utd2GOy+ZdCrmkSUDeDn0vPzBRaxRWGm4sjKkXLZhum+HQG6M84RxpdDVMCw7fFlMOhFBfi54o5N
KNagm9q6fyfoqGmQ+rJ41+TqQVyPw8wFf7eTqnHIWoMOaMITx0o8wxzFhoaZXLW3GdyprCmB3wfr
pmE/FGTavBaMS+4V1Sh7mTsNh6HUzm99mXt06PIF5GUFicnWw3pQXayWyCrinLK2K+jxaEdSYDyk
6kmDtEKMTlQypWvEgh7o3uWA+Ms6ez8pHFIzIW2W5iItl9GDkOoQnARO1neER31brvQTs+lvDmC6
aTN1h5A8ucgHmCbtQcyhkYGlABeeSMUEsslULS4UwRb/QsRmSKodRodVRyyS37kITGLDhQODfL10
lsYar3XOEBgrUT/boXLTHw2ABMGk+1PBdde4oaPmD4fxgkkNIQ9MYZkKNUH0rc46hZW13BUHvRCt
ScCiR3AieHt7zHVyqkR67yXnNEa/ycmS20ES+Mtsb/Dx+T4ggBYBMo/bBHeZvdwNfPxtBx7VBaXX
OJD63h+dJ97VrrgjEVNkXBXKfR0P4PGTr/2OMHRgsDjA40Tu2nw7J7lGZKRh/911QE0PT1LXaIWP
Lszplp+HraTJWtTJZTqfNPBKXUt65VTJ+24BaDWlnh1gDMItjqzwTX+S0xU31gLz6yALeMIm/+Nl
iEa8//Zb5Gv2Lo8kIOUCo3X9Y7dcXmv3bsASZso3DoUHztJkghQf9Kpt2CJN+dangwRzXLyz7Uto
qwe3lSRCAlV+BuyCCl/YzV+FV1SE7EvJAa2/1dNFjxep+TIam37Bsk/WWdUKonURx+xS8NmJhjn7
Bj/N2jelkCucvCwS3o6Hv0i7AQJsFY7OACGfM0oHpdDi3P56UHxXJ2Yvvczp6uQv5eDhVw5z+TX3
Vo1xxMJnGtIT23yJdi1ZJnIqKNjnKNNNTchkCAAbwA8l+ffOU/voFzso1AqUCuOgSCBiWa0agQP2
EN10c3SfrVWFfpCTGZlLHl3bKwPtkQ9FGdw4GfT8o33zFcTcWrkJwJfemtxG47P2pQuykAWfbi2v
83qdGDvCSnWkAufK7szXObtsANIvSzDRSMvXdeBtoDsfGl+kwYQKUL1tDkkHYd6+e1d3dGt3rbr/
JQ7B1YivJRC79ttNqCIXTffZftFuqKDbq7AaVq8/M52Tv1dXmqdmgIagS9KH9NEJR/hS0VjjGUzW
KPW4ztVD7T/rJDsDAkrijP5azcwzOux/GLkDA/1nohHNuMs8YrZkoazGnFKR0GIKPqVHx7PQJH5J
7XLRVtk/tabPlUpHpeKFmNGGSFFXyu6mPtjVgtghopegnQrpvF1ixkXLfQsWoHDx3xeu06UBqm/Q
94I8EQKuK3Tglobs8FHmSIz4QJxsUoetETIrSI1xWhVFN+k23NY8B9NWSV/fRDDkDlLndhY/Hv2H
OGAbp2138i23cEiB637+2OZWzwkLSxRahVcT8KzjZxEFSaAweWAiZrGIHuj22xKbsDlnpzlufBGQ
c2DmGPsDSENRBjLVr5bU7MSpE9StlGrxi5EPN2P1c9Jo2sKRf/aMFtkaXh2wwrTcrxldxEGx1vcQ
IaC0OHlTc+P5JVfLsuSvqY6qYiJUrfTxzLoEWvrV1M8tJD0Y4D/e+pO755+L1rqbsdj2XcnMNMPX
gYGV9s+kC2YnHutgrEt5wC5vJFe+/4YSIHw+QrCRnPbQ97wEmhdIuTT3whsviSExjynfgrHfDeMc
xgnbyjVhcHOUFFjA78vnX1+To26JNfSi6HxcnCT4GQGFGP6CzH9XJVvbqrtTteWiv6jQTGFPzWoI
u1SxcWwQDqAEGUVoFAEGq5g2eHLar1ZybEWQntgcYxccrAvHls2HRPS70vHrqOyPm6CLEy1wn2a1
JJ+1+qOAjxtJbGliE6heeabiDRY/GsIX4W1DX7Qp8wCzcPnoXZpjQb/5fN7U89LeLBlCiYz6owXS
4qF7cyQz7wFPqXvNeWY3861n0FaDK8py6JnrlpodYafs/PBK6NT49Cxl1mo5K5CUrdTzeh48TSah
UWq0bbGrPJF8fFXsCiWKIdG1pUudWsGihKmKAU0WafhOsFfpL445uyCp3SL40MLnuWyMeddfwXh6
SbtmJn6F59y22BiQ7JGDqZFrYY0KNVDaNnzX3RRIlNTihpXXITP7O6x+YA3VRKn6tZK0ge/Je+R3
X526JhaYPcm+HNc1GgqbahnNnBJctKVHhzfQkbNu7xelhoV/WBHpALwNINwf7uMWYSCYz5IcEmdc
XvSREadp0vSrR1ylAKxc50bgz0Smo1a8vIlt48TmsgrjlkAKAUp72dIO5wCA+YjukzW0q+64tByK
PkdXujRO0KjgcO/Qy+uUm8clAA4qG1HMt2B8dO1RIYF0z3MDvfq4KwIdaEHhy7RV0CF2bKPOiT4H
k4gv/obv6rJgd2NSkCotHAWnXxY25lnBRHYTCN6Ke+JSy+fBXEGgOS9hvQ14gkXBEYNuGxA+jk2X
vOhA3g1/OWK7kTMTAw9C+OCkhnTUAQhsngKsv35IRO+clAnHZO+ZRMeB0hhf5JuWadDR5smID2vc
yBTHYX2KWvf06HHvhFU1NhooMl1VGN9hCkoxnXRthleoZVjr645Kcbeo36y+/+n+K8un2qSzh/qj
4VHAyXb6ZDQ8US7eMSMinOCVoYeDG0NzWfDn2R94PlXGx/USK4WiWyLAVTtRFb+N2SVt4ICFTM0C
XDfRhkumecQnmXqqtjOOBRikHz4i7sY0nS7VxWx+MuZnVXovPlba3x0Q/tuBJ8kHaVSe1nI+xpPe
pIMI4pCG1FZVRvcSLI5UfUxLmjSksu8S+xuvDVJs0pa/47Ut0/+UKE+hRU49N68j700yY/3Jk82v
AbOoKZmJVrgjIZg+p0AR4tVxybOIAiEym2RPcoY7Bb/0lVnp1rjFaRLSh1xB0UcUnwVA0VaDj2C5
7yRlKRBO4N9ZaADRaq9XgTPhU85z/r0L1pTEbMHPvXAV/3X5+XzxFLmsyTjpnz2ehYlI2SiEbMy6
aDNKn1UHCzFxoJlQZQWOKmpKuLb8v+obbS0ULUosAtmM7yn6Z9od4O7t36yPAX3gRTPL3VLYjGJ7
zZ4rO4atV3QJWVhdWAFP9LD5JZ0jy6N5CSAorxMv4XSUSk4D2+FDOVm5/fchdmgbh7xC6d7yeuji
cAqaQE3LTrzcC/MrI6subdgGdBFBi3ZowAtnCYFsht3YwY8dEBFgLGpxcrC47oM0FuuyRwET5Oy3
VGRLF6N5+Az2tjSrL5pY+0KIUp/muArl1uH5959odAjmqwgL+RuWXVWLWXCSFOYwAurGLRVTnV08
0ergwDO43R7NiIDMPDOBDPwz7Rike2mDYCT3zS1SO+eoRNmLE4zHJ6zrVcl4viC3r5QjQ3YNNQNF
KnXVhefGvtbJjM63NAcS3izC72VabO1s+ucW4V3fidNI9C8UMg1dd/YgB6fj8E0r51OZTeePIUTY
c11NDRuxwznb1EbIxSvCJi4+s2HO6yz5Us/M8EqFLB0k7GBc77XP5dXjhMXwATUE9D3zomAlqL23
RDnX22cAwAGQ62rN8VvmOPP85La0wU14/JggW/fM9WiIJVFIQ+Jp7Og/WUEOepAnQ15g89t3ScrF
EVQCSyLPk/XYk5tucQqUz3pHSh60JeNgdiDMg07B0XqdXpNEQFm0MB/+Iq3xAUj1dOxgTjtmTuV2
RbnXXDD55PfuxRQrrZ96wq7u3dpKy7fbFvHpq9+Dc02SkX8Z/D29DmdjnCMegyuAbKL8ph19WBkh
oPQGhIvdI/6SDq0VqoJ0fgP36gGg3Gu1k4YRWaRj0h76B6vG4UGd6cBeaZ42ksr54kZzJjE1NXfN
C3Rrx83zUzje0jLNF0IJTWcwSv6F/tqVZqBihU4LWmUhyuESRY5awamzQWdEYM69UC09pdeWN9UG
ylPhwv0MdbJ8OcBWd6vtb4v+gsJTp+3BIOjc7pE9zuQ1uoQS15u/+2Q132oqk37jBxolOcXquNRC
raqvEnaoyI2bZnebZbBMQC1/FlaF7rnCLHxyceCFCgNJh1BZ7MGZpwfP10gj5RYzkhvBKC1zkO3U
MFaJ4VQtijAb3WeXf91tXXYl/xKOM2GLKC9iqOHJF0+411xfd3X4GG8XcF7uVr0+WFHpB8+nVcZp
T43a8LWnxu4qXoxWvUo3odLwN1mmSPVCLfZnXGviyENqWnNb8OiPk3yn0/BdkjiRD8jpYO8wczwc
PtXlqyx6cBk5Sv2H6CeD0sggw9lf1lIuMTLGd9xr5wejc+zdOU+A82Hajpt/JNlUVU77VxevH54i
zv7N3wXi6HFCeK/6rXRvOwQhpJ6NRf0VavW7KuGtqJH6qoi+7WouXbQxFM2xVq2dwq/Gb0nmSTfK
zbex+ZK0nYRLi2tu30TsjsMHCj0MzOz5SCMaCMbwsklQBXON9EpPTCgcT86jYgjfbu9iM1RHFJ4d
D30CljQVtfahg6PNK3TlvuI5TsozunxhOJ5PajIfGnPQWox7AxEevIT4wlxidC5OFpk94aNSbVGb
czyVI/fXv9hEm28MHfeKaVxiwGmtXcxv6yjacJk0w4p74ENWUScul2FN86Etepaf46DqcT5M9rpq
FTH5tJrzDisws96QLUurnTwksensDBaB439YCI154SgdYnwjlp85bE7rIRD0CNu0v3EXtWVff1KU
yUsK1ni321MXA86Jr+eKqVvE3R9mf540ncrmHWCvbrgbgaozPi4kesOSPwcE/jbTy+ZtbzQ3xTsD
600mNc6CzwG5WpERK7DCjp2/Ji5BriiO3p0xDWD+MglF11bD50qHWP1fWqmxfXtGfZZl/UL8Q5Xu
TPCz7GSdjAOX30v06LvvNRz/YO5qMlhmZB2JI/wdJbDx+LSj7ivhbnB2o9H77LGHwxBMjzKKRp2k
03ypY8vPMA3H/mGjYwo+u/DoVaDlamj5+4rNHWd0OpwAhDZBWXi76oOWIEoiEnuwFmJsVbJsoYec
wtWnPEhAXcp+354tv1InpTiBQDjGJZn1BzzX8g/XrNerkcJpXLny087CxAJmFe4OeLUD/fSyXoKK
uYqkcw2cKqFHIFxgMHx02lnWFVWUl+BiiLNFOTk5vAh8Rf5PB2yNLU1wzJp+/O7C7/dcsEAAcYFi
n3e+MEteg6yPJy+jXZZ8/CW6fqPFJNCXjxUwZdALdF7DuFqg40gR1uel1ExCknGJAx7dHr4Lu0Ev
KYhyYVSzOC8yrDa5OWVeMPcgq1vUwgF139QHlpEbDI5ucL1QElzFy2mxtu2Ea271NtRhF7zFp4mF
O5kxUF1hNSkAFwymZKLiAjSdedq7sgwFwI2bhooJX/J3H8/R2B8WHIYqCCprvxQTPcKmwaxMCZEn
RlBEe4jZsUpANfyFU23DuU8Zw7V5WMA6h2UL9u1FO3hjoELLzEbEU4Tjl/f4/OpDpv1ZcD3uqSk7
kXoIBf40xqicf6SjPPBX+GGn5xJHjUESS7Gf0K3k5hVTlsPoB3Pica+fzcixlPVWwFcRkaKebTs0
U+dKVhCLGZZjq4OAaHNqlrr7UHGvLZQLD7x+Sex/0r8TcEuNTF5buDRymsqufhljzM1c/RtALsEI
WT8mIg0xW0haC3IsBLrteZ7CRUbjk2UmAx10Le/cVG7Qk2882jxICrzmLSJ+hmqnZyWXVY3wTZKk
OqoIKq0rx0fmdktWUpKDDBMzv2cQ7xVMKvn63liJ8uh8Tn8OxODqS85FGCjWcItSlKke3ZFlmtSu
TzZTybZVg3SXufQQZ/qiIQoC7lC2atrTpr7PREMTvgZO+t3sS3uVrdcK4rjAPT/237JQ/ipnNhZv
pxpfPTPplYLIa1peAP75IueWjVpFMW57lPN7TTycAkLwsOF1PkwbOuSQ/WLcUEU/oN/X5hbN/TMu
1GFZ0wMwd4NltKqZXvIJtAEAgQG9AnvTr2LgzL5yemFyc/K3wxO00jVpML0o5THQ21KIlVyBfRfO
U2prc0c7lZd+/wWHOdLgeT3iZLo2uUIthiO05cLzEKcU4Zno/0rRcaARNDBxmedUZjf0N2iQ8V/E
lYTb6pNxQoGyB0+4AK/vvJ5tCAdNRwY552717uGGXg9OyFI8qR6h7hI751E1tWDhFDUAoutlBVKT
0NPiX9mu2f3k2uG0jdsvNP6fU7ZBtJMZ5gR+C1O8R05UfOUezhTBgsWDVGJ4qxQOzy8Kltx6mEue
dG21ir/MoIhRhLBcVQsFd8h9UG32nORQP0B97cuGG8otB/X+Br9LE7/jcWnemEzVHE+jTScL+3NY
SZgBBCOA52Q6ENMPWleDrkd0Tx8c2hMoB29WGkZ29rj3nH9TZZHKM01d9dUS75BWL16M6IPcD27J
SrRfv5RMTWgTSWS8XqqCYB+FHYQB3eM1/N1FQNNwq65Ek18R6cmxcQBLA527vDd9wr98XfC1dfgd
KZCcHGE2/p1wRmRaTPJQH+/mbJUew4lS4iXUz2DX2xNzQRPv+f/J0IvIohr/EFoCDKPRU5OrdCSf
OFdU70wZjW52Odzv6q8JXFp1si2pvw5hRE0T1J8q5QJ4JHB423tRZK/C7QXeowSptpmf2av5VWr7
ucMsDC0cirhc02g/iJemPwraShS0ipi5dxSd5PDcu1QlTjuvVUTcCoikN4ADgC8vTXj+nHpqltyW
sbw6JZwCiMKTeWzInRFY9BKlCLHovaO8j8QHrDHAvwDstb4ndNaRLoq+C/L/8V8mpfITEWWhHVN2
3yWYY9E7izz7BLT07lOPDwydE039ONiTRnUq9HHqEohwWQu7oZsprhhRt4Nsy0apXXkOBCw5g2UE
/hopsYCASlIRJRIo0njrqBXlB7jH02JwOa0tIdaOnWH8+9LWlYJKvVSLbJY8EYg/MzJL22RwB0aw
vGyVG4MrhVrr/JWuBQT1oTTZz3ZCFKr6QIE0BgH1YeNur+ej0+Ypxs8UTdD7csQBmwZKUVdbwagb
C78+gsfUzzvsE88C7W9LdVZNo/w6SwQ4h7qVbUTmlKVcTmUY0kuCX/6EWbOp5opK3vOZhKK3j3m0
o0qUvNV2nNVUWbXxwOruOMXlpR6fufS6sZgvUt7ggzAOsRmfMWwpfP28bCf2Aja2/wGuO5QVfCLf
ZG3ZDXw2ur8ALy3MqA4NCOV5vITZHvzwspKCcHdz32TVEily170/F72vxH/x/7+CNJN/GJcHGM4w
5QCNkdiVzzJxlZHWRJwT9BNFPkdJwwVYMtYog7Vy/7SjPwfv9dhYEBGuuIvhddia89onN+hss/kn
EEV9nzYSosJC31dHJWxV0s9Fs9lY+IGBsr4cNXIKHL+ciPTUvjY3Uypz5POo0mpl+qWwSVO2SjjS
QJEUUMTYMB6z7n1Q785PPqbCSLMvHUgCbphyVvFLKxDgjeQT1FL3OY2S9vUlWUuVifvahPMb5JDO
aZaSa9JPtSqGGs7/ORjg7soWDZDGW/SDaDAiYfvCrzhxGPjB8GLrNSxnLJofz/JPJAyEGxWCfciq
PzRr7fP37HqGJ5IvNQvF3CqRgvNM9Ik70QxjTcfsedQZPFXMVjtiEmvwyJSL1zzNvhr8O0xD+vai
JtxYCW+OZCme3Ql77q/gcSyF4jQdFTDWsjJKxB4smYTfB2q2FQ5qf48HR24sg28YaK+/VTU73qqH
BuSmjhISuyKniLI1lTsUZgwju9numArNGdHyoxLjyv6jdytZZHel2WbAIFCbljOdjjy5160EnuAh
J/VBs4sWWOlmJZnaps/KIECmi96Hm0KG6w5BTzuHGJ6JBgpf+5Ae2HOLeW4zNya1rzJFVuKq/A4o
Sxb0rff5UF11E+2u70HFU+Eb7ysGONksHt2Owy0zkrPgaa2bLhPYZ2Aj3t/IEe/09E1/6Undps0i
huHmmybfkVaYs1cdSNzonsgDFEACNF0PCJXD2x71owxEyZ/RZAc/x8yT1kyFubCHW8nNCMARYJHL
Nsad4fAnajbzMomANXNxDRKjEA2sV45KIFr/pf9uzKfrlYjF8wiEUer014okavkXfGpf3YMLb076
b/dqUFmdCQT0dY+nPuxtxe1FM/noRMU9e48Vnet37ZslhUQCAFvzMVdx3CVU7NVi8+mk2pa7EXyr
pPninlJuL05LMA7iqLnT05tDM/9mz3o3UwfU3qesgdrfP7YD18R4B5BH71hnXUIeJKEn8FK/bETa
LKt0nGdxctxZnyrIdGyHBn01+j0enHDa7sF6inJJfzZSJEQuH/8VSDocRb05Z0Jk5ZqM4j4CwsNg
2EyoIPedJV3W4aT6BL9F1SfZiDLIN8P7b+6LoHEYnSl/7dOFFxISagZb0MRgQ7JGZGOqxt+3MtEg
BlMw2tEm+fCSPAAYQbmvNZw1lsqfGRfJUEbqmnPwj++5XODiVTQYLdzgjdpo8rak3FRJG1bcuvZd
htd8DXcoivBL0Aq0G/M4IeT1Vw//0tBtAnjF3WLsllO8YM5FXCWtxwBK/n+Qo7D/ba8Np6+KyF/H
dNEVmujJFKpbvDwhvB7xCKz0KMG+hBFquMghaJVrKOPWa5uPRoxTQrkjsGs5STUqJp4pA8Awt6aA
tZA+O891k6LLgfDQx1uMrZ5VHFwzki513X6M8LNr2LgxJJypBPyV+M5avzuCt0G25pLQMmPgbhiE
plPWT18H0bwiuN9cUHasMUjb6v3Ng0D7MxfESqzxzC1M1tE6wAatbkRjIeM1ro91mseBt69VBe5p
53f5VnNteb5tvj5a9GZBDfckp2ZA8Mk5dkfdBZExO1g+Mx1lXLJIWE48wne2ZJc73cBC3xSW6zK8
zLuBJdm3t9jwps0DTkmGqwpsXrD3DxtdyT/cYnRpCGKVlsw7W953jizNH5cxQoQm5R7lKFRpp5VY
UX9DgjDkEP1I8bJ1hl1HY64yoL+v6E9DYAyFMvlYD7qCewjj2z+8QOhGcn+xYYUEF00Hl2twIOXv
3kTxf2nbzWkrh+iSB2fyyj/yx4NBTii1Oj7Xs16q+2dIo4zveus2wPC24+cKnCAhp7r+sxmvenmr
mBQcXllPvf7lSCLFQ4Eok13DasVh/hOc87M1REEjyrvtZA8C9TkrfFsoii9cH9bYTezWuwlbr/DN
scf4rXqppryDmGTcSNUGmPgakoF4LI1yas19k+dgNRs7g3oR+e4JHrghv0xLR1Q8X+N90r0RnoFH
sMJiNLKjLH1wstkTQtaIpU/eG2duiqdXHd0ie7T8Xp/SBmH5GvNNA8gFm+3Nk+Ctwq1ZgeG2Y1RU
jFFKRF1dlMi5uGATMmionFJHpdTOWgfdKftBaIr+XYAMNsEW2H3ffLSrBHONkSQpGA8SNC54yDp1
59WOY1bcbhhso9Z4V9b5sZDnldO1DcQq6R+33cMCsBiGy4KKxok8/ezJau61oKctxg9rTGh+2519
2DxiFVLFYf79Tqa4jV/n2xNnmajTQhwiaJLpeM+2PBaREeya98U9eN8ziwGqDcAiqiGxfAz42Mb6
lV7sIw4kkFcpooiR0evMwMuUrvZfgReCVgTdMsmV3mG1QuFQk3RUj9ZG+pvW02FcCIGbd3MpENRE
Vx5gxdieqvgD12vobKSzmnXh0VCgk22qvkXjC+7WM8mBu1wd2Vqf4uc7sIhHIjLnYrBogC/PTBkH
5w05akZgYvNVVT2ARVXVu0rg774QFACFSO2HWvKPM3HUmxDQtU37Ki58k4YnZ3CRZ73db/46MRlP
rikoid5uKvGy54aZzrAR85HPvUBCVg8HuiHFBS9T05Ra87Nb2y/vqAZnfI9wtT+EVb8WeMbqM4Ve
Zg+LDYEOlBArykWJws/JDrpeUGWTjcbfwveCiHcix2e7rSWAbrcJAVYogaRvgCIhX1V9l1wDCOUw
F/soe71B8F2oG5zrIpzMsSIiAaQvlionNpg2DEFSQuVWqqB9y5jWXNnipoCaDnF3ecko8zD+muM/
Z8OHUNXEtUsZJOzdD48gV2X6IvPckg8NhiOc/SGZdrNcZFZP3vAjkWH3hgpGcbE9sS/PZZRb8MZp
VMJFJifX+iscyvSwikS9nbjFrqS+HYjayP9MYwpKFy+oPmWM5/ie56RGlip4u6JqxW3d2dwgLQnQ
owCelSxb6+ByqeU8PuNRElJ/uAASM1+cAZsT9jBlAJwPJZ+5x/AfVBi0dM8h4axiOU4rteKaH2a/
I+PDD3mh6x2RKKn/xPb1lZhIBn/d/qjEEItF+Z9AVx6tcy7WwfXnpTuMxqEZ91S4vS5/0ZZI+8yT
Nz992b3UiT0FKD92YlTsMgwzfh6lFrTDquGNIiGmfLwGjs60t8VdFb6j7R8HmbrlhhMpEiF6uk+S
JuB+y2yQxPiv+3XY6aJx+bFwQV762s5CRs/6RQZA2cDFeEb2Y4Qkvc4XsmH/FcP/0GCQj3WdTIYX
s4Z6CoA9aZBhaLvBK6QK5PNZ5F8bybE1ZqJVstDmQvdaHVdaxCdbe/QMSzeCEWOBt2e09nQnigFG
oCSB426/DA5KyN2Xw/CAUP3cuOdr1cvsmK0pJsF6pXjK3hmKNREBlsrY5MKiu4lwwayt14MWEWAR
PVVN/o4/qwfcbtPDntSGAEggvKI5/3IBL/92MlU+5NUwtCF0/AK9weW9xLY0+g9ize/l5est6IsU
B0olO0SUg//nPY7McYFT5fQSkWeZTvv9Kvd75wbdmpflIHH2Z1X0kG+omyQhTWZt+1mX12lNlGCV
eAea3iH/d4DzRxtNSc+bfwesNZ8T5wsxPxliBSHd5R92nY78ne+g/t9FXrx7iAyprpN6UusXKVWl
XmgXFLlL9DpsofGz87BqyOffq00zREeg4KbuX/+zYld662yhQw0IxCQxqcsyc2PDcR0d0Ink6179
8ZGjzmcISXheMO65NGB+uQOoM9dC8cL2qV/dYg52RMeujHxdgesw5chl4wJGqMUMo8DgcjYk58Ba
IGHno+CvfAQmfFmGYDeyPKig++iN838v8gO/bdvggUHQtUj7iIZQPkA+RVOszPQAf3zuCAEjWVwc
4ggk0bTF2K0EwZfQTZjanpXDziy3Q3DUYxmjtmpdPm85nMfkfo1LoM4ggS4X54nHAiGaCD+nhXbM
iXbWkE4EAL7DW0GE/oKeXXXKjOgEh8+wZhQp4GMYYzWGIH34lap3b7UNOnMQRerTDu4AZnu63ieZ
eCMKj2qOBu02oNKbJyoX910O03UqvodnHJqGxFeHnrrCGmY18WOs1zTQGmq4NcpE9x/iOVJqW1j4
PNcKQKu4AX6RKU3pArnc2l7gG6FNcdK6HTEOR0YnUzmQKwN119nqIE+pRlc5B/u5/N2nWW1K4/4Q
n/qEMxVUzp3kfzbIhRxnYMUm7tMBHLPmnEwVrcbwed0UQZE5jY2Bu8u7TZFnOAqYKswRUsd3LBez
5dceYndcQMOdxlP9eINcFVuQ3qFnj6B7VOdYJcd8bZV+5FBWi0LeRNUO1SM88JkaMp3GHC3CUvxy
wit263RELtGRuc5Tt83++Tw0nuXH1TAilTrkhjC8VRadYT35xDGn+bbm60QO/oJ6A56Ie6bPRZ6G
jWSl/QoX3gzPpUghXC/hLHCY37SWNSw5BvBDr6OvBZny7rflSYNTPr7KR+jB3f74pqneYvkwGniC
APGfKLpYSPNuyJ+7xWPoVjPYbzCa5TqKpqxhrRZL8NzoP5dEwqI2UoZ6LEz4pPM9UF+q76BKMJJz
8ogR6MEMi/i3Sd8NjEZGom/4fdFqOdT/Kfyf2K+XEwGwmcIeRf1bq42d6X+2d+eLvrCodwbUFlmy
9TgpymLK3+4TC6tjQz2cJdrozJg2mQfDoCJzy4v1SrYN7hRwtAcGHPv81C2fS/Sivw8q4tw5JxC7
o6YbMo0l75YhvtY69bZY0YCGC8lpMUYZeBWIB7qOP+KU8JactUVs5Y5/UFzz5hl2GuvW1D0+2n+X
PTCTS0440xFdPpRMvy5A0OqUMQyodPYSyzywkoujdmdQo4XQ7GyX3h+bws9bzgbTTn8CDoOxJ5ok
MEkFEieCZw9uVuNJHQ1mGjTt1zmyvuwxjPYNGxHxM71bLg02XSmMyilgSvYicib52MFaySxRHmoT
S4crC0L46xJWjh9k/lZGRjEnqI+enk+kWBqbUpnZagj3LxuRaAFj0meGLg70Wqsn+7RcFfecR7MF
K3GcqHbJX12h86G+mE4Q4qsWj1IgBmAm7SYF8vFXJpaDYizglnwBLFQkYwDBXGL930a+B+7MSnb8
TQV8bR4I5B3ZoxyuzQRJZbk89AUz5lepzb2cXp0XnLw/flgdRW+q3Oxj86mDZiN2wiSameduta/y
kumGXoGSb9IXmYcRWA1N9vImiffVzA7ON5mvzrM0qrbRX+MJZSoi0ViPr3Rto/aFJxLzNp2n0IKy
/GW55drjna2gmji7U5CVde+W7269l8aJXXE6jj5ol1pOOM/7vcgvYyCeNhRwf+7CYNaush7Kw+70
6OH2N4HCQlPRUOT27sqOlpFS4vpBwLa0EW5y6GDpNq2B/L7EHMAuUkPGnsDawmKBfMqy01UouQLI
SzRIXWqAOEhSmOIyiLCdSo5uYqhxrlKzF2WYw6GaFWACkAGzzbqzM7PTWv1BHTyOdsBj8FwvJaoM
NrKyvhQv9y4pQP1lI9bZjgC/uCBHx+WF9ffCeSqwLkBakh/qTzbZhNZ3+VGOGlA68IYeXeajSBjO
Hz6vmChoJ3o58QcrgQ0sspAdzf6WgXftleVCLy0pZYTPNfnhg1YrnbFN8HjMD+UqDT/8ICNoKYCo
5fmECis8MYyVWmwetwMP5GW2B264IpssRmW3Y8wJ+24z1obB8HaQAGQC5G0YCsja3PjImF5MF0zr
gLxWjWXk4hP1uIwjBDJMpSKY1Fwvbefvc/yxQo+L4DNDodtnFcFpgzfoeQrvZscFijesDBW3/LqS
/TK6o56aHbKGmTYxQOO5aWN9QMVY72q47U2InH7UKrLEDLp9NuRC0Z0bLpQ2DWU4DMrjDV0+iVg1
o+120CnZnOpTmFilPkgm5wGlsVrkNP+a6C/Aymp1SDADTHKrf/PATYocx1DSexMXTAcRai6uc99t
ysvrJYlqXqqF8rHffycvfAgcLjFoFSP0IUWfdB7wZQ2DXPz0WSovzMEwh1CaN2gYxVKTxMxytcBk
S4nwl9VZx3AvDD82KFIqcyN8X95L+m6hsXv1+MRuHc9I19ttqh3Sz/ONVD2AOM1ZMfMWyAyll6fV
FSQVoQqfNcFO8zR7wENq+GEbfCTOa2m3UjJl0IDhfeNfP9Ow8eele6U5Syghr13Da3+pkIgFnbB7
4ufKZK8iKSajttfZbjkCaVymxlZRZHkcOTggr7uTxRWg4kj4/xK7W1Hn0/ETiUfw6WfpMb5Isgi/
9/urATrSmdtxoJx+ma1TcTmHX9F2knD2yP/sr1VWrWIZrhW/K+vExutfVVY03/Q5yK9ux2ILkCVi
CyaisiowQIpcHuVQHXGxcnYiK3025gi35b1fCTW4YZ28w93OK8oNZzzLiuT54RL7gxQPCv3wdCId
QfMddSiNg9vgjGxXJ5zEC0tgvMflZEsuYllynzZWEoBm+Wz1ALSw34C/7Ot7S5L0VWEE+iI4CsDm
eklnqC2rAH0GXL22nIgPZEcy+PNZsQxtnfehoPi6vRmapncNF4bWRXX3KAztsF6i4Ns+BM61zAIW
1gQRYZKnJkJijkqRCdqEMPTF0GTiBle4RWUxt7AcgUuLix8ClkGDYzNDBMHcCH+RMiY1bh0zFPqr
VzZ+dOvH5QpCGR5SW+223YPyj1aDe2NB98YlwCveO3OeGvhAUf4GRV91at99L0w4pyVP8qakLMsk
jH+b2CnL6UYLfNvV1NrEAnfe5Mfjp3rgnq6sEslOPZtVyv9iUNsOT16/qcCgCZHa+zSwSrXlzQUZ
GzM4bngAqUKGqkiJQ6L+3Ecu9DROlbSoF0F74BHan9yDMAk4KX+a/CFnRJJftu9C1otnIVg5zFXb
vWE25HCWKVZ9RmZA5J5MhAc8Ek1kYf5vGJ3XcjLW609LRqi7IWfr+HzSZLYQDfzZy98wqr3xSmPV
peKpan8DvX1msD9Aqh27na3VZ+fIfk11Ql2Hlms6c5e0LgCilmP0lf2jE3ily7OqnUdr+G8ZaHcX
esVQjCZmY7DFxleF9foiw9kT8+CtK1oXRANKa+pb2po3D6q08FqiUDbnww7imw7h7b9kufbjMtS3
vzFZjPpJeV8qfSW/V+ch4RGpllGo5nLlU/tlzqtrFYxoogxYqUOqv9P/K5pyON1AilGbiLlSioS/
cI2JFZJuwUWsb3vMDmotpVNa/i3qd/N5kx8aYh71QG5vlTE8xAIRSF1tzIK7R+LRjXppT6tM17Kx
YRIRo8jLUnxHTMFzc8xXf+n1CfvLc3SemMXnalczAuSVgU8VsCJUTs4QXWZhCgmUqPcd9ED8cafb
A52o474ItZzfR10WBiJcd1cZ4/8mOCbrsfNtP6SHiRbgqbD9iT2PLnmCOUUu5I0Zuybc3mZA1Fmx
77ruRBv2pDOt0ixdkpyxWEKaBWoqMEUqfdCF+sbICLVM3KB48wHkonKFnVy7+u/kHSv0IaZvTGNB
OBce+XbT1PGnUA6jGNzx/arz0n/P73oabXckWOcVyZ9cLQuuDSbLrXkgFA/i+tyWEiTqer8cHVbX
6+JJnszai3Rb0IvoRIXQFdUi13CdwMWbEzlX9AJWydGPon5RIGv2F9URaYF3T3/0vHsJA4+O+ufz
ap+9sPwrxHEZJZ5O2UoglcBfaJcTZiBdy8ltk6485nnOLYjQmJpghodA/Gb0Ei6fuIX3KVIrBG5K
QlGBCevCPO3I8KWVlV2xVM3uWRrWMInafho16zZ6nG0WrcUNRxB+Hi7vEOUBREGb7H19vjbrTZkV
NfCcOOqfE6yq3Pn2Pn9od7EBhKiMy++Vz9+YmybGrX5/B6BT6vs16PnuoLdNqSsltMAizROm+QmG
wyjiUglR3dxLvT2OWyDZusWpoiCmr4k3r3usabiFfQskd7h4tWt62GMzJDEiVjUmCH1See5vy3RU
lN7/ctQVPEpVvmalHRlrY6GGn68pmk8mA4tI8PC9Octa2ulT9SLvLqVJ/R9MWw7dkpZ/wkwr1DQO
N+PrnCkJMjLhjr8VNGw/hiUywqIdNWj3Mh7T3cnCSuhsfhnSuIPRW9S9FqVruVoe17RN+7ft8szW
o2en8EAjxVZiMfoOUJbOHRGfoRwka3U8eJKS+i42AEu+Rr/HA3vjbjrLsDYWJI8ZfHYjDSOZLJrm
0cdjEzTfV3xAmn+yZ+HaVLcoSt6m4HByigzkG4f9WkyalB9Y+TdgbU6JDSY4SYMGa9dUX0iR1C1R
j+lKi5vCTSHd0G7hflqFLtaiKD/HNpnUis6gBY7a4FFOpmOvgOvqcntgyDv9volZz5U+hneF0uB7
mU6LOvFFz3E8Y+cfl7CykYdtak3EDLcBHgldo162NCART+jsDLEAaa1381qnSPLznwedAo0gpljV
yNI58S5HKLVI+Gtp5pPKz2UB2QhjkZnkVyEG01f6dNB7lCQl9s0ZbnoKi+/nPGRhtP1yhhr9Xq2e
nb63j/Ilu/Ib4ohCeiEeFQM1AfuV+EW4IDr8Z6sfF7enLGGk42hmKpCqT8a8cuZSB9F9eG+hxOMi
epbVLOUEkU8e4wsLKD5W9rqmhkE8D+7S2pXFkak0QViQh6X515huJ0ukSbPy0rAkMKhOjdvrVdRv
/UYUBtlwCWxJY7UodvQENEuyGrKpCpJqi5nfLYwrCm3ejeRS7Zyeyo4gJHoXnyNVRmJeLl3ZBmtt
K1HfNiYBLVccvnTuVN5lQJxinIi8rrILlvzpiHZCFnDEOsl62UEa5wVUC3/Unn+rhHA0733Um6gq
d3GjkretBmnIZpaebNZmihn9p10SXBJXjQfVJhe6SJfIOL/8XrJTEtxH3GYfFgJoO0v2QooJk49e
ac9YoNYpkHTeo0Sx2jNF/uOZBWsdLugvKC2Q6x4mHgxquyXxsX6rcQVTOWYfcSi23gqQ+A8R4W2R
3RjVfSDIYvY3XhlzYMTpVxwJEyTAkvuZ+7i3UpfgWE0843BOxIqqp5WE8abi2Vs2xLY3gib8d6Nk
G+/cRgscWRdnSVRH+TA1g0VgDKb4m7rd2dgTaTY7XCsdm6augvXUnsdMkyLivyit2t4PTgh6AW1N
c3dnl0okm7s/O4Fol28c7unRMga3GEePPsl033ZBT0EdinsIXOZHZ4+DBS1dyISVzXAu3lyg7HvC
POJCzJbifyRmWRPUbQHvleKF+Z4KulsF+4VY97PSCas1iCrAKnqeXeyCfmatmVkLMvR2aqZFWAvW
MeIkDj0+SNkx4TI6gOxcKIfDWj+5/I8cD3Q3RpbuSLrLzj3K4evimdWZpaHr5jgBeroR3ZccH+X9
e/wmMdZml/+6RldMNj/aMR5mxmgQImLVMYut6lzEtDOoCLTucn+r5SSAHl4alHseikVvG+08ZMU3
Ugmt9kP6rvQKHXfpETKetDQgpEhGvNF7wX/Jxx4Ap+wPumlF/MpB6IIfit1GutSBKF/cmyh3DnVV
NlFfyVZHIr7XQDTBn9ZeMiKQJAZdbB12MG7TEcTC33u1rcbLnQqSbHZaJ9xjHi5JIv9oF0FRfJaC
QN0v66nB64H8aSh/sO0FATBg/K0CeZPeL3bvB8crMaaI0IE4SW4gbc8SWmGZaiu5vzv8fGif910S
9Pj+1MdVS2oPoYUuxMwYxxsDHqbnKNyqLZfeIiGLqxdgbTexHiyDXnvnP4F3Udhd2BFDXSgoMKFr
EnMfta8hxxNUfl8kYSMDe55xTt5zPsPcop6akFq9pkNopA7Ep2Ov2Kie5K5xuaAV2bGkotQOoKxY
0fwMVElZro4VPGmNGjqpkC2JdoI358nuk7PLMF9FqcjtNO9C2q41B/HbNDexo3rKDfV7WdYbOYdD
SQL9F/m6u/Gk08RJr1xs3fbhJSaWuSZzFEBm7rwNFy4L0eEmtL+aQJOu0d46nsGn9ucIclxQW4YF
SAQ+jxwUkXAZGD8RkCALbdYiQmn1z62P99fFPHmad9S4hTa2nrXMdzt2Pe79vOajADU7dSK+pR7r
J4BHf3jRj2P9c4EKyj/8ag8R8Rkrj0SkN+Z9zydvGs9HxgEx5baDMjY6eMRewJvfKoRfBRG81yVu
7kyVUT5sXGDcUjebr/idpVNq7geDHE/6K5JBoQF7LWoHcXsD+PJPkZdNUfoGOBmH5XUF3+oGk4A3
qTpqVmiuX1H/3b7Wm/gjsG3PZOkGiQtClgS1y+eG20f6xnhHKVKckXzU0du1sIP1lnE7rLi9gjMI
bLHxzRd0VX/O5JAHx6JXEHJBbmyh7+tN3n5aOwskhJAK+IhJwH2a3+LsvL0DoWRkAWfImvlDh9SO
OgIH+fjqbEY9JHQJv64Fuef/jEzj/XecfR+FX6XRK3xTQXWIXsmFED2/Igm5a6dZ6GtOXennUtV9
ARKsVZ6zdkwmWflPywLnNknWKjRQJLiBqIsdO7lrV/2usCMb5CCcA0XwMTFBQk94qLyaCnRGkMDy
OS+CWdWp1AOIJWaQyMob3lID16MOmByw4e6a03cPo7L9hPQvGR7h5Us2kE1KECs/TPpRCdTSKch0
f3q97BCXavvB/rVaKEmKy5jKtn3BtvvwzL3zXDtSmRHMTpA6JD0/58CZUian77I/qry45ylOZXii
PmbBchp7blYoIa26LhyUCUswhkQPrvOSwd2g3r+NQrxp6o8k5NqdNXfXvVsCEKX3v6+KsRybKPqa
MQnrraf9eLGxSxtMSLm//b4GUtLwYUmhReffblkf01Xv6vUsposuO/ayRRCVxTtVGtqjNuRznzx8
4O7OnR1xJGrcQ276f+nCmIg+0qiD9x60vHp59/wcYEEWAB/koFQvxtlJRgNRtFB2BNxs2mwyFqNa
roHGG7pnhmU4e6j5RPw9VtL7KtQGPeSJi4gHQfF6vTYkoObmkYh2ZxkK7QJKhtgOTAe8xgKIDhfO
QpkkW9vSix53baUDU2t7VKMlfiPgeAHP1Dr7DiUrNdM08dmsi3MD9ZDPj549wi2VLADaQwb24QED
UWWSTrF5rgBsF48mJvz+ScrT3myrjHG6QKnjvU/Zhg0YPXrzFxxrxyEgjetB2iP7iWxmmGvKlYL+
t/AqE18TNrPsX0fHc6RjUK5EQZlIieX6+2XvGFY7KKoZm9oDyA/V6jCYZVFxGA1Nmq2YaUw5gSuz
78xghK7cliqC3DOz0C+sd5hkSFcjk2wQCsc5rR2zE3U9UloJtoh8a6OgE78cG1g6dXe2GDm8TPoh
+LrplN283rPO9eo5NDWc9RcNEVCCfhHTAJqtZBnumjbGX23DAKj/UfLOqtI2OJlyYz1xZa1WO8kD
HzpoWEml6gTAF+4l8EU6jmoY1uIOq/EDELW/rLe8jfhOmRDVQAhLmmI+OfBzmAZNxmkF79y0Ua40
5lWPRfeYsqSt1Y637W+2PzubpxcZEWS/W50Rf4zt+ONiKPS2AsNuD9DYsUuQ2HTjRGM3XWdme30b
71OYCdU2afM0InAIIdNSxjxNLVbk501GXRMhLfiI62CiU9cr7RfDOiy0RrbRMcPQ6lNhLMzPkdsD
ATC0qG4Sf+XEZDRlbZEv1ve2qVzHZLQGZrdOB81/IONPLLQ9qY19kMnUibxyQusEhqXcvmSVPVUv
6+9aE4ofbnF05CwyjQbGQDsKhQRmLqy/RSMkgWl8jG3KBgmT+KMDpBvGXaB6Q0UX/W61k8cMmUdl
22ErN8UWDf2xT2AkdaKIxRyrqV77fOqZfCPBbLlNmMHuAxDRJlhoIFR/B6b9ZmulIjtZ/HBGWLHK
xKh7ismzbNuD9F6MD22y76BVFwTf1gCOtceFFyQWCgiTLKDjbZkbcTWomZwD/Y+hmSm3hyxqLfXU
H9NdoJCjBkYlsYRWYPbBDiVVzXer6wY/ZPLp0c8zoI8EPs2PHivFKh7vD8eF0R7q/I2iWgKOemdl
1w1cOExGa1Jd8pEExXHL5xjY6yEiVpiZ+UxBh1ShPKiudcofxIPvYzAEA57XY8TFbbidcA9C5vag
u0M9MmuS37jImorshI8qwlDVFLZls1ZnwTX1ZvYQ8s9D27R58ruugWoSHKQf0Z28YY22Y3rBmaH6
9UDYimDxWwtsvrynZ5JDeqQRI5cxl9fOWCZCYd6DdiXcumCucruy3j0GqLKWi1gp8i+Vck8Bei1e
lKEtv8pnYrt5tQmwFapAYQ1nQsvRzWY05l43O/ocNkLmN0qJNfmAwmhaqtQkz1fnqt7jHE5HvKp6
tc7i6zEvhJteCkH1J4Z2r2qV5g5RVXLsrtS7OBM9Eu0WiwgEqZB1vRLGJwCnrKCF0nrLuiH1bOxo
prn+lj6dh800oDmIg8kOu0IrrCWFFXYSWUkAG9KcvngR0P2BMdpRfE6AHNT+WgNKaaK07PDDdcS2
GrkskEDlNYpi2VmhN5gquHTMe11xxkt1+nqFo4TTKKa7jsodfCXReYwNvsUP8IEgswYToP0b9muH
AYRmY7t6KPdUILcCTaitacj5AglTnGUzCUvtaZsK15mQAEtQI38P2CvBHcj3Wd4sBuh+JKOgeGPD
px3Bi9axzaGByAtXsQYfFKrSQA0CYUWvfyUrtIx0m//hlpAOGAHlsCS0VKySidtlT9DTQcnjqOUI
UC8RCQe2hU0Oh/fpxUmC4Fj0GaKAwT5ijGTykxAXETbWQALrXI/G+ivMUV/bGmM/hXNDrYft8Ght
nQA8u4ZFgr/PE3fD9BWgRl8AsYeHeJnpEBfDmcdjF+2DzBGH9kDlMmaQrubG4AZpWFQq3BJUmxYt
8qNwPwy8t59KaBfGVq3sqgBkgbcTGR65ZfrJYeh9oslQ4ozqPiLNhX4t5oVUaLcxZspsGzxHwwWM
7oJYHyMixSkMlCT5MhpXmV0XQRiUISd4n6a51YaP7mAxj91gN6B5xeXbW1IKtfIHhj5eAzmALwr2
ToLP/+21ekqhr9ZwvL0qYhXUE9pbMnjarOADmhLIAHeE7Owz8t/5Mir2loLPKrwOF5mra+BXepxx
7py9aFG0y2K1hfnToM+Hs6hyfp8+n6OAC++LPYrK/by7Sni+o7UlNhrzlGrhctGm4M3C6BkyqjbQ
TbGJyXnkbCc3T7ejg2cMMsGAFAnPKtEQ/7wJse/TRRaqwu3+Gd9X2c8ZRAQJQFAdtoz4K4xlALi0
JYEqMj/Pi+cpf24j1NRbceADbM7NBRBosKba6Jk1Zrdn8srm79dceNoH8Bd5dYwb7mY1Nnh/zW2d
BKpGr5OW3LDuJmJy0Sr/RmeoP4wNoY81DjC86jCyKwv6MtPqZUK2Zf2wFqvCLaeXW8wJn5PeTk0o
ZGs2/2wXK5QV1Loum5G5hDXzctSeKluiNiQCJ/fgG6odW82INF4SlUNkdSwMemLaYnTr9lbTSEHq
GVevgJnWEqE8JE2g+RTG/BAriGFocfWMjnTbRKBFKT++MPvOihUr1DL52gQS59ptHABHFJiDjizL
vqcOP9kySU1PpLS86NXUR9ZrG3dHx+Ka/TicVbEq14DKmph8knPGxaB/VN6ypBeqsPsQ7k2rIVZM
XA2j1FN4pnJPc0xV2pLCJwH187p6kmk2Nd3o6BGbVWGSQ8mPY6cfOcqjSGAlc3rYkoPctUcK3gAT
yvaHlaLQlwgG79N2zJGqDooFLF7q4PtxD36Xk9QmQJui2Gn5ajWwAp/isXaCEY5cn4HaEkInorHb
6ojEAae1wFOI1WfWQCZX6IWXW4WbRqkvsJDDdx9N5eHVH6rYxY8/Mq0yMOGdmOk3Zoqirn+bY911
8pzicn872JkUmpn0tqAbFC3ZYWlsuShlmWjnhcUvukHr2hQXbQkEJS3IZSr8m1DZnJU6SooeCTsG
v28t+ZShSFgw2LeZQ2eBmlaO5Jmqzue+UeGMuYCK3TFiZCn8zskOXwcsWWfGKAlAlcNS+iBuKucn
lzaEiYYHOtc40IHyjxsCDQB7Kn/LUWesTEnPYAV8+mu81iUVWY/9bbK1rQTJd3JzS+VWQyQNLubX
6u51wz1jfGzM1ViQXzL8umJX/bNUTfv8mcnQVffBUcPD3CIH1KVUjW/F/yXEV698ljJ8QrabmByH
iRQdUnX2OuYfv3v4rWQi8JTZlsrEt0IFRz95jqImB8f+hwp4iM0hYQ5/m/xJF/R297qogOv1A/j/
Wm3gfbLUUvXqy4jHjOJMOR1rGWsfdWSfq+ooZhglVP8tBnz+wcuXxE2cYr4FoZRzkJ0syNpvlcSO
/Oe4kVvwyUGlit9psoQ3ZRLMJJg6ZP83wnDI/JYHjgnSg3bYYTHo50xU1bPp2fXDEe/3V5+vs2dH
UqgJqxdqQOa32REarFpEdBJpetzaXlxlutC/qA5AmW7zUdRTrA+ZMiOSmbtjkm2dqsYRypsk5T87
AHbwGTuhVB+U5TApjatMV/TAzqzEmJA+USikbw1ZeZ+0B4bxGm/uVpYrW4yCuWiAalbyW46/w9ZY
OYQtY5g1UL1Q0sorpbYvPOIiLw1qnBWTjvScti4Xg25NsJ+bI553HkIF8Gdq+HX+Q9TFXMdeXBqT
q2fLUSJx/BBJfysBYZKxv6al0Jhrec+rmPgolZJtXXU7W6DNhMS+tuWmZEBwXxRZBuln03TFg7Kw
l0nAhN+lid8P4QtOJ5cNl9vrUgLSZd++nAFdHIGCyqfQ3kVMeI/oiQM+7GZP7v1ecNabHe4Vi74w
QSCqqxlrnmG+wzL8ALSWP4zbHTNi9bTOj/Lju020zfke3JzU9rjkPTvYqNPPMRvgKIS3Is0s27uF
UOd5G2i53CcI3AHVSfRXZtq0zGP9XsyO6G8pvx6YQ61Z0e5uHvuaeVJa0eDLPEB3gyD7OxF+cYi0
cMS//7wlV1XkZl5QYqDBNczWA9nrjacFDliW6uxOWW58KDDuu0v3bEbIzmZ0hkxj0D98ar0inbvz
HHbq8axmIxUpo5LzvMclnATN0mKbY3wOGLREVJmmKy0pxOa9BF6sPapFFZhK63szQlBatFBpswUn
RCij0QVFIBJnEJfYNvwzUQUVx0ed80JF8i3Vfe7dY85R3gDbkNwhjBiVG558F5o4v8YkBxB7iMqX
pTWf+ScIIHkKXXTkUrqyqTl0QhXHsrcLQctXtgbSnIIR9vhP0wOwCe2qBV0zv4lT3cIYu3jYYaR0
K+3CkQsUgig/VkqcwmDtAgTz/yKt7ZVlnlVxXvht/qiU/ZAtjlgONXJFsH3ksJxFwTN5g+xjIdeu
QWEPsWexqi5jHo/zHsMO1fcHJq32P5l/1ZQTjHfOm2UWfkB74dX1i9tltYRTap8HtR/83h2KD706
Asv5Xwxxvuv8B7nHis2/VGhQPmDyc7GzbO6owPrUkKWYh+GBhqunPfcmycAuUYYEjjQW3qJ0l+vW
a2wxIm+lS9wZESNLKKFYpfp7YjEQAXhK8oFkqFSCBaJwZUilNwzNFSwXcG0sQoRTzbeBkMKnMq0t
46SU1Nrhopt/AmX18g/zdnaSC6mPM9PbGmQHEqOFWwQeu+4BaNdFkHa4k7pT072lDELzN5DXYgkE
QuFBCKzIW9T21FWPJp2mmrlfkErikb55xTvBc6wmGcnYMvY7BjX1eRVR/O/LCK+gTMCah1jBONq3
55k/u7MIfekxPMHB2lJZhTnutGTBGC9iNc7+QujPkGWL33NmjjjGjYnpl/sUDa+ML2+tDWELjFTJ
/yjjj6MNF45mc9Wyh4hqEpdJYwP+AQYhzXl3zIRLb7MjmNq1fgGCKeqBNoZz6Q3rBdUpj1TIZoxf
XqNrca/ONEQ0eBGZykhldEKc2VzLVNTdQAcOaWH8gH85523mcJq0KsKc4mPqTqvcnyhetcdOso71
BS+0k746WjEDiTq8riupSvz4WQrLOG75grZ8F4xb0vIqUDIVsxTEyJC8pE7h65xcRpzecUvZJhMP
8ylieOGwLAwXBSRnzfzEh6h99EkubtlwEezPInk3gfefkaRAkqVPKkqPtStxA0t5Y7n6iOPVdXSA
mmAqNjRY6FArbMMYWU0LzM9zRIRNgSMDLKagqDat4AST2vFvVW0fCESYQABYS4HJZRUfLyoJrTfv
U0UwY31tPc+CMhYm1ZB3N6JAENf/qucjQkxHj9ZZRTUBEUZgtxb6nkjV06+eWZ7Uz8/YR2X7TK1D
w3bpFgEA/x3gmyBrREO6e99LL2WlYifhmA/mBdG1PE7nNk4Tx2IqrQIaP59qo8vAmb1UEl+3Mf+t
hbzLOrUDBDx5PTdhq7Pm604f02iV3Hr6d9NMtFIku073GJfFR4nVIdwDI0UvqLemkdR7+jFjg5sF
io1Aiyb7KD42wu5h6SQgU6R9skVI0vBMmujcwYTRdat5V+2xrh0/cGp8bIkhNyFec+/yb86f4va9
jxQ+6cWjysog3fHvLd/YO0+HlIxa5vnG2gC5mSCHqvXN9aBxQJhXwAYlSRiC80MMssX3I2mR1MOl
DqHoYUn8V1SgUBcKOYalXZED63M0826ZJ9MQr2+y3DACEgVT0rj4d1asBF37BsK2xEZPILxxCWWg
gVgDAWV9OQ8nfCozFdrbpIEIOjgsRNrmN+Hm4U9oYw48/FHCvmWY21laZkEywTFYVAVtE+c1q7CM
ooWLX7PJ/Rf0F1+oY4CNDJKM2NCif1ftjnOhjP1ZGPfQYtUriFkDTL9G1yKw4FlaxSBztn26HTHN
02YtU/oj2m9e3TEyCr66DPUvZXaV5tABu8ADSeRLMSgw2vr7X+TTYIRzD1OmO1ux4PAo9x4560xE
Nnt4tCloa8nzvTgMmIzfOifEslKykOxWOsVCbjVPJsgEWo9yP4Ny54YpktnLRLJ8ieab9N7t3Zn1
x2ETej1GkZn3fiJ+6ebry3CAmK+v7IqwzayGeHs1ZJblDNxOQOqY0Xmpy4Df541kuO4xI4PTFz1f
6l01d86c6PSkuL4O/dQLv4xnJyXevD+ITgOOgwL7swEk+o6RfCsoXG5JqFx/gTrta1zYEuhDmvbv
vZelRJ9Gab6ajRlr6VKkhJX74yk+FYu5aO8Ck8ZOH1cLh/ufMDREK4vn7Oy9yWhHEvY4Mpv7Nkn/
VPJSfaM/XCINhGHY6OtPPGsw8cqxxjJrYhHGm9nu2p+hsAhdkNcTYw+k2yH74v8fv3JcdUhC+kKw
BKGcqv5jXtTZukLk4Osb00TJ3xpC6PVd0wY9iBnDId4wBWgOeV/DrWg1trupLEwksZpyJvtlxMMj
VeSb6OcxhEupj9W0Te3biC3MgXqXg6LBVyFqkxNxAaoTExnVVOQF6uLpKMlTilLW2OoPYD87ad1L
G2l2o/K1fn/uqILaS/vnT+Bbjk0GwdpdgejPFcF5g3S7R7hckLy4loifMSkKM6fXPZiJZhx3S2U5
PBVjWpoQcHPymcYKvnzBwaepaoH59kYWDUINbWEE/xa1EJ4xcgVsrJf1NX4bMbDNDaY7hg3hMP6d
pedqfJJx5cnvr+BudkAFReljX96gci9apiB7IAu5lq2G7se5bYBMrWI9O7sHkpVGyV6JSGAIgpAU
/CVBuguhphPJDDuBP/eMaWuPFMa96PrU3EpOxeXCmNDSDsZgxJLpIiCuakAcmAItZC0O6XyL2KEP
QD+5pmXEAwoGQSNlTvHHNuDsdWF5C0fpqwrHZQMqpLi0AHCYGSWPoLQQD/dRJcFILf33eZJIIEjn
joQOEFBns02oxsL00jDbafO/isNPrCizKQUirRq1EeXnoX5lDQlN0W2Yx7eo9wlA+7ALpxEWG4Hk
v77xzceEMx4Bh151qrccgzxSvf24ltApqnkcMrBF74sibuKg5tLZTccPROQAeh1BVA9HAAo6PCwR
LKN6GVmvMyxoPkXlbFqH0doTNLZ2mv8Sylw0v8FvapihKVsi90T3L0U8UFHAAXyxiyliZrBvtWnb
/1kxHKD9kWT2oGtBgcYVT6QxrMlBvPnoCYWuX/ZBhdk+uqE1pKXJkFWQJdu7h9/j305NC9IYyd9v
bUHIRxJ0KjlAK9G81uVXYGheAEpnbb7O0WF4eYK2g9dJwWYMGJ8WC4rf73VbO4AnQTIeHT11AVAI
GanknizFhCh+1OU7AP94/p+YPF26+R3HqXHLGm3O8gdtTjrCSlvG4JTC0480O8QL84MqLeh24wAu
MYuygZgYjkMaevPmH4/94LQhzKoV6EX030b2r9160eULdjJhcZhqmWKmCxdV1Qhr+EYErEgJ2IWY
mBmx9UAJgDTGR424XhganW8V6brCnq7u0H14UMswA8OHfPaoSt6ju4HPpGGVCGEYbTCFQxmYbRQz
MEvhqgZ+ADER3fxA6VjnxSJiDqfZnnDz+h0M13fCT6NkvIL92jkJBh9spBaAqFe3fy7Bx/Z4VO+L
s9Sao3m7ANsefZ4/5x1A4mVfskmUllkRlngFtufRpTfkgsy0IvdHq4ARxxU5AdRnDpmR8omjSwwm
rVh0caUftHOE7+AOngiPrmTUaU0IHAmxrRr2LwGx+fGDUce3H1vh44OXUCXQh87dH6E4hw11lmht
dB7nbA0NdwB1+gGEkx2Tp0ola6XeHhl8rM9ISabedeFZVl/fv0aENtT0LAZ5vvochFAm76aMsa1a
EUyR8xLKRgx8KTVS37ZonhjTo7GvsWzcmde/CxjEuu3kDW2aLTuoWfnz3q3AlzqwBv7O8FnVECpX
g9ua7whlj9hq/bRQi2d53B/kU9lKnw+pO1JIykO6JIVZiXAd4uldqaEXy204om9CxXdG8bUzv341
wKiYBzzXvhXCek9DzaxLIbKAJrASafonI7am4N3ZrYraOu9PdI+5VNQ6dX0eoA0tNh20m8topWDc
Hit7TKfkxKdbum19zXU0ZohPjbTMJZy0cmrB2n8/K8IQAA1o4vyP4z0/B0EvXGps4Sz/PjnwxJnH
veNrhjpvtyDi/ETFxJ+1KVfHioT0+2SPFqQqooIIE0UyR5jXebOLBKe6kvVcThFdq5dFizWvGoED
b3OXPNd9R95slLzschY+UNITzF7RCAbda9/3oHlUmaGi9m5b+yX0symSdqeZSta9HjdA+fXi+TnA
8v7iBpneRwnKkrGjFvUgOjZRxyU2VAFDZiof3MISsc1psYDiSn1FxnmgnI2x9fWoSC/8KuO8JzBS
UM6vc3NFl5xUdblGMLOGScw7LSCL+QLUPe9LpYpdJN3IT6m+BNs0Cb6sUo0M5OskmyUiiw7TPK2D
/RsTLJFs6CTP2m6M/aTOX0+5oOdJLc5RkOZcjqs8/alqwzVROFykxyitYpHfqfdw0izfnNLAcsSJ
MRc+laeBPYhjF10FRGaOBqG1WZivQfqEavggfxSBJGUYAUvSPoLv5ARECbosJvQ2VjLs2Bhk6UI3
PnOqLtwUHEako7l2kRt/R5+MoCcBfSBuZUOQrSMCYIPvEan97qk1TGIO4KBZqBqU7nC/8zQEK5iL
mM+1Cou4ASxcEwBNX27Vpnb4ZH050W8wWxU9ZztF7nA1KvRENA8sY7XPz6s4YZjU+wxMGuFmwD8W
UjLoBFAyS66Lwxwj05sJEXrrDZ9XOT6dWBI9Mvxv5HcJqLQ/zI6SaJy3pU/V387Yy3Lli4R03KhF
yKXqJ4u2sSieOB1YSvYgDHpHjpWcDqXBdQHkSFpKeeJulpUdg1qtRN+QEFdRpN45E1fDm2yv2e6L
lh9yn0aaI2k6hnA1mZTKa5u/nD2LTDM0OizVZeo7ITcevEY0Nrv9AB1HYnwyDqaCqP2H5NJ37fGF
5J8biM6wvj+8EaxWmXrdfHC7ai5Uwi4+egS6KGUdUzcld+7w2QhuSi2iFqpq5Un3wAtU9gk8KnsE
BrW9KzlXYySYbQwRASNnT0HxTz8+AXK34DGZwhUdzjIWINcSwPdA3ELevzx+9SSxXvHHD+dJhMZd
o78v4jDPYhd1cEXaNOS1DfCuR+qzXWOjQfLqOW3nV//jnZxyFqx2HBNk5FKvCxDZqmsPwOkhKqdL
hPEUOZYUXz4+6h/96xLxJPu9zqOqeUzVVRsdx9DpB4feiMwIIm1Bgc5BifhnInJmadvEM+pDsrmr
5d+2l59R4HJgvAALqvy+DWBbUAgEtgKeZCgaDb7br0iMc1AeBtXT393e2pKseYSBAD0fccDIovam
3ZZkx71FgeFprF90LFtsXVIgGiyU2yG70lgCQLu0WpuRdMeNCUFK+WHnueCzdmdbKGgm7w5/htQS
G6tScaYkLtbBgm3FITX42lW+IxQ1gNeO5nqiLjCvoSjrSqilQxspgCV9euVxVo1BsfCg47Pmk1/H
Tgj/icP7W606+UtAqAsmUyxqY292UsfGcj02A3Hh/hZpivvdGKz08+YNYbmjtAh3nqD3GfU9KSMg
wizryisrxWAM++TS+rkKWFzxzRxwWoAapyPFAN3mhxkvMwEy14SNuh3tW7i8Gpg9glT6nDiGI09W
YgkxRUOOHhlyG5pMm7GgOLMS7kbYeA5DB1s2LpWlpfQSq+hzLy8DUVdojntrxInFF4Hjc+jLbyfi
8C2/PNT1OxsfEn8sAbZFnMw12+2fQMiPKOrTyX61ABY7ZVQBD1g6fLcEZ36v6eqFO2NLktbIJUAa
Yt+9o1lyh6FLmTe1FWgEzObmp/G+QiPhxUSAJgq5SEh1NElfokAkTBt/XQGVXSV72zz0x6GyByvK
VuNDHemJsZNZxWZwpT3+9m5QvWNYMdvAngN8dFqeLvVaj4sLaz2jsNI7XJI8rftq+lSvCsP7qJwN
JhSQcqwlB6Y7/vMsi9L1d+2XKFhlDjQRb8ZnKS+gBXbsmag4Xihjv+KxqNmP4jyR7yj7jXLVfPC2
I/GlmD3KR1pu95PwUTT6oe6nhAf3WgGbsj1LU0r5LTZxvghHX9tB27Blp/lvVB50rqD6iqONKmuN
V8bRE2/VYeuiMCSDzNd75vNBmzuAU8VkerWhsmQ+AS4onbEBx6j5M5F/lNqkHbX7GJZivui3V9QA
41GiLU9nN8euLk9QPGdBtrL//BnoFfUcTfeZFXoaub7aKBJLDvGqYydXmSUhXujrUuP8NtHVZMVb
ZdypuWisLyJWyjXaIjkxnxxPE4TiZ0d1Gt2JYYELjSLeXf5UDp+Flx5DrloX8Wx+HLg/uV3WxagO
c/r2hTQT2bJE2gPH9aw1lMSMCDxdlMuJFMpJ1m/SO3mGyOOoZM6rv9LrgvHFZeG9dlLhHep3dJAC
47MnxeLp/q1IZUHOXITmnsafBqJqqIbGDFWlZqlTomcRrDsbrwFyAfQ+JR2f4qPNxbvqmJNvq0Gx
NJHLdHMkDHoktDd1vJqRK2ptSgMEweFOlr6/tOwZ8oGt6AQO5bSdjWHVG1hqZ/RnDK1J/E4Hkbw7
ENSq/vdxJXYzo4OSw12MFPRDDRuLX9ic8pMxYzUZ6+RtfBxgRro2IrFgo/mjYWAcKdERHw6G4hQS
xe09dTsmbsRqxIDJvYXMnKCkGvvct8ObiRO81eql5H3RbkvJ0Eq7mlbOR/iNX7OGsT+DtwucorMi
sxHVmTsxXL23DhF4ZbeylpI2Z2DMytbf/H1QvqVfMBEuyf94c5VUWLGWf6vjRitfTtyc8r7eqG0l
RnXoO5xXzbUod2G/NH+so9kZg87hwwifjT7sNEy22yePoh4JseXhvADBg8S0jkhevZy0Qroz4eAX
TZRg5FWyiWb0zc6BUUuhuEDUYZa6t7qPW/RfySER3db7XqHSTRC4qFCwCyJOlSASwsKqXlv35q3i
HP9ncgJdFT1bRC6QdhQ6wRYG1aetaFPs3isqgnUdrF6n/fDsUOI2CGKyyKjMXBkWIBI3k8kAdAay
RuedXQfqytd6LcbY/e8+XftE0IWAWjVlYwRJ196bysH9SpoxeEUO44fCe5YSMWWLD0b72sLtxgp8
98f7doJwJRyKy2eG111mdHo9htBzm/jLyvLwNZ2cnfQAs88zEbRpHOUkYqgJyhsJL99J2QLUNlBO
7IcDE77xCdxOQJ1x7Qtiqj7YMd30TZ3u+11WHreHNzsRyhAWym0qq0eBU5ViutsAw12DdGYentrd
ogqxbYPw2VVYIEAua799ZSiDWmdDcavJmbBsOvCUil5uLaWs/OX6w8peIfaPWvRmJXC6yTPXba1N
uWMRygPpqMSDAvLN+GL8vNZA6ifG4BwKn5Vtuu8UXERAGF5VH2v3RhAJlHHeNSoIon2EEz7/DXzU
Svl71tLYO27irZtTA4IZZYfUko29IVEacLe4cpxAeh1my08N4VqvKGnc22WXDO7myl7BxLMvJMe8
7v8jHMCiUMUfYfR1UFZhk9M1fNeeULnoI+CwvE3bRRWELnWHzs3Mk5Ks7OhetmW4ojZwnOwx8AWC
fA75FXkgrLS6RBknV94oi/6NivFht9Tgu8KexCyUTRX4XTSm72ZLYcohxe6mw52CKj5JeVRSlkVN
DuQN5dRJTg5Tl7NS/FEqoo4PeG5OYYk2vXiFXWH5iqiH0MEcXFNlmTgV5BXks2L5eUPmbwgfLJmm
jiAC0ouWaCDHc8QZLpInSkitPB7GKCfNdaOArwJ3KA8y0tTA2MUhIhZBUVThWOIe+rIDcY+/l6yr
HO2LJLF7tZj3+mvsEWZP2asq/MfYcWzHpg6y/TxitLWgN0+cRl/9MyZuNC6MV6m5SYiO1hRW5t+F
MejIrGyXHkwZKAoyQnnoSUzmx63wqkF1FzKsq+gxUg4vkxp9mjApMT4b/2yOBXq42n+t2W/UEXj6
sDSeAX0BhHXWsVorxKHdkVEWsryDHAm6BfwoxSRa1ExsZI1FjzF5wSpMvJX7zV+4/7muB1Yp8OZQ
rit4frZW/FM2MXewmBzx4JCkqI5um1R0L4Vdm0oQBLneduOPn1itNG43a0SMMmByedC+29uG7EZE
rs2NsanQcSRkecuYVZRY48nTTMhdxRH+MYGBFKVMx2V53fT5yfBTm0TSzGQw1WrVt3gWQz/1/H63
o/5OuIZw8K/EnM9kXgw/UGVcRbeQZDksnF/vZe+17n5MWtX4n++8ri/Q1FfOmhs1osMsxYkH+6Kw
qCaAmLCk88gvRS0TXkJwDBMJHBfJa173q/9UMgtgfH48/p+r3n8Qyr8XNEbypF8q6xBo0c6usQy3
GnnoQZdJaBtZ/LDBBFxxtKFNy4+H0GTcVBj9bDgHkSN5hMek95lfpowB3lZ2n4sNq09qbgQjoa+5
RrJ0mkqnszqwg2BOrIemDigdWHeoVkft3z4BTXJquw57CrYpTTlVPyXKjkDkHbw8daFUkQBGwY1Y
77fl20jE2cNcAyfMvB5e3mU2lK2gtNQ1Mwxes5cnzEu6cheSi3a4QGE2kehuSyjwDPOVEiA5dmC0
58ZVLFRvqRFzmEaBYxO+FR7Jd96Af9PLxJnbtVNqeFPRdtDzqxFQilsXsfWqfNmLI0CFpUgLp2Yg
ixQdljqKhdOGKEtYk0xNxYDnVqfERicqZxQ8G8l4XJ6SC74II5C49QHPeg05NtlQu6MsQ1jliGx2
YKB9fkVOsT4jAdWc7O7H+ylxJRslbZhxp9r+3ogTrAkYkiWf8qepTlZeflakCRb3YkHP/8nJf1hO
gCzQ/64fd8VgugoUYJmduakDdDty0JNfxWPWeenkF5JRLiMVBiLUYNZuHNbEclsxv4gxLe6nB8Fp
4MKux9CkNltdeCD/mVsb1lQe6iTO/FdRJ8PAvkxmk/8pPRk6uqGUa9o2OBTIb/W+GnDADtlPvblH
rrh+8cnomW/xPrK9QeT9RLm3QapfhmZIVlJZ4cVGD2JdQpCA6hLzVhHAV/8G43eVvk2XRfhOLR80
y2XVbXNv/5g+4NHSJH3QC/r9jFpFqFDi779KtivcqQXnNu7XfLp1Vu7vGFu2UpwaxtF6XoEHsBoi
fQ4tIZ9rW72SvciU+beST5bcKlaKcFjU1ZEy1yCZ03O1MHaokYYyLw4L+ss0EFOy8cBnM1Z3ynNR
KnjjJI/VJ/c9oGcMzIzStBOyKJ0nJlmakLFeUCfl69o4FeHOFECHDfMmTY+KF66idQrpkcUJfyvM
ssy9kg2NTuiZwCz8pcqEuvcspieKF2r28AztQeQB1opXzrk79IRRc8dHFlTlOhA3FXBy1SKdNCzE
kNtHsiwphKqgd/sRFroHwtun1eoKjk8rXgaCnmirn1yQnSHlxchE9cXUUmrScRJATV1uGzrykMtf
WhGG0GzarexrvFgPLwWwVrixOms7jHKYH99CpMegPlVMgx43VkDMWNozH1W8hcba/NlSHarFljNc
7rmeimNMjmNuX24AGI+26Fcj5Dpauy8U7f1QO5iXv4N9fpPesQgMpd+a8Q0VLmWX3uz8EL4DIRne
AJ4on1L18MkZISSE9y5WARk0AM/v8aRdNXfJy5PNOEko9sk/LB1lA3ByUh7IinNimOe8BKrI615d
uaz6ZljZqgzzbh/Nl0NvIfWwVvEHy8mfPqkuB0VXpe/UxY+PoX+PywreWOlUjrIfl3NhzMLzdrfn
EGgtBXlnPaPLlW2615lBxgzOv0SEpEQd/rhGlTf1fRTf+sJEwJ/NtsJxigIv2xqkHZ1ySXlfTGly
Vil0eUN6nL5nVTkKx7ohZpQk96GiK9bnRVAIDGE5XxKdQSBhPHi0smz+UgV+UhbYHPEWUwY7iWTa
fe6aWw9aB1RI+NGQTGILIzr62KpXxZ3W9/U7foZYbnOwRZT3tLTJARPlNPrBnlYFclcVru0GuBWB
TdG8XP0RG90xYJ/6l7rzs/mY1J6q8jT/JoYvNr6Cwfh2eT4VZGaUShclfWHd9tr1Crleh9rTdS0/
UlVM1p8yfdWnsfyCyGCtuB2bzmv1OLbGouJoct4jV9PF/74NALuOTCua7dqf6B1Ea4CQqz5zWcUI
f2KYghSyPgwz1upK8yg4xJNdEahpLD41OHMmqaA6Jm2fk1FeKbDP4jTwEo4VwmsVOfwJ0RA6vB3w
bxL7IhscIk4IoxZiMGGTR49bRm/NAadh2Mi6feyXb/fnEPrZ1qwT4ABppFFNI5YycUBXRMAATsOw
HNRZOVT9Zo/4cRnAbYsu/aF9KlcPWAdU8UJ61xu0kHkQTVLWllTWrLwvqa+nRS34ejotuOxcwSDH
dl444OY3xAlNDrYJn2Z9A5RB569v+sTISQ/hW8g+3QgL5J04cd5XoGO2TVW/f/ysAzylt1EpfQLh
mtACHgcRzmwnMzWR0+lNIDdkAWte4zckLB/vGHU/d65l9cdDyY4KUduYEm/CUoB8945FFn/10fvr
L1JZn1W4DL5oWqd+V7b5Mmdl+Ev2VlnxAJgfGumhMCof7Bt8KNoG3ifap7Ias20M+ufvuqQAgLLb
KCj+ndnxHa364qjW1GSo3vC1FySL+h0mlZKGOIPIiEu6fflzWyS3NMT7WaLwzh4hTDrrsHy8s0II
jTA7T2HXivGMEQPH4QgiqAk/DGWyLYmxKGrmRKqB+bOHZrg6tHh/YUqiqVR25xOYT7VMegwZlgXS
Px7W0pEGuenTd/NdIJY29YlmphxkJ3uCpEBXmZSoWYPkznKnSeFTOxZXC1t2ucpkK2xVLgipRxpI
k/b27xvK0ssxlUOVvAGm28IIYMqXfHRWxSIwYPV/D2b+l4i/h80XzRVt/WrP5hMiwvp50MqGdeNy
cbyChhjtkllQlvSHejWODfDDl1NCLVn9/0uDeRsE+td+cNMInJUaJ/JY4772DgKnUetJ61+OWNSy
DYhqYFhP6OU4wGAGlX0KCzxTvwtphv7dYtvJpsccf8Iwl211a5a/2VPmP2vQYaCTlVdKNdX1Oiwk
BiI8/fCPz5NEQoJ+u8aSYZ4RrPZPqCNQk8Cwjuja/abXqcIUjSrgWmGBYDjRMCdmE1OUwwZ6lYAw
k+H2c+Iu6SOT+m49BNmExljUZpYNTgixS236z07oeXZpOwOfPAQVc87G1Ma0rfhhEu1MlR08sJPI
bb2+0KSxr+mSvKGE5GN8Ue8EiTFLHI0K9aPrYBDuviemrg2xJvpnPgfJeMRI7skrVYa6YK7Pbh5u
XiiGKmPbMxDMhdu042p5Bd3aO+hg0uELaWFCU4We2aAYv5VTk9HmXn/n/419fpD76vKvwYijxfQr
658JZb8k/Kw8c46GHAZ9RQwC1w3vyJjuox/F8JUi96A1tZmAzADhMVzvKPbJgIBVbzmknCVc4tEu
IUp00DmFHZ5pMAxv8RJLVDhHuzcfl7LJiGJ+tMgWkDULvrdB9kHa7Zo+ElMedQom7g7kVyiMfbjv
3V90YhAyr03+qbWv//jhzPQf69UB5YHIKL1Ez3iKL70GC9tKnoAaM0Jii4zfK5OH2bPX84KUFl5i
bh6ZdNu5+mkqBHgVk5piDOzEo2Z8rDBvMKWaEctx7Xpc+zjwr+1dNT5igXUKPZrpXAZZSXtXHOXP
yjU1boHTdRb/X6Ixf/wD9rfidk4jHg6neptm5f0k2zsgqL3aRekNEJK2gcn87AjX7jyLfXW0zpU1
I4RPC20YvIM0o9WDRZlhpFfPA4lCFCC1WeDVj+jp88Fo5I3GDHCj7hceEUVz/UjxejSQT3ibG752
7yfvWZfILD4p4MkV+eonyTmvn/Lp9TX2kccEUdssvGzyP0s0if3WaMk5Fmo3LOr5Wm25lX0j3k6j
nAjkZ7lVyisHkPz/tltRRnJ4ZISFszQRJCfAU2ux9M/n2f1CWO7VUotoRilZ9yCAaeNwyoIUQK6U
6bDAOdOJBntOvGgc6WJfaE+jgZ6v8eFD37v20oL//B9+KwCkDpBQldscjjlWNmjhzQXlIfb7lfxw
DsGz/5kkFwq6HX72i0ikWjopU607/F1Hj7oIGgzbgiQ4fLySggm80pymrrMec0kPjRZuX1DTg+vx
Lm89vLmF8Qk/lEksyGqFWiBkGSOUXj1WpjvJo6PbcJve2aYnduTW88i2Hfrc89ukD68wtaEQdYZZ
bozGZxC4AtEAyHAz6O1qBu+mbvQpY6I45TPzSDvf/jzAz8byJBJifZ1hzytKIQYQWQKGGQI4DIFZ
kz/IXsCJnCI3mj8oePQRFM6datS9jNLIxZPkZ6DV2N3bL/QBDcOvZOUf4ypIB7DkjE/iSmOIdDSd
96L5Qk3hndNFUtt1yBNRnURK/q3xED3ZusvX0x7z2Eb3SVziQqh3E9581fkblh7Eau2nVddTWRlW
oqw8iqGMBa2Ott7FEzqdQkcFdc0oWIkQTeLouW4LpymOBivkywxC5ZkRWJeswHaVrZF9BbYa+v3f
WR4AMAMKjKITb9lwcPsB9LR4Uw+gJkiLLvBM7AgFgcPskJ0gvpeplPfZWHhZF3c6RN9z0q4i9KE9
QsioU9uqvA0/2kN27TEACCFvCRLIrmh35dWIqDJZUXwPF7pOEazSK1aihzZe5TDKvn9kNwb8YgQ2
XIKDj7V/5A1zbWOixJpSrV8L8MRj5EnnpjwoEU/MhvHT9AxfgD3NRyqWoLP0eARpAHYJCM9SIAe0
yS3GBcqFuk5o2ftC4xlk6gUMbLTnOEX55/Bm6V+GYsywr1T4kVHWttogqv/NC/l7/1aG8PonBvz7
0FI2fINQf1WdCzqNXZ4AUpSyKK+kI82VHDwU1ESCTNG5DDtCau5RjrjN1CyQnrkXB23LiPWwK2C3
LqSsIebAtRAiZ7ild4kN9ziladsc6wpKEAJFXYzcvaolONllc5C441ArKKGmRcZnqT4t8Y4E75h2
hyA6KcVf+FH80As4qWlm9PxxOdtLAb7NzYJPTHv+3bOAZaF36NQLavi1ooap6tZTs1H3GlJjPK+t
+AkHivFU//g6h1yoqR21OKi11nEHFtrWvCaF2nmccdW6hDNwTwQxxERHtwPqgK3Uj18dOaZQwun0
pSUkRweOcAeN+84UYxJdI8HZJlu+FBGUHCrRwK91k+ZjeqTTHaSJh0ck0FCd/XbQrudk9lDd75kB
rAYN600fRahVge0UA1B2eOFn8y+I+mXcnIqS4sZ2uz2njJV+Q/oGBVAGbK2xQEGG9F2Kkvo9KY5w
Qc5V1XIM4mO6/0ilUU4ibKuOHeTaPrleCmEWkHJd/1Q8N7fARIVJzOTVKWlBx9B5BS22sI3cqoFR
QnyYhO8ExFBOq+FBPwfe1DxQBOW0yuky+WwSL7sTVxl1ddQHP6NE0+1gsj8i8JboDbqWeQ7iqMQi
ZxDQ5cP97tl++9dP82hUV5Dx/67byihqiK6wsBhz9aUudKXrkSWohcVluzlUFNHN1w9vxr1UoQHL
M0YzWo7tuCS98oURVhhrLEEmXxB/wzbUNK1eYp+yADsUe3JBSFQMRKVSt+oy7sYRSJn/26/3g09Z
hW+RxN7KlUZH61Xh/ja33tZQyMjF1fja5mk2LXjj2VDo3YPP9QepuMS0oDW50UnIAsR/FtNS4UdV
L85f/VQ0gSX0Ru4kJVcIZcqC17TpF7fJfitOoc7ackxCwHk9NAm1nt06hO3iw763pn6TtbC3bmV4
K3tS1zKw/VqewkH23GJAI335dw1QrEBOa0VGrDKWeS2mjOtoB6ydjGgX8eblROJLWDu/Kj9ffqCI
5CrH2Fv5lVyyFF0BnLjn+JjQHqcqKBA0K5NDANvq3AH7w80AS/VL7Q8UrGDuSZ0Wg/f0bH9nr2Mj
ikoXZ0dEABu54tV3ywnIjx8ogkDMBySJudhmQql2XoyxAECtKuTE6QTXuVdlVpPeHDT0TJ0bGjby
JaUlIpYkPrpGViTJU8k9Zx+Rb6o4/d/Vi9r6OekJLxlPj8kS2wlSRYmcmto1CrOV+AUWmyZGdPp6
aoD8HIf+8h5XrCEbLKK9ZZjLLoXpvYj4HhQn74V1fTDnQqvZKvE0cXt+gneRPJ1HlUOQqS7lfdpO
vGtHM3c12x2pTv/MVMHPTfA6mFrB2QwjD/ucPEdPKHjTiKR5CPagBB2zqL21LnPiSEgIaLmM6/mX
UQiKxomHPLx0pwR6s/fT7tprdmHgwG8CTA49ql510AmdVnqijwe7nBSTkPrP0BO/C+WQaW3SFSAp
jOOk88cF601Q6UVB8R5fKwN6Wa71bwHGJ7k6aVDyyFZtvDj+GQItkJwNUjr4XQ/QdopW6nPNrMsp
ilhqzG4tNky71dzb6PF9g3ACmjs7WgWduvdrKW1hd3yKzABUysHYoHJS8FhCJbZNalRDgFjfZpH5
Oh/57TSgW2reapV+IyBazIaa36I50/R7AqId4U/wkrIwlKZLGtLJOuQtiPZqfHiDSzNL0rBsi5iS
ELhOolCqu89biCISzHdidTIU/HgYQ7OV8FVwAPrTGcFz0vq1doyWw/tb7xNANVee2o8dIk7JK+3x
JafwgnXGbAtNrQ/8cKaR1iXj9/h2ifz7Sr6+dFVEoBuwQOHKp2ID5pCK+1Lob9Jl/KBxme7Ojnpv
BmSE4QtZU1p0C/HWPJlBjc0NTyd6JR5Cq2gBBFb6wc8cYQpyqAGgSD6VmRSDUKxjHslH1OxTsQ9y
Jjzj64JOueTmHrd2hzgaOL4dsYrCb46EfsEdTsyKnfE+FZAUmCbgkKuJ5etck4aleMovbEioyRdS
zUVBm08K4JvbapjfXZ4jnM6eONidNjhKc+Hg4DRMqDhwebjOr67/GC3oMByTc7b7FNNw7H8FYSlc
GeXnjN0dvItQ/XXB99VhtQe6Q30d/ovaCwZSMkBDnlVYRPgjI2HbsepKH8kQJeKIFwVHr3N8lM8J
2T83g+Flq7uLEeXaxlkFtWnHLC/OTXzxOZikDjwF0NlGY16uZOT/2V1YVr02j77ARdzanQU9FiOJ
/tJC4IvKKEtlCYORs0WSQNJUY07HkyuI8P56XG4j7AE73NcjjtugBn3TELV8nFNpHQSYTaca++J5
0FWrz1gy3nf9J0Q7uSDnudejeVRnT3XedT6+X7jkiXWp0OWfJg00x6CGHsbh718qGgelAkEnxQlk
DTL/7nBi2xYMpGQu9KE319uRhrRrhOdfQqnr8pAYUHuMYqjXnKo9ftjAR107oSoDkFXJQWJwVyM/
gOuQVq7A4CLXAfsp8wW1b0BkNP8x6V2zOyQ+PaCl9Sj077d04rLiDuPWniOcfzMnBWmm73jvn+XS
+metWFCKsLYmYe+8crKVyrxLWk7CkTMCgYstMf24BIhfyi95wUoB3IYRJqqo7YusarL2x0Ep1E/Q
XsJ6eYKa1C3/lS61AFmxqaH8it8Aw6D18lP+lG1UVyticfALy3haE0uX6uobXnBHek0demRbWcI/
s1n+CqocsGLSpcGfp9WoI6tNd0nUj12FOr3OnC55t3U7uYcUOXfjxtwXRcZeYn2t9s3Ge3f2jVcV
C/yEEGUPuUK+aVfcb/VVtmt9qDlnT2j+ALA76RMB1bk1dsT2ty50lHoX1xGOQ59ytGfusKOLNc9/
WD4CATiNI4eyqzypkOkyWYD9uSVrq2rl37KQZ+eETYl1jTReiHCPUqw7LSC4bXXpMXGjjmyVtYBo
GHb2wVXowyoXVJaicWtV3wQxhaJ0uN/KkffVq88t/w+wrBpdiIcI8nQX4m4Io4VD0B3FDlDYvrvK
9t/6PM9dXZRyFZO2MqSGQEF3I3qiaCE2Xb7p4eHVGTXEO5g6ufNAJKzg2EVnht5q9Y2vXbhQToGw
EH97iMJqwcaLlJ8zCseVyjeMzyi5MebDGWuwc6n8V49IuBmHXuFgXdFyy72MF0l4GmRfnO30EShs
g9YZ0HfIH1uG/AiR+xpfwc3jpl5JU8g4+md9XP09gwcQxOU2E2ZkXy7sGgzzVzjHeaHY1ogGSBK7
RvJQ46LLUaA6gdo+Na0WUk0J/jr1LmhDO4D1vcpobhjDNxhKYTmG4VmTOCp4XnSq9dIUZqsjh5kd
PPIgfpceMkiCa1RH+dIBDTUfkfuddG0SRpgJgKwY5KSWdPavjlQLshEhMg5NG9FPCTbsRtRmBpJh
koW+RThTeU+he5X1JwC+Ju8GX3kC+Cv1uTVFbcBKMU7o9uSLDHfigpzz8InFmoS8mvyEg8qvEHiG
EUQtAiq8WkvsHbbnJx5AJaZxDcLlculwiLd7EFOG99XKN6tDARhfaxPzGqVDSIYUSjQZs3bKma4G
/rMKu2Gucuqa1RcAcUsMDnPZX8jEop4lASQKcpABp1lYLD42YG0BklQ28KMW3fB7g9P/O+DBlUa8
plvZKxHa5n9ea/vSXwh5tO/5Pw8Ug7xv741LNL/FXHAkyaz6//JkNz4dQzdCeEZpLcQ1fj/zuCOF
aXltwoRvkx84MUlgyzw5SkLA5yMDIZcA0GfK+CiiFN2nI+Di/ji46M7UoXPadRUXHCBgi5ymh/+P
s4x2L1reiD/1yhCPHsjbUKo5MaHPMLLWyoqQ5zHANlWdDgSOrjIyCag6uNmNlRxolquAVfP2veo+
cYj+SgnCpPPmqm1NX8A3+DPAzhwxtK4Wy1YYVasGHwpItxvad0YcUySbNq4mzYzYQzE5swVbKsR1
Ogha+8EIySFiSuPyDi2A6uJVkB4U2n2xfpa9+q5FvGNW6Qm2p9XBPvrjhaI+RzHjEh7Dq3kvLuPc
ISHr7uX1cOk5bYm2wvPUByOIh6eWseAxwj9u7SOS79RbrLCHHTEjGivhhuqtuPC4cUFqKakDcaLX
JczEuSR5MlN9gcXNPL3YnA8YNN+4l7Zh7ZW3kg3TMel2+VOo+qSeRasui+ePUGgEdW8A7Q3V5Iwr
L0ysTnB1HcB4fUq+MHraG0YNwkvj4JHcUr0ZXyDrWvBhhz8eT+iEENkqUM9QMHHzFkG2Z8gbJ3Mb
nRFBk+POAD+U92qPfL3dwXUmzarqFeH4q5urtCl6faBAq7WWVYYvFlSwNSRlhL57aMvYYOWakgBc
8rBoJH1d+4bfSwLgJGU7dpVuxvSB5EVCXZ3JXf/1T3Ai3ENoHWhAIwf5/uy0JHMIDw9ukJfqokjH
7fYMiBR3/ab8NnwtFuGoz5xYUIYf6S90MWV2Rbh8maysZ/djc6Bltc44wjYbUI/dbj53wRNQT4C5
vU/qPGmGQy0D6WpaA0gXcYVYsBhOqA220UMp5Fqx2p9STl68iQkOZzLMgH0DqQXIq+2VvogpDPYe
tWoOcOHDqcbJsPQkMn9vXLzQ0ap4WwuS9uYPeRHxnCsTqeIQCb7+P4AuM1FIWo4bQOJzeKwWW99a
5bJRHzqwDlpaMhDiVek6oGzBqDzPBq6GSkQEO0R/RjEi65X5ybs+354AvJswo9/OOSyh6esxBHUp
vhwfgygUk/sivxdG3KQxlA7/beCWrSQh0DFjCKAI28YgGvKYXzr0Vf9pjmLFhKC/sELw5Hb1LUiJ
0dvG1UtWNyYhMIQ1XuBvGF3tTUAh8A9hv9A7A53Ht8d1qbq05evn5opkX1yIBxEUKeLWbNPmUg17
3N7GbjcpjLeN35Kg6esoyD8biIY8w1AJl79j5aSA3ROwF3hCuk+ulBWa1kr9Lvz6FOMo/YWeJIjs
SmnUoP8H1SdljxiSpoGsIQJS2V0knbi5f0OJVK8X/mfLsUpU73ULH+rx/abtttxsYO2QOUVPj8Kg
bS4U0FV6+pzmekm5K8xt7Fe+89p4tgIxDNLHQH9dA2OPTKGLZeuqK682lXNEdA8BEZVldkL6yyvU
gxCUVYgSEBg/9yUhyNm4aPddEGAHtyhKom4+K/pyKYh8lqKoAabvDrfBWMboPwVn8BO7A0GLZ2dp
GU2AKFmqY3cHWQZ5c7Q6dVZCk9znaRa3a83VpaoLI0tQchV0Fxc5KSNeQX760lJe9nkqxj2o1uc4
tjSpXxzcO9wVT+J93/JnLMMoudwbHRV95JrVT8SaEFpeE2OOYEOXauY+lT4PoJiXBzspeIiI/O2S
+OUgSjv8mityBESZwuevnaBUT7gdyZ/cMQXRgirh6To+7ddd4H1BP+Uthj/bFXB0T4LlFtyUD7iM
skn6SbzRp9vHujmzMsdtv9RSIvfX95ly/0m2pDnBhoHJv37CE4lGg0nUG03k8GzC9ezWdrRMn1tD
AckWgijAjicossfXvSeWYoWTjMSQ9skK2HpAuEZTxAGgdDq63iyzVk4uO6thRUiAJxih0xWhpX/c
8IYELPRhJ9Rg8foL4q3lgs++q5IVfsvkPjESZhCqS4Ed6gSsqD5X53IMSds0wmsSKYBLdbNV/UX5
wGXNf55Hu/dgE6t/hVLFb0yJ0owqxCa9A9YvqtEVRzMY58tnDau5kLdyvMaXGWfwL/uaCvtDCRq2
NZ+LqNIm1I7l32BMgbVzMLMQxoCcIJhAbxdRllCc30LUkM0M19cFPIABE9HNqtPoy9X0mxa/v4tl
sKDsXMRuZTsN35Iwown8bWHl3sgQe12FbSIvZafyHUazTWDpdAT45ff4K6UveSNQOVLTCSQJOB//
ukopCc4+3Y2Ssy44QC7yPEpJOcUE0Mt0257D8DCyWmTTlR5StihZZu2hdlit7cv0+ZMs8WquQqzI
5WWlWMtPxoZH1CkaZtfrvcUVXzF6K0W8i1qY0ESTVkimIfwEo4SBrOekwXlblIu7VQ75BgGfeqPa
+d+TFGVuYjBD60o54QdZJx+o34senjj2AjMDMcrmtEm9YEoeC2qGgOQK+8aHZT9tMs09xcCi4BXl
3LBH4l/z5f1egx+FkpZm1W3i/7LqxdBsp3pwsI4KllC/R0Qn8wCesbNcWcWZ5dqcPHesumNTeylW
s9bbSQjllNHS1jzroZ7bQC9XXqs4Z2KM9FA5QQFDdA74bYaGnE7pmlkXur3bLb5Gwzz2kK43wkDO
CCBHhmBNaedxsK0lqpquqbCfamnOm8Txi5sWnOzBonIR71D1LHACI2XAdSb6DcTRW3JaxLGf4feC
C8B8hV37j/6hli5iSu/ncdhBf1BBDu6mbZT2mKO15/+9p9eQAB6cmYodqufukOmJqGEzRLoQch0j
GiKgrcpxE2b/YZVot1XQYistKbf1f+VYT1NnR45R6UxMbPgDF0pxxtu6rq2b3PKytd/Xt5TXvEbd
LRgCyX7zgY9FcMpWkOcCAUmJoeKWCK0gLSKxdurYrgUT/wGTQ8VVe28LQfJIAbCd8FWrm6HLRHoE
QA9NeY3UCTlfVkzAAUa+pAWRrahH16iKLZRcUC2iNu7Yh2PfEpevAYVluktScXNqkgrsrVUNtF4T
rfppCO+w4WRop+j2mY1TKvGbTLbO1sgjJY6Ru+svUzLmijZ8JhpEygKcTDzviwqucOXZQPK4fNxQ
2xDRND0D2Cy1DeJj2G4xUPmYLcKjVvWS6efg1Votcm1TJlLXPOwcVE380TeVVWkysI+6b8tB+BT7
fLAKtrtvMJi5uXML99Eq1ZqbNSTIhyz3UpUeAzcdt59E6ftn64lQr+dgh2iCSxWsyg/DHNovacHR
yMCeH1ZeLhEU/rHUVhyTkNQ9NAa1B7xGvm70gdyQ+lspsesnRF2x8T38ytbvN4jnfAAGWqusAvO3
fTrA/bmVzado8MRq50Om2vPtscTaGZ5y6Ej9kuZMQLyZbpjp23TEq+4z/9fMTyipifXB/jt7r6zL
8bxwxWXahIdJHXzJRlXnweT58WwsmvcvNSXo2NaSbTTSH+H3CfVfmYkux58mI8+skWy8matbiQmO
YlNwp/jB9TIdfDTOT5MDeTm8Xp6wrJ8Bykjpo16ULaennEI4dZBTlcLJC1m7668IvGR4Nzzmfc+K
JGhFZ/PT+rcpzeNmFqekGZzQ+YUT+JJRX6L119ipW5YaK34Ya0efueMMbNtWbFIlglkmYUuTleGh
IFfMI4Xs0WF/Md4ehTbc7w2Xb6ZKXjsstysIfK33aKxECd/va5V3lhC6GDJtCf6Lh0Cp9fYwqh0F
wOCzPVjd2ozRQm7lXagzAtNkg6UnqDeDso+rFz00UZzdyeBiv5FTSjqVwEa1O6MUzTBNEPYs1rxL
f17fc4HKygkJXU1TexlH7v65fIxa6rw06+wpreFMVWRm5gkH1khby6T1m8I8Q7Rai756HaUUft1N
uPzDz6PozQ5Rn5h5rP1oPpIdtr0WJPU5A9B6OSeYC3kzLdKujJVjcKHvWo1nUuIC3GUHubx8lQ67
JkGaRSFmRmjb7Rgs+LZspmoWcx6uDiU7nlf+MiIDP5Tzoq1JCX7qXQ4prIKpHNJmbtqFJ+ruosGp
SiJC4XoUM3ffZESRUTGEDcT4W7ORW2ksjCkROuUQ71MiN2G8hxChg1DTQ07dTZ0fcJl6QhZ1WnzZ
uuB3wmF6PhmDUGPAhFdZzAJbdrDM65a/Hnvv3wmHRcHOlbPwsTxROARUaVgW07azAt6evlH2kNlP
xFvqWf/FvPfvQKRH+Zlkkh26cdi1ykfM+GaZvnwFa0IZ7BJScW/DUvjbn3vcflCl0fTyraUzt3V7
GCl3GBBwVB0zAyTZ8vFPySo3GvlnM7gKxVCn9sLkLZnlFVjPM9h+ULP7ZQeRSVP0ftaQS7FEVeaA
Fr0484NhEfu9Ni29l43BeTQNXIhtwvWxTchQf/Ks1HqFPB02RPQ428N+tuuml/lW/qDGk5S9LxgW
8KKbQ709ZLRN0HQD0Q3Ao5RWqLZ2e8ucYpxuC2bBrpZwRjMcQw92ROqV47ciUBiF2qzeU71r4FLn
uIr7nObMli6v9M99My9lYMzXkYlm8uyDS9C1u7dTXacD6Kt8wB/VGHrPI8arlvQOV+g5Mi+CNtW1
X48egQeNhUSo8VaCTxjQhaWGfmfPdv5cywB4LEkCeVAuJeuRsYOtG2AIxNiCCX2xrfjocIJ+Akbj
M6RRHJkn2YH9WeGrCtOb7QrtXdTisuQjwvw9d1r3AQJzr1D9RAJyHYzdCHWCZjEBqVDCGWiqUoRo
QUySDtt5baI/N14XBbi/nzyvqwnxFqLmZUhBu03Ps2+/ZNeKzqVoDQrnkh/LQ1muciEIf9VZ0MQG
0LJmBj5RhwtIie8qAJE6cUoNkmCHXSOtbk93alNo2ZxLAr6u6pk1RHjQes/IYSuoxxZ9OcB/Z3Fr
yCKiwUfsO9hVgQ65xLvx5a0JTAK3PcWgoF5NljZnrv4TggqfbbuYiWoqKjFfeosmcVjiBrQR9QKm
ud0jCa/cY1H2ynxkc3z3fXTpn5VTS4DX+jC9VJxQnfhZhMiZ+EgMA+fBbYf1rjcK8r0JxAfkr7a0
V/S4I2m1fXHi5g5XpnN6ur7HJhK0qdwcLkGsigLAWjNSb5H3o3iWtjqCFYdLRo8e7Xp/GI0J72rb
NT+eHLkE+DYNxKPShHuA4ihGOCahybznqtCcrPlPRhKUaUYy8hIKn+Shy44ZynXAaxh0uGYn3N2h
UdX4V7yxC6osdNvMrF4HJxQflW0lHmKHpd3IPXQxmz3giTD7ucHvWo1x3EWRm5gQQ02vYZSIxJdk
JR1j66onHapIait7Kz+mOO7DfQR8u/tXsRlBG6Jk65QqYDDzqsJ5YYOdWm0Z61fnYSrCFhVaum0B
LeIm8eu0aUAbeWC7gNyyGoW+ZVPtzpUfaTbkT3VeKyegC45K4NtCWZJ6YMLNGtT2/6KkTFsAIntc
SuJwTE52WZRWJsSwz9NBMtyY5sTPHyTPydzzrCCYXxgRsGWWy8cA0LqNRr2a4+vNlrYU4GzvpZhB
E2x3Nrh8JDpu5yNhA3UIcUN902g7N4UZbWnstbmbgirN19kyyLdoSfaVREeVZhWDOy88iAuFp+0S
AGLxyYz9i+ZKfo2/Lj8qNMwshYTtKXveoljN9/8rLQdIZA/qyizkbqd03Gu19FUzLRx0lrHsZhDj
7TYyKJf2NXdoZQ9Lvi3rIRU/6e5Ztjws7IIALWRY4K43dWTLdT683fQQ4lv4DD+yxJ+FYQpWh3YU
8+MLGDGk6hJzFHKozMLidP2eydXUDeeR+y+jTj+ua1M/GBnCZa1LPDF6bOli4GOLxOqK+hYz8DFL
IGm0rlJtin1M1kKuZoHph6WQTI2tm9fxn4XIuO58vn6zsy2YzWCqihCnERvs7wKnqg92gDs67tjf
I/mAidEjh0RtmGSc5s6KFSSj3YAgF/QCGENg+IDsRUv7vZRhI4Yy03KCwaEJDyWzK0OmiQ1Zvd4R
ymat9qUrAWCBE7+yu1Gy3Q/VC8RgrtEeTJIbsNsvNZrrADAP+SlFAgL8YbT5BqObHWKWqhcE/NMr
xyqcWpvcTkCD7Np4af0YqiMdTkMOi1Pcak7l/kMHIMiWdwIN5mxe7qO3K7Yafc85HouPL8Rowl+q
cQj4eL9/8Wq0LNXVnLGWrHJwfLbuzjQn5WOaC0BYv9upa2QVY00PI2GYu/02SzM0+EmmkA+MvoKm
mCOGlqlSFsw3mO0scmuZEZkfYv3jWZku0BK7573DTuWxILjoSlg30pKbsb1mj7NfkDuioxl0DkL9
aGIyZ2CPCT/hNns1Z8QaBNTHk3c6Qopy7rrAnSrRdhczG5NdqqEL5MWzd1zzLxKc3pRHMpIkMw8z
+sNx+j1cZvtzS3Kf1Blq/tgybYfk0SwSZpwa+6xlowT7wt9D1q7NJDciOQnc3+56drYpAXDW/jSW
Xuq4SB9P2ZaG8UcO0mIzqIwPqO2lG+6Einx1w+Fmpq0U2Vjed3vtVc3RqVxWOdL91x9crnfzfTrz
ocPw1wAyXil9g/fu5Fp6ZpYhTyNML5KwwpikLjp3gHLi6mwVcp3gjSUeFG7pC/bskxyLbG0zQmgb
qLipYgnPzyJivC2Eli2/Nt7KzpPPv3jXmIkkD+61Trx+DcTx+289HjPcz0IvXSoqrcZaSEdXfO5g
feJmfqKaddfkQ6aYnJTquFyqK8sj0rt/0qpxKoI2IzDr5U7v5aaLeMj94bn0I+By23VredZgGPdJ
q8VVo7FSONYzqPsfNn/6nBSOKKPPXT6e9SST5Ysnq6uhMEcGMRv1tCCfPVSOA96npR0SVOfpLlD+
PgnRH9R/pAFraPek/ylfqLV5itKeORKaWJMiQ3T3ZkMh2+6Zs6h3e7uReaJ5wFLTXk4ZyULa7DvE
fBePLBSOv9qznZdTaCeX6I7Gfw887YsU+YE2kePJaP38JRkOjadwB44hlposH0DqvokXGR1jlRiq
hmJoSxpLoE4gWSWJkiMpbG8F/25TcgDlhs+JDBYcarf3ttWj5dxZnUswlSFzyXFoXy8yBvzCNOWM
Jox6oFn42ff0iCqKsZEYGHdF8ZFvryASp7enbMht0CbhdqXWCKugKkqaPHTdoJOi0e9RIaqLRk/D
Z0K5g/vlFUvfsm6fQivkTptkDPNMDkfMDjbWz/eS2fqDC2uM4n2XU3iO3y8eXZJlU01XA42DXzfz
kYTUB9C5eB84OaaBCnq00UKT73In/sgsX+HoHmaNXTBGDryZAk9Y06CM/EMJJEvXU02muDndyWnR
35WHAmNelrKB5lO7TxJrh4LgQzZgH+Gnfgwo3iR/Tv8Y0vukEqzcgVt20h8eEf4HSvcIYeV4IqUc
7GIFYKjCD3+OOxMxJGjAKXygL+j6jXO7N87mbhAeBD+tc1BSX82VtodSKwaJXTWfJ9GrFYzBSMpG
YesADLvV6NKHKjuDcEXx91YJIwFU9EEK0QoK2TCNJxysZrzcJyn1mwY/l92BsnkKj1RxK8aiB5BF
YvD9WIqW77uSLUtrXga6XhtI/+1rjte/lP66GcwlkkUgsGB9u5yf1rpIvkWYeR/N18X2oYFxphPY
0J6Y6o73MU/2Kok68nGW3xD/DdjqPyLfXQJsXlvamTwcfxnwa3053kbUSyyxE1XfxPVUbe886ycf
BbpDd7SQDLJ1t43U29suK4B84FakGtRzF6ei5CspAVmVG4JEKuy1oBuhrgPLv8iWDTX6t/oncKPa
yGlcw4417ZsFGcKc8kvm9kr33Q/od1/ox+YkuGGnsBnMlNwqY07Q6jky3cFT9BvlZlwQvRhIzgTW
kLQNVb98MLfyHCvaHBIFWYf7CGw8qkx0dYws1YK+TICZeNBE/5auPcZ/ZsBovwju1qRZfpJ4o0yk
ZkKZ/u6r6DNZMlwinUpxZUmj2ahIFjc4o226GVoAzpTPu+r8o+nLLJZ1c00yMYWsqaeq+O6SOVJ+
HTQmLY+mhwsqOEiCIGzc28EaLt4FkTqVCSMAwX1Mlwgy+m/NbWVH0n3moNy8kfPd1mkUt93073K5
UBsU7QwQn6WKpn8nbSmBDu4OFSsnXBzwDQmNNC+zx3hYQe4bYZ4fsAPsnE8EvysrNUr6S5167IZ2
JXaMrorDHL6r6GPsst1kZu+7ou6X3n8PK0hh74MWhUBI5d134Cv5XJ8LKfeRSWvraY5mMXX/0STr
EChgekajRIhJJvmCyFPi9R8XGy0+kF4arnQncMDcCoyrEvdhEufWzLkm0BT/+5DVEevJrmJtPffB
FoNKwu8oKACjwDvNzHeOBXglsDjsAQzORZXWhuSc8uoYoWZCpCQiQQTvD6U+xHvW7AOe4iuBwlB1
kKkeZj3JDOQLNRBzIiz2fdJ/R0iOkP5zOdyfRtr5kA1a9U9b7s/NolLUkNdnAPD+GJ1wwsi1xnq/
VfKwOmfO5lYYRGjGu/9qpO2gbP6tzf+w/3xcMJAdw5rTly1zCraOAhLzq4fYBIusmzwZFVjF0XG7
/3GePNb7/CObBPJFOQsEr/thXE79ENMxOUARyE/8kMC1zX+baw9d6eOb1XuuYyeaTv2ERDyPcma8
EUXLiIS8k5N511cpxuIn2rjZTE3I9WQ1+Cmhal3WrqtyToG0hTPg+kx34w4jZYXe3SSvLg1nlChA
Zr/U7mgoiWZQasGA5qLRcIXJa/1Zk9PDMUA2qmgNmz3le8UZWSu1MmcX305jongy05li5ehI7N9i
i8ft268Ne08Rwuz1aNyD/fFaXtE10K5LlsRjuc104AhXfiF4HCjF8Cj0LDh0Srf6cFEt+WdTLvAE
xxdMFHq4cD38Ib/aPtjy4mjrg/jgC2vDWV+pdnuNLaIKryU4eQtIFS4wJYIDLyxvjn6XEVZtQK47
ikd4owgyxoDAd7j4CAedFvoUpZi6rOKvnYzfsPie80qjTr1G33Yjw/f/IzxHey4uMzV+fO1UlbNT
/d/xODWAJWXtB4ctTAUjhl9mNFuOHErT5pdupiAMnmMCO5mhm+wzvc+WqhJo3Smn2l4GXSz6IIE+
UTfFOHdvfwrcxro4xLfWbymkJIgWT8Pm7vJVVYQb3Ot1OXZOB9oObpkvvEuYEeTR0D9BNfMcIa2M
rEbLcXMXrZHai8A70wAKeg6gJxPMaE0Py3L7Lmfppa8OaLn0XJ8L3bkqGjCUr0pXx3nWnXaeDoTw
keXn8v33FKzI9HNC0IrxJbM2/SWpvMxMbN5J6JlS2h2UiwXek1Gjs4txK8HKFoo2nxRyE4pjUgbK
0PcvaYxBgE7xG/iau/gN0GNTiP6DolS1W8ib1yvEQVfTWf4MqFdkIo2T8+BUQ5Gpl0VsU8FXxJHX
/JlFyZtXEkvw/hENCmrb0Bx6yZMpoayy1qWHvpHkWz2CUQs5wUGLulX63dendxQzUuTdsqAj8fsG
o7OLkaNAZ7/WQMmRSWg6315ANWBjSd0snthpnygQBpZfLiwzY5ZqPDK9Yjg6G2stcDoWh8pw2VaB
3urAi9aRqeAdxkKE5u/2BqnvOifiZlwIolOqy75ThIl+k2gOtzdM0jAFJxSAUl3voyDnmPVrtcyx
/ivpLAAhvxOTjLQpBAC8FGQ45ND8lDI9eau8MTDrlD9Gl8rvpBCOei7hikW5ZMyo3VTlbfiHUT4w
ALjv6r0aKeolWTuesi68pjrY0TkRWdvw0rb8UNIUJHSAUS6QhCUMcIFX/Cljl0vjcQwld5L+nNRD
Cx/0ejCqHSp5KDfSvGG7JeldG0s9iHZM0thhneEQk/H4H3Dlz4SeaOEAvRY0NZhBMpWmK/RGF4gJ
zOKYekRhY2PeE22HKSjgknYjuDQ5A13x6we5D+I5jRrE/k5XTobiZBgmvs5MyrT66Pc2txj+XyMf
TXidU6cQDIYi+8M8s96W6tYXZnI5AeoaTln9/Kc5y85lyj8PZQja/nRRt686hHig6Z9tt51083wU
MmAh1KyWepSVaUAa9BsmKalBEBAP2cS7qOSeqjpPwJxqtrmuOHraVafcuiqfLirz1e0QxZ2lWuRa
kTjc95UwN1vGHCdmUzhVF3h2gDcXDKJwB6Ay8Rerhug9GoKo/B0vHYrFoydenFyw8LTPWzcKENxV
QEzJdygLnF/+pPzdNbypHdSyXsCWwR1c9JR79YVNwWWER1nS7+nRgoh9493Bv8STP102CdxJFPZF
RjlGOfMCyD19687yC6tvXHzHklDFqLxq01WMtCFIvP7SK2ev6aTQBl77c7L+u08UdiFC6SIUlODm
5TBIeuKKpTU8D05/Rrx3BpJPK2WtNvsTzsSAU4VI+9rTKeI+f4wjXSQbI6XQ4hWz7Lq7QEDMplYB
Cr5C1r+9t7kmeVxCw+mGo60oQrXQgjLPJJ5JszUdPaty4WYzs68BchTlFC5Dfewx0FvVyLym66zM
Rhv+mE769zj4JTMatLMfX9cp6y2la25SFYVQbiaOpgW6H3L0eMe+FXadFmXUNPJgJBWZAykv7Dd7
WoqeiuVCdM/HkB155zdaaJNOWK6So7rkZH1KeMm9B6M27MY1KUQ3LYeDvIqAVXfNpAyq4+jf3TFP
TP3OZM1zQh8+5y/3XWZ8enCTWEKyeXk+hx4xyyCmr7mWN8bLR2A2NxCxD4ybnAWlI/opw8r4ezkH
R3EbG+SEM+qtMSiQCLqyiGSX2d3YHuaLmOioibvfi+rfncbz1KN5fUBunMAoQeDzAFhhrborl2Bz
P9p0OQBwpalkYvwuP46WV9JATYH1QduLH95GAQz7sOpgvdyQzQ1kIOChCgfa0qiuMmvfWAOhQX4n
Az/bcyTC+wSqJH74QxKQc0TzTBucMcoPl7kpjloVdtOiGjVUpwGH+KeDfxuMByBboyqaHaFxAQSa
Wt3et5GsT6EbH4dZEMh2Nx1FM3h/Tt0YlzPrjjiOAayc4Nz8ABQnp6Dj2mrNzUyAb+CIhKvVb4rW
V+iFpmg8ctY9WDonqvu8U3O7R5pLuxdypxV+Hw06ols8IplWK1iU6sZeqHQgXWDM7shaxHQrxm6M
NWrU+2G8BCjCmEinD6NRQmVPHRVAL8p3zuRZTM0NpuXUVje0yWzI4V+x7J4UAoAXd1g19ClTQVrk
zeYe+vx43dh2ytxCafWhC1r9ijKR62arnFqhEHIWZTOm89xm2Tv/T3sOtXCi+5C5L3VMODBKrSw0
0iW0fE+ixsTH2y50QkbsAMEAXIGIZGv6PhxtZ79K/KwGsMbfvcK3ic2U3WDoBys1FdlVQziZ6yTV
YXNNEd4SipNhcSKCmadCbLHi54nWfW1vkHV7dzY+HT2HHVpPcVtAs4c1j8pnkRgsiAVrIMnR7QJN
90kHWctb/cbk5ms2G6u9MnDW12645H31vTxOiflNPCQmOkS9fYqLoeXrnVGB6VGn8vDw0sz7Ya10
mejwJPcz3CPojZpKm4L5QffSc6lFdddGR5qvhWj72goAr7b9s/P7AObRVVd8X5uk11IKtlw61aeR
CU4ehXTqgRgwj6TlKZ4TxTD5wAtd5oRFLeJGu0jKd3Ks/+iY4Re71gB65ttuJtxrKBMqKSL86Dxn
LE3p00pj+Hj34/9vCkHEZe8wxkNuR1WIZ/D6eGwvacsab7ztOCtmga8xa76F62eua8E8Wk37QKOY
VeTywwxLQ7HPxrI3YZRgiannxzqw26o8oEhWE7T3RyEI6LjkSULHWv9BWfVhuGT6wtK3m0HalnGB
duTHWm2mnSyMfR8tdlm06eAU4yunD6n9I4bwnpaUmFdldWMZNKtVeEn/Tt9Z9kBD5cDLU0Q3lTj/
jKyWXDrtyhVuIZMQ/svDhwHC6RlU2QZTxSnG7N9vS2GPJRDFc28+27gI/Mc5GXXJoaCg9lXIjYsg
Mmjh71CbUuV77saXUOXZP/h3moAyE1raV5G55EMGS9krMj9vw9YV/4Gywpf9ijZINXPB6eqRYSqi
OywskUf6mWc5pRopuL3ZSZXsI1XwQJmTyth7c/3jWkPZM57Cy/XITjL5vF6IfLEQALqIzD9TTu4F
OsNd5MTSuRfdcNNU3IUb32Iiqp08idijBxJnLzB9zy2tvRm343hQwn3eY+bCLXgWlAxMOakv5BM2
pitcvx8R2KoLI66hUVTtNxrP45Y1ezIYWzZoIL7Fiu1/IX39gD25GfXKScci49SAtR1gA5uBGJs7
Z2dYJpOrClE5gzhVzqDyFOEpcG5IrLdhVHmTTVz0+9xKApgcNfp4dDsJZnqiSh0ozh4reQTpKmNM
WHHGLCxtMNkuP1mF89TbBvOWsVFVcb8Hu2RrZwaCGvDJJG+Hli5jjxs31laXAyTDZuBNXSNc5/G7
5xqFpar0HFT+gFV4LOEWJjO5M8YKtDWCXRYSgpUGWtUW/XwjAvF7XPfMFugPpieKmK9wTpfv/LK8
ec8NCFwT4DXe19pWwvSgRvTRACxQylkp3TVcXi9GS2zCqlTjHFs5UtdFj/SBWSmPlpHgMpqazy1J
J8GLGoPsGOefmBFq4izBBuB8wtoya+KDq6nT8dsoSNgBU4pY0/eZZ0+Ti7Ibyj6gocajxEXPv+r2
5p8lMVDSvI3n6Oyu2CvLplUgtny/YQjrYvSYDLWSH5yKW7oHdovoQqVV2wRShupMJNv7GWASNFL0
u2LCD6Drkdoj48qfntfrkv3VNQbCPfFqzl2ojlIUOiudrBlZMz72u0+prsaFDsCqM8PbWVQf6EVq
WAQkSGVxd0OonC8MTvFvVCSorjkPGaA9y5VrqhiUDsT6uG85cOrenEA2yE8MsvkUnXbmB8DhJLDH
UC5p+px0afdopkK+Qp5FAjaax/eUApDhmFmAR67RvYPDOMfXGS3flSXDrb/thtNEgZYlAr/iX8/d
U7RhPN8QbL0yiN67evNk+eFRPptsO1FDrGwr5QuXJRPFz2bsZj9KVlQNq4wIm8Mr31TmLv9e2RaT
GqNUaVS4VzdIVF7R50hRgOoIzfKHSOf9jQ/hVdNviMz9Ya9X6wCobdp0UxYiCDZCemMHTJJeYPbA
/O6vYQD3mmzKnRrd/ZOweEMFS4cKTp2nIh7+zNRJgS5LCDm9zCc8GZyiWvKTY9FLr5NprFcwhlrr
+tPz1IwstjjHLgiOMkoJwl37tCF13eXepXwfQYDQBypD/6two/TSLfGn+t4FC6AUsW0TJ7uopqPh
6Pgp0QItd8IOLhbSLFqiZN17yMS9kxELs+iPqGPap4Obopj1+Bn/eoteicj92Kx5+sWskiDNlxa0
k3JQfiretM3eGqueyxfywjnOI1nwWnGz/n9s/Lzl4Td/W/Go9G/30UMWC2hQ7al+encvZ47G6ghv
T8ogOVNjCA528C7B6D1udU8AzDe6PJsQd/mTYOaiEthLKV+/KGbCgzmfr0WSNliKLLKYUQtt1/Ya
NC59C6R6Gi0mrUWtTGHSB+A6i686L/YPhIEmN7Qy/IAGy+BpXRFFJZs+6JfMV2u5aOygTnyMC0VI
dzNv3UiHlo0mgVaJHCTEYxwo8v628cNiGTocMkwYdDkXlJqycersE3YsVXeu7lx3NbLOq7qaMZjC
ZY+nQETkDO5nyux/H/TXrEK7a1tp2CiMFfdXWEofsKJgL6Aqys02ix2yNFO11UsKgCIN8alsSqCT
pmyluqYCQjcmonurT9u/hAyjzraWY6+/V5xBAOc4AEJbDDYtXPo9vmo+StU2DgGXOu4BB9HtXeq3
O6tA0Wf2n55AAUDgKCoGYmoDzU0Ss0wXw3WITbSVIyFbkOSSPv+gdc7bERnBKWLs1Mrg5Km/M/Ar
4CEVGmCT2bGv1OOhz8jfCtKlckhyM96lBmngfSt2JJDPI0vsW4sV0xkxRrW4zsek/TivWZhbxAia
NSiqag0yv+1eClMr+ENj3EFPlzhb2TLDlgioEizbC6GrnvGx6MPAkBIslRPGJ2+VJh+1UAMDzL5w
pDF3z1GOX1Ha2WHBrXuAQeFae6IqdEdS1BPuJhh14qMirdNJsOT9QxovhnbY3GeQqFitrP9p9d/L
WDEiCmc8gIpoE74GTqZqar3OWoYL4LXFj2vVc7FKLcWw7n3byBvg5iNmTwqXIF0pXb6NuZgJbnV1
iiar7BSuHCj2pEkNkKCq7nhhRzrOrkDKso7WVL75E0gjdcWBEN8Y3IcZjy673jBLMicZRsWQZw3S
TKvZCJjqcuPrWCeuT2ZRelNDIPvePVILWTKskgcMENNA7xqOcfN6BPCya/Lg0+qpOBCr8175x8Ni
8hsYgs8kOm5f4IzaAQJN5NjfTGWXpWNeK2jGIN6aKuzsFelt4+LuDYM4fOcYbVu6Yj49b3g/F75O
uviccOBmDLm3kVeXjKExlnFxZvK9d+KFygu8tFbQkXxhHZ9Vq4dLgT/PxQsh5DHqvOEnSY9vBnjU
6r/wCh0Ff1h2lnS34/XzDIVSmRmvTbRR6eg0TB9O8TA7g/PvhgUflSl7YRjd6QpXMB+wz7p5P3u7
rseYr6MjRsjgInqfp3rPu7k3QZbaNKTiRW93TPuCIozC5IRwW9RIrrPeLtn5nYhKVoRSX08PXqCG
Jzj+TiMMeeCivUPlhbLVc477d4qth1pvBwMCyzrCPoYj36pPXacuCKRVb87FddeCcG7azHyplqMG
DKRJwTE66Y8yIALn1nrbiNMOMIkqlkh2qNljb9M+WJ0wBxrvZEuGIDAk2xmZh60ccfOoLEItGVF1
r/2PucocAVaZ/qZsEjTQCmQax4tPGD10q/urAhEu3kxW8zjEAjw0VaYfEGpb4BAkWZ/IjG90Avne
tB164CG7g3+MdKNSqC8U/7vRK1LrlWUin0i3UuSjN7TjBP2hLnpPF3dkIrh14HAB663Si2qcPKTm
/77NUcYAyvc1D4G0z7Dzn9gYtJtbe3ey0dhaqCG65QxHAWZVk5c9zM4ghmKFhDowPPYGREMItLcJ
qX7l3tpTEvIZw2OfZRJHoRMg04GKOtxq5+prc4XtI/CASop3qZZyvV7DuvOzPeK+1P/mzljV1PsV
NW0MucJ2vLPkaXbBmomKjlkGr1vcKKc7AAo7u9k2h5gRLB/qtfcD78hm4cveLRpTUT7pVHiZQs1t
8DPnKg+w5DooLehl/Y4DZTyIs8FoIBSfy6dhNcHvXxdHMaysh0V0eldjJ3xa0i5g7jmNJshm5PTI
FkIRfBxuGeH1ZmY+ZUSf4JrTMX/W77/GVgH68e/Z8eSPA7AQS03+RyDrvDgH8qVF6KTnKW1i1/d+
UaH0TaDayraTjPvxoOy0bBNDEFZ5i07mkFeRnW4Ea1vCM3geJ2FnU0Y55MznbOrye44h6KImB0aG
GQyh9oCcwL323RopU1SyLb/gH+F+TEo4wt1capna5HAw0zJ+jOgOOXhDUOQVSAxdHn/b9+KqScoo
MiVKZuo1YpldlRhHir4Caa7SI1Jd3anIcqa0Ka4hAF0fHvtOkBHZGSXL00hQ93rZlFRuuBjBthGz
X0pr1RZfH7GWdy40jpVrwB5LekhY3IFIoXwi8XyzOkTL64hWUozCP8Ae7IfRpb6ILDts18JdSrvF
V2Nq8jGEktF0FMlRzQT79/zg67o4nKyBUYNaRutJo4Bs9Gwoc0bWlYpwBXsCEkgC9Gei9GDCj3OJ
iq20I7VE5ZiGTDpgAh4HpDDvIdENm7fIMCtH+y+PEMMg9o5p4iwcHiy0QvBEtSbjiqu38V9cZV27
bwxPnvVbWQzcmDa15/ZKRmMyaBvqcaVASh8NnvTWiaeOgsU/fUa65K4BtHP7GY/a991dvDl2h3yt
C51c8d0IDeD5bFBEAsK8b+TBXjKi4s53UcieBqS5vBbB4iD8fo8F4hHdVds9zzZjS1IB5aVY1dw1
nt7RKWW0cou0yZzMGdvV1ZrKD7qBXVvwCWnd4sHKQXpnpghjRn6XsRTZuMOScsau2y/F8bEqUC13
5P+Sop80vGXIjrJraB/0/wsnDZYr1sLYgckknyWoS2iCReMROeB9lttnro2Qiqi0usnUVfNpAOvJ
1E659FmKAIrPEBpQrj9M0W1zoSgGWRFBJzc6HcJAI62T5Pcsf2WStWPl5O15hXRjCosoMrIYpzRt
/W4gTsQZFZPW/8iDpClMmOg5VvogJrLYtmSH0zoTaK8jxTE5nVWkLaUrcsi85UW2bqO9C4Mc+NXm
XPPcZlM8FRLBQgz3Lexb0+QLotp5YVY6fs6qKFSpS0HD85vd6dDmqF6xc0fw3gizD5BBdQqhkiFm
8wL9dx1guLDKeYGcsQocrzuZjFJX6Z6rqQ2xDIuOCXrpb/xTUzFYl0knFz+BxsU/EpbNdONJ7FJg
S87JOa38FjPOKIvWqGZsYJnOQOoc/PuxZHU+51oJdo6M3NayX2ZgpC+p1QUtygyTXoQ/e0fXuTpP
u2JQDKWZNolaJBR69o8rudk3q53luOJIGmQO7vQkm6a9VhLDJG/s/Zaf6BXcChDDll72jmj7naKX
td/0GN/4018pYImsGpzwwzx/VdFPr6uTiwRiJxln94xVmMJtKk1sK/gurMNnc5r16/4Rm88MdYkv
NcVWJ32BZLJOEm1KStPMlafEUk/lLo7iV1Ot97rapINOs9x7kG+2c8ahx1oRfRts26hFWUWFTAqj
KKOljTtC9MDCghhSidk4Z7DovDpmEbhU5DclEAC+DQZ08HY50/NDqu/GRaDjkwa4eSMgD2HJfiJi
LvjrQIU3DoOdMVNy1IQjYcmHlraBaWdpQ12w0mYB0MpdTrJtJ1eS9+YgNU+SIeyDZWr4wZ0qwN+e
Yf6N9V3TufhhwFTl/B0tROLiR9RwElivBt02GaGmOc74eRIUJUMkOmVxItQRIvG43N1sMNwTi4eT
ufFGoUUABG3JSkrpw/SVHtQtaUJwdmzIRByQiAv8kzdCt4/Wkb3IIqm2/EhBwtsYZlTqu72G+j/o
66SoTcFTdnIcoItzFTg0LpXqG+3M79N/9Mb3jYjo2TfSyyurJ2PtuZyx3CMrXCSANXcA11X+A+vb
LQbyJP0sT6mF6mKWY/YvZHFTHCMRJpBtAXYJ96xjIcjDnAqNrlZIDd7Jl2X0M3yvbmGCKCZo9wqB
fecNhtFY1sZe4DCYfKI2uUSTO66k/MB/WVDtdXSEGXNcgW/5r6brlf9w7fJArU7PkgGi4wWKCBru
FsfenoPxEKT5GnIM06/EfbMw0ZXXej9yE8zYMxnZnqNXTQGqH4G9T/tosTVyt2lvB5Yf7Dg3Ct8i
sYv0D2NO7xEY3rum4UFpffdKhXomuv2KBOVIzlqbiGBte7JXskv8sM23RRpVyGUdXPOZSDyeG5wU
hy/GjfoUuVkc/7vAtkx+tYjkbfkcIk2eDpWlGBB7Dnhy/KWQjuYsrW4bDByJMQdAZ+CJ7qIDyE71
W2H1V2MrYLSd6FTYZHGWZZ3IeUV+viVlaKkp+MLkM0Rwp6ZvIC85a7MjaBsWblHkvpk2aO7airAW
WMxmI47mEmiPuz5n2kRQx4CVyFFvyi78EVmkzsbJ3ni1ItITQJbFMNttTvsTV3B0jrXLyVi4pXAV
YbNCEEC+yhOTacOXHApDJtezG7ACnaltBfcjX+XLH13tfG1AyTxm5jSp0n46HODGSZ+ypQ6kEXnk
RLdyEy0jih4hpRyQz5BJtEnFS0owGkVfjv282OyCMGJeTP9+FTC381We/xx+mQgY4R2aSmkTYiEY
4JBfKJaLSHNXEBKak0pXffwDUODhkns77UraJ611txqDxi73cKUt3wedDhyKm1QC4NZR50T8ih8V
KNbUNnjpUqFjRKRo0aSCW8wXvJ3I8PAvWOU+Ry158BpnMfK/bzKW5APVYqVoY0mdzq7XUwJToHnb
Z1lqxAVFhEhjKIG6EiUqOEGPdh555sJBcCImTEhXR2xahIsoAvI78RLib3oOcHUw5JvlaYpLVNna
3srCC1srQM3zfeHpvQd7qYZbMV/InO0VFzMz5aWylvXDVEOlz6MfEZQkHuCZCpbgflD3i1LbyEzn
hIh0YtlKDPi6fRfz8pFpreyhkUO8Wt1gvX00nsVHPHrnEAG7Wh9s1acHcUSUc+JWSTiJRJFd89d6
GI9uUlSkyncogl9aMVmjdJ/xfP+I8kddB2A8EU7CrVfiFGt5wr7oHS2FwzS2iQ1csgO5F2/AgKEw
lnKLTK6hsi9GvTv9FrIY3HbdMLKN6CmdSjcDPGNFJyUVRsRBHrQ3rA3jaljjnBGjq1whMdh5tuIo
3HEtga159RXvj1Mz0WHrsCBXEhraDn1jS5odcgtGxUVoEkQ6ig7Nbw8Cai4IuiJru9F3qBuLo7ve
A40SVGuKxabAHmb4hvtmmTwYWpzROKdRGtaouHZe96i+sjbsax+WIyHzhMXLDDKTrleTn0myqpO5
7tWYuQgxh7mMdudtU4958Dukn0e2m4kwbSMjIWmwQVeL8Zu433Ik01xYoJuJW3+aDJRn4FsjGurL
5tm9BfwGrBWOGY7Y1VgV1l0Q3FnlVMljGTCHSVRFTCcbiWD+m45fmyindxMxmxucKf4fJjytD3cs
GkpOkmF5xgql23JpcBL8+ETN9u0aoPbd6KXc0D20iQ7THEr/51oG6Cnw02AI6EuCokvRcVxoCP0d
i9KOEtBpOdW7QHf0guspLjjnWbdzxPftkzu8Wb71fzCFeFXCWqci00SnNO8sZw7/36Jqo5akbvGY
tyEWu9Fre0U1ah+u05Hlik2ottcHCCFJZvOWvwGi19PvEGx+pBCXw/huCOWNw5Yb9wF2km7Pw4jK
iTpspvnTZqQB7orLnW5NB3FTaArAVdhWjD6PS/1HPPTL22s5bSLnWmcKeMqK6pNci9uRjLILnnvu
RZWRYnohOH7+1LZMnX0uKLL2Ut60HJirNg+g+8oEJ68pUizfZZcNc5pY1zNdjaZa1sqSB7u29jYN
Am8JGocRdOIpPATOpIvnUdIBn7XMoU4xj32dR87+j+zngvFc8Puoz2He6WIkpBOniXZn6IlDnJ+I
o8b/GKGEiY2hHp/EtzfKkPQRvpYD9AQLgxnxlA+K3WgKuu9y0z1Vtc0iysvvkG0FDHyvTxtVDAwm
G1v+p6F3A+M2p0td/flq2O080d1vA5QBcZm6RKd6znJ+1mwj3sjiXHF9jIMcLhPfvAtN68hi+66L
BSNUUep32N9wcZ0kHcGpXJhvRBRnoBb9ABA+tibsu1HISjxE8JJotGPYC2USwQn0zA9kZLDs4McF
6N2TRZ17IVAK0kprgUPNY53q5GXdBmPQCLZeko8+D7KItkJMyVi+fWQibX9LvZd69IlYdnTp/hE6
vjdjB13R1LnBWoqkLemr6RLQ8XKz+k69IY+D/FFb7A2W4CDBrOMx1o78FCBlhCAzD2n9s9rdZ98D
ONYwq1qAPRBgY2zliWMa3stBH3guG1o2UgsqPbZEUVcs9ol4nDbJ9v76ssB1YOAkxm3Zh4My7O2g
qAAFImvc8ymqKwXSk/3CrvhaSBrJc7Er8R/J412Bj8Hd/wPpgT1zcsbcKvwXGuYxFtxLaLiMHpcR
IdSTG1d4wcIADJeh6O2HM2kIbprtUyK3w2TsX0g8wQj3I6L7zO63rmxc9L4zXNcc6xORo7SjiPwr
yZF2hJ3+L6Xf+LdKIZtHvadt+QEGieqnKtk4YYL+taJ0Zb5sxkcZVuvMr7+j1fTlLFWyECKSq4Dn
2Yuq/yDCs4xJFSG+UYhyH2lD9VLQOsbKs+7XtwpHzGFixQXONha5DkuHlj4CabcJow1R5AMCC1YR
TLtuWl23LEWBoar8h0kHtYbHhbD5tLS9VrrmwVFxekfCtwHCcJRQtq7zEJhE1sVC7vMCHOgC/0lB
36GMbhZxvYhImtcjMO4GhuXJnG8p1tXK9V47LzzNrTnuFscaSm9D+Cwr6T8mVeKDURp2fFlFX5UU
Ic9bLm59KlY9VlSObRDvzzAfRetlme/Cb8u5DAWlfzqkqZuXV/nxeiAIeH+wnlziM+3LwCKba2pY
YxSbiVrztP1OPISIiBlHDq6uIObUkMsJe9aGyBmRfoUZsT8mmLI4B8wSx45ufS/92XHzn3Odk2oN
KqhxtHQdvaBrXuafCsoKtIYIOUhChzxeoY2zyp4iT9bVUBX7bxYVwwIMNxiGqciyNyaIWJTyOBrD
zQW0uGqCtbkPH1EG+hTppO/Mwo+3AAt9CMdHoRqbs+uNBZcwWPCnEvAye4zwZN/XaWteUoMpKmtY
W/FokCIb2bKrEO0z2ILOybFVndiDQelolc6uKC898MWs5wrueMJPWorEq4C64E7KePr7n/nMk/ja
D8vO+n+25nFt99qnxyhbtyzpJyLtll0096e7pA9fofMqL/P5H1wpEoKIoramiIj0NKUfSt69bPod
U7pTBp4WcRbWz7uB88A3LBXz5ww9j6q+2T/bWgBH9YZHmTPM7AeTiv959hfRxpn1IqhOws30M/2/
VjZ368y258vt34IL71DzsVuv4IKBi0qdQ9/rUiq0otwDBET13bA2fhq6953s+zITxWCuiP8JiXEG
YsdyInd29MfK14jyNkJ376s+jfXDQ/wxw1I7J/ZXKwNbJkZKTShDme9FeQ3YgA6Epi/ivsTjvLba
CvsER6N3EqJE5kih+/1J2ICuTL5m4QwpydZYwS1mNaPh7grVzvEtqiKXMbEXbcGu8ZmPI2r1DKQL
ldnzooXVpYWocuRV9uZl6wJnOmObkgFrlIduQRkBXc6re05uK9FryoXkSBt6hFpHSqMokQ1HERoV
OdvPahLHZRzsiNkVdiANSbamindQgimbIqu6rrcIGo2KK5FlbXNUhwQaW+HPr8zojlvsGCLtFGAQ
hX3awxef5K0XGz2oB9GwuKp3EOcWG6h7e5RzUIhI1DypcMnONQVJJUjJW/oqwea9jcoSJjFL/kCt
k8JDPU9PY7vIyRnAen3higaW3ZvNoRrhEOfQt9huYGmYkU1qQaR/3UCNWQCRnOJsHE8df7x7vxGO
uMGdV8XW8lWTeKmxV3GO3fguyK0T37n37plG94hbKFAl5kkGR+5hlFs/32zChqPbDTneaPnzVlYV
TWAvSMStyA0ZHO8NIkkIRoHdQiUoA/EZO+f2eMaW3JxEZOI6o7YMLjj/FaSJQgxT5r+8G6xcIT7Y
OqJ2Gm3B8yXLmkXS/Idj1c0Eve+tk4CIY/7DebeMv2lOrLAuLC9kxLpHS3cQSNPuvL13Vb/ramBb
4ur44eETJ/KQGvCcU8n8KXeBF/44lcmLh5PZq98OjEVAkRFdx5Wm4AhCmzjt4AFgycn/d/2Mqg+S
ZlJu2exAy1JFXJbQoQt+2aOoNHlMLsUegcPHTnqaA0k/9BJ0pThpcbfeZ7XnJmnhcZyXNOCUh9/7
lfkbQCbXNPQ5otfm6kgtYBYZpiQ5vyG+MeR4Sk7kEywTYzjZo4cBz5mKfc7s5nrxFkUw+XlUqLnN
7DHzI/dUXzvYwWu93RYF2/uRl1ql61ISZeW2ybaeA0VW5hVGVC6Re5JQK3hxXu8z4IqlNIW//ii7
/9wgmuo8ddInmimgqnJl1LgUMyalMHzN5IUq/FmKCeQ3aG5JrMPEa2u+VKZF9/Mfwe4eRD378BN7
8VtLmebKxw0M4Y/6+9RUdCo1wAojZJh7k8N7REbcNrPuavwfkDGU9dxfQkaI1hXSHrMnGTrKprAY
3K13webCT3ppPERf8dnjUbdVdU/q8B0vOUcXRYc9EQWKw0KyeDWbfXjdKCs8JbroO40rmIYwfkWM
EnnNY5xGRDIPIQohTkNm3BILjl9r0bVOGhbBhj19jGnU8G17TNsFLEiHhEweCyD8KvRDYQoq/ztQ
YlkMpUhnK041lwR0osEsstJChPGPwv/6saJamPum/r++hmzBYu32KB1fTo25NzOBA03f1SXbO0vg
HXk8Yb1YBCSpieDfzGfMyp+r7ajj17THM5hEspV7sBHmHzebMauOlOHrWrrSHwDjcTw37oX3jaBO
39Ot+3+JEOhq3eICpca3+BsVHbbNgEp1cY8OXJfY16rvtzXHvlIU6qLN2yGXEf5WWVmweyC26Jnw
ARPYAc2ewLZNU0sxEWJgLwN9to8Ppb2hCTkxztshLkiQ/OK8sITHn+GY9XR7dBv9W6YVEH+O9BHP
DJnw+XrGdJLNJZvD0JzP1FrLvqF6U+xZn8zt9xGafTtTumW9PDdoOkMgSmUJm+HHpNVP304GT21l
KGiP4BU91bnOO0b/nNg7YR+hqjwCqQpC6NubA7ump3UhOp5Z4JlZgrxKnwUqQEBpnn98yw5/DnmC
BHMRpHuS/uyfZf6IyNvFQ8ALyIGsFTuiFUPC60EEeMQCeMnYY5fg1ftUlkEmM1dDQ5RAWZYvcE4R
ncZDkSrr6VpZdHXbEBaAQvRUgwY2utut0af0s9vKM+sSG+iHPSlR6fQ3bWihae2BT7T1PevKu78Y
q7puzvhnSRiDdGx37itcikz/2Fn8/BPFDDS4heqOcHzYIFezdW2WEgEAJXldEw6PuWbuVFyx74DG
Ib+4JnjQWsttOR9IfcBcBn+XOIX/BwmoRZfbHuJmWVt2yZKyKsWcEyWonKLc0P4LOV+RK6KM+gHI
rTJqzxKG9hh3PlRRDCMxEuVwe2eM5dKfZ9aLA+FtlyCqhbiqVxTusNLpCn1Jwn7FZ6b+tlTzzTUk
qpy6wbmATnHqBYm/WavmgoR+jZ2//Z9Q02VAZrdGVifcsQ0REJ9Zw1dyi5fg4JP2VnyTQtpkGbkr
VJQ9RyGmme0Ih2yd85XnEXe9X958gjkJwTJzrr0/IAYQRgifZ2TIJpCxVWQt34e1AWaYxy56PhYk
cS8a/6N5cTD+4zYdJq4QnTfbHFMJXeuOavxiW1NI5wooLNdPOCtCS7O1X/zOy0YDbA71KxXhAv/L
12hm6WXlngr8DXh50RexmJG2w1blpXBIlKcPshCcbwIAxoKAi1BpIeMhuKeSHyX4KX+JBekuG4h9
cPe2Pyi+CQqdo6jWS/x1c3tbeRCuKi8lWqH/RzeOMcU3YYUqFJAKfbeq5p60QQ9VrwShDvliLqvr
Wc6yEslXEI1ycpvDdPTNv0HB0EEj4CG9zMmLwYtVhs38gQYxqM18ceC8mhjdxVK/DdgsjTfLGswO
tSmG+l108MgvjAS2U7SzSGP1/jNHoR5d9cCz9onUMhCM8SeUW5eJ/vDhbuFwpMVL21EswXVHZcZt
Zwzy3FvJn3GYzLIeahzw7mIk6D3etuGyBtXJzfbYxFgJm/5cOTz+C8Ph1sr2JdUlzod9VPwurDCA
ZeIkyEkCiepli7dlh3WmOTp9KRRAX0VcUi3q6lMUoZQSvG/XFfBYHj/aVm09kfr9hzhQOnPCT13W
2Y2jwGQrPpL6VVikgN1MJlkAbWHJ85BqVe1rQwIexqexj/5ujyQSQXMDMqGFspTkmyJpMjTBnNms
/3VgyDg9zsQftBPNIS/lQQX/6DxbWMW5iXIAT/99ljg0reG21YChIVbxOjRZFon+25APJgwETSni
ToHbVzOrMlcp3nO+2l/CgCr9xFNaUjiomRzlZQ4l0K406Ap2bxRUbsdJFoyA6hH4XHTaJ5irC7ki
bxzPrR4xn+173NkHlaP1xcAPmov8zWTAkl0Yj7paV5WSL6//5RJHD6QHUsrWV/jesKfFK9Lv23zN
Bpt7PLm9r/DfKtvwjH6tHhBChjBF8V5+JaEy+8os6Gx1aCpliGfqWBFYEW86qbIhYfQCPvNPm23J
80iTpvIAoRSN8Uc17Vk4MZYXvWxxVueYlaVD4j2hUZKIxu2gzPs+LnRK6zcYxpeZTDwfII/z35Ts
fvaq5T9o9KYiyxdrN12VrbOHNFaSlDliDHOWdbtT7DhalNYQQ8GLXIvb8f29tocHlpLumjNJUVZ/
eEk/Yp6TIvahQ3PmnK1VTMK2ZxNYMPsuZA7/WNDh9Ca+dx53krEe3Y4IH6U6nEXMEJ/Bs92ifd99
+of+UuNwQmYiFUIJG8+I1WOMvuKACX3Yqd6Ke2oIFtZlrlfRFUlDgZrcAy23DF2DAIXnzsFRAuS7
Cg9l0Fkz4NavrwVj4ixL8GVraGKZFuxAFumcw9tryhwJtimJOL1Fvxg2g3EdKOUZbDnzlaLbdAGb
mgn7ywuebSkTHRFxcpvIbyKrh7hcVDpyHEqHfj1dE8NzWvNyIuCozd6KJ648oBSaAfLlkYBzQzgR
jC25YwTDwOtNvs0Lmytn2PEwCC5oD+Mdwg9GK3qyfKbAugFoancur/FcSHlj3Nx4kR9IO3+t5cvF
tmlXT99mW2yjRb1mIWqmZffZ/oRaaRuenOMcidGeVJpZGTrYaD6Bj+5+x1i2cwt+rjoyOBE9nm+f
fyXomuOdUy0jUrEsaqZzElLGGgMYXqQNcMiW/I4dlQM/bDAKdW0G13niAaaLm4cr66co7T7YPe5Y
r+XVLFFAb7xbnHkdMWXMrDEB6ssuRrPhNJSG9bsaeKuiMfjeJjVqy3GPp3axzEwg3eMlQsPs9sPI
nxEWCNEiFjlindRSf7W6LmtuNTVob+nQjARbYTFWH0Z3JZj2qwE0IHnURkC3mDwWUmq+b2SKmEBj
5bv6oq3VJifAJhcPEkcG/Fav5D/BKZF3x1B3/YfHS4mWlUYCT5/6UYNX7YFz+xDWyhKBi0OfTObL
0vqSm8xVpd8UpE1dkXZhjZQ7jFLbIlG8R8LTwS/p8sG0x+Ro49JoT7oxlSl+yuk6yOnyp68DUFa3
9WCeHSPJWg64HKLdCEn/O7eR/D9rP8tk2aPwrOwjCofKMCxSHAEH06qNcfwlfK4wCU/qmURWGgaK
Qy4d8XCcDmceoOazIj/W0+NEwRnP6AxmxEYL+exaE3BT94fmkN9IUYwfSXmXb34d8TM4QMq3wkzE
M6VHpG3VQULgCexvmAcK8z0AimN/lNVPz4wIQMyABVtTEH6pyldVYO77EFE8XioLV63IOo1ari5x
/pUywZbgDe87h7bQjUGUGP7QaZO5ebyGs7OCNKOUlt/TLZYS6GPRJYlpticF/dOshYilFcrME1AB
ThGEw4GH3TfqUEXWdPAvQ9FbaW5C4bQ4GEJMp2zga3bcfHqCyQxuj+FG19H8Y7bBUyeIr27FUVXg
oksHBu5ViotFFWKCa64sMR2fyXEXIwjy1BLodqQiXB4Hk6v96GmtLzbTTtmBQO4q1Fb2EgaB/BmP
sa05bNmKR/aPgMGHetfeiGk1z2BBqdUoWGVAmORjrGoRgsDRXxtIPSJGLbIQ3H0rqtHf5EJ87fLV
erG6JemDLi8IbfBYdJWdqo2HVsW7x0jekuJI/WIN34BeQE/Ku/EIM3XHG/pyY5DrSryCypX6ncJz
UjXJmVmtlrYFpH9IxhWrX0upYL3G//XWxys+vsnWhK73ctdiUc/pOCFj8wDgGtVgjHScuHJ4CI3L
Iy0MfTuy7lU4yW1JOLIRHewj+hmUHsCkd40aIMiO3nYjO563faFvYNUxWtm10Zvrm3HpHPHQ0x43
eAwnOv7yOqFJmxvVyewjSkFa3yIx5Ips08NbqazqWvTyVSoehT9x8qrqnZmiVjLJFf5yGVnuMffI
fTXsTmyCMtQUlmmeagsKuuETNBtM533Ms63NRycGgQRXEZzGfGM+btmjFBtRUvbgexQ4jtQL3iUf
524xDPVjoWRJVt0fPIf2ene9VkibnMhSt9oDpYAd09Ly45fFjnZ/IgGCiu8xd+hEbbpH5eTq2GuM
mRNAogoJIk12VT2XIGXl9CbaVGSP8V7AYW/5YVuv48Z6QR50CfDKyo0WSpC0TyzBu4qvdTPeCXf5
asWt0amVorUm5pnrtGPuX9byHw4SSriiPlQuBQyznePXAyjLeVmXvddQWh+otJrIubTweN+vTDid
tKr9U8TuCn6q2cIQS3qtvgTZeTbNK37Ock+c33qny96L2fXLiJ5CDz+1h+diuhCxvxR1oKngJByT
PPJOPBUDHRkEIUVubq6LgooqU4hbnEFWAGRV7H8c61rU+/T1rDn9wKS7Fs6G2ctHQXfsRpTlOO13
0t13vD0nn0toN4l2zJW9Yrbr1T9c+BPMhdFQnXA9O0Fk9uOCVwhGOX/LvCADLWMick06VHtZ549U
qQw+HHZ+81rV0GFWBBXvbJEYJUvEvmg7+NGHw4BN2LT8T2XETUPaLEhj+UBnybT+mJKaKp4HXWEK
K5CUU+P/eC9Xy7dKJjtME6/B108hp82p/WWGiyovEhN0yEtk5neUnAI35z5FoC6yJs7ihYLlJtd1
vo3R0r1cNPKonYXscL4Z6hbT1+sxsYMW5Bq5N0SAhhHaTlC2iBP6VZh/diPW/1UIi5ZZL8CT+s3M
iHWJ/8sh+ukT5ObkoTzbGg8pNLrzTsiA62lLavbFE69QJAzMjRjCMXSsbH3LYFs5vo3NJEtS+YAX
E+CCAEprW/bFnvzY8bQKSbpLM64oeMcJ4f74wX6TCurK11qIN0Ipyd0CMQ+b7D22qaSDGZNs8Tta
GmmnxA5gt4wEi+4qsMYgVG1EI/BWaSKKLVVdFi1n/cLUYHdWHMN4Kr0zJgQkeUASHhoef5305/bB
7QEoq3idH4uJh9ZOH9VFqpoyZtI6EqchcjHCiFwdzFYz/tRRPDdW177r5qGoKxgGMKpyCwvAgRTD
xzd45Lr3NV7fcGtiUyhyTYrQJSj2hHP7ST3C9INGg/LAX3j+PcWEt+hVWfq6hhImmhjkmiaD2CmS
glmvE9tPo0N1utfeTFJkVAZYkOCIGKR/vJJNpBbAJI/mZBVx0pzLaOYSAd9FvNO/vFTFivTbzaLB
le8o9CHlCGMaGpnzAIEsv/0O7c1OeCln6dhPfNr9gzrOjV3kYVBNpamZAaZhpfafIF440nBK7gNf
kYeIitaoE2+OtIYpXFirj6QkcRoe9LpXDzdufnbzCodpRjj75JU5f9/xBLHkBYWATGHWUgS2okjy
4bEJuSuDPW71OL7+b9sM3V3z5ZKdVe9up7sP9daExINu2gmrKPC2PBqNGzF7sRQNszF5PXMe3oel
bmcVTQ3OtIbltn8x2+uRICzpu7JUxXCq/R1i/HVVEenb1PrFCBIAmqoRiFciSRMSBRYq2ES8OnHk
qvxmDxqpkFTCjdEd85sKZIRWt1pWWHzGIsMBSkSfQGfcXomrvWdeE8N9C3kuGV7Y590fEsGMuBxC
VwNGR76qQFiOi0JUlBDXoDJ8pGp4DaxiDLa/abrsT5EsWbE+8bhd5gzio7cKD3VmOPXAN9D9o/NZ
fLnxH3jbBf5C/Bkt+Cun8D8idiEJ6uiJN48nJBV+9GLLhqgexGCKGZKa8LEpee3nZgn1/7XDC5VY
uIZUDfV7Xe4LYDGYT4VJYoHlWO+B6uobZZALPzHWlh3pHdEdD/ZtbAJDpc0bazUEfy3s1O9gyM0D
qz8I6SaCnGv+2zcRSgplLAN5aJJJqd6Grt5AymDbGSS3b326sW4Lxq05cHZC6yz0P/N6byzeEEZu
pxxjjk3A8Nipmxtnmmiuk4FixAKSk+58F5J4FDxjfJbFMzrdus64FqZY60VJBZyvLJKLmvxmC9MF
UUeywuHhmcL84NWFtUqOXOUTsWrA1EHIU/BH/cSeTmvc/57/AR+ebS2TTPGrwzeMul03UMrUr02o
NtyxpqkpMUwG2c9qsfAKpk0EicMDhD0ACmsOyfILdfvMLsbmVcw+JsRsfnVyEJ09oVk038RSvVyq
FJqkcJUBNNr/KqXaGbKzocvoI2S1e/MVfgmi3VNKHw2qPJTJDsQGWpoUEEmGMrBOutlr0RpZ66Ov
xUb/UcXl8AZWAq4jmpKPxJ9cDEoAlQVQjwSvrY5GU61p0lpwlM3IdKoQgwi5I+rYP5KmHJYvNLPE
itzb0X/M2UDR3IQq2t8nc4lD7/bo6nLk18ut2lx/aG4qJmaA0qwYybO6xPB/m0Z78CI80fMl3Pm5
emImhoFwfgP4anqJzLPC5i1sruhrSB3ADuMHWFrfM21x6nIgpOfqemtwX6GY+UgiqQEe2WoCbyrB
dx03A9NE9f+SFJNo/Ylq1OadRtc2Y/A+4QkCYIhbMaRh2vtVPs9wqh4HHC4VhSrOPhC12rmEjdSP
J8uICWctxnmQpeLtzQfnRoe962z7kYIenjGd0cZiD2Tg4TLMJUKzW5z9QaO/OP1A23mC3IXOA/9t
2HoVNoqWU2CBJZgo1r+I6zrbWsSu502uL0fIZ1QhVf1QGUopK8HLiazBTPrEJCVZ8yo/NaL+o6Fg
51GPJs5ApaRWqSrLy1fGB8U3cjtuxh5Nxp7ZrSu5Ar6WGiu1wJjfwYQCbic8n6j/sgpLjGpv4SuN
QefgeKzqL/RLwG3Zljr1w+lu9UHzkCHGiu9UFS6bUbwoLt4fV/lElngfEZH4Jx551nUsX+0LDtZ1
w6oRxgCLdh80znRg/NYKLt23OaB6YivbhMefyUgoCoHsKAJC9tnhg4Rzn6UUGZ21JUZ3ozbEX8hR
wpg++/ovCp7rwG+Vke4tMofHfNPSX5xyalYdNrUUtCF1iftvZ61v56UyVTHGc9RgB4Tu2cOSiWAc
91pw6Z2SUziTVgfAlfz9Dvm112ttDV985N5YA9lzb40CH5I+YwYJQc5+Qgur7r5wYD9zJiJM+v4i
z4XBa3Io/qiZl9zizer2OXel955l5YW8V9iS/dtOqCqmv9bOoaLXFWeQo5sPsoyC/6GMMcOy0YCT
nl3AUJwuZ/rGauHkB5pcYZJHnjgm/pwmu2szsnQZwNAWNq/y14hw4n8sr1ktreY4GCdTYpUPDXEZ
rHTpXMRV5I5ETf5EPCOjIQxHV99q4ifZvGI1JbMueBzaqaK/tLEmi1qfzdE7yUEyWPFhcXFITlGP
OO3WMecz14Tb/MtzwEvGzdMd0JiQXQpT4s121vwzm6payesPNf/B2G9+iAH9JXhCESUZCUaqyjqU
bfHOBNziqCAQIR1YpJ2fRpsjVJt6QNILl8u9OXHBVWE6t6PLUVA8zyTX2zGHHleVJATj14vSbCAP
qS4fF+rhjPEyqiT7OOJfAnNY7QHL7+e1k68e6rFgkiI2DlmpUTCq2iv5DH0A2GlOcMXBvckRm8Uf
cLISiRHUFk9kP2vVLbHMCDYQT5Ebbb7mhavRilCCqsu2jcWPfqAr9IXu0duSTf0LqS1yJt9UDHt0
pO1/NyuKvUIvxmRF/gqOX7au8UbPEtxhoRSWJ+OMx/+Ljdb6gSouee0CuWHqJQcWF073+HNs47TP
Zcgcs4n8lugqop1FEBiBkbrphOglwuQcZj1vsYh9jV7bfoctrjlSVoIX6/mg7rMplS+t+XfjJPVm
abdKmTYyKFGso+Xo6Ix2l6GMsQ46rAF3vOcdYTiqAOCEsDhzTAwPMSuKFaeC57beYVlLcyaxNy+/
FcWiuMaKGmUTJ54SB5OwBz2mR+/7a77g2tRLtJ7vH54iBxzQqyfpLeYO4Kt3HGw1+BJlJsoEdRbu
6jA54gZxfOnINU1P7Tp/0dZY6WsKYRnQMUpy/V0vH9DhcU9yFu3vFpCEzVsAb3ePN1/e96fvqN6F
Q6ekU6dAEWpYzjfRO+9Zeo+nTTeAb8dm9TgwB2VnBpLG5MAWdLAK1Ii2zJsct/Y6Ioez1Do52FBm
2SHKRKeyJv269BeOUsIWMMJXhuIIbNKli3M2rntpYT3dlvZHJsUldBm/clTTbo+HH/VZmFh0PhpG
Ry/bVNMEz9j3wq5vfim+fQlMtdA3VCvw+UA8xxKmOs/vEO7TsBeuBxswgzYczIR0Vkv9wFXYtvME
Pw+STeoma5XKLa4cdACJEjpYFH8QNk4vKKS2jGtWKI+R2nmwpb6XZdtfFgCZi9enUPKoqhjxtpCJ
FCciGRcP8JmdpYw6YCkc12QfBszGrH8THjHUQhAhkunBsB5N/Af+t/BL19ulTcpUrHa2H4+r8x3Z
Vv+n6Df7tg1rOJHQhNbPpsTt8NTcfuZOnuXHBSxMnClfkvvfutL4Z5frH99+vYhm0ey5TtpD+tp5
aISojgxWy3jGbqSz7efwW8zpNITDRF02J6v4do55Q2kBzxLpRIbr6el14XRXD1RZngYlfAjFvPBq
YmcjXdtmn8oDTS/lioW3Z4Vruk+JeenhQSyerSbyUCwVsi/s9a09UsQNggc47J970n4tGVnn0mUH
le/VsZE4qUwhNx15Mk2qlown6ZUbvVnNceI+MpoUeXGVVYDv9whERvjPUOLOwIkNnS2piJF4uE2Y
eSJBnWW+jgMgeITKlDAAZ6a3QZFR2N+urIV/tU9YrOSeOeIgjr8MhxYBqAPrVOLmrjVHmatV1Qw8
uqKXYrQkiI/hBX/yKBsWwJxJTWss68w+9O3aWUIVKIeqsehbhFEpwKiB2vya2zqzSSsc7tN4YN2i
XW0+aegwrDLdQhqQcJF5Al6kzYeywi2kMhO60fnEPu3RtbR18ZL/1XmYF3hhVTmzQyzA/dXodaSd
di53/YYxzrO53OCiQYuWmPzRbvWn+3Pw8DV8qyFlI9DWQyF/EzWbhkT4ukyrn+xz8io0fpoHnOYJ
ob6suVr5yvCaNUSE5eyfByIFL5md+EvBDbjf66PNS2uXfvbw32SdZsMklVNTlaE5RaOe43Y9j6wp
j+n8FA4dojXXjUHc9Y/ixfoTDk50snFh8r9TWXXqC+o1hceMJvXrcKVtkXSV01lum1d+ZeqWf3Ih
PEI1EVMtUi4QgykuUEeZFM9pAuczT5nQjgIktnkaD3UFViWGzvDD/rPwwvPyDfQVXiT8qQxt9h83
nz/3Eg1gLFAdD9R6ULrCCU1+GD7L/A5GXRxvpusLkp6++SndCEtA7HWuYcL74buLdfjdzWsuEDee
luB/B0EAatuhmOcfw4Hbhto7J8NjR5q+tsOU4Wa07d5y3uziMH5hDThJUO3QMEL02zbHiWT6a5GG
Y35E1W2zIa3yJBAwVfKliYlp9qpFeJe1JMfTfNdq3PZg4YjUVI/PxaJcCNfNnZNr0EYspJclZHtD
2is/c32RX72n5aNW9BEUtee19PjnnTgLE1YyrfSCTq2Y3quAfga7zxUjV15n3OizVlRCiQomjSBj
mjYObsiSEQKr48REHXWA7bJRuxsx4kAOsI1ETzU6csiW3IBX2Tu6RnYAAJZCx55DKqmIFGSR+9E1
AL/+IDr31V/7tQXiM6Yxqx279m9bftxutxkLFwe7mXCqbpj9OSj/yUrzcx9TmoV4ymZFDUImiGAM
VI7+NhAWb4cV6lSBNJJp0URAeEb2MDEyk58zuWPLBFQ7hbK5a2lA/LdRwHYIFmATE9jf/Gg1Abk7
VS2MIzGziAxCRTZM4vdX+vH24rmr+TV4zjxhWQIvdE7v9YoYnBy5J61DYgGDk4OIgpEHpamZvmLC
wJH9hit8ZTdUqm0NqoEI2R5rhswZPeWXbbFC11d0sxaq6Nstmip0EFUy0GJym9M5iTUz16rJIQ4j
CSJKZTeViIQb0ZRJJbV5p0a6/XAc1ERpvT1xf7plCBgNUql62bmVVj3gaMzr7an+GIwbldY4xFlm
6JVWGtyH1WNk2sn2gxoOJVZtXrcTFKN/QOa0zWA8NSXk7z+daw9MbNUOieSRWYGjTLKGkx3aqJcm
mDbebT6DZQGKey/ilhVyE58FXJUI0WKnCEKx3HpBGbQ+3VvjJvHT6ozXmfw1+yTLZjWa+QHMePkn
urt2TDOf91M0uMraKH0qbr1aWTe5jsjQ89Bwxf4g28x9ZrGofiUuqhytuHm8NthDI4258g8MloOb
1QJwPeK96k+8L5tikqFlqYfNhKos+HAInYgIlhavkQ17mYEzIgOlmbt0pV5j5CyLQw0TPhQ7NiZ1
pn08t0Tqt/LctTKy8PFcNERD8wJX8FIaYoDPDKkrGUfz8ArWJNdax3p1grR8h9cjGRv8Es/PZ3FI
EOWLWZQ4Wx620Q4tkBPqfk/QWeJwT/4WBfqj7YxS3m2FSKL3MeLYO/vBzU1dSf4ORFIO39oEZu1Y
EaE7l4f9PmeyNbXzuAp13fwU7jvllC0VLogBgwujZlRH+j//ShNw9by37d+DSkEnqSVdx196G27A
iYdRrKelSLTVdTb46mDKXCOY/iBXdM8y0DZJkdTXL0Q4doAWEwJGCAESudTBZMx1Rv9igMA1E7IF
8KHeVnnEIiDbDJO+276QJSkbHSn7yEGTiKhMzsQINZdQnjtTpgQMyEEHjNGBst006erYaVvtUZNr
EhPsw+V0vcdhmlK98ELXiFB2JiEdbbrWEBiIvKevpuii8WEFZ5wgC5hGFRpTQy670x208zc0QhXI
wJEzC4hrx7TYVjyYIdqh6YCpMqMrM9mkupfEWLB/n6+bNjU4UAceYKJ7cOo2+/TzJsPe8gq221N5
3CPEQgLv+9fE8YLpbJVN9/X+vAl7K/fuezSGhFEW8jyggSzUiEYNF8eJ0zYaXoZb66Sr6rZGlUf1
qfUu44AWFbrcKFGW/VAL2akXgrMMfZpbunGaIwNZi+1nNZdItJ0J3OfWKOTYMkx+Nt5gSRjXLTfL
yAOjLGfQKOjUwYwAG64EeU2IpWeBgA90l7gjHWmsZjQCBPMwXUC7OxeQb3Rx+oLOb9hK5xg6Oxw0
cHjyd6rpSVtwvA8wLKLLW6BmMdh+HuumpUry2uXxjZjp+BUjika3fD1cM7FYjvmm78UcaNuzDl7m
XI6mTHhssPh5IbomU8TmskvBTrtNXVine62z41Ehuv6fhYZMon0zvOCFbrvmlmZu9/9HfUFRlz7y
MUh2MYalRHgr0KHjkC++OU7wTVVNxfwsNHtWlThxCSgIinl5MyIqPi+gU0wRrBmx1douqoTNqi7G
TpSrFFF7xhNx6jgJOItrUCmn1ylOfE2Qbvk5o0F9/f1CXP0OGeW2TU8pzmmpvjR3gHasLfwaK1mZ
EZjSXCCsvBNr3C1LnPSKSJqtXtfaf3cPreHjIjx/QU+HxTGDDq2ddtL8KJpgKIV6cJYoU55IKiVY
7zhsQG5itfBF3RJ9+zNfZ4+/bpwD/1ATggTKW4/PgMEILphl5beL/oNN6v4TN86XOXXUtLnyTsbv
CrQ0kJ4jhGMuTQI7CzDx6wPH4WQg9lCbJLKuU13CClLi6gOW0Q3Q2KTdmH9vtTp8vYlsEMEaKUej
y5bB7MBbw4D+Z91tjtJj1eQ7kzUOjv1D57cmVNWdpSq1dVBbqalqZUOEgA7VoJGW7T/9GphMkrd9
jtakMQKspf7XDYWUeqzi0nPMMMTt/eJygE7Lxl/+znSB4mPaACRTGVJTVzoGmTCIZC4eEpVIbljt
EVs4CaRbtuD1MDAPREKLi74X4XhRSUv00ZworohXWjJmFPKwHXPpjulZDeojXFQO2NujIlKsCFCA
vaTh+f4cZNTvBvWoHCwyPZ46B/XzLC4OiRw3We7JC7jgqoMh1B+wMHn/ChCswHCzU3gE8sqSIB5E
GozYI4LskAWJq8NZ+mbBNMhn19KmyHDDCx3ILexEqsueRMSTd0S0q8057BLu2lYzxDPn8ziCTi7t
0pF3dxx66LYJTop3vxuOcCAJ2QFeC4nivurWnB7nGAnYuCzcyQzIjvbRt2DEIG8ddOxA6vQ3rhxX
yv/w8Tx0vcti/9KErdQsYyUVonWtDlWoROEwmbkBJs+P02sYAEHtzl9HEupXUebzT/xrAVAxxvs5
zcYwrF0GtAAve7950cEY9oU90sB2ehtpYzpiSSm6l5EL4ru7oRO8M880bstM/IaD6JIXL8C4eHve
i88LR87uGyqT0oJGr9zpkHqI/vR65pmiNPfIoSfQr15V0sm6IZ8+VUjTiGl4wGhx/0qBD9r2By9I
BDlSfFjPcyvu2CTHoegZmou6zCxzk9lVjOMZjS05WGl/j4RWjm+ILmTuxak4lwY4MNFwmNnPt0k/
HIK/wkjZWyFzPJ2nlFLLxUjaYeFKRureQbYNi+Q0dAt2LNpOOcr96Tl8ldXGeNVAoGWwfiS6JoHd
13THrM6f0oQ788U1EvItBQZJUDUAQRzhVyHNkGHnIeXJmP+CsOrgR4W/oG2vay4fjqyA5ynRTZ5f
Wy+1Bg7NPvDK9vyR9ogkOd3mZJJhy7Zm1hxsrzCU3VfNqfL8i8tntWKvi8KGDLSGcR2SZjfQVCpk
cTMzxxLjV0oNBFZkAXW0lllHXSmo+QdNleHP1//nbOz6ScWSgmF6yAX7uqDMAVnLh7MlhCx9TbCY
xpVx22/elMELkSRT8mKCGMMnZ3C3bUDN+XSKx9B9IioI5Swk4+9fIcWDJ2K+hbfGZ3/A8wdJyi9F
ADZp5mW6vvFhtH422m5tMj8zRKsZdid1l2zVyxUm757X2AAH6lgBA1kAJI5FA7K/EBuh4NqcJT0y
7KLxQzhxArqyodpMj2rp8TVj9v2kL/kLe0si9Hd+9HH3jEkn8jaoD1/H9CNk8jcg1Ui6vmdpyW31
WlAs6kW0i0hBclrtHNtxZeITR+t9lLpsamUHVV9P1Ha3bQwphVaCIfzJxwZlC+Dl94o2Rk1CbJ1S
haBXPagoi3nEs6SfW8l/kDlDTbrT4MKWrrjgeR0RCUvTX/ukQLDmYwOKp8pZxb/iE5vqTKRyQ0yP
Qt+WrfOMMILnkwds+C3TCxOGabtFNFBiX873qS+kPkqVQUdzd9+OlbZQDdfYdPl/f6DWqYQLpfQs
6LJQwiOTZqaOGGaYadtfI+FxkovOidbaBpc9PHkIK0o7jkTB6ryRp3JcXzhEekNLoEbrdyhrcqPR
f0ivjz1qAeKI/TPyABx8q9qg0PUZS0aFxOwAro0anENFv2HWM3bmZrU9Cqo+zbld7RqeH9s8CWEo
7dsZfNtPVc7PUZz57RQihXr3jCD3F25dK7zq07ojB4xNaFH4A6tzpp+TJVZZreEPrNmprkwzVhb0
JzaMSnQGegh5oDqpyI1nclhwtlRJ+eFZ1o5MJtMiZyzvAA09/gQQLl8ECaFWPwtAHwnR6KLMIu4r
agP8SdupIGXA7exYWrWmWTnXPMJsaqjMLQN4X3a6dGa02+8iDa+Yx0ISyzAtNndedD21o+09sxjt
prx96xFbiZPzrmbunB1ScGr7eltiKcpAdIui+qyZQBx2TNODRqWg3cCjVGUROMjg0hAuQG11WSGZ
Jcrwf9DQ9hqTUiiwyWTYutpbGhgK+TX9R9oyv9tufoozSua0WPqB+QGjpWJ9WSPE7a/CBMPgtA4b
KxEOB9ovl9sA8snrFYbnOlxbEhcQOO0QEg+VxZpKlKYw7eJaJ53cN1qCMrmDacvN5wDKNO6iQ7jZ
fN8J6oEOhNGkCZYJFvE85gv5F1hLQ2eziTMCUiSlqUOgS4NhLP9H6Fv+5NGFou1C898ZxgWeWh06
SNgGi6gmmg1y6SoijkPYl3LRfiexzkxrgvoEDP36jROMnwOlXzNVkwrlMQjZkkghXdVpwfLT5JPX
ODVMJ1So/uHknlMe8LyzDUoPuWlVi63eMmtJHvIdznNOEcF7xQfLrqSFEyN93/yA0pewz0lYEb1z
4mTKuHOVFhfrMt1d9uNRj6Ej8HtNVTpDqDfmDmoJsdfYi1EdmH0wtGokSlqHesbVdB59UXRbsZ5e
r62eP+nKaMR4s/Q2jWaP+ltB+2q48YirCcs7uTO3bsbKdgz5Wbihc/d/YysJK+Ui1K2DyW2DDDeF
Csouj+ST8hUNb69P33BvOF93DGW498sXnWcNtkn1Hjl7r+HRWnEFgOIQ0he/86MuZBAJHxBKP0UZ
qHfhNyqVl9BJNsa7d27mLyTQEs3HcFk71XoL2bwkr8WhY2+YU08oAAxV2L/zLf4zSzq4qbV33lqa
kXdPDVCuHp4QwVoUTK4VVz5ePZ11wtmTwfIxS13AfH5YarQu5rQFZ5LvrUsRDID8omTLXPWKVfju
vbJUD81CroEViEnvsvMBIKsPacKiZ1X4UKx5nlg/7M6dHeMEJ6sWjmDfO47e2SwzeXrBD67mnKzW
xG5QDCv4rTXPIaOuGYZ+z7vd4AQKnINvR4r578d5UpnH6Ecm4EU443HnzNl54m2ekjzDlUVzAQkR
Woo6+BA37l5Qz+VS0vBEhlffbIuwKCesX581T9jC52HbgTPu1sD+1dDLA8dr7Bprj9M5E6v1iui8
RASpVxnNGJtMis6ZkyKVpbq/BriU+zIljS8n8g6vJJ7U4VQ5yDSmu+JqI3Ep5Ho5Yo00CwgmahbL
abJam9A+MbSWTgw00XHefW7AcRyyRUEinLSxdSmMHtzEhNxsxT/3pue1A3nuqlSbjxoT6ZQUEOh8
8q/jad4AJ6DtzJ7+bNjMR1hoFyUhFlY/bhj6n0dS+TjB9bReeVfFA9nDdn3DEF4fXM8PuxqeY2P+
STiIE+En29Ht8RnPryLIKtxYi0UlsFLFHypuscLzt8vhO7I/2kD2ph0NGiCNsddjw1zyFbsyhxC/
elryyNQTZWj+O8hpF2pY7StIw+Opfm9VmGZPiYKLiAAfl/yNo6NRHSP2Mfb4XgHbfLShuRUISQ9d
HqCm760oUI4EKG3TRP7roJxAw5RO4D3r+eCdh+s0xCeFV6vjpziO/xrkElsF5LRwfIH5BBYnAplx
VzKI1b+A7d0v9ffhINYN2UM4IVNLRpcPUC7yBhbwxAqbLxwQVQ6IN0fr2Td3ENuB5OuwSdw4LlKC
3x3mym9MWtGNfU3G3D5E/MkaPUboG7rOyIT9KBKizdCbPqemDkxnMdFATtJxjuurr4Qq8kyAquk+
ymeYIDqzCSPkHMR5u3MKUWib5a3Fuyte96Y72o+Hb+sOAMiryR09CzWYefhfk4fx3kMBfjJps3lw
IDU409n2rvXsR5grdcmpTAjjRKB1yfKjVrSIpYg9K+GQfcucupzS8eKrAU85BBOC0fmQp9/jqUcN
1eKUCW15JZgsMtoJsec99Nh8P/brZgt7/eoPTFx+HJYdMhvR9k7o8NywmpFrhL9c2qjLbYmPlzdn
WUVk+9XESLuFMKfj9f0taExJaZi97+SXF/N09DNYgzCsxXaxZ678dXCA7R69ch7KA1qOieroCYLB
UNzd/+3JbINdHxOgqiaM+6p8sXGM8EwmBTpj5q4ZJ58aQo4F82reOeSsIgzBykd69L67enzAWZBT
iLM4m9VosFymWLhBw940ZE97rlFlhhMSq07vuCwncuYdKzCXTiqJeuyObpSX/x9ye2+TjBMGP42Y
2w5ejQOzsO+lOcZ5PN6M7yiteC8lM9fbqoBvJhwJlWfgiSZCDF9JFhbqzta+eorOeoiBPK3Gyr9p
a5luZvl5D0yjaMH+K/cF5+22wQ/OpuOSyVHuO12Dbvll7O8J9oJDfCgbJM/69TaisA9BhyA/Ypb3
xvg6g2VnrqH5k/BNI2bH5v+U53jS1pNyyQ3jsX49XKuQisbJPNC1G5Q/EZX9mZEiG9jZ0zQPiVpn
oeD2Jz4/vbJ9pwh+JYOvZNmuxGIiE/ZSylkrWIZD1KPdKlwohZCja67Foo+qMiNbAgRBHHWFOOKs
H5sQXVRAzoVHZ8f7HbpQ6ZXDfVgDty8xIANbmFHnPz6c0VAkkNt1W4B5eR5XYp1Jhi2niTPDqF9Z
1Lm8ff91vo+MhiK+QHWYvneiv0446oDqLej8NRaO0Xi7A3eulZn1Ag/u/kTR/xczpEDv0mW0IS31
y+31bOr8lV81Bj5UnVzprQnHAd1gGzZQHpS5KHU5VABcvUCJ3oG8qPDjyJ7X73/+NKUKbfrRW0Ie
ErgSjzs9hTIv0xDAhyEBirUKUQGj173zg0wqyYX2tKU/opz13LZiYaLGCcbslI0m2/u426AfGbMb
YdVcIalh7tTR60WWSY+cvFR7PdXdvRKa5TYoUWeCPfPozQvLLLdFzh0VmU2kVT+q+oHbh3//Re7R
xYUZKZLyW5Z71DjK9wt4JaX7U6AdxD0ZBK8I33W3XBZi8YIAUkM7kWuXCVDMaOesYPa0Fvw2xwxo
ZoVamGBj4maD4IIiF9WG+TeJLN5cBxDsQoc//uMb0GKMmp4KOe7Utz9wRaZ8fvB0HUPYaZRgLgPh
tMP0BiRlZcnHL5jMW12yLCAJIUh+qiMW0A7Vx94x2yOhwW27BR8DCmG446Ky74Mu7cmlTy0fN71E
bvRBqHPHOAxK1tk3UNETV+VnA2CYt0AKc97Ttb3+kximrFhqBqFc1gHGjPi/B7DN0WiShzvFAuJB
I9D2X9iDG7F6Dq1K6BDngd0sRCI8lJblGz06JA++Rldl4Ymuce1796zhkFnzRiRQmCCIe6jy0qed
s+G/Tec9CmS0ZLA/bQnMEsF4kkFoBO2xfE5t7DXb01ljCLKLo46vYDm6ZrD5C2DwBxFjqe6jHz6Y
iFtbORuEFAgJ8vCVJPezlPzX5+RCJI1Gd/kY1mIeuLjm2koxJfh6Bx7/0auNF8QMgydML+6ch8MY
Z4CXgVXxn039cAvB9fNHNkEwGLHHvc8GBonYYPmBPzlaqgvW9uUkT8teUKM5fDkE3pfQqGkryMMI
PZbptbFnnezd9mPg+uyUzkxB0kuZHAEKvSiZwQT2oPAwgdY6LvSsaAHU57BzEBUICYoAh+lBFEId
V9ESu2sJX56jdyD34pqr50qxNKj73c282tiMB2vFDgVJ1b8h8VykB7m0J2s14DL2mG8gNcGt5KG9
BuDaW7OuWrwH4dEH7p4FP0KZzqoeQGjT48AcCm2EbkfT894z77RD/bdCi8U6uxm775xjJ3ZPfnm+
3Jh0pmqtbQdSFjeRYXMDGpMkRl5Ml5B8uP4SC8Qa0GhFnL+tGBR9JxEEDJ3U5sVnxv8UabeP7Z+s
4xF6yUArGTgeZJ8NKxqLlO3yMEe1BVLnNXI64M5gGR3wObIeI/MEY+OpJQtvUT+yf03hqIeQqCjz
kOTg0xr3/POMZ5mOWcLUIXaXWL924QCx1w4JcN7vjJtYzJp1sRZ0wBZK+r9YcdXXpafGR5NYDXCT
i63htUBdAO3El2Praav9gM5Jqw3iNRJUmcAsOiJhKiJ8B5Ht6yCW1qYxsSimVpFY4H0ekZrMeeT4
qPAil5XwgQzueAGzB+6cwYmJK6SZwA3PyeQkYdLuShkMTuju+IQ7CYMP2Gp7b0JrsFsFFzUwcdeS
K+wZWuI8Yvxs6XmI//mrJuz1CugLr29Q3iN4uOgrfG571tSlaCZKLpNGgsJGjPrzH+k6Gx1OrHpD
cF+1Of1ojfCidj2nAVpiqji8oTHYl9oU+3NOt9Ef5SlqZo6kcIX8wT1On7Wu9wmmjRO/be0eR1LZ
muS1EVpLPlcXNLwiEkb6+KEkwYlEB4QiTNglwVXPLlqwecURLQcdm0QAacfD/qSYPw+0mrF2U1F5
0KVIVU/C38HciRAK5Py5FkwTcRnk8aHdY1BjnbxpSo2/tMpPOXOE/shh3OXdkvoRzOaUvK6KKUPS
o4fPpmsTOzK1ZUo/AqXzVwnsvGY+6AIlWpeAuUv15MP/kSgBRluquzxQ/dIiFnjqasFk5+w5bEr/
4D+l0TIBJZEpK7uaEumAK1PYe8GcTCoXryI3zYbXLOyWppk1A0RKsM30xD2gELz+rXB6llXtKU6N
xGLCYIPUb5qtpT1uCX2nxEWw9lJl2g7YscsGu0qBY551o0l+Xz7BH2rKYFT/rPJDXwPSnsXdEG0E
GvHFBsjEmjF7eK8WBd8nrH93cJJakezg2MbakARH0PPa3gccWtBHbbgiuiRtXW9Muy5AD/Ld8uEU
iygZWWdlZRIH82i3lLj8gBnOcbbgUiH40vjh2t0p4B7ErsTlc5P8akNlOrHw6NyIRqbq87woQtKm
bEzOASXQ1IW0bveWfIy49GIpRKlOhTf3jpxA5mIiZDXnvLxTQvQTNDXk6ZUgyB7niiGU4SCqtKjR
aDop2Inb7tY2HY3eIld0JpV3h4s+LjYcH33oBZatiWZToksKvamlAsYvx74FvBTxnh2RKX9n1vQa
GzjynQ55t2jwjKLrN/Q6NstXC4u6GSPXpMz3BmLwXElCTmJavs8iLDRTsaNESzpdGj5Uta3WH14s
c8j1OKApWOFmWLRLE37UOfKQAAqJPyE6WOfV3Jq9nZ/gpwiK0etnMr52H3tL8jDhGXg7Rz3L/fPD
mbfrrbPaoj9M5Ph3L9zs0EyBJPZeTpqTsQ+xC1y9yEk02a1ZaEAmiMAHEgTXS3vlsaGp+xblBFxx
Su72motHmXZ4z/njQ0FO3oz0iA1g5u96Eb+/GSfLrgE90yUsmEMhDz4BA3wUqY5d9fJoTDgA+Mut
JNke2xOIOk0HCD5cJUQSA4dVMDX9ycyx4Rl/KjAGfK4CJbguVQZR1zNJWtrbS4Uj7ClhW/Mw32yY
+uDJzLNznzsBFTmLlAymJjbqwIA2cWSoykm3mKsYCdfxw87+b/5uIcux4BhOqQqydRuqevd/ohL1
/Zq+pxCvfHNSCjGZokIyrjcAiwfErGA93T2ElvgCK8tT5m0nD59YJT51mLE+UQ3GOpsVPF5Q4XDC
6WiB1LNX34xIFJF4K7nRN5nceQnxtzb87WnqVqu3pJEU1UUbfBX9ARLhXRtfEvpa9gznyRxrs/WU
OBg0SUWOL/343rkq2CQiRVyR+cEsBZ551ME2MVwk8VJYbFcdv4ZiHBTUMup7xZEfs70MF5Uh33ih
TLZGbW4b5ul2pJyrDNFt3MB2bp4O/6SIy5KnoZ67KkmC986I503lVjkx0NfwKfHtzbo1GBi5stXv
pD/yGX79t2sVuZ+NOnEw+t2Z2nmYvMQL0HnVuzPUWDpkdy04ueuX+VmBunKDQRSLJy4iq1RGAnTE
+xS52azIAv1P2ptg/k64K+PVlJwMzGKKAteZZu7E8QOA4/g2uPryfmsSCA30Nlx245Rk/RogTzV+
OkW5Jdcb84GKsBjCkpJOWhwWINuiqXF38BGjLubBvibWCUg9B/9y0p3bZAO/58fpZSRSp350mOvh
D2w33s5FL1OLv/VJ94zwliNbYalk2zy4QpuV0e19M3HS2oBgmdhki3/wasYnmnh3i928kopjNobf
mEqK6yp89wtOG6BLm6erPDqJox4zWuNsw9iFD5BxG7Z+gw5UMSyfdPOFWvz+9+jx8O2Db/ueQCtd
Y4jy+9YFHFCT4GZrsj/sC4VPOnJQu6CLpCj1mMJjOiDrPG0HkiJVrl2H6tl2Mh0Jw4sEy7q3hDUB
qK9qfr5xu8fEmVDzLeAHZGtUZZNWBjXsnEu9jYmsC0ppk2hCNeimwKV5LHiM92MNdtcO7+ElFp/3
uVvDQSr63+bzkkygNDiCLV+Le8GIKzSX7hwDqHu858YMdoS9a52AZH+TKsmTLdduKUcy0ejTVIJs
PHTXXyWiLHGEJORXgFeXt6mGxPlgFlMK50ZI00yJnEBA7LrFjD6lXt+aOeInVYp2Zcox35ol0OhD
MnoHYggDy7dDGKk0fkUmX0Jpcwm9wGX7qLSJa18meDju1l3qg/Mz66h3Zoi7+HhhExG1tqXwWAEn
O2LdYmJ83YV7RNy72PDSGw1+VJMFpS0HtqAz0HUqoP90jADtm3/T7XEEYsLqtX6px/FANSuUhNbK
MXcoya3k9sOAOruJfWTlJqNpGdkTdoL2uoau/U1CXQaHoiQXLquuK/kgsY2SDl51JxIZLIFTZgfe
yPdVsR0N0Dv0OCxcFng58AJsecMVb0mlp2QUxAVLc5pmFV+3ULxU80yntnAxk+E0/AVaFaevZdzQ
OC/0/nU9tuIQUp2CFpHdVQuZ+qzbLDoDiWsl3xP2cgfnaGNUaXJIdImErmqLTQe/PymKICW6o6wQ
KGoBAm00XPPEGN9nipcOMZpAqK7/ox+ClTp+pTfaZAZe0M/YDWmokmbOFFHQNLkXh94Pf3aHoIoF
id0ivJJlIZQSe4TsgHMej49mlr4x2LAptFylhzmaKaBVM/4mZSBiQwdm67CubXlkUCjsFgTxVqJ6
2rThybTHDSEl6j0qxtAo4fTmW8cGE3yvrdj7sx+EdWcjHhRXln/kNj0skuGMmYlCj/gQ68Qd1rSq
SU/pSC+z8I+0YgVU+KWg3ShmZ1p+aqJBCTsmUiGUfN1PnABXNROPsvX4V63JYMsHO/xOVcY8e2ri
CX7hI72R0Ald7/0VhXdZiRp6KGbBzLperm6GHqzK/e+JF8o3n4yzUp0BNUaEbUCwkBtpi4H4Ieja
2sS9tVtfqhFvzyyeunYOoJbPd6PCIhRYlEhXyV8cztcIb5s2TT4+NffBBv8nUSzKfvRpwefKoQFd
3Ix4fwgErkKto/sjcJOtjrV/rUoYmboqSnUFNznZXlWHzdtHD89nzxvqNLsf35zvllhmvCmXsRjP
FSeLId6EBGaMGbA+laf+X2VJI0eDGMmSgIWJ7/DCG2QONS8u/gqobjQexucTVDGM8Q8qKyckDZKs
UGl1zwAloCxLsJFahqXDVsdBnz7h3sNBPbTjfXUpqIIahtdXOnamkOp1rAQEdX1eSwCNHfGJMlKs
LwYsuOhiCp6VJfH1HkvhCg5Mjfs5ArulJPKGLSrxjm5FgJoCT5NCeDNBmyBabo2qNXwQYmINOVUq
rdIb9+0peMJbYNRR/rTIGXKWgKgQOZWgIOD9nrcW1/OftCY1JOQkF8TfOWRNSkFGHO4dylMTisYD
4h5Y/vT3hPo2SJ3Qt1mxeNPdRJw9B4yhN7Ksby0cnN/LUZndWzZtIeqb78EeQ+wgX2xNpv7vf1j0
g04Pes/IdMJaE+TAsGmjQPwZfhVavbnGAO1WS7ot+jkluvVxMA7xAn6hgvAjCpXS7uiqFG+ks97y
WTN3iWq32j4AsX0JjXu6Bwf+n4Yke7ly0uJ0cds5rd74i8S1+LVv5MiAlvHz96GV3upGmPV5rdSC
bJZZVKb0pk7jLk1TY45E662IDQTYsmgoPxwjVIXiBRBvYx5djHpmqnSZOK+Nbm/zUyESW9xVvXXI
UD86LNdRARiE594+d/VVyYMRfoc1avK92q5aOUlr0mRlc0pqsAiwosluQ2ZFZxGc3nYK0sMGPdgF
xljMUsDSvonmd5za56qjN8kQocFIWOTOcKYSWgKxAQSz2d1JoSLDYzW2pfzO91v+UClu+qLCm/GC
3NUbnDYfYxbFYWG1pPcGCFRSA5qJFFP/EaWxtIq+AYqGTljyFWDYgL6x1JSvJAshoKKpRN/c/lrM
aKJBGuxv0oo8G4PEi5FxD2VWjP9cHAIfrdhf8jaUDpkThwsZVgOIUkcqIUaC7MJohavazrKwAkaC
2UYKjP/ZraTiTCh4L+jomRCaVADucS/5LbrEukLmfW+Ia+/6iZ5EAHDYCQ6AInRyyG1sFE5QUfTu
1Hu4VWv95Pu8h/zFSy5e1HmJOIIZPEsW/KNQUfgK/+dwgI8uK1bpUltGBPMoLeFoeEDJF0+ADKh7
Q71xliE9+ZZWhQI9euw3oCSEESjIVUAWtZBOrX3kZHgct6TsJCBT/HIQSLgTVPuOBO7gLtpEtOVh
VLHQwzgMOEYUtRjlkreJXtdwn7RGvDIbZ0UaIiSL5Ls4zLXMPgi/uJ7IWP+9OOZlLAXlawip9O5P
gYkPhXS3qx9c3QJ1JXsgCcEAq7Nxl/i/QJ3Qtc+nrWwQv5C/bVZ9Su0VcXUrY1TVQ10UNrtefJW9
UZQaS5dGRDxdCy8DMcJ+V9tNANc23RYWOt2dsRztqnFFwaXTCNc2riM9M4FeL0IJA0M5JQ9+xZco
AdjpmYqbRBleq6yNkg7/oM3I7JpRM6pE2tLZoaBJ4eHYcW76wZ79BARVddEh5y8F7ypvX0NUQfDc
iXWa0XafkcVm7s6OG4OhbfjJuC6x+L9i1/ILqb9+vzwFUlf8Ke+815SKlJRYRo/uzZ8/HkOapH2n
as4MHZFZNpYl+cKJw9SKVa6y9+xXALCeLsrlwrEe5cNWyPJf9TrkzWcHkHr9ih0TETgsaWDW9DbZ
hxojlji9rbse820pLCbPnZji+VLqYhrRf7yOuVrYyKiRiE13TGSb+QAoXkP1F7b33NMYttMiTFHD
oVMpDOVB5ha7FroHS0tgJ+pcPGpn1hgzRDV3+Kj83L3E2JoYQOvD/w+MFcnxlGe/cTb/gUjZ/D1c
pNfNbZOZZA5qY7dXYMLPF/a6Trnlo5c4nuBqf/YWbwZg7c26qNB3fsz9hs5TCD12E1HKuTrhr8I+
NEVZqDkRSxTw3AZZL6GrDj6PXjLI6W7oLOJX+LWq9N6QotXqcCxZFe9riKRZfztBc/r73K4JhlYG
1Y+H2N15lCzpGHk/9ieUiYk7taGzMjtWAKN21b6HbmQg3PuNNXTZ+UAiA6Cf6hrVtzOmM1DpNlfH
W0Ucs1ZBVvGtpX5Pg/kZ1GQMD14hCA6wgYXH3fa1FK+m76dLEbBobYGnZ+drTyEyyLlvaYCzxEEb
EZnG6b5UGD6bXbNQ7YnSSJa10R6z2uDSz6EXF47/Q0ts3454rjddqdSnWot41svgCcAdje0aRPhF
ThM1LQX5/SIAFnippDpHLaMJdWceo0age8SqqXqUN2Cz9hVBJCiqqZT5u/0CDzrktkktZ8re1/Fv
z73YWexhqetbTKnRjuEoWVneDeQiQQMBUmZLrcCuZSC8MgrkHHgnkGqV3FtRkmxIjmfspNf93zUV
xWnP20/BM+jODCmykiBw5nD3oviMEekhXIQNIjjejzA76Zp0GsQISP39v9soL2L6H7DT/4E+7kbw
Vz+YC5QehA/vgOSbj+OIgAt9pJKVYgflXZ7CaGzjyx4aAPOAv4s8CQLlaN5OZIMBa1Sq++I32BcN
AWO3ZaWS4+BSzBcuUTPVI1nvrBRA/OSmeDXRYQzRQip1Yh27XcsttlWcIILoeUORWsTfmQeFh2LG
WOflwMpgLUBa87rJVOACCGv7Xf5tWiRbPBlfF58h9cd7Jse0GrVBrtzPcZF5ekvIZwfSkqWIvsIP
W184icHTAHFZ7j7PpHpAaJ3/94g/Ak7NaVPmjPPQ0U5j2EDaqoifAz+UDj4AA7ne48HUlfq4QZlQ
hfNUcg3DItZ7ZXWNTXn8z59Ryd1NiYzFSwerfbjYdB7a5uo7Kxjwe7CgEOaifjYv673UgDudrRea
6r1z6nektEE8X/nhC8IXCOY4RLyHkOsX/OrPpApH0XuSVKrN17YYWkDr+xgSjb3KSVf/BngUnGOb
WDK9ocwlRzTFKPyau/R43NFXnaOmXvLaQGtUlYb3YbRs62w7lwpvGL+Jq1/1PghXdyv8Vih6Ya/b
7Rm9aJKKrK3AVTurBH6UZgIJlTcP/WEvPfMGaVGizDnr00woBRUV9qkw/OctruFFVAHIPBCaIZnf
c0bir/COd69DY25EYSCqrkwcvGqT8Ds5TzSgAD/NTMwwTIqW41B1X8e++Q8pJpOzF09Nn4nNZurd
ViKyd+InHkk2kKqs75Swjr5zCPIv2AuPn9WkNqplM0kOrL2euQASGT2XWfyAnCfNQkxNrGHlRzVE
jyrOBjIi5ZFEL8S0Yy+RHtTYlWPRe6E+YWwOIZtY3czeh/QjqPNAa5skApspuGVGw3gEsNtEcPwJ
/XJuDNLgUj7NFFR3eE72DFUFXFVCZHi42nzZGuohQ3NL0ekibWluT+Qh9QK6u+5YWLlPyXy7cu3a
k9c2kiEfc6jyJ+L3ppQKtUmbf3FHDQ285b/ku2KevMXX0N4+BIV5jVGvcvvf104p1PzPZZg55OhI
RJ5b1+CIbM3BV5YDGouCpsPAuK0wGmhIn2MAQOSFsaTAW8fMG8RG1z91Q7I3AXDJbB/vCAqJA+pw
587/JSZRDS70f9/Zf2XbmMLAKtbh08CC4PtavHbN1DiMd+1N89M6oLtFpnAa59poNGJls4oGobuM
rN9L3CaIQPloE14+7utMeyLjE9xRC40kn9+hrKXDw+CPj95R5cCHAbgfaToOslm2cTlIKivKF1HC
l51KiEqLOiLjuSWbkv7oKT0DggCF+fG2nnJp+UwJEpatEJEgyyxSvVRCCc8/Z2w6G8sqSws4QCzy
8jpGj6I+DEduE/R2kGOrEjl1RM9HD+0MhzeG2+81KZwAMYEq861BQo5hqRcxMuDpxdJ3NIlxsaTN
yhOtqLXUw18sNZsWEB2TYrxAQmCDjM+SkxKSVcfA+FWSYDH3pLIAlBDvjGjkC4AzhA+9ioCwogT3
mdrV/LWF7t+vjk06rLet/Fo/tqslSr3lJ1RxDmH0MLE8+lpP3gsuoYV3sL86HRsGwX4rcXF6O3IE
hf/DnXNaSqsO9eXePfhhvf7Hm/1rjngqn9R5u7T98rA3eQ8GNZQH99l1oPDgGW7pMsuSjIepTVY4
+nOt7/ogZ5f9P/xjBEtfey8OoXWenBNZWuzyvwA4SlJXKcEpHZJPD3gKdBqGZb/Qi5o4UO8OHaw2
iBPk2VJeZTZfq2T509JPqPqvYbxD2cYAeUbaF7yxidcKsJbAQzQP9eDZxI5orZevoeJkjhevoyQo
4402ubGEmvKpaCZepA2k5D/I/cnIFritLTIAirJemrF2cWwl3b5jWOse7DcglvLE/l3WC0bxAn65
VMIESCZ78vI4d6Eo/g89UX9nEn5rKIeHnLwSPICnGcjJ97SGVwKMxeaE/w/FlEfd3IIvCqArGaiE
TPEWSajt4pp2uMQpVyCp6NvsKYn7+mo66YHhJQMkHNyi5uC3+VFneMWLhCCujOJvWi645Cr10Y7C
Q0e8lbUHgWfijYjT0NWEDGWiKcFs/wGgU9B4yWKk5uopqevH6ABuEuI89aUJHmCObdY4XElYZ6ow
FmN7LG57hZKsz3olrLcLT/UEs4T1llurEz4Cvg3a8bna3ZunDCNKdiYw6l3rDVxCcce4cqxKmQQG
KTM+LOZa7WHC4cvTFWamAiJySWADIbKxzj8m9uSRvBefNm2e1pQKlVIlMQPP+4vf78l9hhkEkyco
TICs1MkF809EpJShWH0nrmsgMpSl1A9HSw4KyATp4IB1cX3fKdBMvt75Au8GazNM+nincdeoGdv6
5p5DCtCo9lVT8o6ZuGu70lmfF+KxM/TaoMpCN0Rel9h24j7ApMJZCn9F6YyZqERMoBVB2/qUVSSx
K+8k8fwIwlM7JDSAdRyG1LT0SrSSlAaeexRIwqipxE3TzJnxcpaoYiH11Fa0HJS1I7JWGQ1t23+l
b0mSSyp9sHVuuAHhwr9ZnRn6De4Cz+LE8avytrofnnbxZtwzTp5DIDdP8S641ClFTrwCVjHDWx3p
gD8PfRNdVAjWFUW8sCW2fDTWlfWIk3b+GZDinRazKByPAJEjDz3eEQrm1dfmDAPOpdjG73//6kQb
tLHWnFi+vOubf8uRq01tfmU18iHio2pP+oSw9xyF2g8QgFRoe9PNXEKzLL9IM0Nc0qDgqW2cIE6i
tjNUWW5r7ZbSL/nU8pJkOSP3bHOq14gsI6QjPySz7T9UIUVTQZLIDa5a41lkNijXhBAbBxciP5e9
TYIlS06nZIMzDxVK/wjEuJt4AginADCgK8oi7megJUMpaBVNoKPOT7tA9t5qQYqu7kbj/hxb2Uk1
4/xNhq+ONQtv9eYU12pUdSjWfKCNrArHPzP4ABQ7P26zm8Q+G6wh6xiVx64M/UR+aeM60NV938ld
kds0dfDcbMzjwKoOFZHM796pEk4OYphlw88/IJKts+udvMnRfiaNvbOJgeEv/LtFhjiKvd11G2oX
59a2f0spziao0DpuQShLH9Ivpv3Zgmcwj+kAdUBWJGKO2H+GMfu/9siIuJMEOyoURnOGcurYCEeF
uT6WpDMYnXpSHAqF/HNOm8RkHaUzC29BwDPlDTqyAZ8k1v9UYjE7zfqtPvnOBa6+6aAl6DfFP83A
+DExNCAK3T4duh7XY3GqcWmdb8SHmf2kiTmdaI1lez06TAPtxMIsobnlz3dCA3Tj9tk+N0VKuWTw
7vT0mpH/KUyE41ExquxFmvxtHmrDUGJwHqOIc/BSCT5CF1ghwaprvg4qivp1MgOF4Dd97OLZ7z7x
Y76g5qSDmO3ZxW9PN5Bba2y6Wpcq7MSXghf96lBU++uvQVF+OzNw3TDaoluKCapW1yUDuq9KnZVt
AnbTtgKKrIVpZbbIBoEDB559o6OebUyX/G+DDHkFD8F47SDie7wONf89dgb9F8PKojdIgZMpe4vb
AfD3g6hRPESR3INeKnWuinWKb9Qcrb6C5FJwKdXaiYmfuti7YhbCYkepYIuNMPYfUQsILor7et2R
q9bF4+yi46jqGOdc3+aZLoSnsdcfQoDUxz0rniVY/C+1xXzVZZK+fuujrVAZJ35wgg/oCo3pfPyS
RPbtBlTWDHg2Dhv0XlGMdmAQEE1g1MmGuUx3JnhJVymSFZUxyOMQQpem/30q/bRaMF+KbIX0YWvb
km0/tT9NmiZKRnCyETqY/hM4bsKTANtglFTn5wOiEkrSbt2OA6y/tcd6OvgfP3Ry6GZrKF3xg/qJ
s4elVLZjvWVMft/YvH/rIQmvxv9WxgeimP4jWP0M10EPwcYZ10cSfKOaSdwBdGdx96heqaZnw6eB
8CPN6zqLdMazdNKb+U8QXFN/MVwPNi7jFOWrLhOL1n6xswliJ8AzucTmPfviz5+/M+hqatr03A1b
aRQdxMbuh6+rwSka+vWx+VEiR5HbO8s1hCaPI3qRbZdp8KJDq3KnuazzlNmug7ukChDG6itGncuw
46GDg1B9qEsG8kys4pMH4MZkaqgFxMKwg102mfKOeIPd+2LVvjI3wypo/pnSHdJdWaJMgBGzAqO7
EHk3dDZg73jmWaiirYWfoxd+MY1HSvyWEjgbtJhFrc7g0DeG4YGKm+xe2aYyAWO2yYsP3154LqcT
3MXAUoo+9FGe/SaorAyc91jYIB5EgUVq3A24gU7JdLNkf76sZ6ctiBvRHQwxybEuQ9V6I2Gtjs3/
s7qyaraDHcL5NywKlImL4NdBtzPov65r2VA79vDuPfmm7aUZZ4kdu0XoOB3jd7UZgO3jblz+fhDd
Gx9BA/NaN4vRa21cZQNaIjmR/kg41Eas8MRu6f2xNyM6sszVoMk+de2hFdPWuq9xiH95+eMKNnUd
Kt8QD4DpXgiywGWqRwkCoNHoEJEPkc9cRxNFk8bl/A6O0NKly8g5AbbABPHPYsdfwL9XAhEZG1gz
he46Wo9vixIpWM/oGya0CkquGD5rF3yjdTPxGU2Uxp8DtiQWXETvWli9fg19HYobxlnMEImUWMbW
aYhsXlwGey/sOdJufejzDGwOHqcxfBiT9MASLtU72+uGRVJvGlsl+L3JdgaS2xkOLKci1M5+9B+Y
xSRl7FVf0vSw1hqaUGX3ClxYzLq+aUljmYS4zIxreRxeDqL2y9Apfi8CndigIVbZDFfdXSIjrsT3
Lr3jdIYapC048zD9t5jTQHJymyiD/6jeLzF7XKLPJm/hukSSIYLAOMe8GV08pqdn2eNXQqIKZQta
eEW+uBSXg8YzpLNomuB/T/kH51ddMAPYXWVaJvZr1GqNKpe3j/cbTlRWqzSa6ogWJw4Q2MoXutlw
9jFqqRhPmNk4MAJzXw6b+uOpPmoi7L4JucJJ4yqz0zrKdg1MrHD9v//ND8sLS7X1P8/NVdTmZYu4
tFaKNHGH2LxooTKBmtZYLv16aV7LtoRK+l5lglDQic6V4FVpZYW/ibB+GgAPxVmxDjmjTsZtEzqE
4Ff95McKrwCZOh8pK7d18Cwe/U9lvkc436a1EPE/QoKI61I5jAz1p/pEN0Z9CXbvL4BRTigaZHph
MdxaOzluOEAe7sdIypzjLzkyrZL5PRYUl45YxToMSpSRhIuB/A+TlrdNnWHnFhJS1JBLJwZYRsh7
l2Ry1rEdAnb3Qq+S3GaRjgxV8Qp3Ij8zkbOhzXk/UaqAiE4OcTNC7oHgtcK77nONTrn085CcwfEb
B3cTajmwyIrmcxsA7FKUfsjZWHXJmIHljB5FUhlKlooDxsM41bwXWb+ITFes0CV58NOxHROdn9jg
uOoSY+3GOLBRtI9IOUEOmHT9iEZcMw+fBW0XSooYA2Ef0UxK+xwe7uCwa9/qNbwzhll88vdZt+Rb
EgtV7/LO1w3dkF0AxvSKsf6j3lXWtGvYjxPG4a6vtvuJ3xGLaLYJtE3H4TVEeEexX6fFaa6/7cXp
yf95HwSk6dzApA5+TQnjrNXWui3tVeGtUY5q5CUvAm8Z9d3E6DEcdn65GaogGMUgIVKIt3bVAMQ6
jJ60efyfIjQPuDAARJDIFDiPhOj/j0y5lpGPKVYdI8mjlFQRUim2ear2nZRQKG1d7qd2H/kNFf1P
M/CgncEO/SWJGjioCt4hr8lWwjrL84Fb97OcFHnGpsqWtUIRXbvZvidxuxoRuEWssCpJrfs8Z4Fq
ZERyQC6X7JjiqawLV+WwF5AaJozKdjJSVfNHn59JulEB0o+AFQBbVzGX/Ey2Oq8D+yx7yZEVukX9
eaezmw7UpvHx8rZSkHjeCOQSvwcCpugVc65+bHqMMTdNwCmOblFSX5LJMzoneDtFVm/DMYBDzflq
vgWxUMGRXpMDSynU4tW0LWm1SI8g1TIYoeCCMS3WnPcn/z1aYlXuI8xOmtr3ZS3jH/prCnK7o2CH
HRDpv/T/wntrah18XIQS7O60KfMg99vqvPuf15qo7WbDWgt4e1M0HhwV4U4ndi0Os/TsmB0U/rKP
835Qx69ggIdBwIJPakQOvAACkd6Hw31g0Yr5XRpl//pjThLhGxx7xZm1tlyglDRN5BpOeD9D0VwZ
mVR7XHEatCK9wwtvA8J+3rrZ0K5xjMiPeL0yCBmiWMpNV5S7GcMk+uH68j7InHzD6WIbXW40woFy
Q9Iq8djbQIwUZTtlpFiQUm8b7lEmKQUKMTypxRArvSSOEt2ciqxYGmu8GxH/QezGSVwIGUlQW0ta
lzxxr1qRrNkyc6smm4lMrpYGE8j0WnKv0U/B4f8WW0QQV2XfzVjctuhLPom0/ViLrHVrrnm6Rc2Q
K4mx6/PE2rfN4lH5JjHGVBopK0PZSDZLQxZ/gEYd/iJiowjhAOUpwSgVcvI8L13AuEY5GmNy22kh
ou9cQuBOdgmb2xqqZ+6kkEMxs61PrdRKBhEu13YxuJgZhQu1AhxTQ55ZARSFjxt3m5YwZ/dBIK97
A1egk1OtB72TuL1zlp/h6hl8Vb77DeCLyAYwss134bV/bfe1qSe0Xq03ztviAR4VIfJXy8LnR85X
zg+PM0243TfKKD0lN+ySqA2eq+v0+iSqmZy0/R9SBh91cYvtU83izOfpIk8HWxmaZN6a4yZtLRxN
HG8Wjabj7dHcGUxhVGbC5qnKNpUFWuKEEyLN5EDazFOEBUtXKn2vR9YGKGGK78Jbfy3KdG6DIyYx
sR3uSUqHeUw1A3RdavKmF4wp97+TcDJI5GShl02rg6BgF+Ft94GRJPTCJDTf62Sc2RsAmmHfdLp2
8Cv0582TEblRc++nQC69mbgx8nlYj264sAywgeX1cvBYryjLq7EGSQEaTbHdvKa7Z97y5o5noKiu
mw37UqP7yUYF4iRtuxAU/dWJLRWM43MC7hcTraZU8vwAl94ULiuCJn5VhC+EzzaCH9HxxaYgowbp
1rVbQe4CIM/jUttbD8hO0Se1o8OyEpSQ0Y3MjoturTdjtP8+fHVlCqFalsoxHpRoCURZWOzkMI9F
fq2Il9ajbTj3w6EWyKgdpHWUsQpQqBRexqkVGIRDKFehHsQjEQIY3qLPwanygF2fM++xPDbBDApV
1IpcH7xGfQrhwSEpHGlcQZdCvNcJuItIw+ZP/DJUHiuMEmh7URxywwr+SL7sczXBc5ZPDtQT/8F4
vrgbUebPfXIdeWfqZNc0jOiDSqlFtVfDKkUBSVRch8JMsNnDY9gi1yrPNEEE2iROoTlmsh6Gprdf
W92Zo/rwZRXJYn5FBLlEol5eDxfo9MfHY9GbxfjOBQDo6p1ohl7ICts6CiyeIFuHXNrP3igluzsv
RygT0WfjFvSFvvu/4BgDfsldWLHLDNCuNfZnlm84kfdhLfwVat3rh2cvNeVbIH7RL8bY4W2h1jIU
V2mjgM3qVUnv+VFEPGs6mbfB/nwuNWUe2ntp0PgNZol90kMLm6jtKrfxNxn0xQlNatKdcCVX/wg1
esgNboDQwGGbwQrCks+DL9Jxn+iQ1AYPcAH7ZT0HQkUIxL8gXJz3FuL/3MJb1OlibmaUeI3HweEc
rGMIrkR+lNT8zzMjQ1aLAzn4sqoP3axd/oUJZ7/F2+GSj9hlE/IJjysyA9VpaBxKOZaUVpAEVxnS
UTOHNj4ZLbddASV2Wp2jGl/khMll1vz4P6JQDRkNL5w5b5OpZL6Bo/XiB3K4I6HNzr/71MnWqQlT
qCtGHVZwbigjBSiTAkiwVs884hI63KxGDoc9eXfsw3EHRHwrjiPXQT0M9y+85gGXVaxTOP7Y4dD5
req5hYbq6GV30tjTm1kD5zaSYV355x8g2CyoRchZq85ritHvaKx9+BuejUgZegIyZz9IyVAm1IVr
EctKQFb2VF9ocwB/X8WEYvqvKfX+LynxLSPwVrQs9s+ZpVrkEp7h531Vkm0epZyTfn1ss7I/ReHT
7w9vPFz6IrYj59yaxa5EP6qYCXrx/Kv9mKD2Iv69IpIo1GhMSW/YjEhCnljH/k970mnbyyGkhxx9
3tTGz4dDIClPkEuLBLqohX5QyDkQZYoDHW9nRpkwOctnpvFv+AHR6bIkxkb6Co5EN7rC9xwFGsFH
lueC3HilzQjzU9c3XuptcQcbmqeEY8jqu36eA8Q3iuO177h1lrS3+e0bP8A1gu0VEcWSneDHowiS
bogoX9V7Y+TxeSNdWJsCiw8ewD8YoOd1xV9yIEc6zNeOHQuTM+h3gwDsbncLHj4RgL7/yq0D4OfE
SbUpJ7YPlxhN5QGwZBTpInA+5B/u8h3v7OTqgcSPlApAL6ViDvA6yFUUzwU0EHSMPjvLdnUTsFzN
fK9rrxu4pcN4tRdiTOSwryJ/f6z/vt6LEjgiW5G5r9tUQGm+o5Kdwl6MQL4u1gqCpsE4NH+RSnKt
wCzKcJjcbNKe6cfIWVLf6EFpiDDz88bOVRsvVht9ZmofZeuJgdm/FNYU6+epao4JdobhId31Ys0G
HXepRyCSQ6b5Y+bPyDRlicrSuz5zMWf46KuZ/QAs/KAMi6PIEYp99tyyTjmwmwAXsCA2/J1gEr5u
v5ecfw8xIzJ3On9hsBZ7WVxh6Z65eVGB9xX7Qd6qN+Jj3jt4XPf409RohRYJPoYY2h1FD6dHBorA
W+ACVXInrzMn3pYSCRJpoRIOx1JRfDVoCr+x97e8B9bfYlM0PRfO/mL/q/UZJ7gyJ2TVS+Hs8czE
krcs9SJjjI+gfrvdmLP+00CVTGA9T47KPB0u1YvxhntpWRhTsi/A0AYP5MQh6AnSLLBwrtCpFLqQ
3AiSbEgFTOiguy5SRHHmETrCx4ELof0hQSlAkVJglXbOjw6j+Ruinp4+4jV75+kB7BaUo26iz4d4
NHn/7OAJKAN7WOfJn+NtZPz7bh97+aPmfGjSTzaTDkfrx4A21tt2Yg07iiSDKWr9YPMQw+SLLZy+
MfPhHlU/yx4lFOQtOzPRoL3Zf1jYz3SCow7dtQ4mMBGV/BhHNVjI1Ls1IqGjdIXzIY0r/IZDTaVW
FU6x7gJ9+AU99F+HTg9dH/VD3XhGqBV4KXhnmI5+ufMLAFV5nL14D2NA3jG7RBsEpTBTmsDohXG8
g/n4LIPI+zX5xGO4Ca974JTxDQn4IOqEhzFkz24TJbi42mEK8MpGsf8RIPcEzp6quLN1CPcNxssj
ZmWfQ5gXu1qy8gYg33PRP26FYxYB6J6s2XV8gAcW5qGjAMqaHsydkSyb8hThEIidXYfQuyPCdhKZ
NKzDjZExgKmdUvLXm56yPfwXzfuGYnWSxA8s6SYRxJ3mstDNDT6bUtp/NCTE0eUthDaEgtImhnO+
StJrZwmNYqZHBdrkv5TeREIndRCcX9HX10J8gl5brClAjJBLnTUaQ7P7G3E3kRFuCdcIwR/SP14Z
TW1jyQipuNDIy8/KSD6lzix0B95tfqmpbGNuSUfuW+6Q2j8JA1vdT2tr4oKB/OneI4/1BvVTEcNb
pcAkUtXdU77Us+cv7Efy352G3cgU/OtQGWDXf6wiWCX1qk9xVAvnsZl2KCfQLKl8xVtHPakncKED
KUYXfsHuzdV0S6y/0p5XG45KOBws382kknDzwBoXsAyLcIfMfefUvrFEj+FEDnlaBGMhD0D0rMcY
yDkkW7y0Gidb0SP4JthHQJj14oEOwOGy1dQj1Kj7UQD52RFfm9q4cqDz4xRG2J8t752GjutLXO3N
0K3GKdPTqzzdm92XxT1M5wv90w9Zr2tLV47EOQJlwm4Zzme9P+Dldcgeda2GT4k78D7HseUhT1Gj
qxTWyFbq6RhKNOuV8NZOXhbxvt167QEuivEL54M768lwKJr2NTP2apJ7z5LcQ9kuKbmn2Fwspb2e
K7QBDw8+0FMTUVz1nrhxccVKGYNTbb2xt4LvZpB+Rt9m5Yaf9l8R4u/ao+Rzt/GVZK0dilrSL0IG
72V2zKccJ1giAnmF9iyCB1hozG8g4A5QN65A0tqBf4ZaaRRcF7aOWSVgNcpywmXMlgRrwFun/czN
Zhvjf+Jf2MatjJHjAvsdG2enY7WJVSWhmjGFA5Q1lvC9+GXgL5RKXffVABfrXv+3kplZjsmPwU3R
/din9A3k/nXUMDP0Z+hGONedq316z/k1SL6r7xy0lN877eEsnx4u1RDeR3WI8Wd8bM6xCdK8uzar
TUkwYdkUuU0OI+OybnyClkzx1s52GWdNKko40kjTNkUydSY9F7j9k4FZlzolhY9v9H4lDnOvxZrd
VHi7xUgv1ADFEPnhKt+atBmJ2JjAHb5txKvlUqUrq1zouN4DFSTzg6QftobEB+3GhBLqtUnRmmFw
gFNOpzsEprYE2SQnHFA8gdmPx++RQWtJTgOx1/nhi+eWVLY8kLf1J5PqFHw4X0BeccbzIKtvlNk7
SQOgfze/K518YpJqqnpZKOyMqVQuSQbWSygf88BK1lGU9EGlci/CaDdRXMS9pOLLbD5xXzb5FKmD
Nu8bSYp94VE7+4VCjsjr/5FYJKUlh9K7diafluI8Pzi0BHO8nOUYD2f6GRGvoPdLRV/HWngt4BWB
XOoAbThtZpyCTil2bwYr5vNHoctgjhfN1s1c7Hc/3G/QIERHw/0RvnnPWUtXQGq8xq3Nf+F8u5wv
zcyXKVVESbDjZSLImNqAirWi3L8z7uRl/CX0EAh+Qqq5f3wbV21Ld0CI1JpblV9NCh6JCVYPpPgh
9bpI+VPfjbEReKO9oNR1rC4JYgQRNLWur9AnCxUwOQYMmX3Wbp/nJDLKDMt7Dl7BpwnlF4OPlh7Z
gg7/83yKCaC4chrYY6pyZHhwz5yGP3/ZJSbXL54dEeDTuFQjyFluLBtUS+5gK+MYQObmtIVjryMJ
S9/t696k5eOGn+2gwsXsNJQro24ByzQ57jUS3CZt4Y0MnKB3JkWmqhctGdlw0gBwbVcmHxCzvQLL
jZWZcZ2+BXMZGMpD6YPqqlGcqUM3/DNty/ev++sXukFo/3s4Ea3E4GX005TVzebpgaFPK73NlfjW
cVzP53jOD4ZyDYWWWSoaZ0pn/ZRoF+RKVPW+T/CpZDoMtPC/VdHwJtI5BaTfA9B1b6r0sJn0owkb
eWxpu+UQIWcDHdwEDY7zzrllUkHbcbsl20MDiEDsJAjQJ/xJsGKffOYvJv8y7DiJuI9sfccUVhJT
Z4u5qR2rf46BpvkWb6juEGwZbIUVfzWC85mukVAzSiOdMr7TVvNaZttII14Fhh51yFPR1S3h2v41
j4gtNx4xXg7YBzbhiixWUXKW1GXaiXc6uz+C0IOtiadqHcwN2srRKeE3sKuTHNHZsIiStRgPhkog
tIr0ZMxkoG/8KOK43UOnVXEkHa04Qf6ZJMD78FlefNqwtwOAhECKIfe5v6pL3+JeYwj7S9/oBwyE
ATjPiNzs615Xi8/EXNjbivWH/ZByhuZ5nVIngisKTMf0TIPlk38qdcdCRMZbm6wnSsBcUuA/zAPb
mXpaGlvO+gs7pq6qmrNHFJM9Y8mVbMh0CaURA2b/eKtWON/T01IBBVgLQuwZTG3YnbVjaxRTlSSJ
uMlEm8nGwuw/sHhLwccEj+9mhA/+GoAz104OREmseXYWR6VyzpaXSXa/s4B33o8kdv1IvdGMocST
xFxw8D5lmkFKq4DYyr/JNa26qGKfvgnrKnNuooM1nph9LY33kjIw8s+uJ5JOG0IVMoXbf4a9FzU3
yWzllotWRIjktzCQ7Q9vy88dSznBJjR3BOWnzL36F8u9tuMASjooRA8zTyif1zap6zvdAkaL3JNB
pN0kdJ+uiJFF1ZTuAMrJLiHSdyuWJhU3wqxoX5sSe+EYoEsMEgT2krxoHQ0tZxil+j+pW7XSxq5o
QnIato2jDmMZQ6TEwFfxYTZAqgSoXCF/s5+MuIinMOZX9vVn8BQkHU949G3xkFnIB5dZpTHcRQ7w
t1gJKh11Xmg+mLJR6WKfklqGxEBbMZipw0iUPqRPQXf+J3lR8dJqq8jAgTW2fzvhHLIoLICLxACg
004yR3T1+132mhOalypkoto5VP6QRvhQKevVQ4LJdHkM8iqY8ZEpS757Hiku54zklZF0bRsnL2bf
SLDYnMvowJTVKgAXvglaGxh6YT62vQuQAYM+GqunttFani1B5riJ+LXA0PGqf/Pw4IwpZg8Y8d21
+QhybEnV/fZitJKlkb1ys6w6spSRZqrCn5he7D4vaQ52xiU3TXZqfi6g2Z0v//097hw4OCUfHEmY
QwikT4W/6K9ZYKJK8NuZ9Xb1OcrK9FgumGBMJBGlTFP1Vj4dE5/HcN84w30zpXCLNiptB6ECWi/S
FomPgT+UyFG6tWiHEkz7YUWipjhGjMQXKibeRld6lZGTY8S/J2A5yl8+Xn6qPbgT5H58XYQCIkBu
SWZcpDAsoZcnKJbHNKDpx9gA2tND001t2/gh1EvrFCyQvIwsWPpN5H4Xm95Ivsd8btX865J7qMju
tzmEQfLlrYpM0o4B8QYvotOclrSNMJ3uq878qiDws46tJienmtwqwAmg9wkq913hlgyyTL7R3Pr/
ONm3F99V5DEarRRUcRwZRts+FO4/bW/633PuQsZpnjDyjecgUCl6EczoSoHR/5SyVMofGyF8VikZ
XhV9M9WzBfQhXgIBuYyixce3FHTcMpvFrNFwrpVqS7XgdX0ZcVk8vVq4jRrQsd7D0FyoiWAlBBVk
LrGsTwNKfVnFQQyhs0iylfpE4NQbsJ0xw3qybgK4LYJKR5/+kTSqmJMKytjn/3oXGVNHN9TuP2OH
ftmuRG1euIh9YeAdOZTsrmS40veqQZmJNpFj3o2pz9arPcX+jgyI4hE0fldONSQzBmQAjLac9n7j
JqpPHJigMwAcyuYSMe7N8mXM4LDGESDeQ83Of2FSrscSnHm98EjoF8zbRx7etU+QZmiAeswE6LXv
HpWS3xuC8yzH6F2+GsJiCnAFS0MuPa3WSrtO/V1bX/f+qTMfOZe48IzLB0ODW+4jRuuXxKiJL0ov
TjwXTTeyXRRfFY5+3lXTcMAqmtfaokw7C96Jbu+NyWKU0D4xx54fNrtkwgFpSm0bzxZi20AU0Hzz
CPnrNcCrXgQDpflqtQvmmkqE9msQXOSVkCgDf8Pe7nh8uhQVZ+OEHcWZwo6l3OkKl/o6b3HNcKq2
fzM9wPF+o6d4TKM6a9D4guSwKlIxsGEeukqc1e0L7rwuvCQpnfXljizcCWHB6pGYzHx8NyuVAPTy
mEHkJAP3zwMVaC0X8zMY5mmYWp6D5t5czn2E5TncpH7UPKSw+IdrVicK8tQ/BaZ1eERasTy4RAdg
EAI/UnHMFLgo27U93b7vsMBW5iLvFO15brqGUJAJeAOr/q4/KULLKqdYLhv2GVtw3svaWsfALbhR
r0lEy6j3F39JyyQsPk1h67Sj3VUkg14iAz/2m4NbSr/BkqGi0c5UPP3ABGLqAuzAGtU+R+XGCy8n
+yiyGLqosfruxCdTyHmPHXFxNWBe4fpdUDW8h0ZeBtHiArfBjPQRCzu6p2nKxiZnMAZBPv7Ro5Ec
iC7obYYYTzwINulsECNNyLDOTh96rrq3IEgU8hU8tyEaTlrm2JkggBuVyiBUgN5TREqtRCgCJ9SO
xd05D01CBYUoCzdlGw5lC8V/LUAdHckEhJwG8q1tlZfj2qckmWNaxkeoA7ABRrMiAWdELrzgwFp+
OwgwSm9hXabRCleqQeKXCTBCeTqhn5zVadNn77EnaouZ9XnmL0xZbpHND7wT6FCCM1U8SHjXCvje
/4IEs+u1rlwO1/vvJyxKh1Yx4mQsrYWt3ozXe9CfFTDv+WfP7XLaEK7ZieZsRcHl8WkfcrnSL+NN
h5z3xr67Px/RNHKUHL8WbJg1btBp4eJiLA1UVprmO20pkvxHY61Ldz+sgzFr9MKbASlBcC1334a3
H/NvN+1F5DW8BLIGIY3wSshU+HA0TdOqPeznVRCr52KrSd9Ydyhaf3utR2+vXEmt1XpoT6GPNvzl
QyX+YRhx2sWfOrMx3//xyOzHqBiWG41cZjDvDAoss6N/BBW8wnuebRsjDsKoSy+NV4tpsryhNl3f
YsPyRDgH0Nq348r/42fesOQpU+lXwBO40gHHKV9Q4X8zIsVKsQm4N52GaH8u/vujWkmUUkz1zWx1
6oyYrVP6eYjt/v4Li7FbZWU2JzYwBSsLWoOXiw/sFHNKjN+hPJO7hjh1v+nq7jid84NKznlx58rt
5Od8Jgi7TG9XTwdyXacwoVlY2r8pBAjkIwlFTW6xFUyPV6urewENoNqZxFmhlFpHgdd/+FOYJHEO
JJ5vyZmDz5Yrom0WdCDzQKrELFA1EgWyiyQmOAJb2LHxn7VD6/ARk2FwTO5AQVWJ2ywblP+7yxj+
QacogXfCeabs2GwBPbr1tTQbn8BIe1MTy/M4DunxGOjyKC1MvPl3kvaGTvH36khN46WLtFgtqlw+
sOfnnSAOn9d+xFq5QAl/h9M+nRLQVVQvyC/21cm+RA5uJXAfdPsm8kiKWjc62qYtr3eAUzCctXxW
MnEH480r9LJqRrP3YT/r9C/M5ANkmDphrn9Os07qfEOw/Mbh4nWcbPZBagsQ+d/MhLAf7QU5E4rI
ZCVKpkYTDGmMAX8sSwM5mS6PmnY/9GRRklvcw4GFaLNPx/0ofzbcJhqVnkIGtfcRmbW9VT6IjjRH
WutEavYZbA+r+1SyOxznPwyAuABMiBBlsaAAejjH3HE1Y6h+zFQNAB/2rd8xnu1X8dKrDmP4ABLI
V6s8iqh0bQNtGAul9ZfvjBGA7GLSDfb2Hq6pVAYkRLqlELyA+Bn4eZvVdYgdJCZpncoN55syuUZD
7XX2oPTNzyZDNDHkYE2dTAOSJ3aHoUhVWub6fnqPiO5fnzIxIy6khf6fViO6Vng2HUxFBKFN/pQ6
0u0mfoIUPv+EZjaMHun9bN944cF+rc8VmnsikwnOR+J8IWGL6IzCQeGMZVSDaQsP5VjMgcI5kLJb
ykgbe2wqtUsFaMBAIwnxxgWXj6FToQGuxLhCRXdhGzAuTDJ5GRAdHuwjVNwEmWyWd3VkltUbwRfT
AYrNa3+1332wcye9MDD+sZxBGKy+9h9mFV3CbvHnUDnAsB97yB0QvS4RdKFq7NYIrLGDmTpV3WcQ
TNwXMv4j3cW2IQRuKWzJOQ2SRDe1OE1A0gQA4sj9Y5GwtXUQuI1mVCZ+zxi0RHEP8Usmi8oq2kyT
i1tv/HRCrG46XJyUYdPDgGS7CWbahro4SgXiDRz2rMz+hYZE1pqluGsbnsIKcu+h/4gUQBQ+Ycbw
GmY5sqHTA5NYMRhA+Ifye4u83hhF6bwkHHuebS6vCEcXDtU1iqtrJVHGNfkAtw6r4kFSA0FyQVS5
4I/rSaEJioHMelVu07lF+sTGlwIKUhjZiCel5UXjUKRe11fkVChDbbn5DTSEKBHk+DEaoA7+cGbX
OcZqqb35V++mGhDuQLYmBJBGUVo6b79r2kSHot921an4vgNThoSBcPoAUzCG9au+EB3x5O/2LqnM
ZGW6wq44Wl9iZcz0Flaxbf3lBUCeXr3gd1f6PJpOGap2onCI33DxaU4uVuv4z2el5sXHqI9TeewL
tEBtv4tXFnaLQhMdMY1ATswBuSxcrcqvqxZXEo09920jlm7zDEsbZwqUlM/JYOvER6oaVMSBtu8I
ND/X0ZzsVgpcsl9hg4HkKIn44I6CGbRFm4aktONkAWZG6fAwi287D2MaBMGzq/jwJgsz3RqEuQAr
uFaffzupEUojncizqRQZ3vyRjMWX8V6yQcVpqv6K2slWbefiGBk8RXCbI7h3Ku/AdGXdTMzqpwTP
y5+3RssddFiIUYeE72Ln0XJiiZV/nblaoSbqE8jNu4fOa+TJfcFhPCHu35CXNR05KBXRktDwl6E8
NUqAvUS0CIxdfMzesHgarcu3wbdBP7lmniQ/f7onWiBGKEW93wyKkWQ9A94+wMiBheRc7HvIdFtu
Z7bbHYUzmkenfzNILMn68O+YjxKZTIirWAiXrDtGQwbHOA2NLLmpmOw43gCKuiNwgaLjF0iW50F6
mn7nnw9ZRxNv+u+VvmL0k9llCeKVfA7NMr06YMYIo3TTpFBOK7LVU+RFCwWHIPbootTCRdQebfBN
3sxraTw7DnLlnmODRiCfR2ZySJIQ4eXyvFTX/WlM+uIi/WezbQEIaK+hwOhramg/lOotE5b0xO+y
rwBGLVD7BglM35UnPGqmhHqHxWp2pJBcTWz501YZeewrlorregnx9KUomrkMA9rb0bICBXH3kash
55ROePNTBpQUfAjr99hvk0YNoYmGNfmdDTlmGiy5lDSw5nT22Nl4YPOBojKCt4s2nCSm+ZY3M6Tf
gCaMZw0uFyNgnJSYFfBsLaZHREdq3k4LdJhvkD8Gzat0xe73Yli6DEpfc+6q8s18dITh+UWBXrZw
FMfxGWswsL6niXTPJpoYuNlzozdrR5OlGqQ1t3JsY2zHpra4AMo2krx6JIq8O4ImeYFADkbfqrLJ
W6xCFTTH4Hi/bPWR3m114Ssj6XR+SAGEowywThs6nMBU1imPKNaHRRiLXtyFBFgwXFJ9TJ3aCszF
upmSzd7/tHGy2UoZ2geUsopLT2sB84Umxftm8eW5UNsE8Cg19JRyuVvWFLFCJ1KrHMLc84qTx7cB
rYuvEiUQvt1JEq/xbgqo2hfhYZB1pVHfcNn961HIW8Qu2bB6dl1qN/wjf8Cc0a87tfIBYZpZOf0U
FMkbIm8GW9UZxnqUQHcYbrT/uitIiTiNZczg6Di7fd0OBCSaNjVPluanW5rft/d1DO+JxXw+u1xp
uDbH9CUzCJKxIm6t0GhGFtFifehshIuBW8f0CTPqaFRdlNAZt9VEefniHZ0fpbIb4DQK3a25Nvy3
1fv1Av9tVFZEXFBCfbk0xJFkMTMoe2hplpziCCvsQ4Vmmp+prgCFPzZm3N7OGJzX8d4XQZLDXMFg
w34cdlVPLUR8XOGuzIBL21FmPGmCZz/VsNY1KhODzxFFdLrJdNKDDEyPFBfvG1avanNL/alc//aW
ogOWpy07D5dOHEZFFecg8eTPGcpx6xMCw0d3s7LsFulPxcoJX5nYrJNd7ystyUpL46j1hgk6kPrF
wtYae9YWFH/ZNNtYlbiZTP0OF6PjeecFAlXrM/PKBOfAatk4YkXZi61TPBoEZekn1D2Ee+PmJA17
9q+Sh7kMeoLjHJ9f/Sob8K37ufvzT3iHeay/1IlkS2ztP2+1f0m978+xGETlNdNr5Fm32VXKefPm
gZ1j4f+/2R4+rtScnth9NDX3lmGYXGX5bxgfxMENSZtVwnfe22L64ycaWazXwPm4486veTBx4f2e
XEBSSm4AT85anZ1nQReiDOojWk6JxuOJt1DMLrtNL+BunVSQ1Ngb9K2Dk2FxsvW0ARtSO2gLj0q6
vXN5EarmlFUiqef1arWADGuf6cp2CF/w7xVtqQaMFkGjiUmhcY1eNfzp3CxteYJN4n9ph00bdVMO
/TVyxa1oMgQj22P/hyWT+uAr5ZD7iVEU4zivN41/KxEaH5cN1JzCuCmeIvY+6n8l6SFGdWHnQeFk
ZXuKYSV86OqNQ9WCJXCEactzVeGZtQUsDziwE+hM5zyuE6wxQ06kpAkLUn0osPaUPjN/zyUcyX87
H7Ca3rz8H4ncRFhPqk+esm+zVV60Rg0GsSLZtNjSm8RsMTWoJ+TnLC2zpl7b9FMwta+z8uCKk/y1
ukZXbSBdRlUPVTQNo2A9zN00NSaBuDHT23caZ05/iG7IcQ8RVrarXNwTFXKfiwzs8ia6Td/TVKWh
k/QOLlQ0OgyK8R5dnpP/5TCahVwW+YjItZXofYkroqzLcXl1sEhWlISbd1mOxOLjC9HVDZSrCeT2
0FYN5WE4ctwSHAO8mYqiAPozHRtZS5PxCpndg2DTYA73isa79QyvDKqm0nDon+b6rFkOH71/VFYl
qhJ46aL6FP1vaAMipad/QMGOefJ2jLyYCrZbH6FtycW69mT8c4aZe5LrOqIQGC8sKPMgVgPm8iHb
87p+zoUKtyGmH9yUUTbXlgJXIXfClxJBWaXytheDzxKrtZpRm+LtSyHUoF8puMEDT/gdTHMygCE4
WozHjQK0mDkRKQAu/aCy0bLYvcHjMD1u4TEd5gkkdYI9FwSlgL+xTm/DETrt2VR4+A3kznl4auHM
gIXzfbrVLFSguuykX/UlNONAXk54JfY07GA9YmBvWgycZ+cDms3JTB37taVQWHwZxyvYbr2xCxXN
lqVgLPG68RJZvttf/BAZNgwKRGbH7VVety9DkRjveUcXs+te1Rv9GiPlXk21fUSRKisiZaHUzl+k
2h2pSEH0jtDu9KfFNLFpK5WS6wgaGz3a81phgzpE6WLviQvNxAzdipoqPph2A/XgMpsoZl95ul7+
gkyx31aEgmIV2zfei3DGz38mE1ImW8AynAGHluxxCwQqVUNvh7dsMjpUmaXxf0wNjzpRodaOwyhY
f5RRVgYlXktyhY6viFqPLaVejeGP2Q3/cZu91fGKC3TwEtmJXskncYx3tUaoNhO1ub91R9e2b+ZQ
SFOxiDlKm1j67czpSVQmLR2pgbH9dPoq3l0AnaobY5OA8ih80OQ+G5F0Iy3X3CTBCPlJuooWNqvJ
AU+FfnccJ6q6yZAmRiZCND61d4tSU6QRqtuSBiWDhW/qWBXR8IXUAwovj+ExuTUHUvWQjF1b5vvt
u/FRb4ClTGPzK5n05A8T5hk6u+BeTKLMqg4J6FtzPAnwoloflVjnX0PE0gIy3VjQjJtqtHkcETft
bBmNrmlfP9E5ShUTv8vpcb1MlZfIV5zOev8ZRvH3K0SsbfW/R49GZ5lK23NyZqIb8JMKYzCfq4Y/
K7VERVd3H9h9VdnRbcHWwLSXhRaWp4IMMQshfYXtI/z39OCPuJLuSquJMWOitW9hn72MC2GMoRao
ZCF73c9BryCUkdFabgycdhdIneOIH05pE8hFooQkoOM5ptDwKPJ5nBo8ngxxMIDTOg6W1OkYSo4w
qOs4zX6wejEu6EYCyMA70UWnbKvyByG1o5Kfjov/M3fdtyZdavuXMnrPgHF4kgIp3Kgip8ljmPbV
KOxtclpimZY3XsHXvV0Gq8+Y4qmwiE1SmM93s8pM8MNxnuWXx2ayYhrRDsHSGZKfDq1XLzW3P4ZU
82rgrVozMLhGah4/TdKy87peRLGMHqaVh3QqffxHwI+ffknRtmiu/0d1/E+74MI0B00PFDssCHvW
x2B0gDpG6S6WV+sS33pMIGUhtprEIhF4T3k629MJWGy/M6ipsIps0qJXvK6l397v8qE93cTjhd5H
+ls0elAW7N/RTUW/NdHMSWbem2unkNyQ/cUZZ8VEgK8uG6BE6NptJDfBq9+B83isZEn2wKEnCYKH
MtTvBVaVlkOMOL50gsrS31TWyXv4DSdWyrprrNFvIo6ZZoFCKJSUtzdVCFcI/uSgZo/2KpcB+c+1
M9lPh7iEE1lHf4mDDEUwtAYblyKtUWnhWWS8bkS36J/U4AEu/x9wCZJT2hTFQp7OVI+F/ay90F4V
VtObL9rf9HcDzjNNsRgAMIcArUNTWyJueF4X6ZxZHW35cjEI/fbJt4A3uNT93I2EQ2tc+WDPMPJN
Vy5ynCaXajyMDYmitHfggPrKIgO4jAjbi+dzXbUVtfSjU7p3ar3qUGXU4y5z/Vg/wDwgdqg7gyCR
KmW5yWakclmwDGF9zd8l7uvkun60crSLCQ3ptxaLWzo/JL6Fi8PxDO6nR4AC1kHTAzeF1N1wYvI8
s0iSpVmXfHnRV7HfOiofeLlSFiR6gt5lJpfqvovDZW/aWtm3DPtoETKe528h6W3nxerVeFaVA2FI
+qLN1BhZPQ52hzBWevHfPmuGBxX7mzZmmDV+OTnsZa8lE5LZiIbpA9JX/hv+ZcelzUyk6Rk9Cu+v
DDihpRVrVmyCRLVWkXEI3q1MdSqQ6RWlfgDPYSC5cVNv/3Cg3gvjF0FPg145uIY7JbsYN+a/ebte
H/NuJFlG8z+8jpiZ4ynoZhyvOrkotLtgljkN49t0HgjrVviYzcugQPvv4jHHU5R8hGs7HuBH6ded
Zftfn0lf8dIalDRWjSpVV/yw0elm6WD4BhB2ZdrfD7Ie+hcdRS1giGjKgtiB4Wfn1VqWDxcx4Xnu
DGdd98s+PWylykJL05wOS0ESucDObJMeKj0AjGKL8ZQ2w7yWrtZT+ovWB71/OivN0wuGU417/V5U
eWPoQ+cdajYxAsIDS4UG1fwF4d95B3XV35Bi9WGEkW18CnKWOOUt8+ZA2pFRSWlwygKkhLn+LKxh
OpRtWiiJC+veD/k4GbcRVvv7EuSsyglhPm6sZAzki5F9Z1fsksFypM4jGQzmURWE6De6tM4suWxR
Jvc38tN1k+XCcwKVHnHnXwFH1mehZ2kq2S6m8+3WXFR6hB6SmiAFFmgIZrd20pxukF7YXSYoIg6S
jFrRXs3+cFMo8CAnRY1aDw4ailIe71lo6h2rDjukW47Pq+G8nuy+UiiAkdf1hFJAZ+T5mTo5r43E
TqycT7CxFbaRUvq7SNAOC2sOiyOlZYGvhDPjS/PeeXBEz2WDtImO6KjEqIjHVzePEKrxcXt6/acL
YkRIoz1NnOeN9p/oeI/olj4ozO/qFyTtWxUiP81HVenOklxkQCXO7lYzkwbWFA29krkLN4H48fcN
ZWCzhTEUYfgzkYePWxuEkw2yDMhGFAfKxPIZaccaQBD8DHyw75cmYefMWvBR6TdBnt8NGGeVefpe
Udlaf5K3YL2hfqEVgkjwxdHDKEBPh1OSTvkUuPvfcbnbdoMW3A0zlv4algvMxXg4sQ/EQ8IjMQfM
YKnZ/MDoZ8OhvrNlAz85BlJkZd3dORrrT07Fo1LH8F0V5q2Ue9FN6+/CDrlxPtWpiuKxY6CyZBJN
7Qi+cdrkxsZRoMM6fV82Fq/lYxM0Fnd1LGx2ljJSlCsVAl1rLuBAvy6ZdvfTcMZoEd00xozadc2f
yOLNKknAQ+Pw6yp5yzY2nbY/Srbl6tFFREhoDq+QOZpKSIBdiUTEVW2r8zWhAe1+mFtNpw+wCRgd
kg4J1TOEXBnFijutHMH3Vfm68nBR3q7hr4Ibh1rN0sLFdQgx3rp5M4rFcCW6lSqxPONJLMWyB8ut
R8GRJc7Fw2oz1EWb88y256Wis2oS6IrGolsIRZTz6Ofhpk20ET2NHUamYO3SGy89tW6gCxpO5Spy
Rv2lCKYNcZ8Ex4PYOulZqzm41sAQqLafDY5163ov997GbB1lgKoO8gIz5u72UwpiTTGc7o7GWlCc
W+jV+J88XmqqFU1N6LzOwj3ZXzXmDUxBOhEbasjScZCeV0AibFQR5TGgE1gh0vrhmSkDa8p5SbPN
0sDPLm2FtyC3Wo8oHuAZbnEK96dgHAhGViQBUeb01lyzRbjfcULOtI6x9avWYbtXuAgmnmd5NYp7
tBrl4Y8npa5rB7BFxIW5mw26Nd3GUCp8hd0rx3lU2onwY1/0k4IvnsWowEIQ7DWNIbCvxIhZXl1s
KsXn8Z1dJ3XAd1Eqo4Tbh/kdn9EdCE3T84RwonmxEYUM824AbQwnue2MX2vTR7L8BvtpINXNlUcp
7Q/p75EJoaCynQA5neOD5saOjtd98vWv3MxNafiboaLB7FfpdDZ57Y7b2Jxd80miDX/4DTQm7FtA
T6M6MW/LZo9JAKPUMKsZJ9/c10tnNDsodow+roANiQswh+Qkd79034v3Lf/7NL/ur/v+7waeJ6ot
dMgYzcmhuq3+QPKpTmYyA6W1wPVm07H3Ovg9jJeQKjPDPuqr812eXbH07M9iUN2MSUc5Jnc3VZXi
1yxOX0WMa2MpB3l8ShHRqyYzfxXe0FqhL0S6r9ZhnnKxizMn2mcmBS+j01y4G/qVwYSiXdP5CJ7y
vhhksE01ko/cIpqdvWcl6T/0NHh804911hsQM0JSoYz4dJat16MgXRUf1maNnHozOgZnU4Rlyce/
mfLR6HIb6WJtZh7Pim6+6l1I6hbNJO5qB+31wIbSCI4ujPGJsrkeP+9T0sylxCDuJMdBYrg79XD5
Heskt8YpRfwI2CGWUJ7k+3/qjYQ0LZ3bNoDsA1LuOJoW9nAUE5A8i7ZXNWEuEgMYfmD/NJ5/PuNl
6+YB9ouePFBkIEgUECk5Y/dZm2eEaxe7uAU5GbvndOFpteJLmDM+Rx8g9TyIVCA0sfOGp7Ku5IKw
KcJAN/ZLjaO4HR1nW+bvbsZmu/eHXRI9z1/88mIKi1LCuIHYRaN5ROX8W2p3twKpRf9FPzSCsehD
2cEaAYmO1FkEoBF8piB3Ux0eG6KT+a1vMgmMJRilGid4PnsVQsLRSFpzQrhnhFgXTkoXt+wFPUNz
/25BYNWMn3bhmGOLzWRaOtvLMvGURlQu63l1wQNPLHJSmsEfC1+6c81MRtnxd+Gjm57E5g7t56TW
Er+weqSqGOkLIzn75TxLG1ZX3fgNRjja1JIPl2oFPHVeLa7RIp2heFaLFfyu4K02gZGMzEDaBC8t
OzxXH24pin7lVH64exJNisqRnPG+W7wA5ugElOuC93WYJSZGBbVgWb1kYEFZVY6T3prf6ZDQtYsb
+IHTBRsiENUkoTxtRAopLpezxK6X9raMbUiywDyYSepCCUL7WZdhTZq01qPKGkY5NKo4PHBt0mMx
wLV5vfWbKqV8gHvylRPqW3SdqB+be5fbDvG2bGn8x9Mt30SqgN09SX8KVX156rGfvDL2zXgoTV2F
2p7LVHoNWd05mg0MsYX4py6bfdyn0O/0WEs/5IR34UIBcXD4p58+UeKliOptztqM0q8R8PDBxqko
3PmwfBXYzuy3z0ELrhoFjYD8FqYTEogBmbOyfEHM1gZlKk1jUdjzyCi1ERoHEQmfGiEpFLNLtPQd
uvbV2ccF7mmvByPwC+KvVwy0zrHlVE783zAuJl3sd4+z32Y4mfrpjFPZGg8cCWIA/MOGRzm6XcXY
ls58eap6jwndcvacqxPkxArgFFKTDGvlqStDdIxVz7cfbcwXwV7FFkr2YSEZz64yj5hUyX/y0+5H
E37QxLXySKVuW8bHcCoUgqUUnueA02gx5ilaVFy8i2AO5meFBwFi6mFhtvLlTBzKijJG+rDTCN7r
yqJA755B7UajehefnWXAQuqRt7wuFhEVagEhopnheOJmQrUbTmGAg+F4Rptb/ZfVGA1vbkegTCSI
k+R/9LsLUeGOHuHTUedqKcwzJ4BxknD9GTcGrodVsFs9YWaLg/R8PlD8Vubza2viu9HSLSmpFLo+
HsUMgvyE2SBj7ukTgajIOVw+A09jygSNyacM9ErDomgp14KBavsaztlJvn9S+qvibszoF1TMk3e+
4vqMXR0poC6Po9oLfAgPzeILUOUlZqZxGxXaQ7C9HxnfVPnb7eD2D9yJf3RCOrPFulcOaF9zXqnu
Tels7GKZbAatQ6cUQaMglua/EVJPtj2p4AwCTLAOfxh3mnU8VQlC9jkOenb02DgJdbpwdyOA5QpW
8/SxTpyR0dHxv694bjQdgELlKS8vJo/GG2TDLaWLYyujsaKv/KciozuHMVEMXzcz2asxCd1o8tWS
cH/g4beFafqw74UnlJqrCid0Ci9WeAONyTyClqGJNMl0pwZIUJQz0mdtZFTEBRnrSLRhCu9/+xfC
lwuo/KWGVrO7UgapmWYiQFO6K16PpNCo244lDbs4DttnWKAY+2onVaT6gU44IVyT/Lp+YqCs0gpc
kM6t2HiQ9tQ1KiXYpmuR6clwdwKosSYeneAIl1NPX1Uubb6BfdOrIYPcMlGFYXW0OkDS/Fx09HiV
jie4B4H30aPknyT2jzz0R7Yzh+2dDqGRhLsdp67m0xkzHjJDKmJ2h6Kjp2kl3va4ftutQQkEZiwe
hAFIgGVOdHJvC6WjGq7jJNIhJExgR1CXA+ty5dCzvkjjzssJmN0GuHeDBuMXSxiwD22wg4NG6tkG
j6/BkD62afjd2tXkPrANOKbBqbIIqB0pZdHsf+3D3i5eEktAQDmesEZcDgdX7gtZAukIMqAVvqKj
VJQuQYHr/z+GExHY9rQn+/v5gXA/EA/ox2F67rzLRS2rrlQMFb4SUF9ddfiQm3Br71tufVip2N8f
vphspqhYT/siScP+2acxvPTkVE1qLdXb0jgwwbYIdOzHDjR1nNoil2iDnPjRc3XDl/rgxIO0VTyW
vXRzP5fg7hpX7rOkpMQQ4R5in1FmkWy5+K42NEhWnRy2bENk+oEil3JQDyFFZO10CB59AZzLTPKA
9fdnu9v68U9j244ZbddRDjKNVdM2ZSjOJC1B3p0dPDA06hTCag6tE+AaceIFDovo83dUzswxqTvN
5E4YJMEVA1MDLWk+acLQSRDPwjPVx6zPo95QCalH4QHS3sYp9bgDXVMOOGTmnfVtjEnrdx8HZP+S
t5WHrs06ap3PS34BNL8xXR1a+fsnR+I8z0Cyal/531wyzlMUAzKtAkAKMSW1qXKnbUcLe0cDgtiF
pWRAbrSGjqi35MIo2OXNqlL6kDIYVu2SJpXWrMyC7uDvzrbjHLkeV72jOBPf+EgkjchDF5aGO1+/
3o1X8Aga8oq3cNyn5BiZxY6B+yZnxHTS874o2TWHQJocFfHf7181YnemkiwHMIvh8H1SAQFexEEz
KQMNzpgZIH3yT3rd7lNTg55njW9+cOStQhdqAb3F8PFC6U+qxVQVoVzIJbzQYGp1VHtHWSmbf1L8
6iCn7ekdJL85+mkg0MFx9pbKkAXTbMtzWN+H8RjjuuL3K41Wcm8BZZkE2aoWn484LYUndpaf8J+x
X5iAafNTeHtneqVybWmdCmZ6EeLA6tnH5/Hmgur30MFKeAtGW7UVMsaX+PZQidCUlF4TeCe6sgwe
BrJ6+B6oVMC3gk9EHp5njH6QUqygovbDlMBx5nMT92redZbR1cXzUDGRsAUhz4GYdTFz7ETDz6et
zjDpSpNWQ3tFQT0sFpzOHu6KMAAxMI+CLMXiM7/DOI+HwvG1Jup+wG8sTLiQOMbHYeW9Q2mZ+ZSQ
Wgjc8Lzw1mcdo/wvyJimowMvKpbk3VDIK1Z1Ev9zspgFT3iS2Ak8BowP7Zx2CLOB9Z6E7zSojj1R
7r1UWIAyQLSIcGIzW/UH9gC0YgMHnvfA5LCMQBZxEqWTLncVmGhUotVaIfF5csb++LCOJ8pZ1+ya
kJI7Y52BsdrajttJ0votP91FXeMZXMt3y1VAT61CoFaexZkY0S+TNw4MQJs5R4BILkDCvMsz9I+0
1361MAmq/zpGeW4CCHXKN+RYYSPtxi+oHf5xV0Er0GgurkwOiT4DA7+xNtvythmEoMWl+ymgZ6Q4
BqmakFCRtRJrLRs7RNREO9U7/GVl4Q0iAdiIZza6wsn5Nfk8I4NjIsbELckfncfOKpGO+BhfSCnM
7i3f4g7o2ySxQ1jZgCIcWSnu7iLQYYhXkZsc0VJEoB7cxT/eHc5/Wb6jtzj1IeK6EpjjLuAFbPua
B8MtXXq/FhR5CqvSixlhxKVxtgRQYrRwBZzw0hb8z0zwcFK/hVjMK5o+Pm3Mbr27m18OTCvX4J1f
nXYlFynneTHp+pLnKqBqXsUVa6aZ4M5rSE5jzMenhEzCwSvzx0FbNCDhKD537VLgd3Wm2EkS3OeF
VEbSscCNsiYZbtgIs4W8InJB52Wog+/G+a6+aAlVDf8aNQs2AfnIVDzBFlJrZy5vI8crWpaSK3QM
XuGVMst2gCGI8Pigii5MwR5DLifsWxCK0SRpGogADobus4FNPagyOxdCVzzfs+bmA3eiriI6EPt3
+0i44R4S878QlTmsEJVcpKzNOIX8KpxJT9xlYkFIYjg+zxBIaTyMzXQkBZ+iUMbmZSwz+nJE7w65
SHi7OXdaurgAihAkdRUTJ/MKscZdlRMPmC0FRhSdyPKDMKMykvPqZsndtR6YKYaBaOHYeqk0SgJG
r/ycRJAZHRZFNm/hBak8dKMsBzm/TSZedOnvdZ81iCHtKqWppS/JZqDm+P1tPedV5xRVxrzNbZVM
zfTh1BrbV7bUNSfPU5eXpycC+VGtvDfS4mZpZW1na52lmwPG43Xu5CLe/BvYngGpR6MOYwAyIPnA
W3qMqXSKppin6IAn5LcNjI4HAjDAuICk94ciNKYkzXuLc2RUCBX7PqRNd8qW4+6hIDB0mQWOKE0z
FwmBJaIscAbq633rn8Jpl8WcuNnmwn3FINvL8Izz2UykvDrKJ0BivZP0XT99QOTgw7YBTdrsP9Bu
Arvjt66XlKY95MsdcKcvZ2HJT8lKROTxcyeHAe5ueU3WK9snIld2SyQtfr+JFjVaGsXHCthHOupl
4R03V4hB44kipp2xWd2YP9tAgqdkfO4tpVU4SViQeFNkHh3EAYfELnWJsDRBrB3XpNYKZjmmoKjy
92KgUarHApkd+NuAE93taV22gyBWZ5eGwJPtGiOqq+aFdzwhpWK/pLPBLEHOm4xSTFig5oC/eRG4
I38LhG1fsFQCRQ2CDm4eWnZWQ0HwV6lJxd7KeA4XAPU+Rxcfr+PFzhg/mbvpqBJJvW64KHsNDEfQ
as1ImpqFOCYrWsAociLFK4Rcbqx3shX/8GD5qfh//ghPLSd+HmxcUgukB2yYXgIVCCQO8RVd8kFI
Uboi0ltkzZ/OcmNXP9omv1bHqC9YX7VHUNTjVI3xhTD1KjawBU5LQUjojQakB99Jxm9zf6GmWEqc
UdsonL7P9SYpLXIjfcU2m0NbesbasAMlUx5ohESctMlQaqmZW5lSx9CfQwRaPdtgk6WMCBNZQeFq
lO+zQxqNQh6tPW3TxFQAPnMmeZxt5pm2TN7kHHsmf4IqJwps5CK91vr7ot72gVhFLD7TpOdtQCSq
owht82wwNHEQwHfSxum+r06bGYIcf5XKOqxTUb8ETuUUanyhpcvV9ugbNh5HsIhRNLC2BEXtTaOi
i7ob4rsaEXioKC2SfC23xRN/WHcfr24S8urXQFoeVpZHTkoIbVejg6LQhzi8CzBzopK5oBzoAAoY
6WlZ0t9moliQSXtw3yIEe9Ckg2yL5g1vYEreDuynsLkEF0R3adIoK4JNWWvS7TlET79ziv59Sld0
pIngNjMAMVCQaI9ogYCEdw0VFBS2djzgDXJuI76HPzjmmgn9Fv/bn2mJZH73pJkZcQ+ugupdw1IE
PaVeFAgwLjN+oN0TiTFLMFhY7hAy0Ty+3ndKpked66A3mwQJibXSN4hdFKwrWsHd3Mojix23wTX8
o2WL0KBe7TT9/FhA5DhvVv6KqAvdAKXtpmnhYLi3fuB7jp+GeAgL6Dn6q+qEqbqMJmEg5XElYeqa
kjJugcDQ7hygiw8ya6D1Zbaj5Vr6editWVv7OqGRfVktysiwgy8DuLX0hDKFobHeMAx4CRgr7UhN
JbhWX3S+4Xpy9M5SP5oAdzfLA4xA+diW8O5T9pHFaCjFwCJDPDJgO72LfQd0INntJPL5Or3CSldg
RFKoJh6y/qU19Iku/GbHObZbNMs5gk89mn771efBfZUINumvGrhpDbt8pLuqKSMUUD0kEAYLLAhW
rqgd3wWgj34iemVB2HzZyXyW8kI94tNytHiAAMlPe77RgioyNuiw+6yhTpSFfW/qQCMWiNQCrK6g
ozyS4StMujQdxlPGziDuquyjGkAqFk7/kCwTZh6MGPJHbxdBn1Q6FeanDihJ/wdKYsYuKJ0yPHKK
GRWth0sAcsKN4mvlOpYuR2L3zIx8qy6dRPZSTO4010GtGmMRE6ByVnnWsHsIH8Sn8/AoxVihyLNB
KWz0K+oBj1WSWBEwUNSt71FyEDZ1vLSMT7+Mtn7cjLje9Yq79gdreM8vxnUXIvhb0AfX+f5IjaOo
AYNq/3Zj92g4iAmHYkSHTR2oMsVJs2wf5lsESP+f5TVZDyHsygf7ax+atZnDx3eBk7JjOH5Op16Y
00vVtpzJUfkTgfj2LbzWZ7foqmBD5zo1UhWl+iPXgKg6NUYlZ8waLb8KYCVPYELHd8DeEk/6yUF3
LrBTY5qRV2lbU3vyQw1CFH5HUgDShZGp2ua2znwRMI1zbln2TrbDw1CsyExwjxtA8Ep8prZKeXmK
U+jGd2ej5+TZp/T8busmWoYjQ2rKG/o0rTPXShQt8sNYq0zCn9e9ctqIg7cdc+zO8zNyOPfmZGM2
BobKCG6jhqd0FjL4ubBDKGTT9DGpAb5vz32Y8dfcOToWk/3H+HLT6ixQXn8m0r4x5sOIe8CoSVNr
F69FH96+bkXydeg0sM41G5qudNHFQZ68uMZkDJFLHzORPOLS+KMq+CfFTBJvF473TRk32N7o8276
1bESe/agJvuW0uleN1s0rH5mOimOfTR/Lxt5YPwrx6ll4KqSRepqdM/beIH4ndi9o/2wrg6tTU3z
re0rUBfdYALXOIa83/eZBvOHbsd/cxBKhJghY2/YFhUW/gEW/PS9iyB6nz8EL1yGMnPMr4FB4e/P
xyTkrtokGjzmwid/1gfHd6tes9CpB789v9v3psKEFgBXhYHBGdUrF+g/2tHv0bGFnt6lGwE8fQCV
Je6kkPaCb1Z945HH+Uy/qc2ELxKidPPC4iTIOJYhCVnQyuN9vOBMPTahFn8jVv30V4RUjnSngA+6
7s6CeYB9AAIXxVIeJe9QxSMMY1KSWTmPS+rFL2GNTW+6Q1ye1k0XghY7DKOHXq7yx3/JSbdxV+Ke
vqGnqcUW5S3T1RPK2roSWLzI2WCIBY14DO0yq01rJ5xxpKyn0t0GDFK6PeNBwP+Mm0a153p0wxMn
xwZb8l3PfPJvBFRf12aydWxQliJC3xc5akPECjqmxluIQEXMO8ITeY4fPNkcVuBcUAUuXMrBW787
0t+zrflc8FNBjVFYul2ohFnMy1LysQwK8vWAp1UyEW/rLaxteOyaWtr6u73PdCcDtlwcYA5xC51E
E6YQEShxb0kXrXAsrfcDCudefPAbuYXzRCVQBQB3KuzcsT/Qwt73SbsGWWPsMEJQW0Sfc9g0+LBQ
9y5bQkx7oU+08yHiafDN+9MAQsSrvM6bB27Eee7DSTdagzeC/LVM7Ti62IH/ory8+2i+YIuXUutx
g5WdGCf19e75yZ9YWe/i4/8kPnsoox08Xadx4aokdRFAzXGuF5DjZwKcUmiou7OuwYiTku1fFRW7
J38K85R9ZOTHV9+nQeKIA3W4mABGEI8UKkq7KYcXF/zqIRypW4Pk5JRO/yesYXDbPpBwdfrInl3E
AKWsaJjZOBoP6BZhcyCjxR8vzgLP9s/TgcEzhidumwAAShXF06ehv1j7wsbdiV/gQvtGuaSMFEZb
xQlazxt2M3I/1wSxvW4Vxr5zjtFMnDhC87vEDtCfzNJlfInzCEA0iB4KjlXvyvddMMfiPEDlHPz1
1sfmY0aGKHh/QQfmGFRLxJ5WitcN3AJaMhm9qlhSYJjHiF7Eg3+rxFw4Tr3AYSPsGriikr1/XXhX
Sc9l+pjotUO84hj3RO15i/o2Za0RTuey1rc3JkiNKeJTomIxmR7PdCxJ7+0Z27tMBiQhJoZNPLOy
Vzhbd/m9g5L+d/qKPh1Wt23vG+EjqB18Nz6A8N97XGR9FVgRL3KKLPgguhGjdegEJSsdBIXOjFuI
kjDixv+hOUcwBqLd0YmbTyxU5ahtEx1k+KmYKjhMKH2SrrQ/0TS5P6rH9wwGQHJjJyoO45LYh3Rf
OmO4LTIQahNh/SeryhazgKNxNnrMVuzhoQGvE2vaK9nbvhK9OO+l5PMIjYHkrPixuOlekiplUzma
UN2UeUpRS3dFoyAYH4bW0Cy75KiA5MlV4L+pJ/LFmObpltmvAQrxsWwv5aQzRf65Vcd5ZUwr8yfJ
NZbFT0ttRxzyd6dFCVnV6jBJ1Gdb4FR+/D/1OrE68UiaiHImiqoWC6xwL0nbaRkZrhBjPZlJPkJM
BVeZlFCbKLAJvxrQKB7sMlAQxT8DhQjFr6bfZ32ThQ1geJPgymNfVBqVT6FOxpERBKxJv6bMe9U1
S5L2HCKfq97aMIYpwj7R/xB3Jy/u8oW3vqrMzfgDqRwZ7k39k6BT6mDFbcru4t55JGxf4lRvT0T2
4l3DQxQS0pcL/cSMHhpy1HTCFMd02JWLdDFFjGn+rqnxbFaGqaanXmKzIKGJXFg/2vUa9jjFyhK9
hpnMpxSQSTTBTHNCEcR8WrDxxjGHcvB3Z00KSVe9PA1ORix+GOfa4W9nVya7N8He1wArruibHWTC
3zIBM88pHjrtAwSg8yP4nkIDO/EX4YUCql6IivUidiktrFHvv3J4uYUwiMxGJurUcAO2cDUwEIHb
8/NQ1sLFCZ0xYN/yzuYNWgl+GM+RK8BArulzPbIDYoNOprDZAvEiQO23WEoKKUY1rHVo52cCAYxm
Y3VRNX/ttw2SqprIHzKLuibjCMUVW3EZjM4+Q050rrSbiRPENGSMJRlSvQ2DaPooJSurpaVJoCLu
2NbNC/jNj6Y3E302/Rv6L0sAhmHoLOHuFbiR7611s5SwP+d3CyQPtR/c1/QSvF0873E0iw90A+hn
IFeZI/AdH2I7zQ0ODt6JJDwTAdKCp9MfKeTWUbwmDsvHvx8wy3Gh+wCli+78gT3q2VbUMQew50hO
zqf+PwsNMdZRaH5up0DbFBKlfSiFH5dkYzFr+ibWKqbo+/Nf9mRlRSwCkdD/gjzZMR34zwf4OK+p
uRG0NgFpN/e48vnxvS5qEi0nLe7llPf/u8kkEugIogpjZFtMykdabCuDPLW3W5Tbznozh1KK0Tgm
sxOxrKFWdt4VX+NqWjpOO4QG7p7wLcVeVa4I0nafIB6h2Udj8iE8mklVSIxOPU37gq+dhHUkGf5X
TPFHPFDFVAsVrVwglc0IBRawalhsiShMgiPvxEYGcRXkrF5b8XGRoBFt0gGFdZnVuGDJNugaleyR
sZvkX+KGSOzmi0anhyrwL6NrX7oZzqXDRWs2Jea9L1DvcKkO+Yx7+btMrq3ZZsuG/12fPgwWyfqJ
8TV/zOfDf0muhtcU8Qlqtf42dqgcFIzB/yParVEkda3etiGG7XMVC51F0sMCcoP/tg8sNhsYMMbV
6LCBBGMnYTsinJOup6H40dXMPTGnQ1VozKCo0W68N4n8DUW00aGFk1DoPWkGYPisqNVy1kMiLHhx
lUfmZRSzgkuNzdcK1kYZX7Zda+oPEd92pDG85YXPB7dqmeVTiR04SqgEEc4PjphiWWjQMw4s+Tcc
ADT5FyngloYlMgTzlnHFRRpFXKOXVo56j45ClClUnnDeoNjXrCqmoxVZIBN89L9uEN/9/M8I77OG
DMw5yK5mSZDPCWPxyCZpS4I7xNi3mmzLdZfjKCR0hZFmsZnzKBkg2w4akBcvNJNcaRrmc5P6/q7m
SKLaX8NZPoRDtNszt0dxD6o4knGZr78rYnk4QP3sSgZMi8+ZGh9ZsYU/dHgb55DsehvWS9absAyt
2YBTE3FRCuNE5AjN7QI09GR6gO68Bg/N39MB4fC1dZxyYizQpawS39F1N36JfPRNMjxnGFFBHEoF
EIH6KqMwpiY294/s4FKqpahRxZyfhzXGL00u597c8IvErZ2g5G2KJnkdNHELTnc3fIkaIIKzQ1ym
G0I3exgiG0IVOj6U05xbu+6fBLTYiwf0aX5tIxBR2To0L6VSsm0P2M5qtDT7dlBopz1aTAcgz/30
t02uVuS7vwxzqvtGsneAAvQ2dviQKaWVgYXPxFLvMxJ+yF2+tK30H0I8yylYMnr4nKYJSot66iTn
y3k8jpFqdgDLolBATMTRVFRjytYbbvE64+eQhEQglNINKZZHVYhBmaHf5utHuCAAU/8giXVnEfym
PrA+Knb5xqnhnEQYsGnmun/RYksYU+veMwGsH7M9tJD7DT2EVwDj3CEddt+61YIZUVBx9Gu7pueQ
Wt4yZhMNDgP/NIVRlsAuwdgGtJrummX9tmK2AY6jZFcTATiFzWg8VP1Hgg6lquhDFGFLmqip+seB
guw27UJPeKDuvXiDo8RIGhPBTW/jLEftCiRObRjgBTcB4AmLa/qUwo6v7V9z/OZifCqp//wvJ1Hm
MP3e0x32CIONki90AMX0tWGHDSqIY6NxIwrlUYBytBIamHAYJEdbp+mfQr9BsymI21m+jWTE7ISu
3UbyVSQlDB0VNLSHNEHIk2IOp6hdpVz6vB0CYIcpVQsRCXl2A5qg5w8Z4vPQrOLooMEB5tLz+PcY
xcjow5YnoYjFCbwiaRETxEzkShchEDi9UoEfJTz3KXXe5bMyZSK+qQetruIwmzBoKv2z3JIBMs5u
KBGRqTyzrpRcWROFn6hfUIyivA83xFaUqzScKkoZUl7iV1Z6j1o2IYDI1K70liUsaJnbqispiOK+
2WbSMN22ppHJ0ssLLyVDH0mSJitWw8gM0pIAPJ0/dHCrcBXMiEmbCD1KbIKMwt7UGALGe98RWc6g
9dTT1gcKVg2qcbX1cBwZYLja4FzphEvdehTA4YGUuDr5wXd0dBGZKcB4TnKKY3p5+cXPT6Fr54X7
3WLJh3irQ7aWvis326gwPJhN6jTJ5gvTw4fzM0SZK3MMDHzy4uTW6Sk84aeWxVr/yhMwXzCrIj0O
UIn4Pfh+c8QCDl1QYPmzgemQDZ/S7l8owoAINj5XZkxZD8Rs+KSz09XuE9CY+ov5exy6urZn/aoK
8ax41WuyKpRO+0K4FU37rNL/uUtUkaGnvD4K+1HMEizRtQwiJisc99JHt7k5wpfbQKe6iF/S6dqq
GcYx14+sXFYAYK60cVQWwPtCwNjE6jU3rmQkO8Oba67J7+ztsQ16VyMNw/Fb6sC33kExmxWgRq8a
6wfcHjc2QSh8cMcB0P69/zYOm+QLslSpQrfc9uibiAkEUzIlNExvwXwrgIXYoG87j+jsSxdyrv0w
QdpEiPYyUaXuzz5rK4u/+pgbCJi4D3+lInedlG+jgcKFeYpEIxI+78u8gl1YKT6/cnBPDrXbLorV
LenZ3KFpMKDxTbcMPjfTmdwfVMKWfxWew2lwuddBJnZHXfVdV0P/1NnNyyqEC+atgwMd76b9/uZ3
egdRxACVAK1m5sqOWM0GiHGuzN/dpKqenWD2/75vyesasuKzZWwFV6ej0/1Ajn0T3TiFkzmFaGi5
fvXnOtG9H+dG8nDBjszs2Ni+pMbZLGDyqXmv8fzYiqDIYJ55biP4rRFuBfORvjSQCsgG4XTNRWwZ
cgo/v9pRoHMm0DZSUdcUAD4OkWoWNzeQxTGvyB325FS/ZATAhYjbzN4a/QHCtIcPdsI6OnefwD7J
QTeNlkyYyK/8P55pCxPup82etFaW4j0+6jsvoIwYduz4KtE11DJ+NufdoUf0i02iIqJ/KfR+e2XO
iVwSAlyCkkvHpcdiC4gEyTqm/CUCgE5h+t9Cbw0DuoQL0cAYC4i5KDDEjSqVwp08whvZ6o+9T9BD
XLiXP/2grezZ3L+ayX3q1ViT2Owz23xYiBu5HZ07fGoo1hld8GyUR+sTmRBjHVGY2/c/bYUChZa0
QLNfnS1BmfKajNowbtXYE3mm2YF4tKDdXh8yOcEQZAErelIh+vqeOSmiaxR1XvWK96p3elJnt4FX
eXdRVI2eg5e8ftlCRHgRiQj4nOCE1ot873bGBUdhibiivcPaQAenzCRRgZk1eQPnyhmKD/7UnhKv
QJf0Rl5SvtzAiIiNYC0QiAeTro72obL62ZkWOiEKg2dE5iVY5I3Ubguw/3pga/Qr7g2jI5JcaA/I
7S2VaEcfP8a2hiTnZQ2lQ5CqcLxtM31dBZ4a9uZfUyMusorqYxrQkDCsxEtObkDSLGrZTnCdjZ4d
OHUafhs2ThVJzilC+rCJeLfWDcvthPEqf+aCq2PZgBNPa+drPdSbmtiPh4HldMI3AOiexDOIhgru
XajbSGsbwTWpDq+JsuuJcC0aKbOLarba0Md/eHrcIp+l9a6ivNeSswqn8XeqeWPff3QVA3eUhjNm
XDBEIL1+9quXiaQaoqHhQW6SFz8ZivjMDv1ZncvgPU7y/6c3+N0v01oKG2aFvwz9Iy08Jb1qyMmG
H7OscRyPoDYh0jBsusMIqPOvxNCS6Kr6qm+kXVNZgaNcRKqY3mjDHwixc6hzd7vsMSIpfZazzPWz
1r2Gs897i6Lx00wKSc8gx1/nHpZJJhqtj2U+UEIlpVOGjo3Gvu1Ike6PgClkngisuybIIsaYEC1/
giL6HvVmP4srHtn0lBIVFtS8r1mo2i7PMc6gfkujyi2ZpbD585O81zmK32+y/BG1WkJX2iV7eSOg
bckK/bKzap/kQqZC005Sv3TcI2SwxhXQU1oBVw+KsgFRTus8t+r25TTMU0eRr5rp4ierj4yEnuWg
roDgtcMANAn5AGZWUyylXOA04QijU86xuvjU9ljY6dmAeEkPh2ihQhEJ8r/wGPMk68rUBhJ/Kk2H
1AY+suyQZ1o6JQfDjQr6v2rp+zKQXohiO1aIaNjzVCrN9fk+6Tkn6A4eeeA7Uac7SZKvGDfkNN3u
mdVW+11bzF5Ryt1fBO7PilbLFQ3hpMFKZLGCv7doWaDYkkKk1fFYOY08Y/fMrvPUAZDiJj04sl+7
SQOTjQRqDBS19S5v2Pwy87SHiQiGv2mfnhO0OvXnGgVuf/3Mc31PGA1B7X6GCT87Cjft5eFaBEpe
rEZgWyVeqTJBTuBJwOFlhu/Tvks4JZ67dbMtnXBVqUh5HH2AAV17IbBgPbwh4CZWXXoHVB6XhejC
vTvaV4yCrmUh+aqLO+hmr3ELFJVoNYaVJEJnIEPfaYMSUTFJD+MKRlKCorq100i/nYkTfWsFtiQC
2s8iwXkc5+J8mjAf1vr7pFNNCKABNUbWadPSVo13YXlQh4O5rA6781eSLiDlR8ksSILMpwHHmmH6
BF+gpi8vMvYq61BnX0w9VxVxt7ZIMVjHj5Kk0ONtDHHYX2Pg+JLmfqAM9XcdZ+hRD6pKHPnlDtSE
fYXQb6fDLV4fvZM6JF9vyEgn4GvffhMj5RJfIKF1UDXJXznh2+h/ydu+eflrWOzU7qoOq0bZbzei
pfGZYTyGu0wOy5wmwfT/fcf21Ik7f8hzoXPqU8EOAAgjxAe6ohsD7bOQJYorCR1DEZRj9M0+UEM/
ODzWx/tXX7+1mSmYcbKlyrQM6MCybS3AeIJhjE3RL9gCrPTIbRLZ5FgcFvUV3KCTtl2wdluQKKAx
1HWGWAZMkJyNSMI0sNwXY9dMB7dWV4ZUtjWoa1ypq7Qqde1YpTrg33sTA4b1fN9zR/m9tvEnhRVV
oH5z/UPKnwVD2YnTfSYjnlsyrnAA+QFzJI/5W2xKNBJ6oyCiAJ/skfJhBVp8Vhv+J5dPv6D5LtfT
EBrjLwUxqi2njFITuPn1SrYoBz9xvT8WuMgC9q85ci9iBfnh1T6iPhc0xoqpGZa7tPSqXCl+dgAV
bobp++bFgNQMrMp5vyCdeY15oyABz0sBBuii0N/p+Hn+iOGiTKZ4+Zdy2YvfYtVjoKo9k1eg04ud
lQzIqpqqvBJSw3Ed8wx4CjRGdKuKIMVM1QmdJvQhefW8NKiJPNRFFMjal8Xxs2+0fJwOPBON6hRj
B8u4WHuXo9xTnO358hZDaYCqQVtHu/N2UYih9uw7rc0leC/NAvtJ979mC2byi5r9qfnSnmo4E7wk
+DkzR59ibh+/Ofrj2lSzpnfLDagqWXdLEsyiFWf7HPcYu9/bZLyRAs0urfSA8cXI1FP0ZOJbTi0+
fWML+/gZnCoQhTnp5Qji36knfUWZR/zOSVjgpEX1MFI33qkIuazYKoE3FOaI2SFXvu7NCG6tFTYV
VkRjxqynFTOGmjouTxLfmwMNosTnxvJnPdNEMMMzVDfXg5o6E3bg7vRXt3Dbyi5hGrTxA3ioiLB0
T3Lk5MeqGBS5nz19O4eXUK8rGJ8mXc8YgQrQdCs63+eINSRwfuPpIelarmRhsGngzePy45HO/fQR
zcQYjWLZBc1F0i0336lnLTQu7zbLlqz7hMBUBFGFQsLgwxHzUN4rqw2tcNoGdXfAoIU3+9mRCgUZ
lJBLUwjmR2pBM5qmXewSJt/glM3RwdN1ohRzCjqrFKefLsnEzT60X4bXBNyayrqtn2VAf3HT5AxK
f6iuoFxjed4Ro9xAuugGQeUK5sAqEeq30TDexHWopAy/jGYsThQ/JgqU2BRaxHMVlLIyOOG3OXwc
TyOQHa6jEqWGOsAxO27+sCZZ1kGcuOyE21UWM41qG5MbZf9ECZj5cUZzHkjbxDB+MhBFKB9CmKXt
2vv5Np5sII8t49GZJSMoMEDUbV1EfWg0rbzSbWf+d3wMufUEwISbyyXl9zpBRf+pFAw3jZ4zGM6U
ja/ifDuxMrN2ZPj/GP4CgQUqaPF9NXFnOU/PFVxHd/FwSgF+VLLoMmY7J/NkN0zlTmZ2mFsBqAis
9MeFaAfnF74jmXi1LdySAzCXL2o1o1ezTXMXQoOAUj2+O3q4hYTxiAbfCMxZ43+c7jZG/ulJYXjR
75eZbv1ix7hajCXpGIW0+oAkgWc32mlEOoc8ZVBe6b3s7DgbhVUoR/ebEHqA9IKqmD0WQZ/UvWyg
P9t10BeCWi8ozBz8blkNOJveNuCF2F1EUynB+TcOycFl8h+ENy6EWrmcDLomDlfou6HnLyWJ0Fba
Nrboinuv2qZnaj+U5Y4uMRH08N87Z64mIvmN3g2CAc2r7ySsyVu+lvNn2a1nxPPBzU4d1WcXsC1J
A2e6RA5P6vtP4GRgdgWBiUBqYCX0XhwIGUDkCGx9FYHMxTrwFEC2X6BkLORyT5fhMMgxf3PkCi+n
z1e7qbQ+syZqDL/NRTdFgL8XxG5pgyUvm0F6aMrAjbRKGzWcLOAx6J+kNo8+s2ASeZ6yrALbCygk
f/SY1Nf96rgsosaSjOwEvGAtEz17u3vV5BjcYXUkc3G4M4Z0Jexj7E0QXQ1DUpAZg1MIKamvQPnl
I7wyJxpX7H+ExJCsmG8pGs+gscXgqvJufAOA8FuSISFRW9B8LjGbqvTJkMj/vNP0mMp6OyXHz9v2
PzsWxezCTByMxP0Zhaqx4OhwYXJpgbRp2qVzVyXai/ETvQQ/2V6iCWpZ8Yv4aVV/V0PnygdYvlcR
Z5XtmNJWdEu/8QM2cLPcx3WSE5iO6Dq+j1AhX6uSAsDpp3YdG5V6lVQazF6DAbWtj5T4kWabAy9U
5Lus0m+rBMZzPA1W5OqbtmQ3RCrCS6MTWUYcgjM9TbPzh9RuR1EPYUHhR+YpZnNmfWXD33NBFFkH
oN4byptguBFgi1FwdhcdaHxL+Saw1Hma/XsCek2lwdOwfXcmvE4ILC4WXOYoZ8PN7XlKAR051PmC
NOCnJpDFKdvjyYNkMWwVVfAg1UN3tJR9fSPLcBRcZpYqFt2J4eQwECsJKMNdo0rsfh4B/HEfy8S8
8pSvLMfdXjx1JNRqD8vwgcJzJjgtsfp7zb+K8tjn2ZvQA1wmD+KeW+d+3sLT4/daZ+yx8L2Hunbr
bJQaAh01ucYQHo6t0CsZi7QWqL29rujhZYemdoEZkR6A9HtJ9EVhCzc+LHafjbgUqMVaYPHkgj4F
pkxblgoaZPQO2zP2lioJlQyGBVdLS8vXhPhkiBUd0cJgMlmf2jqzOZE57/S/9r9ztsA0TUW7x6KV
PZ+yhjcr3/7ovNAKapRI3VQbohicRXmRyqGgEvAPGAmYR8sACWDLSefo090lFv1UaQdOJNSULhHI
6xEhLzN0VuCm4ethW2qtEjthkx6753zGSXvm3JpL1dno+w4P8IEeXVIxso6KOs/NBtWHBHksaWD3
2vFBc20zPcIZeTqi6wYfYZ6SG/4AJbV7jNOAJWJ8sneISiA0KTaAlrJAPny8gaV32PnJeMhtcpw5
xqdkIp8XS7pQ9tsMCS5jKhFhHDRSWZExNIpZeqsI+zFPW2ovJ4Qh3KQXwjRGOaIkwXmn1Mdz3zZc
57mnL03x6FBAR7yp++ueBn0+taykQ8lX7iPsdw0Wa4Pc1Mrthj1sNa3WEIZkJ1l1yKr3vcIYe6OL
7JFoliZ1/2jWW6r9oxwy+pIc5oA/tiBXryNxAF3tddQ1DGzcFuFhN3FbP++056nkqcJtombPRLo6
R2tL9J5151hrzZXI3iTgdx2ElZN3emL9M+tzvq3Uhn3gSGixlkhW+TzPwhuOLjF//DB66qfjLaNs
rdB4J+j/dccCCSdJ+Z0l5LAzp9APOPzPw/mmWfvGbKokYBdo5xe0h5Esb/opYwlyIgCYa42xE0Sm
dcCG4/RQ77lZi5RUxoD8YtJfQtTbQiUhG0m6+p95mA1XogAoEPUUElMMsymlWklKD0f/nHEv3tQh
KdI9+fj6Ul2KlKO30e4kzkuhhjzcjmiRTWhOU+JEdVYlWqjWAVyBXiAWF8mKa1fIeBPDAOp3XYDb
hYelxwbmvJTS3103Awv7mvzcW1FfEF2eJdcJh+Ub2GGdNZ7TaSoqh1r/le8KBq7Qd26zDk+lDuTz
ALfTFjM1VEExM3ixMz1xC+N2EDc3gpNCf+8lkmFKqdB99Ku+bQtD1KCsiYeb7wx+z5S+jdo6BnW1
EvSsNFg+BXBrDg52xW36n/eFJ/4xTzowHF2pcnUQGmKK0BrYjWlqVZQtIUdNs9Mvt3pu5Vhj5PHh
bMoAn+yWECJryqYHcNPTujJZurEeaw9+612TQWxiewEdxprwkzqQkU0+UQ+TzHB+CQAOf0PaJY4v
OrvaETzmAtvkHftrf43mm7OoUY6IcWhDCSmUjYtd5UbiFbNZgiEjGrA7kiYCUZV4D+JDLQ2lFF6R
3pS6rmpb19BX5mmjQVpvLo8ebtN1C7IZhpeYl3efcOq810/I0hW7VwYEDIn+YjW21rWxlpRFWRCa
A4OqReWZ7LxNslhAaDS4G1araMqx5P17C6yPfZxM5PycLRF07pZfpmaFsSuumjwm3SytmWq8UIFu
Rf+NPKQr1fReT/N64y9jchsTjVYn9sfPWyIPBpXL8lv8YAPH6EFpQNyRaSBSKm+SdLCfBRzejOE8
Ycam9qOqknn2tnj3iGX0/Vri4hLiVYb6cmgcihI2ZChyCZUfCFcfNPQvc0ODtpMi63WPG17YgiJm
8nMynuXVyWGzhr/WRMvPZy3En0WzZatUNTkGJ7s8mKPerCNUcp4JuXMCvG7BOO+Lc4a2ZEqEK7q2
ilF7Dr2u6P8rLixNfGWiLPHX9s8z4JcGNJ8zoxfnH6vTO/12hzSJOsgsoWbDJA+yf104Za11Oovx
CeucU4lDzUqYR/n6BqpZrfju/NdWOYgtrkM2jSix5WLqDoUeYLnR2rp0PbQ57u0PJjLk9e0bVlwM
3aijEGu3/GSevJeBPTeu9paCyKhp6FFonb4BBOlFrkpnCFGCbSMU6dgedPabJ46IX04+1pc2k22t
eR6D+Z9wGrBojTGlj5ojHEii+RB+5z3ZROP9r5imklABhsnmG8B4CFcmHd7VG5QdCV9QdPKQkBVA
B3uAE44BJ5cOOEzZ6esEFM+fqi0Zh6/KS8gNq3zgvpmSlOsLCTnrEEjuIBBB1oqEwE4pKkff+u9y
pmZgsF+8U8YEbs+uLRJ/nnxr+tptpUXNakYdbIxLMpR07ffq8b2jV8lMtmrU2gJLySiTExyaQYc1
1qoz37F42XpYwWEuxGpa0FqRyNBizgQJMSnU5CnsXga4jKVr2wxJT4CiwjWfaDnymLz4woYpMBCk
mLeBx7pJiIDAjH0VkeXvhutQd1F19EBsLJQxQmmT7IbAcOPYO3N9zvGmtnhLmkGibryohMBmj9b2
U2ZVQwaQhGpRNUajiBKbIe/CoA1vaJVS6mzMFJr1mh4fEbI/QUMzthsU4gxRUHktTPh0ydx2OUmy
bPjr847SXXOq4UrKGreaxj2jRhIwLqiNy0xjtcqZHc2eptIx7bXlmHyfrB1vJZo2QQI0PdGdj+u2
8adAl+0Ru8XPJgTisX9dr91oQjlM2cUnfBFUK+nPRQUm6XDohIlF8WIFuykGsS5N5YOEakgT2z7g
Q4UyxJK4gYzd9RyOM5EQObVZFME7ledWpcAmkoRnrtuJxRHff7K5mjUMRKXPLFXVlVKnJ3v5bVuG
cCHVO0jyS6Mge/xcAjSyGH76/z4B+wNebzBfh9s8+5wU7ox0GT5whYxwQ4RReAStzrFnJVu5i8vL
aM9GqtUsJ57ZDRbC6+mWKMNYo0Sv61PMq0kf68z7/9KphzuEvr3grCbQ7G5qM3SXQr3l/WSs/tpU
Yywpdq/gl8pNHCc6WUUj+3HbQEBXNap/uzBYQA0qiNrEh6USxeW8Oau1GfNqWUuHcZtwhwbiOAeE
6QcbUQCZkicv3v+PdVfZrKwcAza1yLZvCntqUrznd/0zEPQOpPvJELNE84J5u18NLk4EBzy6Lmnq
yiwagzMNRFeFPnpQJVzRCbsCeoPL2l5P+GHt3txELFoavNMpACS0bhXn8o73s/MYp3OONiPPXiPV
3PFB0kPkKQMCUmiQu4WPQyhWsvUjJywD6OGDV96BMnaDuk4DR7weApCYqb5Yb076WlC7Bvbqw2Ti
snJq4V2aUiEJgecmhX+DqyOQjGOe1NB/fhEAvmMv/+a82uOEkG+kHeWyw+QblOABW2WhKr2qFnqI
gsM4wDcDG2V7wI6Kmr8bVooRnn4ekZnYELxkdcrSJQgeL+Y09amHsahOVPUB4Iy0vlFFV0jsFCYG
HTVLA4heNyJSNTQ3pMPZHxwPDE+IF8kfd7qZpgDq7eG0LiRL5v4PYAZq3J6qBmUd8E5j+FK8K6te
6uqvFlJnUCkkjt8x4ygvxKyw6T8EAmBfpWEAbpNGNPTRHNfHZkWxx6Xc3i/8cwCiCfG0wmk/ngTm
RHmu6sHQuvFHEMvNu75PYnYo1Iq36zRCiZYg04I0z4lKKmrLjURp6O7o1Hr5Ei8+RF1G5t9BwtCP
WfAMifhywwonffAHJ0/3cp6l5HPuoMzmZeS3YzcJLaVYRHf+gqCxwlU482lbrIGrz//OdBbRu0x9
pYWsgfa8dWpmAl8x5R48cYopk+Msfc/GSBHleSfsJjQwRfpymST4n1D3UwYBGzjUIUl+aJPBdv8L
UggyiK3r8iAYEO75VWLDAqTc5UZyk4UU3cyy/fILD8bP1mIcp5in1zsHf6pD8NsE6DgJi8W3KyqS
sZYeJx9o3gFVobC2athJzOwEn8x5+Fq1rKjRjum0VfEj1WcmGB9tNw75mD8LVHkivZXPf4dTBmTl
/NCOzo140NTmcVF2Fmks6Wbrne1vyLlbhdETK1JDhv2KHPXjImQrWROQfliEImxsGFIJ2VlmBfH2
eb1luldbOLS78OrT7eSLo0+7q+SUjeKG/twR4BNNBCw8Ha484lwn1rhYj1UkofBuUn5MY1MdCSfr
21KokPt9iZKjh4Iy5HVRLtd6c0yAXtSyUsBBprgSaZqRdsPwctx6dyaLxB2wyifwLx+RxGRSgwa7
floucil8yBrJ8rQDfQHjCEwkr6zcNjYn2y3VMZ6di90ZvowgCBwz5jRzU80sLv+ygxVqAOI4YKO2
niDvOPK8g2XauHNJQElI4liPkXV1IwZ3p3VrJ0na7TvOqIQ/FWuhBzK3NEEybuiytq4iiOkFczUk
hHI39ayB2/iDyjmg0QFhyq4+SPnEUp+w7AaRloPAkpLVHKJ1Xm6cYhqt8LrGcCgSSpMlth/W+y0w
wq8o+N7mPb0VMnR4pNbmj+WaOcIHVVNYx/QI1wy8PTbVc9/x1+5QVethzgT3dAFQMJ8PRqPTNkas
7PSUKvoys1uv0G47AUMLqY+bWIX1sLAoMTqxmdpt1wAL1K41+dkxi3hzRwRmMWs+i8P3iQaaj1VN
R5bW5HTW4QGq9wu95lC7VNCXiS/mV37w0GBEui72yynvBkWt8RZETSoLBTWHbpv7Ch5lBrXsjt12
+4WKptFut66Iwr6arZD/WkEmk1jkaEud5BodWBfc/+Vr1BZk2rNQyrHxhuBANS/eA9vBBWXpNju3
OoRgtQLOHoqkD4q1GDy5LngrFbg9IVMxfIKkSINMm9qm3mk13QId8THO8fyEFpHik9qvfluMCxtJ
E27ZxhJKtY9XojmTRLCLSK92MW+JffCTqZrxV+8CiGO0SG8BA2nEkY5fy5f8ZUX1Mjlax8y1GWdW
zaJ3BFyXfCQcMfzj+A52v3HJRP06Zz/YOHCCafjIsyx6PKfdPb3ShdSG4Tzzavx/zk07Ce26wmDl
Wkmyw1v/QCt7e0DGu3TQB9+XPpOOk0RIu7XldUCxWC4Z+r9Xf7M3otZpOmHI+BkrUM7lR3N0Gx4A
9HdeDC7ajfhYPpoeVfICtLCs5qndZJf2GqbRcj2AAMtlMI0T5mi58Rg/mxAmQynwe/SkyePbM9Rv
E065ap1ma8df3UryDItYisVNoFAAoggI4ttbvCN5D+bZhG4sOWFXZ39KeLYqgX++Ir3JEuqmoWK5
i0MN9pagafYSJVQ+4qkbj0bbqqj0ppzA2S19fhTC3aYpoownH2eGTTaJn0QSwo8As5fczk7vqe9I
WSV0Bbv78VLC0yDp2jMDnFwIcRj/kw/n5FImXJCpLIKcDVlvDQTA13jkIsk2vzkRrm5j9v9A/9OH
wl3tqjDEmK5BbLUbUj9Cr6BRL5ysEVVf6XJXc2SXdvopeZsj+frMJ1P0KDVDgZkOnFpP/kbz9T8v
AYmLeZGt9G0k3JGoQB+GoXTNCbg8IOuscTcgtzXb17dRk/FcNIIln2xvgCELZpvFt3WgL1BG6b+L
e+dIYHc7x341zeVe7E8pbG2AKEfGKitzc5FXwwx6xMgttsj31VKSR6QpTfroaZNNpWTrGohAMjK0
v9m375vpTW1RdE/rAcgRA7o1pqaR/nTtz4VqCL0yACBpRYXhJRsfvMWwdyQb/Ijd+vtzJGUqGaET
U4P8DaU4AlzM3ulh/3FxiTWlPyz0+z/GetrhW0qep6J6uTfym723tV0bXy3y6JSNdAiinxGUbDWq
Ey7xmCWyFnOeoGvHeCfrndDIUpM6T26OMuiiG1ueSgrOapdu+4sSORaIDmOGwc43it+NrSb1Rd+q
a3ER3pT/38Y2wINGwRGYjeQVQbuT2nHBN1G4l4mNYuGPwsLq6KXE/RGAMeCOOUIkKz3ROkyEbEhF
J+lsKTSgZRBfasD2Kv+JpuQKxmwzjEZR4hz8YsBN0pE7NY1geF9MwVUQfkltYDrZE/PtHUWiRm2W
AURNjmn4pUlzeVT20aXeLw/crwNag9GOLLNbHhBfJBMBTjohPLES/iWkeESBABsmDPPI1iVdZm5s
wCkujgyUjZzrHKlsvARAvTHWcfhVbPOK87vrhTsDTPOBk7tpWEXXHuxXbPEVN/YHJhuWveM1TSQ6
LE0ez+hjekZZVyzsQT1uUCdzBNedUinyC8NSz+zycKyJhUJBmypAUHZjcYCwLSEIO/eE+HSG5P5P
9oZQusuWtyBvKnSgUBk5JgJnwbLmHvopy16nm3XylYEA8SrR7pO5eNgULk3f+PTcTfZvNkmhEmwg
lbLWHrslnzchk2lKt0oMQoTwJzRybzlaExqKQTui918xnpSxlix89UWPIjCkgYbwtX9vfeRkyiE2
LYM19ooaja62Kpql8sexCL4YnQqurpJghYD18/Zi0VeNTSyfd9y72VYk9mpcd90Ugek0CVCwtydo
OQfHbDiCt6att81izJ79/EzYHgS7snC+Akau8Cpqh9y4S7JiDJJc4VymAUbU7dgFpnxJ4aaGRmia
/0IpJntT0QtUJbu9rmNGeb50eX2v+eoWBs/fxmA47qsaLppv3Fe+YlWAnSla077B9ZlgT6myK9mT
IOY64whrNgREJ+0N1OujkP7St9sAImlsZe7pjqHeoJttni8wflijyK71Ewc5SqzBAa70p4QdVbp0
+YP62seN2bRdsuxjSC0OEmV6Ts5LyBk8avCLri91gOm5cDBM87jFCAcOSQu8gYG94Hiy1bZ09fVf
mAnAxs3Pg+0PlJwzDjPxE5v0y2FITh60SGAeYgheZsxETWoEwc+7WwJciQoHWxvJxecIVvSQ+aW4
Xepgd7rSISXdewpwVNwJblwNewvjRxRK2Nw2UwPRX8P42Dtq+jYdHLOWOD3WpxyW5ePLJd1WRhId
IkH7zuKx1Cn3UM+IRI0npFC0X1zJ+Q+iIg/UpuG5pIW+mLPNemHxuxJJYxb/5s7Wp+lnrF2O3cBQ
iIhSaZdYLoyph3MNXmBIik5Hzru96bJMdQc5rjs+q9iki+3zs+mPavBd1oIyn0R6mLrUitx2EiNr
F+8dyzFonB55HbwANW+ISxLIcE9JCTt/lgrY4vlBae2pc6WGObuYVLhtSuQBk7Ap3vnx6MLr3ntp
0A9AzwNXNnt4a63EJIF0UflCoHOnkryIIMYFluzqVJK7ngIemSNs37r5q0Jf7xhjMudgs/MOO62E
1tMcaiax0nfXXXAWnxypN7jVmxB4K/nMeKvGf0JXo5rj9V7MvH/Qn+7EyFxMd0vU+lsDPQ2xMnqq
Zg7cjFrUV/EEuMTcXGqHvQ+EV7nP0n/XC3AIFrmcZHEA40NcKyNEjvWWIQp1FLRaX1g9kYio56JE
Yp7HGItDsO79L2AbgHGi3fqHXUkDozvqOlPQ59oWjo4hiBgyy+c8V1NEXwp5+kn6NJtBhspCF6SX
fmBC7JZqEf7P+25ENEctmyPAFywNObLzXLRq1nI5FJFKQ07EEnNtA+WB2a4+Rrrf1iFWg9fIx9RO
GgJ7q4Y46nCC8fnyvfIzwFOAsvdcBuMVsC/cAmIh1ZD6agcj7fEt2fIbAVtExQaEv6X77/ZMAr44
Uz2mJkBaPDb45/p0aKwEWB4Db4+NNm9tBLgJWSlexVy28vvjxllZg33TFQArEYgcSAhgvQgI0mq4
0t+m0EQYHDWWsG8EaBYCNxu95xxIez8bolnAKyfzUQpmI1+X0rWC205rm2nCyRG6gXOwn5Arep2e
XknuGDfjBSGCr9RB0+G98TgIGEhh+V/0r4wFdv7sEeYoSKV6gTxktqCIbyRzmd9kiS1et7/wANKY
2GJ/Jr2PXTjGPYybSGIQAFOpGsC+B48bMsUD2T4tS2vGra/ahKMro1mHdfsTh9DQvJsPomsfzAuu
fWZ3UMUxMn03qbEF1Q6gsgJ3aHbV28FygwvHjvJagiyuUHwWINei33Ql/ftWEeoVdd6AJxfg2fuy
764E1rEv51dndd9dSlBjx8ssKIzk9CtV98lpASba5mGHp2V5+AvtDv5SyQUBtIVNuW6tPzmpBKrT
A3NIqLNojoXsL9975juFcyA2LPOaBnDEYi6HX93mAgc7LELIVwgON2zHcTOvFMIoei/N48E2W47e
ffeXKieaccF0rqHG8KpP0O+hinCpoxU7EFRyiK3SRu65MQ1hgddgMNxFIkkyuHyFklDGP3HvNy5O
Cw1Am35QH7DOiZMPpKNWBu0J1cV1Bd5a6U2k0rgDMFVHMF2AVNeYSBdWrye3gOAcMJVQ8xNExspZ
/+KtkxYVzpoonoj7ilaBT/al7baMEqklVkVLCoLBVMZuBWfOn/aNn5QzFCFwMySvrYSHWAd7cb5I
xU8/0lciI1pyytZM1p8DW+wPo+nopIFlRgDMYAWrLYCPJDwTYcu5Sq0zk6a35mxzGyyKeShXHLkC
GeE7yTIBzx1SobvUlya996S/siH6tfO8Ub1Uw5qftJKQnG0W0FNVro+E0oxNTNfUGeEebNWp+pua
0h74/TL8DlCcVaKfG1Toqga7kiba4/QMLyTnVC/gbpx9irqIdhqB4MkhJYm/HesVkj3VAJHMr9IO
2BvZFyHRO2mWC65vph5NpYmnvAWAmcDPbrFXGsFbHSyzmOPfAW70gXx61qSC8njiNZvpMERcP4+6
4hLyDebQhgcXjhTl8iHQNFG5nMcVpcJheVv4/aFso2F+bzZTELmG1UWJIi3E8AEqIE9T5f4Y6yEO
+nTATXxd2Rm+wGSWpAqUx/e+wi8qI7RPmcM/X4EsUFtaBlL949LY6Mks1r1JkyohFG2oAGNn/JM9
Wdsw/UOOhkE09Uq0tHEBb+DIUHSIILYM3oVikPH77YSp3VU8Wworn6KieRGa2CfCZvFJo6OLJkFd
7HloFY94I4Ut+SauGK4Y5sUWqHrLS8O0m+3IfPmnQlBYoJ4Q8e82gENvo9xtoNf4pgtKc+b2XhWz
lz7ICQuIHjSZ/2NHFX5sAplJnanVmwJuNsJa3O2DhRji1DWxzqwhAeg8GYMvthmnHZPhxI3WDj9U
S4aDJltkZKQE6HYkp51Z4XrvpfygRxVddJSdghxu8EqtQQqO0BuvGNRnT3GNjUe74dzOU4ZNunf5
1Adj8D6udIoGzAvdg5s8pVBw+ew095bJ6EORQFUwKEZJ1RJ5MHx1BK/Tu9UK5/pXtcWVslfYsAMj
fa0ZGc7SdjWW8B+0sn0lGT3mUmLtJXforOTYOZFotFO/RL2J86PKh1PVUevuYz5W5JCo1FcEyuPx
BhNtv9cBCYwpW5zDwRU/QmrwPTuIu0txpZ/xY/JhgDPXheJwCBoI9iknf39MnQMNlK+HBZlqWZ5G
PqiJi2oUAY4xqUDvtgL6UUO/r2sp0rqTVN3L4xB/WYiwgY4XImHIKg8bYITeiUWayKBg+S0yEPHe
Z0q6XH91OmFu/bRy3yCyKZ90jGMbZTE1NcH2Yl3wcTM9EQsicfMSVoAQioXeFrg8n6+bpaBTM+m3
WamStkgluF5OUCt7ClfhV733Hyrz6cpl4pD8WNB9sfDJV2/uKLMjdcRN3fH8JRsLI2zqG/SyeIsX
fXsRwLsYajYYjulWj6W3vURT4rNdHhrstqA3mlgaaEo4UJs4zW2lwekn52EexT3qFFE8P04jR2Zn
Hgr+qRdkHlQrw3QUILNQNf3UcKouAmJZdNdIZ4FLbPKFSgoWnmWXY9jFWZbmuAuWLyXrQIDpBbu4
W1C9qwWODoEGRsbYhi/8ufg7OQ/3g2IFMqleWYHY0HcLaRa80XwRndMO27rHg0jNxnq2rXr3JuYF
SInS6FbbfG/Dlh+uK9DYz7tNn5e7Vozn8NUqeK2J/Nuid/oEPqreiMeAWQLe+YKAEJHVfcihaNWf
MGdk7i06Yuf35SLOW/ytRjn9YMLiHz9fqDD5/HCJvaTxaKv7iJfaHl/prQnvz0HW8oHCpxvhZerO
278SBoSIj84YktBuyN7wISYMkPPaqaZsquvKBZDQQqA/PG6zBGXnXlUaRPRSIInO93F8HjLBd1pp
HcNkxFZfah5RjilFTpWKiN3FrQTdTFjihwLb0+LG2uGNIXz++WiFA+SJfi6v8xW2CZxW0zuQu3rt
MsU135kJsI3KwYW9W9OpZLFkVJUIihA05kNwJEjUxEZsrnRqsBMuuYQuIq37bHEA1vB20Gp+/VEs
G2NMOQpjlOEPGAouZIEBC46lfVyIgrsTtKQPa5i8eW2zAp5GZVTvLY5bOdJn8ENaVfK9b3pcjccZ
lp67/OuF02qvYhv4tiHrL3bdnHwFiVwBQCsCCPxa4ywP8t9xuvz4C2aHLOO9l1HCc/ztsGmmNqKQ
NLqyF2br7EzRLelquJI+mgee2XvbK9ySr7H9d7GR+zr28GI5JgOvvgVhObFxJxL1ZCTvC1di0vYl
vxY8JYut05RueY1XRYNXp9gOm6kvd0NFVSUrr8AFfNbvp95RgEfRGS43avAzkndYorCyHhcK26Zv
a8/Jf9//u5blaZXxY280WhPJovTZPPH8ZpK6fE8LGsS6a2r4gqD0fxtDLntbbREf0qVI9NVCj7+/
FKznhzTeD1WYQq0kjsI6E5hpMIm/8cf+1CXhyhAvAltV99IvbEAu95AlmoEc6AbRQm22EPKtPZDN
nKuVGLpps+mVYccHppiI/wYBBehuLfRUagEp+TdC3hgjfcGPCA/BmgrUi5TvSNuu+zJOsKbHGQLU
GFcoDS9eL8sGOYIJl0Zw0pO+rH9+975ZVQFSBnxlgweurYH+NTRgKvgBFFA7AQ1Pp4PbTl92+Bgm
gVqUeNpeNf8B8fZj5XO2wU9dHQQnWKFYvD/HCkdXa4Y4Qg5sgHZ7kDe9yIlHGPAiHdbgal3rCIZC
Vd1P+EhScivVhuPdENCCeNxfa8s3YNGyy1BpHcfGbLbMINjUhm8xOHt467WdTAvmCm9ULbYJWYUg
6JXnET7OOYligr50fG74ZTU3T/DP7RdIhRKMrspP5Eg/tEtyFEhLmH8vklQOAuxmMpviniKxSwbz
b7qDcjeMmvEeBS8MaJOyUUCY8HKQ3xDhVblNFJWnJvGITTCB4f4zjBmvaPvHPa8wbiPGTgIjr+PA
lbM+AVBSeqlKArIuEUDjUQ0nYD2FB624JKDhREWPgwepsqkhVgGF5T0B/yE5FkvWojTD3lpD7sMI
bc0qmgorO5DTxLm5oWA9CTMCJzAtxis96EhRt7LYjLXiNZg+dp3Zh4H3c4OtwtFqG3MdH+DFMSLS
sTynMO7RDSP4jSBNTjkL4VJq8u/t6C0xvJsNVXDV2JnRJSQ3meHP1JZnVq3eVr3mGKTD76TrwAR4
5pg3sqo8eiKCIeJ+SZcD95YRTnUYjw465ZsQU2O6P+9m3htAdYVwxJiJF/MRx6xe54P+GHHQxe+a
Q7rwFtJlTqj8kTNsyASBvPzYOO04Uci3RrDB8IHjWD+ZqNwIw9c5T1XbKSEfIMtyE8FHkCGMQNIJ
3vRC+Lm5MGphH6V9lSYHUPIwJA7QkssOea2vdKO2+4LN/RjZ/CvUz20kYqmWne1nqtH1Q2eXL/1Z
ZLPxRRBo/yHz//88427TO55E/VKr3dNGNKXGXJUe0zG2dXlQKTnTc+vF9avdtIhBSAO/ujVgQa4c
gN49rTATC9uZqGgRBOvH/QZMBnYrKJ5Q2PZkIc16nQ5LXhIBqIcL69V/sQmZyHc/3rdPdot3aLh+
CoDQ6cu99TCw7HOe3LUdgBIwnIX/ervuLMYlAplAXsE0T8v2lzw8hJtf2XRv81dXbmTrYF6OS0jW
9BcfiLb8UFFOVIDNdUQBmxBdv2Czi3oVGqkQqmfNSihjEjwFq7w0WwLPrMNBkRCv2o6mrnOU/SuE
+0H0/kfhWsKIHYpZh0dDpTYUwa5kF9hYyp9ypuV+3Xp9QmfEUHsDpVD2ygEt53C0oCnsUhC9UAUp
rKN7u9QyttkODYABg9NN+KCNa7uXgHOaRpi9sTr2j0RZFX+lj0Lyi7t2z3npO1y1qc2WddaQfAIU
JKKsNtZ2pPYseIyz8l9JF6syUI/2xRxZ1hcK4lVbavVSQRYfvdXzuoyiMuZ9vOC5PmXQ4My27n2R
Ky2FKjVC1t6xhnNxIjgzubQfhGwqk1xWROfj9f1EvP57ZIawzejkoXZrXYsdRFrwXP/uvSlwDRGa
0N9aAnRLqDNfqyxujeqUrU5NMJn0yJf9nXoK3aswNeIv+93SSfZVRcxkNDoTwttkQ0NG4bFeStlH
vhQVPoxOfoWkisyY/IVTIxUA0K7GFRFTGKVRXqStT67IB8FDGe7/w+CpKeodXMZykDRccd8slVXk
El2QdfysW7myKQHU5KrOcEgi1O7NpPM1Q/BsJ8z/pSAmFWYtMH3LCHlFwyYAmmyEnIbwhYDWm5Qm
NqQPBIh3V1L9TeNmmYNfLd328fDUJWtZ/Tqnqsa3pVVu5Lug7FMU55vPr8mg1wYHE7rErH/lCNbG
sW2NQpky4uC6UC6GqxEQG2IH7r05Mk5+KGD34e+wYxJGT86A1gCkfnM5xzGlKxOLZPxFGCJc2xU6
5cXvxNuKXwDP4s06XNGYOp9wnSVQ4JK5qh7SuUnPLHS1UuCNraC/foIMoL6pqk4+/3HcgYklGTPf
i4vAYRDLXTHGRhOJ27qjXMEAUGh6b7IOtFHCH/z4aaFaZKm2mAS287zXjht6pSeLHnWuGBwOKwya
6nM4kdJy5RLaX5rrmxI/l9aKzPMkCPKMCH6rbyqtcxApPtdpSQo4J28eWXcbo/7mDZpv3l1dxH9W
kchrbGlG4zcPl/T4fR/q+Kl4UIAmp6kR8wXbYKioKprBmuuoA7k6omb27Hp+7zgqT3o5n4q80hBr
5MTrcsniZBYecReFqb828EoimES27eW/dGfjT8K8ooC2BraC/T3ESp8XOKNJfb3y1hN+Ktcv6h8P
wV0N4hNbZGsOKVuHispaYBTb4sroX7Z7W7IWDyyCUnOiPZId/cHkgv2G9CILeXWDXpLWrT5RS+fN
JH4nLGS8lJxdIL6zMVvfcuh1clC0yNI3SQrZ6/2P2+2ctORS4Hne2vaQAZsUvoxIP6QtjsVVhGi6
nWmnJCKd0/naKZ44Qx8Oh0JxzzWsfs0Zd23MKaes5KMUbVKxseYOKzejPgMyBRiCeXv6buTRIusl
6rzyUU9/Cb0YD+TfJt/TGVfvy5//ux1cN8URJ35+ncNj5hEN0t2Ri/2aD61cLPW6Pwp6PiwiK3g7
JAHTkLtn6AOSfoqOmNJovrsHE8mnRPhBP0q1l9RdYygbtCDN+owz1viS4HVZN3xG6MNvksETT61v
fQ/lI4EXYew8PXuOQCKcI7n6VJ0LkfbG0qTYQT5X8uZ+LgjUxaDgmfLn7HOAgFtIeuVFAIS9RyQI
24mJkRjJ/Rmaocgq/u4pIm6sDGDkSq2xLuQA3sy19nP2M46V5MLS94fgcqFWBP2dUrKJM3aXXSCk
pjP5NUxq6GatV3jPCzjXH49lUgWGX4wSqazcntnvt+jAKp1AigFDraopFbVMGlMB45xeTvWbIVJL
DsSEC4alQwbqu4wGxJuWaM+Xx5D7x8TYsHzGngjqwOwmnBNJQOz4Uz+VM9TZRhWxQSxGNmIb3TiL
wa15SZgM9YdkTHVgoG7S1YIqzCzPjj2TAaDGWtSrqaTaX0LYwDIPjRPyQSujHcxYjkZLJRXwzemU
gDnAZKtcTOUs4a+1MnJuKGYCP6nWSfoAboO0Nvu4moz0TeW973VhzMoY+3X1Tw8ymBpBesU9r2Ih
i4lUzB1B+u77dUwHGTr4DiaFoLRU8YcQRDH917n1jZpnlUn7JAQ1d4XeivKFUPR3YGZHxj2gc6u4
wenvW03BmCiP7ln/JsCW3TLJHEj133Rg/XeYXdRPvI6dQpw0jWtvFGmZ/ehxwTMY9LlSAmOob0BU
qymsVL5vuP9v2phsq3H3QxlPTDICem2uj/OqoPzyyNESazuWVdxt3R2D6WdAD76SL1fQabkA9vHg
1i0sPaN3LS228sF/Qt2rzZHBGLLgIi3lYF0JcJUzbBq/VU802G1XyFZ44ZU0s5TfFzeC/nkWQfQX
idaAP4S2yxkICIaicUq0FmTY0liyFsu/rDLaFZwQyHsjxbiHSIp8s0+nJIbBoGZXXJ2SsUHBkfB7
b5xCfLdNcehaoboaPksSsGVLFYxX46hleCMVYF0gPvRM+7aKlc5GnRop14QdKA/cAc/x089yWQai
9VE4eK1ev7ARq+ypGkhe85lFh6z3QcGjFMp2iguj24FgoBAQ2y3a2iKRc3L62t3Ts44AHFHc93QN
AATSdQcfcg8ujVupoZiqQf1qtdYiFzAZSJn+z055Xk3NdzsA3CC2cYA+u9W2brtu2W02O6/SzFjJ
y4oCCH1SRnFFvpOyI28q4p6VTQ3NNhdWo+315IDtr9D6EsVpC4B8jvlCG37b3e0ECNr810kXoV/T
oMUsT8uEYwszi/8Hot44qPK23HRtBCBmHL3AEthWFDdu1o0RP9PAV5yq2S/6sCUu6+6dJF8ZAve+
KPdalTz/Ps3c6KBwywGHKSnFo3GSiMEPD4v9IEmvzGIN9AI4bGqiKpn8eeSvnKY34Q7KXcesqq7j
athk7UrhZZFmEaCN0FSACo2yoeNjLXi6tass8MqABcNePqQMoqRqTpqb/nwLqlujL+/8pccUPHM5
omnmZnGcWqlDFgPY2be3FpdIbiNOG8QM3cE2jGp4R2HUOlwDd/e3j4enAHvkfetoXt5u8PTzklO6
miKhlBSh/tmaQyHmVPLIToHvshcyO2hVplyq+PVDQnRwSvwek/KDR0RPLvXEeBE9Xh0XVArbkUzb
g/rGh9EZPxcwP4XcT+vIvaUSKAlIAtRZwb/YOepSYocX1skq1tfFdg+d7WY41CnliXINrnWNIP19
cWFGvCpjuaqmrib020k/taZ7DDWIaiRiokB1pqfRZ8HXinWG6L+MW2OR+j/qNaMYyz6JnWvZDYBL
E38A2TAtzb9w+Zp9n83VnuMFur5aaIgO5fyFbhjtW2UvbhWVt87DRVshiqQdT2rSZZkD8LtYw0Ng
d6NFjp7fh0K/+2gdq+wCYA6IcSOCaI1VNCaVr79K83lJf2zuLurhadClApcwRtnqsP/vQyhSRZPN
dhaeFKqnNwHqWiUjAKp0qf0jpjSxmYNCDErCf5rR2d6lhvLcm0HHh4Jk/7fKpzR7gjoy25MQc1cO
cXZismJ8XOr8r2QIztRgmyFqohFZElnQvoXlllMcapSpECY8/MMKoLa4JGhm8pGnB+iy+fhg9/fo
uAtlSaLA4X92iHYxbjMD6LHLx8CQPVJSvPGgDZoMao7tkOuaKem4QUcIyQ0nRrygWS7qqfArI9vv
0g74BDs0l8kLGw1Xi2RPGiBan77V92W413/TFG7ylalBcxj3Nq3JzqIWFCAm4UN7laW+YTUhk5yt
TBpcpxUynd4wQFjMEYFOtyXHUBlw9DJ60BgSXhjlAljEDEuCpCnXxLcg80jxVl+29kPNtm0ED1qT
A+kAciiyAFGHpIlrqRaTTsH0Mdx3XpsFt5rSb/PzxOM42odvgG7M7mb7Wo48gMH65j9vv5XwVolm
g3CcKmITw4u21wsRpsNDfSkFRIBr6Ys3L/AfBaA1Ufh1jzzkusATvkz1YvThVYovRtdz9SFGOytH
PodvnLRtF9nw4Iake8YkojRMbbryB/y/gZdBDEuR2/GjPD/oUGcilk70H+d12B7fKF3lIlnwUyns
7ubY7spxKHtY1ufynhlq3/rKiXOosNu9lEZM/nB+zUFWR66fH8UAccKx3TW91jE7HHJ2oJK3BdFI
o0RCRQ+gTicFFO/DLMm19lqnozkF9Hht8/mKw8V9+jsmB6kwiC0E8eFD1/OhMVGu85hVCVzQ71ox
0GEStzVCG8JIbJl4zhE1CqTop7yl0CE1SppVgQURERiyihnxgyVnnsUf5WPaNO0Qx2JbXDbiWCkc
8FNTKhd2NeUgwMt5Itd1CX8SQvTl+WhAjw1xJ3tdKSXLD+faMWoC8qV4WYaSKEFxS3r+0B54m+d+
7rkFBCO/nwWcGCXOirc2P1KL7GJeCJPBkzL8kAyFce7106LVXKxORynUwSjEE/q/w59yB+VzyQaD
DePiJ5RDUVn8+23BlMAocTpOy+x/5gltpfFHCKG6L/UgatXV+DzkzYTiNDta6iJsuH9qiF4/DSMF
d4DTmdm/CcyJp5JHXNLYpv6qhqps6OdSTuDikevzB6bT7S160q/UnLsy5dc+6rEGz+uaNkeTXKe/
0Bk/5Y6Dfv6crZIxcfOoeU8Asu2xGGRrkEXhKjyPO5d8cXyb8yRDdQ/BLSMY0ROma13X2h6mH6MQ
tLQ+ezS8Ik+qlJa0eTHuT6ux1RoW0pzJEQqcEC9VvXKun63QpYEurkPhl1mvdQ37rsr1dN52OqSE
RBC001qdir1luLVWfzVSUQEoNr7AnLpSdni+Se+SUB4kGIJZut7uG+yudXKHmnnmPHzowNUItrqO
XcjiAerbpuYVBqcPYU/yVSrMuGBBCrrp0Y7xr9FviGHcljH30zvn9B77zL7GeVBNRRItrSpgBk7N
Ova6spdshfYz1CFhCbub86Fiq/y5iLEZyNp+CV1jtSu4rPQh/fTKd0vDOJ2c66iWEJYU09+/76RX
WaXWMDtGLKZXRif0Ci2Y8vwmbAAJLJtBIU0ML8Hbm1xVAjR6YDOg+6ZFcStoy/xvo3eVZIQY2/7A
4aeIA7QXKTB4t2MBT4qHf3oWrWKnpwiCx+Zn64osbQNTCNSShCFW492r9/O1iM54cBNSJZAvqkVh
eUn7NJ2b10xFJ5J1MgKKzjUjvuf9mTzlP9CRkn8pBO3wD91FrN+lnV/KxPfyB7/2v1XwJza6cZ+2
9zFwGpRuY6mDUGqKgwzhIca5TdnOfCRhkLmk4UyVLa5Q2dhc1cfGX3mNYcuymBNmm7a65cPOUi8/
rGla8IoA+bB2KoS+thZbvxV6BVi+XDvXLqBwqbllcgOG0JmJbDUAxcI0j2OSTYPyxs09ANBXDHJY
xR6DYJ++Ycr57UmAH0y/KVPaUAg0T10S74hWM7oV/5RKqCfxPqtJKwwvFL2O8wudf1dk6uEhqrDR
64PIqtgyXRwGLk2NPi3Y3x0JvjH/fmfkum/puYPpXj5ZCVZwvYTwx3ZB7jwy4N9gcZAbyS7pgAD4
grzAsoHXbD8CxaFljkd1iP4I8v8AJKQTyFZ4GTJyelL0U7B5FD3oMPu3oV6erPVmpRZm12ha3PDY
lkC07rDz0i1m+gFroybMKpqIQd43UrYpasq5LqYqFk2JCsP4F7uquy0JlvY2EbZkptOoXAAMtD4h
pjEaUZSN58A8qKHZpVMdwVjU5DzcTDzIdD/SXvPT6BxOLQGeO6eUyjTqAGu8qK3tUEMN9/hnbKBL
LDBt6zafAyZ2hayCq0sn93koaUsuXGdLImy9MUPHF/8EISJLEiweXQutFHaKuu/qEONl37la9cLz
9lrQGcql0nt1jLDH7pmwnWlzjtf+AIkrHNBn52znO8KO4q2X1sqlAvLyDjtaaLTKF7RIxKKHPsB2
gjQ8UM3GOUCmK8Zf5789sUitCAvjOebrcfEZw1sUwwBP1vw+gT2UxE7YWF6QDPLEhonawU82DOWi
LosZDxZvGQOjmlR2lYeaWCYkmM0f6N3AlHAdxpeN2nNpV7oExtOS6cB8IkIZiCv9Cn3Y1FKVJWv2
M2b6FPQMZT9kO2Wu2cPLkdXIzrz3uPWa6uKdezyGR7UjazZNChgzzjmPwkjLfZD2FFUOq/qj2TpZ
PL5BC0ccjFUawF+UKJTufg51VmMCYOC5avpDPP64wwjMDR4Yww5b5dxSAaKUtvER3FdMuJoQxUSh
MmU+jUoPFtp69ye00Ak5ZeXiFpJgSwIi9TqAs2wIJpmTxjuE60HQYsta1Iu8f+wpKmRX7m01NCnv
COxX822ZSkPlf86L200BLNa6ncNjctpzcdvm7EAUgL5zycDOc2qzPYUl2D4XgZW29BtdEsUQNa8c
csADgmNHT7ey2rig8qkl2AdODqCWi0T4fb4qltVkV88gqNPMY+eg/ekObRkNbpt1i7te/S0qSC9Z
05lXcbdq36Xg7fwyG32+YXr22JZUG8hzFBcgcn6DzSjqcRhUJ9mpbwrTSo38/2CYFQxQ0Fe9+a7U
aTnzNqUsrBhKUEuwIvQS6okMjMdESlEDuepsfmS6wil07mDrET2JUupTscj5L1dQG0L0lNTo8SFF
9Xu7E+5CDqWtay3cokPwjAGGn6Azubi4inFSuSRTRtD6m0bcN3lyUW52u025iDdGnQe4SW0bUenM
rzYOYNDwML95zI7u2DNHo1gFz7CcDC585pDw5KE/Qvg7rJkobpWjMSa3ORDg8tJ7aDOeXHjlPNK/
y+/9zoZD74oVbPeqe0pW+o9M8huNn5QKk22HZAyojgeId4zPfqeqaCWN5USAf5B7eYn3xINiyR9Z
VDY65+sRDzmI+ao6iH0K+8b3DLAqk5EUIml2hnzU1jU2fgN4o/QGgdxgQ4elmAfua8O70Fp8+njX
uCdW3MzeFD0o3aM3vt4mTNWUqvccAKs9wVgux9XqGZPNdv84KuYiI3/i3RtTiGxM2iHvQsRCSkE3
HrUiXWBB4UoMUrZG+gsct13l7hvJQJHbjmqxFT1mD0C2wzk74a27w3Z7j0W3cVJ4Q5cSx77Hn4Xe
mbihvpOPQCV1NzJm57Tv6qjnzedZTgKYJxH9I/DOjKN4ggNo25eX82XcLO6Hu9QmSH/ObP5k+20T
jVbpTYxxCKU0XDvoUsiBXcqymNlC6ot4Ywur5P7/ZM8cW1FxaLac97FtNzxJEYw3V5UL8yTG5OYn
oRmh1JgdbyEVGUJ5vMppd0JjSfJTe2SeSPMpB5lGhJ3a2NZ6VNXENTLyqIQQWpn8AuVYQlEnFtQD
+OkrqI4zPYBX+vbhg7OOgNYuPyF/JlV7ZDHgJobNKG/N0Zcqjazn+4xQpC2wF3TJ5A/egKqSFhOD
qVrqURzr+SAb5YrrwN2FefiNG4tEkEOdNFqJhpod4Z0ZIsiC/0LX/QROdEzUcJIPted315+JSWQg
6iG/o6zZR4Uwl0vlw/YJsv74KfzaTK4jNn3J36/IGabY8bggPtX0Zqfzvfzs0HHrzuFHSOKG47IQ
9zZUEpQprrvdVbFIJscUOn7WW9sZnQsf5sqw/hjsUQuKucZup507PSy+GYkR8WeIM57vPw2SHiHH
KbuRXN2O0ICDse4dl7k51F/9Vjre+zGnilfOYGoDglpoe9NCATIAWlNH8zBH8Ej7njBSv+t8DnCG
g1ip1V9YAWyDOJfjkdxfhQucnRfI8l9V3Y9PHDYmCIO3fIvzfjt6Lhq6Oot378ifQyrJ8yO2z4J4
zT4hpE2Y7CaqSJ6Yqwp7jMG5XR2CP3BHzl9HaE0bJd8jKdX+nYlYj5zqzPqxKPcwZWk5M/M79NQV
C6Beyhx2qKBfp9DPcECb5Ylw8PsWXRCEg3PZrQC3oQzRxSle8fy1o4fgzzm9dA6iYkXKSK9/NMKn
kBajXl51Cn3upZ8ldlCBN/MOtHgSVgOfsMA4r7nzvLRQgO6YG6209rWUDT2ADcujutxp7Gja/oBs
zHBAkcQ1z48+EvOL56hWTjIv3AYoRtWO+6/vl1WAHwLhETZ05lJnGhL4m87r1aE4XNoNLbGNhEGS
obhhaORa0KUK9e/YVxd0ozhto78vaEb/3WuCqIwPU/FGAsl8fFmbE8R7Yie0KbSKh7CjMclP6T1g
WCFvF9ywBUfWoHsBNLnkVjbQBL505UOqo8OxlRfmBXkw0XDm+uR6S6yp7lTAPKfu+R8EuK+cfvlk
myEqNZS6ObVk7ljH754O30k69TtYyTCgA5fshf4mBcKMF5iK7V6HcRJlGrcLlES58kAHozIMAQ8n
/E4P2JBfNuMy8OPnGTY/XmC+RWVn70a0GITcql38fmy7JeFMJJI918XllDdL5ak4Mfvf65/ZRHU+
J/VINPeUdXMHbmlCUJqRCv+86wKXwYnYxuI3DS4zxNUO4bVYE+sUl7U8/zxnaJBCM5Kbzndu/H78
ExvQ3OSqQUE3A2rEGdK+66Q/XwyyLB4pIRof7gNFwrpk5Mxhv3KOLr5RIAzUdvTZ9q36v9d7GxQL
0xwDuXv3jsq7MfiCURWks4mKnr1duRV8cDUXvwCwdTftRa8N2RlbiFRg396usbJmC2BfdKTUxkCi
SB/I7HAJCVXVt3YSdVawOgqaqYuMswwzKAOE7ijXNoUJkA6nzFE3+VeMSFEZ7OsR0oFSCMF3iqGu
JExRqmflu6fygDY7SNqOBQEcgW/uyLCThJH/Cj068m6J80UEVQZhDeFbSAfyjbag/hB3qHjppqUh
Phx/ghs8BJG5OTNMgJff2G0bxzSl1ripYkRvCjucgwyf3CkuKz9+b1lV3him4uQhOMDAcJ2O4O+j
zo3j7syJDSRKHGdzfAQ913CkbEOFcaRZQs2O2WWkQXgw8aY93YRS9PpP0egRyRNb06myKETWyDGk
Va0dmbDqkT0XUfkS4gst3eN0PMaFItD6d9jHC4yCb06YnFoBrtqDkKmaaO5Aw8+8m+dh3hdbA9uf
PEwdMlCxH7pFhue5H72oU2lPP2zkOkTqMVd32cML/BLfHYvzpkXnYy0GjpJV2X5XxzU8R4WAe5pi
4Hcrt/kew31g2X9Cn0YvE6cAONBH8CHiU4uWZ1Z8oCC5l2v3OvRQ3twrXDVnH/megj8QB/fYJhYK
kFA1W6qBrCEX/vxzFO7aa+JWdeyf0KXED4DcZb1znFDKjuxgKg2bcsz7s3USSOD4HPzNNGzzOKSr
tjqGjrRfY0M7BNZ4H1OQlUxpi4A+yCIjwPR5yce7Yg3J1i0IRnTlk1sVF9uKOOKbd213n0FgxD/L
ddYsBmoYppDW1mloQ1JJadbw/Hn/6C4ou5CY0Wc8Pl1DBDvTzkhRExqZxc2uPyXwq+dwPU4ohKWI
BXi2qpjLCFNq1sJak5EI93XYI+/AdlOBucEUrwa5WAZyB34hxNMpAYgsvlJxhf5GNVrWKBiLV4/+
7K2pp0eI0ICtV9HbMqbxZmY3YdPQPyUeOpZHETJrXrdS8WxdOBSWT8BpH5fgzqvocNUcL3A5EcLL
wREqpqaN5urrJJGNGba3FuhVr2tARJXL9oWsWG/YSOKBmyqwfm0rddH9LUtVpAp4DBBrGCc296B5
pKaFVEBlW4U4anlAuoAgRiGVuE0VSLioo41r7YZHD3ePgEUGHQlDS73G5Z4h/5IHVNo5ibGbQp6M
G1r77clOEJinLAWFehFku6fALPcRflZG7SxLfMVAsjly+BN72707rrERRq/FmbtOTHKOOUJlQ33D
efPpNPayM5CtB1tMG4JyOx4p6Z+2TikKSX8WoH2I2P2WkhwQAYe8k6dmLIybFmGQleAdUrPtVpRX
AZpluDtdJp+Y6LXW1M0DyCyM6QrljQIXdTykFID91zhiAd5UXR4crZbSN7mghLitIrOkr1azQvQd
C1C0TtB8VfZiZWcVptzagYOJSxbsS7vmcQsJl+Kfmv/kSNnNrZ1YgfDp5IhjrBZ1KDIzTcL2LgTH
vyPe1JPWBxBTkIcSAIkGRGA/y0lSM0lxyfLGuulqhcsVbTsvkoAlYG1lZIkC1Oi3LO6PcR1LzGJA
AIWxjY9LPLW3kSA0mEAPO7FCMbSak/YyvjILzDxI5AaN3enp4W75Y87v17imTxUI7mc5DXRekPkJ
qYgr9DqWEYwjeas28yNl1HEaSO3RIZIIopfACpNLY9/7cUMEDj7g77NMMyhexdw0ELh4dw9e6VPS
QQMrHDH51A3W9eU+V2qyTH8ZQRrhhvWFQv3PuYRCjOAKbj+X0HQ9yZ6nLmQcOZ/7eTITVcSikxfW
uvzhpB22maygLLPYukg42elgZjkYUQ9NEd0QEDiISbfqZXyL4c1LCt2zl7YQDD/p1Ygl5sjSyw6y
wKEUeUCp2vPQjH8Iy/E2770crEvbaIoUsSe6kNlz/V25PmCUSGTpbCcd8+ylSUWwZhpAy+8YwkAP
ZJPJSwsY6r1Ef+jOc7X0MkKelTldjkqk4/ajhB5NTzUkLUqHA/o2scw8Xazv5xh5wwRjG/9qfTFI
fciVvyKApFEfpSg+pxrp1cjgLXlr7iBbW//ogYCqGgx7wTwGnwxzar3qe9YBPZXqnDln3e22nhUy
8lkLCb7VHC8qmVbKZ35qQEgevOzw1p+1iGu/vSRGtzp4ju8D4bLewUT4uUjRhpeyUoKBUc4zptc1
OglulHIMhFS+7ZRwQq31OSpyww+oI7PgvmbRTTWM9mJiiXyIcclnOYZhQiCzrvjV3PTlno67ecrN
UQzXL4dBhteS1Nzlxu7tclqdmqTjZduunoDJ0tqbXJsy4iqKAqnJayeOOo/W5UrTYMosr9lt7pGu
pwi6Zwp4ghg8Rpk6uLTQagkI+nF1XcULyBqZwbR5iqvf++pYNbVZQopt658O59YaPkT63u8HtFm+
+G+pKDbl+UMLRnCdoHgz6PUefuwzdtjL6m7wwpSrqEfBOXaaYEP6vxKSYudqrIyzQ80i8ANXnB+7
6kH+zQHBb2J1ymFps8rcxNG3BLP5TE5XPs9Xd8Tz4zIVYPvbcGiwOk2hGmSneyy8kMiCDW5Cosfe
qrvTmoSZ3BK9x0bURLM0fPj4kwDzgoJnIdFsuQ+kGOZeXVC/Ch1O3ZVbh0/XRvNeP9sHgPOAyw5U
XmWabDNigfzmlJXZ8wf43im4nhcNscgShAWiAWD6j+8sG8tefIyKKG1vUv/57Z5HLMo5psvjsYtN
SplqKmuEivnIDXPOMaCxK9iFCUImbJvu3UANuK+5WZn00gOpdiH1vTWaijz9wKyo6/ZpnDBqlLnm
Xt5VrfGl010k55pi0/o4EIm97mK6h/F6dgZSnHDzqc+7St1akTIqoLQEU/osetMB2hpBpGyUVgbD
0f+zjhnfspffOk3Ej06cdTM24RGUT/8gwjyk2clABoCp7qfRMziMGOI8E3BlddozUfSwD6074QSk
w+URSts8vC+GBOvAb1okgihWVyvE3pbm+OHRYa7Hsv1t7idf+2IjXJEoGW/Q4UVKBHb/6nPleTdy
SlZPJ+dWKAjKU8QNzzk9iZkJOoVrO5dVO9vOjHq5It65ctza5JgxiXrhz0IMcjoXh4y3d7gWHTH5
iYt6ZMZlYJ60Yi7PIqRbrHkb2m91+rh5c7DfqN6jnJ7k+I05PmFt0erdRC4YAogtAOOSfdsV7/ag
eEsR0Hi/6tqKZtlvRwaJc1BA20rp9PtSmlpExVRNkmZHT8nimt4MjQpSV0UZ0mAZyO3YLXwuQ461
khS49bIFBathoBLmSLIZCBnHtdvfd0hbnZFRsypEnwdShIQsRpoT7fNSRg2ILi2PEXpL93rBP9qk
CcL4q+l/tzwnCrNk7eRMSN2JwRA0u8QobYzUiqlY9TA5hPAMLJsUbC4QqMFWJgG6qyQYFvADGm2I
HRT2qPXwnthVZA/BjkzZQewg5mokjuqg0OooS5BcFrL0UfCzof3e3cB0MeD6owl/BuKDbk0GLsJI
PD3SVIeQB5izWnPAJTErkpSAgWcfOsbeKyPHJiWQhZs9/1v+sac+4BZooThjSWbaJ2S7FzoGx3wz
wPjrVbEwX7AucAiydBh3P+BzLEOnoiXMjCAP2Bm7xC6p3IrZnqV5Gv44mU7MN5nhhDXFG0Uu5jL5
VLSulaw4/edTnImwdVokg4U0Q/i7q+/+ZEXhKra0II+HtvDbcsnpEbWNXIq0t1K/V6AcHzfHLP4g
iVh0uf0yVTrbxdUQEkubVDtCAjzwcyj4+Eu6IpFkTbQDHmrj6CDjAWmDBaj1SvdWpzhGHJtD+KFx
CevdTHfRsm0hper9qCCe9p4vPIwjTrSzhMnXiuptWDn5S1Na2Y3qXubJ+GvpejuwTYmlxXNUlkNX
2M9Yz9M/Tx9NyiYPoQMXAZNDOhdKMHHtrk0GQFLgGGTsV4PIpOtXZ3GSwqSXa9GLPgz0ye482vXF
CtH08qHaSxWkM7EdTN/3jCgpd+u4gGEKvd2pSn0YyLzcLEIWIy8tuydsP6i1QvVnh5KCfDgXTA7e
Z6/kqPiKjLjVVftqtAxPVrDw48d88uN2SKTxecTZY+OgDAAgiLDHCPravp4t3ix3Q7xmATcmV6+K
9mvgOiGO5m3igw1QuSnIYRKgB6V8+CFkw+T9/FZjoDX4VAQAJFQHNZ8FkHel4zkoCqItwueDW+el
AuDu7Ha/LJ2JgG4cKuxWleTEhOCIPkpMSFgG1iHBrAPdqCNiu/TiS5ujAFpsxIuOk9vmRJ8Xels8
nGx57FLzNRooAJE4vOSph7BahiBLtmMp10AO0uaJjaorQgZWGAPjFHpeDhWRy9OzCKsmM0zbZBT5
h2IYPDkc9MrrgasGU1MfKi/w+YcDyI7URIswlYUSKuFOqHoNcxxqiTZch1DY4OHEX1IlwFdTu01I
23UwvWecp7YFHXFR972OYnHPo4j2P7Ko3KrehyfW6Vxg4POmIDhNZ1aAOgLo/ijSnuuwJTch7Z4O
seM9uFeKx8us3AVrqDmhHxmSWSD8zxG9y/HJ0K3wUVjgCKe9OIHpaIVhH0QMD1vIHBSfah29FXg0
9H1GeuLqiXJc/vx4ILBq7fANECoOAeGmygpl9DEXm1Uws5yEzmR/r8mjMxsIM8C24LH3dJ3gOM/8
cHEBGqgg4xUoHeJcg6U50wlJ7vru0R1/Ra2nULr+G9oKA4wk7lg5QvkNr1x8SmjSW9GQd1Lin7YM
AXJBMFspgMxSB8wn3Z63HYOUZEhiYSIE7Y8NJ5Bfo4heiIpM1XdHByhXlEJsAVkrbyrtYekqfs4X
GIJywnNDfAULbYMkSD12XTTlW1l3aogzwvm7rEjE1Hkyz397DSoiSvcd0Hn5PwDjzmxPk1tk9sJT
qxmOLBLwSsFOgWRRlyvKlcNnFENkQf+U4tcVPnOG1PpU/41ThhuKs3WNiKItTesJ+EYDNTX9eTjg
OwidNabXBNiTGsnDgRCsESXFgKbe2AHpLpQi5iFUXMcXfvDUUmb5kkglOriov2np743ifLIPYA58
AngM0+gxHgFw7Fb0tRedN8FKGWVN6ROcMTrem6bMQ0xYBI+rjChBE5/ZtZB6ygL5ZoLh4T3uI0I/
U68hd+byFol34AKX1j0y1AbQIvT5ojLLQ8aZL2Fs+izQwETB66iGe4o1cM/GZCYxpuRxI0uBXWey
1Kb57OBCBmEBMgLW1DtvlqD51baGMVs8CwTJJ8BplfcosMvgJaXkGee/Yk3eMgdeNU5AShJxz92o
P+celrqcZB9NbLSZTPl+nSJOBfCsK49AmfCdhNKgHfTGlWGd6UTaSnasV0NJ4VqMqEE+Db9sgg1q
okOv3VLLQnw4X+rga0826udnfwW7mELOkxljAddWlK65LyA4I7miKQjwJkZai5GblJJgVZ3DMFlL
x4vyO9XSDJaNIVHYSbp1L+s5fOU1ooFad2t3Pr7NNERbafK8qvluzx9qoANKg6BSOXYGETYNL5ru
Ph7fUpdcsaNO/VFeAXtNKRN2esgNCoIy8LAXNSJu/17+wrHG27k3dvhfl1mcNg/vdX44pupd0YFy
29tLydtMLxuWHwvQkqsSwRgHherpyw1KPrDuTCnzlLTtCYIsOYct+JfTebyF8ram2pdhlw2tYNwj
QFhrLGCDFqFnyIASRrrMqfVnYs9aeJPNpuSWtM48Bhz7osV95Z7x0T1t4uEZcoEac55+rFdPNcoH
6v+u9n+1BknsTiqjayv5LdCyU9fGOL5pJRg5zIgD+dGkYBeEqMgAyfZau65BA13OQmAQEjC+VaZC
zfEcdnXqtKzEkmD9q/c2Yl729QBwejiGDO05wPD4O4N322IJl0/76k3W+ysky7DXQ8rdCq6hGEz7
wx6aTaLE+NfSVOZVbD4s6fPTtDf9kTY4wDkl+oKGFhbPcThv4fu7QfNKC/U0BP8BAQlDAXURj1Sr
rNhWBINEKNnhgqJ9aJp6mP0pZIKRHfBGEXohLY4X1j0GlCyl/Fvk6VtU2Ex5XMcV7vSytXIH6Rs9
fkZr6wWkIy/SQ4TPGrkvRTsGgGEonM4jdNsWo80Xlc8xun9PwnmdbR//E1k+YYcHUPvo7b6xjh0y
HJ0I6yIKxUVpYY62lV3U2gYh9oJazrw6OKYz85ro805TshwwTbsPVswkcrNlGW+yx1xCsjBZlrCa
NRcxRnVVeK7YJfG22Ja8J/Uypf/1/w7giopmDxsl65U8ZZ1SGmbjvtGiyXf0iDL6fFMv+/8AMh85
gmngx9U6tg1/MEJzkQy2lgDJeb4cP1XDWCoAIO5T5S/RrKNm7hWwi7fsr/QqzSgCCu9gFFCDt8/t
zPcVhcsghGZg9gY9r+nkjiwhYeykZFTkIaJhgIPdE8bbYKGkKfKawbBg/45eSBB1gI7FAc1kGfid
/mpknJA7nA9+WJLsrSRwNWxxYRgxi8BLbeUt2/UD95fq06CuttxxOxllr7yztoKIoIx9lcsh/Dcd
JRyjmNzDLPZACpIW451pVYSR3AwM3sjupqr3EshfHUBYzM0C9EjsAQ8FoNRrWcC/iJHnWthPxR0l
AMxTLNzqCirKunBhprGh+Yn81tT2fCaZd9JE0bYrmeLT+qfy0p98JlR/BIYavAaGjywLqsnCa926
Ie0I3LM8jdm+cVwpGtAb3CGaSXuDNwFm8TI8wTNmxRDUiyjB0vzHKltbD5kZfkTHog15mfY1rQWq
s/6Ghh5aB5hA0KyxLEd81b8rUOpANhWt87FykMh/GPnbi1LK3nn0SyDgDbVsSNfnvgwRHgOUeLHF
Pkm9KsWDoDPblrOtii3JDhlmG48wU5DBQIMCtAwyYhmJk9Qs3vFbaDBFEHiNIpaP7aupn1anN1+y
w2+dciH6hMKk2cBtN52Ts3YcnMJXmDQy/9Jhf9Mpp6X5AT/PEQuFLf+hG9e4j012BAdgD5S6CsHF
jncdY/yXZAY3OpxoXZPhU53LKlHLP9vBD9jfdm0OkdC6fZ6YZIWPlL27ZXJOEQVHgAjkdx42Lf3D
MeT7jm0f0YhBqN2Ddo1y0K+leJK18iLYrvxxnyzDQf4cRn5gPcMJvwKD3kWsrm4oFSoxlzY0mOBN
beT0utLddcc7eWY6q+xj1ndayAXFKSWxCC0bIwFS3ig70g8n++E5jD/X4PU8BMwWDtJU9RDn1ACd
abavkQpw7OOd/3MSg8aMZWGpZviYjAMEeb0vkWeNzEBE56ekY3Kp/V4Kxr7aWMbCBCJIA5UHBRo3
gZ8wLg38iUD6/V+WR8VdQy/YIs4abSL0o2eNYFrVT53lZ6r9hxN8X4/G7AoWQadWADQnwPCKQjiV
Aewaxx3+q5wm5eYOydC+qhHqBK89txVk8FiQ6aRtRyz3ME7nOqFL3DT6hQSzteBSec9GUaS1TnMu
cJ+Hy5AzcVu/USZNT3axa4BI71Em1bNSgZw8uY06mtOz/uPiawklZpGTvS+EoMQLruOKH0eYrVex
TuY5n9Xqs6H/Z6x+g3ICI/4FQw95pOJsig0LY8OG9h/FVb/ApdmEm6z28de282+orIpmPINHr6cF
tiU1ogLbOppF3n+WOZ9sP6LRt7zIT5QQMVe7S22xqC+LHsVQRk4OMLnTlsSTpeYK/QUFrtP0cxmR
7OkM+lCyxx/Tcb4HYYVr2AKPRBhsN+hs9YpKRD/112jUhvtg8DE0FDvNtTgyGlVXhiI1ZgQqKPiq
z1iHKk0MByjEKd1pfVgDp1kHJmbUqg091gpU4kXl76oCzyzIOUjcdgGKpRLfqhgO4OBqX3OwruxX
gcyGEHffwKqVTpmIfMeoJ2wk39VaUyYxD/9x/AVtqV8e6iDfdv19H8NUzgE0sVplfDEb026dNdXh
xVAxU+87Ho31wClU9hrHCP6pozb+12fHRDp8w3lrCuDfTdN3YPk/SYWhycyy2lF4TSQDtJyVZElf
SbaOvlL8L75uFjvQTGFV1ucWNqQpISFoipr5onkOmCtrLw3XPyAvvpaR4T3bciibDrUAmIEpB8jo
XUT1qOl6IiIxkBbV0YXA/vflSb0kQBMfbym/G/6zZFIPpoX8N7Bi+sERsPW3x12OzB7A1f/bGrmg
065UWdWqKc6yBEQ4tDRY5k0V2Rzbn7vCcinaI7AdTt90z/YDCc3AvXcuTCRRBa5xSblI4Vi1hIg9
DkRfMPxmcx7RbAnuGpbm8rMmnlsq4YysHkQfxWWGYq/CYJLGJKz/5D0lFAPSZo4Q27P1r5qYvuIw
ZqIXIcSKRIFEbpgbkWzjArPbW+3oEb2NrvI1BQeV2pyWpOsFH7H7Vbfhu1+QCw3/oWbQlHekEEiU
g5Bb24ipZIvDAbCSd2/wNvBNxOFKBHqdnfBu9t0yi5yMuIAE0bf7MOOD8J8z1Hm7Isd+E9ntLZPN
bqap34sU7Z7RPyR4JcZUeTBoRBp88Pl9/BUrq7X516X+DEhQo7YLI8nhpd7+3Xyf/M2LAWXMYHtI
WEMeoN9u63RnaxQCEgKEfwGjAsib+K2g5Ed7XoZawZs3H+LFTT1sGU0msIp5m7DenQRG8y+vIT0h
U7SFxjmNtVIvZ8oIaJIG0yWD+4nC7vRfteLialA4b+ZyXQdnOek20DfQDaWtKpr4wvpObDiimche
/tx8RB737K7P5gmhrJAiIuUgRsf+g908vLkjzT8R2SWaTG4LSd3qseGA7RrNN/vLoe2kIz3bqr+X
U7J/OQLK8ZejEDpYESsBd+3CtGAWQUXgtNrRahxpB+oJ/mLwCI4MpQpSrj07v6JGOew51A4MlOQs
qQQ9kQ4bIa8oEoZfcWNOuvfT9+/sSPOHIN5QzLNv+n8WI8gkeKnFiB1L8bTE0xapQ9lGA9P8cux6
7eUlIx5que5GXZTDea3y5MH315vh0GD6GMeCSOXbiE+Tntj/iOFnw1UdQe2uwoKVJVOZlwjo331R
i7Vt9O1eJnAawmf1mx7hK8p46QhWX1a3t1mKwe19JTJOKEY2ro4i54P1TYRyVg3mojsrHTHpViOZ
w04wXN/clb9TPL92EM3eyTfQHC8fwJe1TB495nV+8UyHBGPG//5G8+uH2aAvwGDnxaV5cWU51IYZ
HnouwUhwFvOmGWbN66ECiVRtWvcktW/G+F3C8RYS1t88sVs8QETkSSdFdXt5MjOQq+ve3lGETafM
A5WPwNyIFKJNRXEsthWZNxBDG9l+73M7FqZqj6v4+AKMWmG31ft3ny9C6CdR3xcUYMZ9Be73U80D
lkRj39GkRI9fgjsE3anne6sU6zy7pjvkpkH3hM2paY7+gwM5GJMqGzjCxURkynjH+RlRwH0dC168
w4+w1R/K7QL1kCYnDHoatJ0PDpdpVQnfT/RwfEgUudouGAJGcQFMJoXbJ+e9oAjVikaNhpTuZT5S
VOufPy8rrI3ZYrXwDpSwY7aPPgWC9wwwz6y0kP8srANr0a9CH2dn+5rpbTxie/gDvZA6hHRu0SkU
28YchQrNXdI3T9BTFLV7zmhu8A8l6FEmYxYLsnV4cDpCRrriT8GCwHiOARJniN8MGm0irVOLi/S4
4fyMVEh1WT07MTVVidzBultfejjGPQp7srQYmLabw74chgsG+WOzw4hyLPvagn9K6NqBFm1Lpig5
tNnvgO3OVi6LmjkBs9MWgva8OUnonpYKocVdo3FmPS/KP5mhcCPmdY14DShor1ZDch8u7cxpRBlN
gjyM4v2HktloDyuIbT7Wz2zXVSgND7+uoAGbdTShN+fd9nDs7XS2CJHyGkdY9Zn6pCO7tOgK2I7f
NCDKOzw9e/HaMUJH/UMc4hq9x6r62NLkh4IlondPkk4g5pFB/ETfqU2KrR48c7zpOirN2588zUFV
URSEOUiYQM3g+oEzX2/FogAiCBBzLJnJgOtlcURDhuw7M5TohYgQAG78qluDlCXP8D8mM/EdUtIT
jZiWTqIZZKDFkIbxkzB60Ca9zLG0u6cf8j8NzlTExoB/xNlh46nvqEIKUGLuDlzRL6o1iGBrYKcG
AeiVIUhPMOvfzC7Ske1Mgg7ed4xbsrLpv75ZocrVYxLx5hgadFoBSBm1AFe2Th4Y3XNewJ+JkOzM
9GymznBXXVi3eGPN1nglTvpGr0mFeCK0sR/JGnAC+d6tmiacaG5aozU6cBHAW2KO3yvuqnH9ZlFq
x/he1D4pF6qp94pmlZE3ADUtpzp2J8phKFcHcScia9StpzvjZUH8jNOONYDqkoRGV6DZEd8fZoSf
dXAh+miJ3TUyQsPnEaofyr8FYgzcwX4X6+gQ/uuRxgBbswRELTeFIVqkD18AlLh/HNNmtScsXEPJ
RTR1eQJHQJAuVdU+leLz8KCznYGUhSJTVmgypndnkRZLMCl1DPOVKOA2JPxQ52fzKLMLZ3AtuKLX
WXZLnoSIkDgsUPyFfdtGadNhfhYyR3zAvu1zV3AbhlqXH4iYZYXoj5DnCXSnjBAjU/rz90K312PM
8xRk5wxPntkL2fS4wbyONXJHLVsNcfTjIrXfnrJSU+ZkJhGlAvuwxr5pE37tXL8E/zDQ/ohBvAiE
9F2v+bn+EczUmFpQII1Zhz6wSoSvxmma+jzgX/kxeTlp558BB6rZJxw6EC85QbHVR2NTHD71ai53
T8YV8DDgOZsWJfPZa1z7cqEaO/zOVylaeSNLEF76TN9EeHwtzuyZVIpE9r+RTKIEOVfJImS8EH2E
+YnsoySICaEwiILozVwI98vzs63QgXgpPg7oJc6HyiGwHtr9f0Yk2xlS0tT2+yFfvL+IANSP1Ihv
ncMnhEU87BY2vgWDxoBF+ePFffcO6HZUB7s/fmQ5YGUBjhq208kpXomkUUhGeesvXY0edw/MQi9Q
0FdOvXHh/pMCxWS5ufqD62RZRGPpYziHSpl4/pFRk2JYaUGEkfXUzHKJzXs1wB4WisVJ01L0Pr/y
bBZfHEwdJ4JZnpd2IqgjeQb0UPKCEpc1fBpwM9B0A8u9NPjhGpgnKEVXxQU2qAx9tU2jjqOMgtUk
Iyqo1SZUmxLJJNdypj8t3DofGIjkvRjW0aQzcR4rguueMLssihugrKdKQVW+oOEwN8DrQs7D1nFv
COKktYXcCNWYVp3MheU0snpvZh8Aevk1Cc5W3GHVEHaWWYuHIeC0/c8TNuX1a9bwPfi8UfDrBPJc
GM0M3zbCoYsyAXmwW1gnxXk8FSMdY1qZIoBQ51fEWwiTCZ1qBR/EfKi1TuJYHjV5haR81K0akeft
4CaGsIpAebEd5OwE/kb+jNJROADmg8s0dig5uBngW7AEuuf6/ahbkJWBfDSf3TNuQW2ZF4Df0+jJ
KsORKTPvIE7UnmkHOrNzcbeRSnzJbRnTo1KqDtNVCPGwsnhRg+0TPlrMGRyiYwvOwDkYnG0Ybgr0
4hd0t+hiLdiLJNZ7OdIA7n72FUmoDyHA6buFZBs47UQu1QH9Ctlk9cFOzoRuYHiFuoRVeivKNw7X
MkTmBgzcAeWC0ZOjjdS23Wx76hSeRiF6TJ7vAYKvyhwK73y1Qbq7FccxpSt8OTIwAO9OCdMcjnxF
S/HnPryKMaTukAQVidSdpvGVrMEfUadoxZ5TRSjrCeH4C2FORaMVns7vkiS2RAH/Va6mz2AmDsrW
6BkwgIf7VN7citdAadFZZrnQ4MCBXj3cfNEXY9XUkZdFbRNAS/UA6KiZOJ/VMrzeuaOScpt3sAqk
t1Bbgcvix8AGwrS10/KEzYWR7bR1J53F+lDikWF/JGF4YXGskwMGgtgAEJfmKQKyQv5QLSfOnA6s
f7CVzwYBJp0LJrFD2AD/W09LZlf8rmjyGx7bSjqMK6AfhHh9yq1oQJ+l0VJN5lmuUSfYNslu114Y
Af+zcwTHOuTUAHf88OUXPEd8gCJVqcJZZ9jQUFDjrPJOlHdYl8jPnC9xvl2TryWyixX9WaFYLLVy
T8ThlF4lmAhxI2pC2vLTHcCo+lHscpe4XcjfIXewjDS/Ch3OdYKo8KX4aaxGpYkl/UsvW5WD4Oax
cHOPkUh+RjUCKGcZGAO7or29J4cG8KzVU7cfqQv1AlCdIUS+B5s0rJ+8SY2wxD/x96nKnLUhZfGF
/PT0/woj1SjzzIwS3CxnIbxU7BJiU4G1w79EPKdOhrDRpwbZviNs+C7on6mBkh2BvM7enWXHCeng
mhqAwGcjpoaS6dr2vsvzhvcyzoojV+3HN+5IoTJozI6SdAUQJwPL6sX0mFHHLjJdkiXK2j61nXlJ
dn2b/Tv9rra9RLvAge5CCml+rrfHDsnWxbmS9a//2GhZjc9oLg7JLMJwRZVs8qwuHGPv+zXCDMh6
T0eRol/9EqKiHnXzdsvar1UVQxRuGpDXQT41V4X9qAlBOnc4YWEElHjwe8wDKExcs17H0F1Atg+D
XtIMHWffUcfzDiEpd/Z+0sSiNnnTpoQQGL1FdvL+j6oBCSYKA91FjB/CK/Gyg9lzCHJYOaBVhSNr
LDHBmUYu9K11fnw4HYIB8U0mBuThxuEMw5b3G0jiTIhOum2gwBtp4aGEe7XKlktQ2bIRtiCkz65e
yHzL/imznBNNB7xl/85D3lNOX1A1ZlLBWny4Y4xWBA3Er8NiCaqxv2GY/r6lg/RMXRHKpSYpFHjo
uvru0Zw0DkbDXx+0VYsrpG3qTSC0Ocs2DQFWy+sY0uGM7reGkgbcuCiCq0NHjespWuxS95oHS78n
sMFkQwuV7Wyr8DBC1Ag4QUeOd7p5yTWOJQ8ifuMR+YMk5Gnq0Uo1j8MsSfHfz/gE+cFOX3cADy8c
Z2nwwNsyiUBdAVvlbgbxFSFlnCzRvveLt5uyy/GGOrRnRyX9qO++rWpiDin20ryhAb93joqANYtC
QZ6KHwEQgimvZpMYXKEcxRUKrzAraC4uoR52z1iR8Q0YCw1Ki0VfFve9WEXn/ZjFzb9cm5C+biWP
1TMgnoobgJRhQa/oAE3KEKVKvHqxRD8J4DMO8nEgO7zz98Wlr50z7M9qsJSlnuh2Zzx9Dl5AGZGv
D9vz47RDTyxvGquY4YVxm21SrYHGN4ZuHkjXVtjfkBf4vEIoBMOZnMhMqLp6NxxbG2aheFted1vc
D7PfznGg3ZnNjAWmE6XRbijwwYUZmXBXx+CGVltD9c+n/7WC7UxqQcvk+EJnYDLTXJ/tR/+pNJoU
NMiaenQ3f5eXbgRqOrr6kaUR4TPBe954juOVEm8oGRmv4d8QyFCiFD7GT5rc1sjygAsYn4iwcBow
sRJxGWUfgp1Iq2DOF1zQgqvlXGRYTiWIkwnfZJRLNBDPADH8xhFJZxs9p30uB+bhTCo6l9nzGrwp
+eAJwpbipw6nzhOB3suc1UZ0wAyVHjiw0hTb+OV2AC6G1F6G/kkpZLVLj7ac+1Pltz0PBVluqR1w
qOgBhIlv8fsaDfhcTYU6qbuuvh6Jzd4r6U/6GlpjrfqwyLZwbuwLXYpQJ6OMGXysrcZ/h4wv7P6F
lUp3dF+U3jXOzbVA91KfNcDqbdy8/Jb9bsMCT7ZDdaR8UCpmDx1xmsDaQqo8kY+SSBBPZX7gbdo2
aiHl12Meb9SHjagZLfNMToJFdSazLKMOM9WI2FZCbB9f8m9kmhL4irHBSbJGGnS+iXeSuPoV0Rvc
cwTAwc4tXsA/j2TIJxEgc/IyBoqcaACizyeHpwN1oZKc7xO95qUMtTQroM5hBjgK9te0deTVADhZ
bEOsOqmtAMZx5CYrckJZrSIlxUPulgOo4KmI8v7CLSRjoxFC6ZAeOyeJO91oVfah4vq+TV/iCOjL
qDWOALM1KiURH5zpqozK36bEIUbuQyRUaij803wDsplkcNfPSR3KNfulOs+kReUCNz+f+8wK+gxy
PXzcAaL5Cao9js1wvRFfkvHiI4X2b/2MbwZoS8p+wWYLad3f0QcHag0Rex/ixWx+ku4mFWhzsCiq
yh9eqbRukYadnd31W0lRR0TABgy4B7vsNRm+lRyQS9FZDKQsDyKOXiaHD2ShTJo7ByYjNSXKAsWu
/h4yy7WIOTGk+Ncms/OVRd5TwYt4GSBAdSXJxG2JNiRe9/YY6w7yfqdzxRfqP8+mLTkOzN+waaY6
7XeY3UiQhuIsnXuw78lAzcV5Vhjdhyr4A1gsecWE58Gm0Va4p5uReI4Sw4GDdI6UyFyct2O3crUS
kD0kg7uOKG1+hnYhYSDVhGy1gOYE5WkYxtkr7Ln4B1hCPc5/qw/Xy48qkfcytRMFwsb3qbwJdDrK
ea8YtQ7DQMskXA0qQ1Nxm0IJQjnL748nQwCT8BFjHavSzJS/a3B/qvY6EmTXs3UBvZom8keX1Bdx
7T/iMCG8ASb3uhDV5s9KwdeHh0p1ZTSErqLc5sDyCv7cFSdywTCB5W3LxZXilqIOmAM/awnxuA7l
XdMi/l18cZ/YaZLX3S9Z+pdvAOs6dtp0ct3S72FR1CJuzNwj4HrBD9sgnJ04MPrDHVWaTB5YwQV+
Qv5y/d0cRVb1eRc2uFK3zMfEMVjXZ/mAupADbGX4xbjCrFqzjN4pTRoqalTOkD0BYViyMNnhBEiN
AgeTFBb5RxXMBHWxSri/9TiQrlAmfmgAP1zSeWzeUaw8N+9HYzxdjOq9I4WEdg2VzWFJMhKCRB5L
6ekod5UqBKmCcWCbFESSFfLPH0QuUASnpT9FW+zzTlQTkq5Zi3ZZVRfBxOru5KEvpvKdxc89xWig
1YsN06f2Nobnxx44A3Tx1+Y2IyCbE63Zw8RYWDncaxDQCV9mbwta44swNktJFH6dpS695/xtyg95
6U60hF7fynY5l3J7EVi1wdfPPXX3Vfd/BLOtXd4PBeYM9LIVh5pZi4k+wyoVFwD1HAdYLG6tze7r
cpOx9M+CGi/qonozzrYNqJbCnHbmNYhhPaaBH9/tCNMAXHy6khlHvYbv6y1Z+iWmItuqi7Zvzfj9
L1ExN3p22rq6cXur1RWkwRtx1bO7TZI1/UXo1fnFNhl4F991llfYrGxXyc7IQkLkG7M5y5Du45R1
MxtY33a9jtCwX1sYPk0x2XPzJyoNsTrOA+g2ltsp0J6fpV1OdNk1Wv58mSkugIe/zjUAM1e1f1lW
wnsnWl1zzETJctFqpTRBM0J5zc67QgFXwM9qI+ompcZhGVnSf0bkiaOpA6QdLoE0ARZVNwFYW/oT
zGlYuqFaNLmCv3E6XABpIPBh7b+aB34/esqaICdY+s7WaXIWb16TxH+3rrg9NLbTfVY7xYoFs+3F
squvzOspzJATzlv/YEjXc/dGNzNN053a9umjtdaH7WwoSmj2TcCzjyWzJHrgD1Favo6WkPJnhk20
IgeHmDInMm89Y/l2+rnzcMusB9bp237wVViYLA5QbtKecg6p5pqfWsnCCSlQO7O2bsNkPxe1bzIN
hT3zrnAX0EHsUF6rhbZlXHXxQ+NnjLb6KU7vrz8dieypS50RvVbWEK4bNTTkXWoPmBuXcL37bfIr
6LIXmfqom5CaECDlX25mq7jZru5KbPM5y6vzuC3IOSaANbQXqmWr1zrqAeF66gqW+xCBvWS8uz6h
WCV72UoUGiyhE08s/FisGOx9YXxZg2l2yVb/dAcNL46gb53oU2GVOmb0c9caKRcheC2pffPFRtER
UVPUkMxyDXTeGTrkiFR1ZikhMH5Ah2MIxzOsW7QeW+TZ6ftnwr8fSpJBGBmu7afoIpnrct6/+w/k
Lu1LWKr7ZUH9wOaZAkTBKpTeUYcZkrVGMZBf4va6MQpijCbnOqsVR/CyxQKSFuC1CtnjcHj01VeO
BWSPmiFTeasdR2Y7Z1fPZIdbrbmTYYGByJEpordXHIGOGkDubvFWDg/jnFoCtdE26tNDPK/zt9zy
PLpk/OclE2KDLumWTGg8nFmmsahfdOhqZZ/gd7Xu8IZeLefVUKBmkMq6tF7LYSAy8OnWzYK4fnw/
IpkZo0vcdFcq4ch44/rTMqSphQ1F+Lax+RmBP9lnAkiGGzhfy/JjRW3Ei0iDq7k14dhVFAUmMWnr
/fYnV7F8tBUZ87ArdI4sRXVPyOSrV62BRWCF13L1gXGal7DZgLlzIZUAApvRBwjjLPmXPDUCq6I/
odlUL2ZHuQmy5sK35IREsMrMd7bbzg+1dM6n5s3AZmZVj75FwsiwK6oEIqnMYknpyDRAGZmT17VG
xB+idC9fwu6w0Pb8tL4ahWUKmy+2y99x1a3BvL6YXJ+LUkqlPjsWz8pCCXYgg42bh6+bIqD1nz6Z
FKn5MbXJdQ05sEPuwSFJ5SCLfqIlMRQc3VM0rCjZC4UqrJfmrhk26CnlZdIbmfodKZpS3MXeAWUt
TO8JbTLT1linEbpCJmTURbNHbpuUuU00MG2DrX79jO3hCgYxALyf7L+DQdCr56oBMKMv6ArS5x2B
9JbGVO8glktRW81JzeXIAHrCJevg50hnM+v5KUQqtUr3n/279GABsU6H/qwje8WwjbDVv/58N7xu
zv040aXwokv10/kY6XDRCpjqOX9PKBuGBqcU9HnO0MlT2BCmOC8aJHuZNjFZaDUlK3lHfdx31QG8
ItYicNoXpywglApo1K1FdwlRVKo9nf0safCVQxPLOk8k11d4gt4EC4vuvgFdU8o4jad2gjRWiCiW
mzhmsuy8BgbU67fvyviacBw0NDRI4vaZxRL2D+KCTAa6vjKTk8/mNGljlmqbzl/ZPHJ0zx+FqZlH
7+YqBhUu67l8Mesy9yseiOtC+abuBzPoblAbsW0xE229q2fnMnbEeusKSKscKS89vr48J0w5paYl
gxkCSHKMQ2kLgRiWj6aDT8AuaT0PtcOjRmxg9rFBvjU3rwTB3HZLLg094c/agrBIQgS8DzjdMaeJ
PT6TrYHMIGiXNj9pOc4MFGHWdOhFMpn4Qfk77XxpVaY69sZ7MUy5cP6HQ7uNoNu3VKaH9iOZp6No
8SKCyLf5rH9QYHOTDTKT0qpAlSx+p1hemTdDGultEeYR9+GVgbztPESqx7SuPhy5OlyUrbW4ypXe
B7WAGRDalUhDKN49oPiZ4jErtjs9MidDxeDiSaMBGRUbJ5ryqqysYFnRFaWekggQ3yA64ZfH7i+n
JWV6gl623cf/q0EtT8kBspEWiIPme2dAgHg554HMuWvJk8L3X79hzmfbRheOo8griKONZi2/OQCK
f4ukKBP91qhFbAow+Frsd91gOP5xbOqMhDlgIzywIRIzzUCFrcw3kiOTJH6uaFkixQPdbRcSXVBP
eKyxI2RdTBpH4jugjqXy++wxpvAR+AumXKkCfYVs8zLFQ698E2iHv4mOIMECd9KDNdbxZsNcHZUo
CceQASFn+Mli0iSNXqakTB2g/lajOawi07k6dWXzjCThTyzDc9/+lwUAk6CuE4f9PJMMpZ6JGd5U
lXZ7F2Fda53dUiqiB1loUQoj4cUqXiFJ1ogXp3KGGxgzfR+BD/PyIO63PKBg+F9t98t6M8F/tQcW
1Kw6tcfEOo0D5To1FxSUblrZDujTKw0ErM6XRej+5alOdidPwAUtxBAQkoCphRQa1d01Vo8AiDbI
0yCPLsvB6tlY33sOAQeT8Jk7F0qwXbEwyiK2x1m6L1aQxjhvJm6uApvWIQlZnTrsYX2EQSa9W/W8
5H7Hh1pGPcHHkC6mk5frCHkGXR1zHR/9aOF2c41jxbcBh8P5QgM/OhB+8PyUkF2v+MHFmmE9OifO
5MsHU02dAc1X/c7iLiQcxBojv3Y9rZokIen+IzXG02m1IkR/lr56joj3wgO3mY09KUswSvNL2iu3
YtihdZZ+gsNIhC7PWvCCe4ybywtkY9FWr9ZQoUNN6Pv7FiKmyRiL1dNFc8TS5G7iTvwOY+LRMToS
xr4MEyGgObXvIhspTx5q1MHhOdJ6UkupfqSZGsEm0ZsURNT3I/iNr019wUOebTJXWrg+YFtm0RwT
h3IWbTXnq9b47jaLYMNQAHCPQ2zV87eOvDOIhm7/Te/Af6ZuomR64+1kpNvlDGzpTDyE/Zn90NPI
B7hONNmoujj/joehPjNR2ErlXdYkB7PpRL5RPeNNqeM3K1t/Xz/4n67GcptmY5t8DBfidIM70fT/
JacRvbyW+2jr4m6Nyjwt/m3Rl3WmjeQXgDjTdg2rtXf2XCvLq1xb79zFm83HREGtpbQu1AzuOEjN
jqsl3yMFQzY1Rk5B1SGszhklO79FHtmZzCxaScNQFrLt/LEiY0/5kmXsHVw0FShls2/vZ//MTBcl
NmfPoa6u95kWQ77nvKUEU0kAehZRKLepo1g8k2yQeiFy1x3YedIms7b8Vpxr1bF0MGPbPWQduPz8
u4JWZoaeZwY5j1jQQkCSJoc3OPWHmjfBrRe8v1NOWE9JKflzMcXUFh6SGpwJ+nol5dasQbzfv16t
tfLuoiXkRvYqoMeksJU9lhhJoCJIH/8s9fpGEhKXJAiFj7iUhrEjQhx3K8M/FgTg5Z206j0AKUY0
rTstKtMKqdMml8T1GmZ0lXfuRN6J8k+NIR6beuLVAunIT+tG9cFFr3PFyKBJt6WnQvyf4dWO2Oym
qJXalHj3xGrZgXTHXxlNLQpV9RWrbTULdVkmjezpkTzmAXtHaX3g0vkwzj0DWWvpAO3dbCYwe60X
1otL5zCwDDIubGNU8pdKpnKUC9t1Ma7r6JFqR5iiofvHMjd5pZK+cH9kja6W9b88TRym3uYKr5UU
/d6hQkDIm9HUM2ClBvxkbmts22Z2/nfHBNuF2WBRoryiVXYzTXKL10GgTOEeiroIRTGg9XRCHx4X
8yIiwuUK7fAsZTCY6i3pXIvaFvocMALMapxX8SyL6FpUl2CCY6suws8Vkec9+Ke72w1o8CAFXtrr
LomL75l1Hfu4l08ogWmBaHuqcNEAI6aSj4cWpjACfJ13Xe0yL2oCqaDjkWHcfrnAYOaGAc6DysjX
rhYAtGAYN0mBqaZov6P2d6h6DKlQsqqJ5dcQZop5hnGtszNAfUp544H/3cUlnmwWkBzR6YjWRM4T
afirko1o9I9O/Q3vUTeo32udQHBeylHlwp+CYMBGoKHDRb8kFGUVA4svIOpoVHsVoWToBQfRFzgz
gdCjoyw6nwYObctYywm3Fkk/bgihtmruDibcMowjIXnFB4xx4w7mPIMZAtr/bgLiIkIR0i7URpKO
0tjcqjzHw+HRV+AjBuRadGUfnTeGzFqMnxqwumARqnt4YkaNiIUMA26+AX7/S///csZLT+kXtC80
daYtPjmuPOzBHGn/8I6kA0wUFCG6KW7MYMgHA1otuKhHT3MEeFyMoxUuC2j8ct8VwNfWzotS/knc
E8AjyaozNu5LDsZX7A+PPA8UCMaDXfosBWIa2lBRnCHE6a/oFiMalemLqcOOK948M68uAzTL7xO1
WRPaC8xP++42THkwb0DVc73LMhZf8vdjR4ibvz2cZXIkAMm/3CevbpwkZV7xq427A0N1eyLSNZaa
NTbIcrWAeAya4+Ud1tjDI90BUYtXTPrOCSYvuytLpYBCe1fdPxAT37xgTvojLUjuclqVO/QgKHw0
F/ywWF85qV9HJZP2pXBFG6iwuWoQsoVExHva2GU5mXCRFhLK6uU2W/HvaGHnT6vraflN3zmBfIY7
WfN9wPVePQK6jv4WhwxIge1cUCBgyXuXYf3kKORC3Ks5RObaT3tYCFc8oMgIJHDHItBBgVptTN8n
5JZt5AFv+xMVxKIk0KukKEo8Y5/jgaJxXivCXa7LOy0Nwh7AJCvVAOCchBvlW054+a8ZA4QaakWw
LzJ9dv4qrBUbaI5XAwjoo26oHn7apdMgjo8lpIyr5HyPTdNBrkrfgLex5FjNKaWVmlwNSQ/3DLVN
/huZI0QANQ3eZP4MTcxcXrl0a7g4iCsGvtQ69yE420qziumTQbVyJZoGOp0Y0c0jog/7x0szghFY
fg3ddbfnrT6WGrIDfHnuBuEtQIcwS9s6MMi5NPmTHolAPrPVz2e2nxjhi9/VEkqYfd7VVn+ln8Ha
wMhm+Q8GSPVW1YSnjZy3JIY1eV+akKMFtiWhCmtLCpQMYHS/owlvvYl4Jqq6a76RS7Aj9wXQ2Sx/
tYNz23YoAFyCMf5tDX/m3kGY32VhgQMbxHeIlToaavO+X27QfNYOaBzAzmZG+hNO+lyMmoAkvP4V
QAQPK8fM+rDJOK/Qr0+pnxWiNBh3kUei0kHRQ4m1aPlZDKWP/qtqNLHm2Q0rSGzwL4YVfaclWwkO
e8wK3PX7pkuCq+im6V6UdhMkYV96T1aw/XQVpe7rG9Men/m9g7E711LTBWKi+VPyeBqTHGr/IgUk
Zx8hL+0nCegpcU2FKvm6Ny5Mpli8StaNCKYRHc1EcpJ74CSgPiNARX8naZhbC770hdBrXW1+9jgq
P62a9Vr5jI8WShNB8mgKNeUNXkqcdenfvlRa7G9+g0AXfIMGvPZGClLljRFt/ywZEXSnTuK9StwT
QfG4Tsf4nsOxeO8IfTAZZpQFB/+Xgg5ebz8QH56E6X+5F842g8oB3KqGyXTJ/994eGew3ysVtS8A
7miqe5U1l43Wh4X2UU1pbK+2FtU+la7HaEk+8SJaPFES3T+rZ7lYXPaky16hv9JwodqOEXiVx6gc
Fv3Vfp4NdPFBvAFqyQGoSayEnMHvJ4042QyJvNGkneAqY9RTe/VMKxpjPULhcJinM+OPF/rGol1J
INHtH1561WqSyeiv6V59UUWKF32fj/mWVQF7qNQ0aDrevje1nUMBwuzTZYLG1A3SmN9/s7abkTvt
kFU8v8V6DFmQKwBN48sYFnuadMgvE+GVZQrHNpp2Ml5DhLXd4ClNQ1BhHaLBs925IWj41lUQ1rhk
Pg0ZZm2GM0T15SHsbcukVdbdcW8mZjqsNNV3czIy7C2wN9GY5YOu8ZrU0SUMclH3fIqdBt/0FnEr
tHcE+I8UjDMI12dcrxTI+i/yQRUhOnOUGmZLc7ZIG0j3DQF0JHfTn9LEBNtwu8a+L6KhLT+/e025
sLcc6tbTRnCV6zz4+Y1PL4hVvaDH4sWJBdof94KCd6BLCHS0Oqpb9bsM80iJpKf6Th1tT/oSv5kY
HUmQRE3IMz4mHcGqjxhT0ttFNz1IZd6iATWXMR2uvhwMGZJ96hE2JWwKY/umYrGVqX+eE7i2EG0U
bn9KuTsud7PCk5v9PGDpPN9BhOmtQLozKjK5h+M5flZmYEABSqsG4xyCWJXls3uhUdve8EAtnIpa
jsKtZgpdtgyftYMeR1ic3+nkomJYC0SoT/5nhWQkjvW/8vFMuF815SNn3/QQITq3cg17TMlbJ4j+
o/sFfwXY+TUaqEwoSr1zfDe8A6u+BtUHPCOJVwk/YiKGfpBiE3FtfDoOuhq1rDlFb+gIT7NNA/g+
LBmbfpPi5sLrj9KwyfKJzUTuJpPXZJ+jZMkzAE93i8/HYlbNy7rmtRFc44WCVMjnY1qzwdz0vI9W
9O30yzdttKq5Mogf0cMMhrh7MBSVX+3xoqHIkZVR9g9qGeMYVHIjkyRWlAITpUiXRDbJ21yDeYWR
lkbD8n8+Y2foYHHoQuuO0M9VYa2cywaZ5iT5s58Xb9SKaROiXfq1Fnjg1lreOe3hrRhzqpKyF9YL
XE4HJtxsPq5xxu5IQjl4Ca0dVIMn73boKHpwnggYh0h4BINuYKc3qDRqLhSGGY3ss3Fgm71HoLxk
t9ewe3V8NORlHLK+NX30mYzrDoo+Z71SpeA4ce/4PjdPe3ghDeMW1FVfd+rnZhNGBFHNH+j+Q3VE
dXXGsoVAJ5LU/MsCGu215yc2/ZkTToVt0BEgiAty3xDzUHM/yaiR4IxgMPamt3ZJ6n/4JYOV7sbc
EB0xNNdvr0q/aZK90suc9VyDB9mYMQRwynUhUQ8FV6OmbBhY2GX65eXAcGMmte6MMZACh1yJFidb
+WQDuhASREQQNveKiBgvBUVNXdqN4wHN+ghVBoz1Okl+vscssTwUuld0nG5iJjLUnz1fSRnYSdSr
AbC5zJWelGSapJGsE9GaSMXFNiC0AeEGtnZ+ZsRUi3VV1c1udr2Xcr1Xhv2310UWqpYYFuPIAFeJ
AWihyOLWusiyEYG3Ts+WKzi+Qs8COYrVvqOrJBhe07WDJ11Po+DE/iM7c05QIS5qNndwuuhETQrL
Kla332ZKLoXo5dKc828CDBwEnCBuiPE5jJE85Lf1b4HAn0YKhvsY1rPvmLPxZNq6UOGQhJvm7IT3
yPYtqOGLFZA7vbt2Tn0M4o0N5U4xQZ6v9Nick7fpGWp2fvO+r0dkTxG+7cOWtXwCrAwnXsKBicZ/
tX0BFdIJGzgga8h3VrfvAyUmjGQvraEVvhyaVmDXTo61OW7gMZEGWmM4wcbgmC6oMiVIwSVyHVS8
waZIjIldwnXzxWUTUaJgm6Zbbs5UCdKYGHz9r+HWmN2HNG+3m6pnvn+pXbkhmWWidbvDnr9zApOl
1PfLqfFXZEhq41n1+1gxgfaStuQWX5HXmjzFUwLNzPruz9peUp+jp6XurtvxHr4Uj3hzP4awsuwj
mynRTmJOzXG6ix/3pbv8ZxOQ4Tcjf68+hFJmNyiZkOp+1p75Uo/SknNPZO1RsFovnvyXqD1uQsEr
JeoU0MO6W2kina9kW9iLx8vJpyNJZIlbgeGG/RtuPiKjKDKHo6pHUSaQDFs6So4X+Hbv0jgV+k3R
jrbalGbnGre/MFxGGYI3mM1fSWjKOAvwV3T+SXtAoE4girM2Kjkns7deQxrqdOYAzstupMUz/ikN
rb1aHn0Qkr2fkvkilP0oAfImHH62fSgaaUHJ3lUGvwp9A1SBtNferUCR5hMWZFQPv6ftSTADNz1N
/5EYs9SBOZHRTB+/3TkPEsZfAZho1EoBF29qQ5DvKvPUrSBtSacIi+bXrFhvDan23aC1QbHVgifj
0tNcS+teHT5rq4L87dAC57YpFp01cs5HaJeBXuUjyFWaJY8q/YCx1BfKSX8GGIwlHUNJ5jEyWCMj
JpurCnZoyFRu5Cl3hLzQYeaYIQRgfsekfUxq2V91B7vCJDWJhf+ngcq1fe+4aoN4NYQFlJRMn8G1
C7TE+StIf+X+CWD89lVWy+DxoaoPedo4G6EyhwOWmVw5JR26QWmW5m5IT5Fj2Thvjwwp/V4yHCw9
Xn8WYQO6SiPaI9ILP7cxUhSfClCCe38xjNmqvp9mxe4VjUqjGixl0KtriZlJihfja19Sf6oBiCSI
VC/Az93rMvHmFZ88M3OFusWaqVdG4EFmO0O3nw0kl4jXhz+AGzfStWu7GYPnOuF+z9kuaGpgthB6
48Qe3sMuxPLxnEC7yKQx8OJGdmlweqiZSotsH2TGbJbN5ZcXIujNNI80OESXPBD87z6k3NyaOx8W
me4bsuvWcQGgsGrNR9Rc1Wt7g74aV6W5srR3vz4Rnhs2yPr2D8SD0p1VB+CZe5RCXx/WkYmweMGs
bid5JTC4UL0ThpgeQDoQyutuCCdlwOoTA0pGmO2KNjXwv7EPRxHHzc9+NnqaHSqDK2kiEIgbLwX0
YV3EgY80/8BQ8uPzN1MHjOp2x5fLaraOxuYba5tlHzkDwTen4ivDR+XlaA7ey0XAQUsrxquf/B8c
B54H84bN3wyk+9UvZ3zMy3EnFzZXfhN3dqiKbCvMTADyOvrLRGA393DsiboZcoMbIqac0USbcfaJ
XU6fNKp0UzIV68PlPMYPWfOMtC/RXapmSbHdTwDuREa57m31tNExhbz/PGGvoN6cE5ZGVogjifnc
PQOM0HR7fcQU6cQgZtA4UPxvQN2vmuF+Ij/xx9VOqY61MDizfzeg9q2PQJaWXweOm8WndLA5IQ7r
tETcx2tk8ldZ0MWNnIuSPlT/xaj8E6oxnUdrIx2i9L7j1GzgDp1/8uIvY8UIw26imFRY9jPEfG1K
BNCcifKWLVmy14RXVMA0ycWruqKiSRZOIwNFxTyl4RevygxNLYKQEVK25PKVcwU5YoSwAvkA9eu5
9Pio401Bfu8nXMorxX20NY6JHVtu5mPJKDgUvdpoQm66w8vY74fzFYrD8CGxeERU2aDvW9wxa68t
fV1OVBXuyclnPlQZ3kZzCBBy8lemcydHRmFNhmPCtQn2qRzTRg+RZ5jEDXHr7egOSJpitt3K5LBd
I1rEyOXWtk+JjaDCx3MsQ2VvBdKz7y+J7p2a+712WxbCxQm3IfbRUdlybLXKJy3t51uSO62Rqe0l
jdtnEcN2hFjY3eMOKrN5ocpEN7crk1O3Nh84EoS93saIuqfDhyqXgq/hCqV/lr0Scp7Tr56hyJx0
aueXSfcpm9X/Ta392DcSd3P1aD9jP4LSrWGvsdP4ioijwIOarjfgmv3cbHRjKgeoUaBJiqUqurYp
rcW5vALDLVRYnqW0HqCSGjoJMRHz1MOuf6B0uw9QygVwqI9pvCDqhZUEuKusjvxKC+D6is7vNbbl
9LxlJlu8Oxen3s8funzrT86WNJeSDF9pIIzik+h1YSkAY2iDVsz+TD4xCWIeA4YL9aT1+pm7k7QH
6TbPBtBNQLOQLfOFBQ+D5bPs3+Fvmg24BYSNSZA1JPvsauxiLwOq4jPiceQxMQrSKU9TQqIXr+0Q
Amq/Kyu910J4tznAnW2Bv+cDRpnxJFf4LxaY6190H/PJg8JKUKS5bAeWUy0GSmjeYfU5QTlq3dcx
FyMbIWcHIWsTYiWjnvXVq9L8AjzRlnIB8sVlMViLDkBKYDuUvmbqAQkfx++2Zq5Z3Kkp9BlUed6H
wGOJzCT4iBI4llsTQPKuWJ/sYZ1+UKljf4tC+/puErEy77cpoIr1h3A3BrggyISoI3ed3OU0pdBN
rFgvjJ8cC+Gf88OcqTlL9Ffr9XSSmW+WDNXcYByyPTtq4zb4A2irsFr+/HRhV2xuwqPBef5X4RHs
gjqN3j1DP4pL/eH4ECsxZu+iusvXFiXrcZe5PRK38vZKLKOpvzA97csqb4sjTgi8V01jOSpA1x0x
eXZU3FlUc8XjZN8AWR9CzdPvtj4cky1EWoaXidWIOB929NuBHfegD+ZM2kZbRrgWtT7NKtI8dZ9A
HiCwd7ewJ1Y4QceOVxDtzE/rv8pdwVnEcTIWde4Pnp1kGIfdSEpYqD7Bpa04zSVky1v/KMMRtg7B
1gH51WqM2A3FUpda1K+FnwmKHak/VP+cRAOko2vTLPsPnzdK+39ijYCxc8FTZGRF04XqhpryCgXP
SrM2idd6UIzKqOrJ5cNyNXlqSqqzGMb4pvFe39dCl2gUL/JZtdVFxU0zBZgfTveHTFivDgleUqms
J1C8W5PR99aV9IpgWFVbK5IfBxbg8i6zNQooAU//iSTLRo/r1X/9Mv0rKTcHUvcdkjLGHDp5aMhV
U9L9G7eyMxHUS/3szH6pFT0cuogTpUWXeVIO1ttFCqhEzQwETtyjsgbsDCKGLH+aYDpz6gNCUYNw
YdIII36im0qkVpx5tu3GYMEvkSd2Ar4pJj6h5sqDO2amYqdzSSOg03nsssf9W2O/lK/I/79CxskS
rwG3IkLCDIZaBc8/Lus34FZnADeKPyLN8k3jQaZ/8Rs6WMh34POXWtlhI3/bfggc67DKjW10HUkW
3/ZJSseJdPU/PSmW91YhDRw44fwJjPw/dR2ncCj6zFVU+NrOg426/LQZYRBikAnMmDjfECQ1PhUa
hg7aqXQhwLuVa3zDJ/wXKDTwBPsFSmnJfvUaBpVIgaI4uh9DnjJ/j9oq4aguNPOC1WvL9WSi66Fk
N8LFHYS++VTo4dsfpXRcJs9R12uIhNHpM+QzaWEAb+1Q3RYAqZ/9M6ofsSPTq+ZVHOeThxZOpUfa
zRxYTAA6NIz859ER+hpYz3ueCkGyfMKDEmgGh+d5tGRWHrkql6nxb8HF5XyZCKP32SnIzQ876809
0QZB7rDGk59EweZnZgj8aTeADPnRkvXXiQYeZ5g7OV7CH0mNRocYoU6t4Djmjm19SQDLZ6J4pu4u
UAOdvWGlt9whiQOSar6+j2rEscd+4zNXRYoiHaQQKcO1q0afdfaX5nQNBgfkbh/dJs+FAaS8buOh
2NPBz54xPToe7F/F2iSCqbxexch8BmpEGVv9oHoOYysjFc/ZvDouwytMfQHiphcmJWHvY9GAPK4y
vD7+icPuuw29/wKxSwLlGajHBRpkUQJKZRXWTxmoqtJPrUAG/l+pqeq2bXxtWNKBhHgIG6T/DMXE
v5rwcPyPdTV5CjFZ5/516l33rGWVlYnV4SY5tk0PGKDtcceqbIrwWzvDW1sRJHKQFSulB78N/brf
gdv6ugBEiWCd0RCNNSY7V8VhqsDYryM507u8JZZd6rEUA82I/WWJHzMOJp3S+0W8O6cAq2llfjtS
utpmYpAD8MIVBt81oF/gT3s0vYwuaEI4CPVFZm3DYODh1RUU8U+kk11WEPs0NUUEWDTlFXKd0iiT
lAy1cScFGopW13Wsyy1V/W6Bx7/QaZbGV8IddCmBaRat/uI7KsR3Q/I5QQxYlrA3Z0mdbJF7ejos
7kTUPJqp1NL1PT42dKXEO0NOKuOG/5DO4Gh5BpWTW1WUJtpeV8ZMQEI3DqjxHKRbIWR6CVT7OuJF
M/W+Q6vqkf9GHC9zLZRdIl65y/lJWy7bT3MdBw6J13/V3tbawSCl/8afATc2/NQ94BjhdtcMaoD1
r9e+YPJ6Hsf2bhjrn4ucv7bQv7Txnenki7duUjbSJruc54PDa4Nh1JXPbGe5mK6DHYHtU+3Uvx2J
umu331vgbEoPEIPeRLBpEHPB8a7Zy7r6YtC+3jTE/+BGvXAQWzdobWFD5Yrt4c4uh58OuDSLT2A6
mLMNMN4nTfXE4M7p1pTNyEkJBqzWVld9fZCMWLZoxDsvMZuWXYWp63jA930QM7RJ5J6Pd3JoZYWb
NHadi7rF514RJdIhYtGbflD929ii0a+/+5PuboQYAmnT8ecij7A7i6l40Cgq++OF/3F37BHIyryR
mXB4Cl0zEX3W8jR1Ue/9AZ/41wo1kqERChcu4u1FbE4ndqurpMV8A4jzBv0LhpLpPy/lswW7ObqJ
UgWierRIrpy06/N1CaH2EFH+GY2z0x2y+cxkDQ6WqwJRFirTa1E0e2Au/lkGbaQB5OuEicovZOSi
ZL6KXog9UTrjkC6H429Bx5jB7Rea7ZfGzuVKily67KYG1LLHg7uMLnEGpGK5vvh767dL2fqXdbcv
9RhZK8173cJdAmWCragNf5E320gBTsVBAqLXLFjR4xS7wfd1ndWGjqf3NZlFHZvzRQMfrYCnvGOt
u9ZeupfNuJhCu7nw4ksabMh5rgEHHhwhPCp5sZggW3UBY+k46zrNaEdKHZDdycP31b7Uscq8Zk3P
UPsAwEG2/QjuQLeF/2RtBXNOg26fzg170gLB1I+bLtDP0HU58236vMacQODTF5HmQN8OEUnZrUCA
X0OpxV5wpOXWco+XwSm91GXnG3JYPjGNulphdMrVulYiXcqOUm6YXGVvCH/QN9JGwYvozdFtP5st
5C2MFcxcwd6zk/IICq7dKJBPokFg3fjTkj3ZLz3RU6TQhdOM3DKt5R64B00J8E48XZzz8LDNw2Mw
DDvznMz92rBtuTFtJOcTfyv9knQFvjNgC/tSYHGod3dHisVbJ+wLSpRBDTN0M8IpbI57MBgPc4HJ
YIty8lTsXVbBI1taxMj7HTSBqk19+a19+p7j2ro0bbuDzxQ/0JPaj4bQorDEOl2rLJlFCfO+KIhB
uQO8TFom8UM/1NQu4JML8qagsB3OUJOrC+a3YsviCVRt5PA4cn7dPuIhm5g4EsJi6hbdDoBddwoR
qgUx03pyo8zMvE5RqmFfXRE5zMV+P8ruRKgy+9AeUDFrhUbdnpk1tMOG0VppEiby2SFu7FpbEwRi
XnI75v9Ap154MQP2DjCJcDC6GnvoyXUCN2nmia/VnyV08huwwOvfL454UG+kh/WS9FzBNVUjsoSY
e0e2jCRN/0GqEXPDOT5CX3gd2M605R4WfCeZWPhUNY7/MS0Mp8JzzEZ1eiYOPL2LqeTkDm4HH50v
Nr3B9NQAKrvc7PZgc0gdAFNq9kGr7MoewH9rSRvh0j5oeyvC/hXYo0r+42uCUTMXkcNeK4isjZIl
LtAt8fCzNXolzdtWnY67Yp01QIHbvqGzrh4BgdY8UWYTxyOwiwo0ye8TgpLkp33t51TiF2FNCtKx
vePOqf2uvdmXjqnsk87Z6GrLoGTNndfD4olbs6t2P83OK94JDK/tr+7GaSulWuczIcAdRparll4R
rfjBB0DIx4Mvp1ujcHhjbOZIQk6bARhCaumKV1n2UGABGJTPYNCsQiB6rIfnq/xO/f03bpSM0Pv0
9PMsIJppiZ4WrxAcWcsLc89IDDGPh5fUGrlUKRsm3YbTfiQSSMYd5Qd192GXDnRonq1ahxn+6fX7
Pr+46IHxePsnL2ddOkP6p34iKQqf93qOWxaJKolsTYlJFcuB8Lyn29grJJyH2uQX+/REvDepq4Y9
Bf1hw3pqVmNYCcOkQ2BTXOKefI84sMT6Ze3JRrr5bY4dTTeJM2ZnzpOo7NWkxU6cB/HF7JiL666o
unUVf5Jt1kbK4atbgb+5zr/Ru9hE0x6PYJPRRzUDVR0JNsyhj26A114AcxalLNT1WY+InQxSDgT/
Lj1tZQfKLCFjlsNGEWwAmSLG8gEvkpPTcQ1kYqgAEA7adNatnzhmJ6Zq0geqaplIbCBnjRQ5NNsI
4bEI6cyKv/3exT59ZpE5VOKuEt27kLnINEs5OBkA6sJ2lFW2Bjg9F2rSDo89UJq00RtCk459L5Ma
V4rT8PUrF9SNWnIFPJdfMFYy5EdWJKUUdrvOLsc5m8M7x5SO4ruqxs5vfO3E3tzlsqpU2tXyGXnD
O6goJwGzmvioKt4+yn2a0HktxjV7YH4SwAZuxlR08MlsNHNDY1JQQdKZR0yMn6czq21m5f/eUKhI
6tTkUVHnAWxwqOqp458ZV4W3v4ogE1PYazz1BoJgsX+i3i9uMYFPwM7xgo/geCSpiifbol5hl9Yz
EeJa+lNWcl3kuf9wZ1TNZaBMttIIJILpBdsok0Xtv4RGcWdUdH3TSpkN2AtfVtzQPiQEfe1Kzs6D
/+S3alKcHVlKi/HMgo1hAKjQ4FFoq7wmx9TpfCHP/YaH599O1SsH7G4O3UBubNDFU0orPatDaVPx
7yraDRbltwhG71wSGvwWMSpWWotdwPftI3xCtgv/b64Icu4BvXnPEfgrp8b5laCj9zHk2Wf8ad5y
Ntkm5Y/Sms0yJzHpVOIcaXN6+g2jTeAQNVkVKuxLRQh3wAHpa4P0nnwsWXuNkkl/AX31/r2yfVO2
E2Y++7ZgzBQOt2Um4bJR+nhMV/L4xnY5Yofd95OsmpTKXtI4RJDbFo1Xfnfldiziboo1ujkeFg1Y
vqf7pbCEbuS9ZqD/Bc7oboQdlwuC+W7sseC1qksmFB6ACUvrYBuNEo4uGNCAKUixpCACreW33KOx
8/YcAPpalQvhJ4LiXLWcKlaQoZXm/bumUGd1dsQ45cL8QV2GwBOB/gxxK7uhndvOVOZpP1yxHIIQ
+uyRy7voBO02kyAUzyDWHLpY0bT8I4i4EtoimxNf/v29nmiBOnqTkw28LXc/8HC6upexYSMfWv1D
KzBa2RbtWYX0rig9z+9PotXnXu5yOh4kr2+5cqVX150Tml9jSDIt2YG6qQv8lQ77/lV409mBqqK0
TKtLFldRcBdfg9YqDITUkyED74ytzqc8W1YcaqB8/Da7PQJfEQyZH5eClrYMWBK5T7/yRaZFR4tY
pJ6dM/PnIBLCCMdcJOPBu/BVNvxFIu2yntnTwgAnaP42i/9uL+ZZDgUHv7vMB+IkH9Bj0sdFsrlC
1BvYa8eOtxuqnuCvQrFnV87AcOjqeVncjYFvPkCgKTbICRc/c7VqEYCY5E6g74/9MiCCp7W7AGk+
0U75BqAHADd4OuNojaVwnVGmoSFNQ39QvIL994bPzHedTtmFI1UzDTOV8tvm1g3pZL0spcJSTWGM
M5Fn2MsmYWpP4jRdb2a8MsNPOSKIc94JfuiNaHo+/eCxnyqC34zeLVUsgQ7dhLiBoNlCKfwsSGk2
FNRxtlVur44Yqub1/QYBhIf+6oLLAnSAlRXMXQ0Is1DHrtxiFTb0UJrE8PWT9dwbiqzQArnhzgM8
g/ENpd8mFux0mHfkb+x/az8V8oyGqbYtJOoLf0esEyAoCsuillQSUHKOp9xuDWDR7UoFtwNv2rWa
hnEJKmkFrVnkMbwcW4oeufNWugSnfFtK/AjeKYb8EqSx6pJc15KRVpp1ocu9lbK+IboJax9f5Yyf
E69l3o9JqR+TyWHfG09hZ5YufWpLZaF6B8WSxl8IGNJfMX6W/Qm3/PhVLCdoAN5NryaBj8g1x0/W
zcMY/dbdRUVaXbZaJljQP5qOVA6X99GjgOaxg94YAIpq9XKj0ak+yUUNzkpVaaV9pIPwa2mZ7236
i9Xn44Hzu+h4Q9MMexIDXHyUoIYKYlC4NUyu11RQKMWpUVIozuAftm/bpIhKrHfJ6tsy8PBYbvDj
PgbRjmnxlIPN0AdWgw/utS0lsTp69PMTEU2UW23tXF09v/fPj1tqA8eEzeAm0KaAkUO+qJJuxau5
yjrNq4c8vhI/KCqsRgLCtUsKPMyHeKGigQfUP5/MYMLUOJx8S2HslYSm1eoWW5Nczjl5ZghRod6z
EMQPPnOIJ/A1LDM3qNkr8+VzLdS3Oxoh2cUfb4oKQBSaAmORqOpeZtH5SGl8eTZ4EIB1vSBhVsih
pBhqf5QfmZfCfHB3gVjuHKO1+BlU20AR995+4ErrzuueKaP8D/eXHZXdsHJ4DE/g30W8l14Q9Drv
iwqLvxUq56MP94CKpk6IwZ5W2A39TuMyDI4kXlYl3QkEfhUd1wKFKL3XbWa3Bwpc7uabb9rIj71f
IROkD/gY2p8keSlSGMAtNll4rNWLkijFrG088qIlXzSLus+DLtDGfdoENQI1oBL8Ga11HF852Gei
APNqppENfX6Z0PZak/1VdJb7PPlKJrbsBlza1QVKVeKChmjUkTG3i6zdvL6GRXe31Dn0UlbpXq2p
SSxV6O4OWjSWC+GUi9ZkqSENSRDAivIoZ+aAm//+0IprOwnHD8/26kbyNgNEN9qSSOl0OJmRkiHn
ajJ5Zc//hQTLt9nPRIdXIvmRrvhuSxShYoyVe49hAJF5B3HXvxedeGDKrPP/ME/UTm0EFOpE9FcM
dhX03gON9HcJZ7KEeP1FEIbVV44Zhscgte11bloL7Ic/XRpQsFVplywNSQwOVn47b3OClEMmjSHF
puyZFcIaRK/O3xwWf/GjZDMqIS27s5UDvYxlI9dgwT+F6MMGX48SF8/QVfgUJmKONbm/Td8YrNgf
reAYg8MrdswwPUb+hnNUUqsnZ1GMFZaFcBkPD0qQRWFm8pQbmWXYlVvHO2OF91/RHSLQvEXdlaSv
qOakgxC0UYnnyKwVzEkqJtTVj0XZaeIQGOx60PSn6QxnSUR2Z/0zyN235VI0wIeNAWsZ1dMwM5D2
MlOVma0ruarQ0+fzF5eRH/knPElhTo01PTxGZKHJc0u0BUjphNf7csFVje6gk8eLmF78HwPj4OkT
V4lBodC1DOPJ46dQFhqBuMUNfN3LA4C+Qks8m6JLd7NklKSWeBw60eLF7LI+5gVB95aYark8C88j
XelGZKF4z2REePlhuP1yAOaCLwoJq6wVS2bqDD79Kg5DNsEggaTIm5C48019ewzhjQoCGu9RNU5M
/Z1sBsj5BHUe9Wj3FYI5KtfD31OH59wqKBRdT2Groo7srRjuSJ1/3a3OwOf3LIINJ8KCxgGQzZjB
owcIBDf2AnxLB3fYRkfKQletn9xCNpPbWSMtnSYFKkpidjOgi6KTXpNTGujvom6qUA52clApZWO0
GI646na/1WX2+KkLtPEJ9vuFzgBxOt5O64FwMpxmRJYa/WHScueh2WlQpcBj2l8c2vLhzXVzl7RO
grNfSFMexwyMtnaWJ/i/VBXCsARPNyRFY+Vmn0e36teGTPfpp2HfR1uC2H5csufPE+yhTuf0WVVy
nbyNn4cF+scTBx2CyaKtl4/5vbRjl6BcpyVms61Oe0T5T/SefSauYfruj6l43ZuXC08DXHhs1i8I
Ln+oWeS+VWhFTtztHNC3sxBjm2f20Ysl/LGR5KZ2J+ffMiO3serYedaCe5zmd6djBmUOx0fTduz4
p2K+5gPvqBjY53q5o8sjAouVOChNuo0eUI/q/SJFE9m12iKYKzqSfkIZ9GaMmdW7YBo70j2Q+ep9
w8miilynbUfY+yFN5WvxkWnsuHBJseUdkr0AunAztKFGy8KB4ewaq15W5ZSoXDtdWW4EqmElSCeO
a1wtP4GAlOxDzSNNxJX063hiYi32qpf/ye36Y0Ig93nAue43rf0aArQcO11DNc+92BkkJhE/FTq7
YWYhEBd9l/7WaDhxNC0uZrjGk87zw9eoQU2hVXLzx61lVLt1ihGx9sk1ggkh9fYmtkSpyteSsjQ1
Hc4THPRJNh9xAB/MDKSmWK3IT0vVHHqxLnHpyFj+LodaeNkrKyzd7+fm0KuSOh8xGzCLoERm1VnZ
z1FxJhtJ0Qy5/Ybc0/bgk6au9SQtsrPWhh7eDJCro01JJY/DZqp6BmG6/FEJQfcFu0EftF7WXFRS
+tLSNXFJr4CYZC2dKFDIjcUyZ4gODs+NIET57Yxavz1+aP8+isg3LXzfAjL3UWCgmy4GupicrVMo
8eo+LTU1X5sKYhzK5nAagob/TVPBadMswAKUn2R6BxnQ3dQ95ghbvkrJ0p3WyuBjIXXvan6LzNBK
562t4ehLwP4qSlMnJtWtZyVcArP5cKOBlFkgBXB58vdjfvmMdjWNna3YcPPLPM0IkMYdv8b0sbgH
tta9o9cC+ZprOELX1OWtLy2UpI0w4HDazBfCPu8fCEnCEK3a91nH0QHO2bdPIq12fdiMn+lDXK8r
pMsIhnnVw7ZZ7aTTwouf07GiOk+dVeqn7UZMBX9BdF2N08Ub9JmzBshLOGNi9vrxSBvaW0GCejTk
CO3F5fcP/CoUAhkCMFEUyBHJUnDsvUrRa5BT6QIzM0GRxJcW8TNIMq8utZ2eco1F5TZGgf0rvpd4
IMvaWiBlo4E9V2hltjHXWXnAxVuqAD7sOTFkHoewioX61aiOq8lMwW/GYxqr9GPJiLLm+5q1yaG7
cWH56JtgU0z+7N5UUCp8JwK2hNKbY9NDtIi8OALbNrGd1+k+3LltiBWr1lp8X4vGCOiP21GFB6qA
dkk8ZcmxWhbC23Sz/fsuTrgbzEq4Cgrfvyg0gHbFCPtfQTTemAhfmGhog8CZG40nXWToh70lhZqi
fL1PczaMMmBewm3uzRQfdP0DX056zckFZ4t2OiWMliOleORHlMfSR19YTvZG1KpLZezHhJvrqnpv
ID9E6/g0WfpU0fhTbAbOveGu8Psbd8aFXd9UmScqHu2yA/yAiN4RHegAf5ddIfOQIgE7RfoWtqmv
pfHyiVaJ5K8OU9fSrgZIHlg0QEQpFq4F8Ob8lfjebuNMpevUHXGtmMdqLQTkK/fBP+WlHW0Nd3DH
3u5j4zcOemddOWi7DzbD/9lZL8tVUs8/X1SKESno7D9MEIXDIZ17rqWuU+8UGdLEtrFBvRC57PZi
UXqxYitlZOPt05IWhfIFtqetLCiTKuSHuZX1+MK39BchbqSZq469efAnSw2LdIKN5n9KcTGrhtb3
lejaUGOFFgwk5B+B/mB7+TwINN4lh8H0+k6xKQ5C39nOxw4AAT/obRMDHwYio5hhbdJt+fd1kV6s
Zgq8JIs0ODzZFnbDkVA3A6F/CKygi1csDUXMz9S4+uU4gWHXtvkus52yGKakFkYKbyyOnBDEKwgs
3EpoajzeFCpzimTjz3G82r0sK1S4ElfkUAw6PIb7rL2Fr3wKwNFiS7LQo8uHZo4NwCQd7s4ePfTv
4TFCqSDeYEnO9rlWT/P8MpYhhMIAloEThfMp5d8xNZf4BH4Rm3NTXxIGwa6IAbZ4c/XSKhNzIfwO
NwIfjGyJ6ieq+CFw4pujkJNQNn7uh4x7gOlm/AOy3VoslBusBKGc1FfByX7tByyhBGivnwejpWnv
8aq+kczmu/uqm9a9dygtA2v+VkMLi9Bz+qYfnGVJ39/fqkdXFYPznay3J4fou6x5eTGmSb3jzwbX
b6OFTXNAgmX46oJ+7SxZmyoHlAafqDZHSWNZMw8WEz5Nb95/rtIGnEqum75xP8NhaHXnb3m2Xkhl
KqLWBxh6AGbHebtXoX+E9QRk/0QUV0/2ZxLldxOoEz0OSDe5qkTNbgPxU3Dy+r/TGFVNpwxIZ7ef
vBqMvAGGbgmdo6Yl3AqXQDN1GSqQlUQddFmpJa3NHRy1WOR96Re6DBuaPzCoxOyw14VnNh4LwBaz
oTeDE8dJ8gTiTk1vMirBb49SXLbDs3CFWc4+wygIRTw5Ejdg89Y9vYSFq0kiSkXoS67OFPR2YvCf
pW0aHkZhScCk6KDa7Skfh6Sr9bquQZwInDouCkjAzodBNygAqkb73NYZTR3bp8qgfcNT5quKTR+t
uetpgVijeNJb3Y6EAkC530ieUo+tK7leLUPKmVDqaVEPg68sBcLDAQ7EiKq+1Ave5VnWz1gS9Yzj
EfGkjxk8ecbobP0sKTlMPppawoFGAR69b0GMl1a0V0KU0wTbSLbKd8L3Xv08mGh6WhLvhHm31WB2
Ni4kXjKKlZZnru03DpitDZ/20IeS3oEDBnKVeRJSRsnHE+66UNYi2oJf05SeUEMOrtrmslQ0OQyM
S3yqRI1znr3riKjsU4RucSNQ5Kf+29PLIykiTtFGmecUv8jLaX0cvL+plZylJWwJNjvUPrLNwrGn
YsYtvcsj+z+kv04DS+Gagzh2u7b3g06e60UcUlVDIWl5EqeAakwFiG7fhkEw5bVopRbvOamAB69L
/u70ghsRd1TNqt1FEqn/BhnITDNEhqf4QRh044iJo3EH0H5k7DpiFzQ2L1uZ7v9ScJ/LwvubS4vU
7DVVhCNk7rMY3caEfmlq7C3XkU/MhJ41Qydc+CzIKpicXWaM8l3H6pg6HJCtvIk+/oO53kZiJxyq
uKjwNW0lmMpwOu4fe0r0DzoB8NtoF0yX6LWmBZVIRDGeE1daMQw2kDSR9Odu6h2QajoAaenGyoxu
cSIrfdFPsiCPIqGm+4s67xlW8tjJL97xRXuqw2I32l7AKPtJJ7Wc0xDnfV3172zDzNm2X6Zjmplu
jyDOjS9ChYjAQnhZ2CfCxiDJ6u7noDJcKy6/fH2Sal0hJwdIw3ZFwMk6RdpjC1aT9k+fqm9oLdJR
Z+Kg1jILk1+7GhJl+5/Lj+sbPHULSS65nfs4O3VV7yY6KZvYjcQmkySCK/SMsIFknMCOMaxPb20P
PYPYly/n5DykDNQDoQ755OiRl7VYwZ3HFcxatcU2Ib0y1Cjsm8LgqaKKdDjRU24QwS5PStNeF94g
DFlG5C2ftE6nLo6xNNeyh406Ad0Vu7ZVhYarZRwQqDLvAqvXycb/62E+8DVg3TYQLBvfKkbt/0wu
VTgrwrOe5uLqEJ9oohiDSzoXqHhHuL6+JYIdx/c1sC+oJZFTiJ5/Zr/SWRuBjlPGUQSI/j062J+H
L0UC8rhcMC6YrJ2GbCiPs3Ef85WWYfD6tV+f3GW5/yk45tghkvFnvn8W8i/4k++My0+B12TD2eIX
gSOeH9y4GSkho/UbuN9vOiqHH4VCF9lkpSxU/SrXBIGDBnkKA5RT8sH8Wy70HEI7FpdCpxC9P54m
sBehY9mRN9Eq44QO2rMen0wI7q1x/zGS9oUrAWEBS6/I63A6sS2Ntu6SMvKbV7JZyXrLsoQTnT9/
hz8eGGqGnfvqUXs7UnLJVbLjHgpEtAYxYcIHctQdY/ptJKNSDUkiVDFjK/AJvKcRlz1/vsI5r1Bf
dzhk0+3nAhfh6wYFcgyHLkgF+EwgcG3LnuppnymtQfvH5fDoHsMsob1SnYBWgGfMBtUBaevx89hO
93EI+6cMPMGqSk4Z94/NxArTZMGK8bJye7AoZHLXJPCgR29+UP1UZJe+9DXoQbsF64Fg4jkirnFZ
NW4vJT7kMQG9CYtV/dUgl7Ybk1fXv2LtRUaZOJU7CvcCs8QaVxG1ZWAl8if9EA8i0T7h1bZ+D0VC
XrdRWQsi1krI4rChQLL+5/OUmC5fVf5/rggjqX61+TpU9jGzZR/Ke3mfhCTMUQcd4yxiH3K5O7o2
BJAhGtNz9nxTMbu0DceiZ5Ej1qPM+BAXkItmUJf1hiMNEb/JHWgd8nP/lukPNpU87qHYF/FWq7YG
xbuq+eQm4zr7DHOWRsXdKux4/AUf1eYTxF2pda96uFWneAhz9mNKZsakABzCpGMYZvmqRpv/5qhC
y5+nqdxz7sci9UwQCyNIRJgGC3aq3OKWtjxDnb0/Rin1e2VoBHjJL6ijqw0Oqn7sDrBiXVSzijjN
Ld1UWJ8ftBTnETw5eNSx85sDqFVWn+cSymg48aal97cmqmGm3Q5wgOT3BgU+NYXZzKgW+HzhBfnq
ybGny7KeVU9jfKHhJboPgCGEFg0FydbEW3OIIeNcqrJiYu+s3AHORMVi5Y2GRQiazKUum8L/fxVp
PwDfTHGDhoMDG8P4EJRc7f0XI1AxANzRgM8P15dvO759o2nHIhi9w3TZFp9Hx5ohJEbXhh/LPlps
zqzc1Nhh0FV4OcUEF0Z0s3GgfqbJfNn9hlWv7zPyu/r1ZYZX2XiwcRwnQtoHVHDHt+mTHbEr0jNT
1iqAyeqKwnJgdTODtrdmzczigtBq+hRamCYeI6FGAFYoUbvQkBEH62kvuOigfIoWnSdM8JSKPv3u
sI/8i2MRzLzjEpCi+qLOcSwIW2+E4uRuR4ezgZlzqBiB/PBsmZ7po54s5R1vpMr7j99qta9Cc3Mm
g2j4t0ALI6AwIhrXPIqMWI3MlvjUyXk6Wc5FX1K2o/m8wNrnM29WNBRDaN3nUFFeznh7BKncHxlz
aeexj5RjZgGKwJmZ3c+7QFmkYwraU3yTanniQRJ7E5NCjhnPapE4osmN19/L27jD7wzdCTQQBjHo
LhHtQpIuW/tUAvKtu4mIZ/pH3jtGxGZvJt3CJUxMi7Vty1QtLHiGERwmPOm+ue8eRvpXL2NRRURb
p0erHBbL3SyNT/Li+UanRX0eoyzZdVAmQAx+wrlDkUFX5vLkwgW0EL+dGQ2hjPCZev3SqNtwXp7e
Qj6y4mqu43tJTBoie1IwerJDINx8m3lX/j5QN/LZF0a3Y9SID7+6ahQIAvbLRj63lPsOdcrP3XwS
a5j8ZfGt4uFy7G+mXJNPHt3Vko+l+ADP9p63RELaqTga6JBnKxxEMwj2FYU0ByWTWQQB1XYl8qXT
uIcwUVfVsxXfpaol5iIZD30YA0AXzkt7B13I8A8eX5QUP/EN504gDs6n43Hce/nNygs/KQXhkrjn
iMrYcqoaCFlVlo3P8s9rl2l61WNft4UsItbdf6ylUIbX2Er/oeWJt4kVe44cc26u3G/wPU0D0JrK
ALknhq2opRgh4/1EOBQNVDoKVIA+qtzkGUpGvrhlhx/5RvlBIXpys/m7WRpqTqK1h+hFt1NJFFuf
V4jU/rD9EldPELz36W9NroFs1LejqM2+7wccpPo9X0wVdXfXaHb17p2Li7PfgO8qDFlfqB35MEIq
WfhZ7+xNdnPDP/JDbKjY3hb4Vm6RnqYgyygkx/1pp4Ou4sFnMwG5VsDkfbKPyZmrFHPg2ElrOIrO
6NlzSI7gWxWG/GGaXa4OA7+bovc5rpIgwGjL26uEWfbMN4LVghC0GHpgE1JFU5HGpJXFR0hEqrRJ
grip/a5K0gDI1O5Q6sNCQG9/ytmNz4lq8KUHHqyU5GxBnarsXMK6CoZpshfBlfAdVRUunnu8Gbc3
BzFsbFmUQKTIHvfloFYLv+O2mhr6EZwGoBuQ60CmPubPBr+f1BLw4lyZLKYAx6W1BwB0OxC3U89P
Ty56Wvsmsc+GTHLUK8vn2phiJPgfoGMtNrKOuV7ubbt48CspHKaSNWrktgDos5SyJtbM/5QzljXz
KWBElhCd3KTgsbL09lX7rfGrukh3qjupbAHw0XWkcqan3JGn3JJBIAboyc9GiViNkuWzmKVAGTgi
3cWGvov1HqsO3g5/HJJSfetCYTQ4QGmPjMKDdsJxKj550ZDKcfqEnnhvVXwFv6uAi1ONvsyZyzmp
bpNUXiyN3dSEYYbZcTr0ekXmtbn6z5bigKKdyLlIZB7Sx8HQ7AIi2UYnX+OHXUPZ9u3f0Ue75E/T
rfuCFpHMKIwTT75j30TQRJuVRET0qPx2znRl30mEyMwhKgoQKmmo3dnidPyOMuA9UfMGHHnOrNSJ
7TqNtspizL31DC7iizml63WnFZwQRd56jGCOjkjqWKuh9i05vr6RZGg+YPaSryppnLSY0sUEpAaw
ExWhCKPD+/XVzyAOPaNFpOl8ImxH/T0DnLve38AWpe8hVcfoBRLuxyBqjD967EtjKpDpNdAsFyEV
Je4kiwDhCQsAHT9BTleZRZq5SNKXQjN15Ya0gHQe+v/Fwp6Q1TLuu8/k72TFbFB76Z6ep5F8GzV8
8RuOr3t80TfCIIOLVvKrtOcU49j8oEvT01F1aKocc46KoC+AI5QjxREfitVJvhNP2pC0tnp0fLEy
1Dzkt9x8a+L4DwSYtwoDCaVgBVdBAZMLIyjmoGNQoGib489WH3CZSKOTpaSRoN6/0AgbhK5qy4TB
VaQXd6AQsYIsjYl63x0Yfm6EJzuWncpxvGBrFO0qiNRrnBewUr7KIjaIjdQm2OGQce7sbSFK1ew0
4pBco8XJFxbp0PxLgFglFDbb0jyx4kBgi8LbwM1nikKY+Ik2CWnWUmC5QB2mbikQfeyZaypZWsc1
uSk2EgnyI6LAjTuMHY4UJFJwLTpKKUlBoF3hqB9WxtB8u50yVdwvoAdToe+E//kq0RkmJp9JDhge
W4J3krfjYHBVkvR0tca2unGtqFI9598RCjKpMVptSMibv4CbcAcjUZeo1xtBB8geMG93CIDwWCC6
cn1vj8aGwjoon5UvjEPVPj9wUfhKQUCqh9dBVx7JEi5kGct+rJ2M16Ky65oKBsfSZJjcdkT+0sm4
Q5AZyBxm4722YHAnQPYPbO4XayF1UPM2piUzNL+rXXQDk2H+uBhk6868gcU0nnS9LFrEeimcdL6L
qcdD8g82jL3jvPUnRpP/HtOrLESo+c4XS90nGAAN2imi5xsTYVUoGhC5NVAFQbNi3eJC/YiMl9D6
StqNKptvXi1HKhJiZQU3okrlGbDq5xHIdzIMvJ5Eaix6zbOXWTnAs0u1XaygdIv5zZS2bZhylO0P
++GJozSdwKIKHdWEF9q8SzkJl3/6lcXV9Yq/h3kAfNWE8lWilat0i0HhrB04jxDkiZEl2oA6DKky
H/bTe9gnqossI+/g6RkmCdQLorx6vNtvAgOnsHHZ3UwVY5+IhA95MVRGNy/uxJLhlCh57vzN8cAx
6WJVKeVgSvD6hcO3RMf8Fpnhme5Bw8yQicufOjJYgtfX2PomEYSPWfJBv/pbZroWSz3qlsgb0NTN
ImxH1PW8uoJwffRDJXqXA0BRsYFB/aqNSzyZHIemVRbMzwti3qI2M6cmHH6WU2J55Gw+os5Y0tWr
J0EM1alF5AONdiD/yBcaJVB+rxmCcnkwAk4lCy9QM36L8y1Qf0S6rDF3ZAuH1160zAW4ogcXuXw+
OQJxvrFjzBeWwMTBl1/n9d66ZA8J9eKT1N/v5pbzP7PkOVY4gKSZlNqJ4iv5L2tcG2lO9aY9LSxU
pCbpA8B4snGLKAarSbxu4lSW8f3IN98zqByRgw7YwNum2ExoJpSYtRk1yqY0oq2PRXbas022rQz2
1vji5MQQHUhMtnSXWfBO4DV6o834accO4eJNdFEJzip9WSytVBS5ywjgCtW59GL0GXevwVfAFQCI
t5SV+amrwl49AnSalchdbMXr0OEGXVfPt2g7+bRGg4H9UFnHKs1GyOqtJS3dxzUhzEsn6lkcNBZT
6AKoY7XzlWZSPAZSr1MVWclq+zcEJpeSRsq1sCRIieFUirAsTQzwX7UnW9wTtHgwFewI124O/kZ3
ZOg0Hn7Fi/bm2XNx7U8hRspKkbObkIqDy+6t+CqAuTj2frDEi4EAWtBwS2edK7GYvXeSDijr3hRm
tG9fx4Cp5zst1hx3VlxT9AL6c08Fuc5XCOxMYKJsHdkHBv2ycXyETDwkXd6sDYhYJNPhedB5n1Bo
3BL0En/t+wPwRjjDUhZ4dP8Y9XnM1UcgRNpBpBpooLGjbTxaC1KFPqM7fImNPsXNGnkWNVhr6XJK
653MADve5pdLo6+Bgr/b/im+lamuXC2u72CvgGQRxhIgie4TTh0w6eU0D0MyT8eO2oIiJy/YXV/m
VVaet4pjwukXAqchGBSe3mCtES6oSKVhaRMIHNOwWGEcpkI9sQ4X/mJBcl4cw2LvnJYEpHGKrdmD
H4/EwR5u3zBKfbBJ7Bu/5GxB+RhP/RVZWNJmj9VCCp66nigvaI2iK/cD80UF9BoQfLkViUBOe5Y2
Cj2Z+GjyxOwVM3Cx+4NrmN1QAlsNezZqYW5WiGHfx1/xFmkpMAtQPxPFDdN5XBo0kuK5ajJmooeL
5S7kYX5qqTEfCYUp51OPvdTXxCAqm4yKTgaeVTJgNUVde7D0h/GlFXYW2xwfRJzSNgeQUGaxKHFf
JO84wLiFY9asQ9dNJ9T60uMCJyEVG0YCONv/bbkkX4xTpfHfoAKMacRDSNpdwKS4ZK2j+0+Q/QFp
ZZvt7yaIQv4TWONOGrhOhJKkGgoxhEDlIw5XCAl8n6zfz2P4UCWtX3C3NLP3tCUSyzjT7ABddzcQ
hL4vxoxk8hzazfEQu6XyZyIdA9jzmUnJPSkGXCi+949ttPGDzA6E3iZTpU+r4x9Pne0h8s+dA9hz
NxoR0W10STqpRlb5ixNRTIqsid3Xd6UAc81wMC6JtwQ9uTvmhSd/fN70JRtpk+sKdtVFp459dDcT
OAOs84pkZHl3gAW9Ri3aB3fxwM/2PmZf44Y3i5ZOB2nBUyPnzhTEEE2nDjmjm+FylyIXn/HbRle/
CzaFZcpmXzc7l8vSR/D/IXc4EWVUzxT9KxWN2YevC/FkDjaXGrVysvrgxd+lXGyYzLjov2P4MWTF
Msw/Fpq3BM36OPak+PLPR7XDYxtehb0jFz/hrDSt6YXjLfqPKAIWbwKSGWQV6LFrOFW25xkL4j/n
zj2FcIt6X8VbN7OjNxIgRX6/0BG8vdes4e/PO3cAC7WYFzK7XgvIZEEbh0tihqpJty++EcNSZxha
4padCjqDOhokX0LM0KgKdKdPbEM/+of795oDYgNb46MFEs44eGe5pspQWXjkKDQ3BY77iVBzwOXp
RTzB7xmwwpo5VP39IxAqd0l2+i740bxJ+cf1yUyO6ojsJuBAI/okf6kNbjmm+4O/2Ngww8F7yj16
Y0WjR2J5q4gcFoTlzbG2TYvM97HxtF1cOLqm+NxA49iW+Be4NQi4mUoVX0XRvUOaoTGHHmS9ZFWH
ZJNjz6p3rfW+yMqYq6/woAN1OdGa6qY0vcM02LiRMboMEA4fDW5QofVaP5oKR0/F0f5si/P4oHhI
RK1NFR+xOGb1fyoIjTEcAkLc1QNzOFqaus+/9GwgFZQweforUzPL5j/ToInFYmFFKqV5a2rFvMmX
woOHfCQp5aYudDZ8fQSenPJXlEqKmuh1+OgLfs6553BAeTu4ZJh0ctm1/EupHzFzR+WDOV3fEh/x
EQ3GTk1bGOLCV9fqgs7tupnBRGUwJNgKJXMyGaf0udvLE1RXSrv+jyG5TpvW4KrQpklpx4SNcSdK
HCi+3hCwSyEnhkOTMpdIuN0J7qSCjBvAU5JzPtZI8YfwFFCJ0CgJrbtwaW5waLSMIrVUfILHm43O
2BZia/44I76YRVtwpx6jfxDQjofg0EhufC73Sg/O7iR+7UUIP8BuSHMkzfEo75OSmsZJN5tt7giE
wh5+cB6I8Fuzm+V3DHxSARwAnaeMAyPPuE9tWM74dCfNwJjj3kyq9N1jcDyF47u2pnYe0go5j7a+
BrIcBcFjGNEBe8+cL/yWzKEMnPrSLnuhnFhUZhc5u7FbveRnc13iK5j++qarGNTFoJ/gmimrtt8G
tF5JB4/s/g49pgplxmj7ONhWcFc59bWIwLu5KjY/gkhShevSvC/nEB6H2PQwkHo6ZQgBE1EfM7DW
NK4/v4ZQ6C9J7GwsISVXbG3WK7BfW8HitoN94xAx7QN7ru1O7fpfs2Je2MaaQTWLjjOgP2yrrfIB
pmVTuuyXSrJ5XojSZdNsDXu+fuhlqJLYdx5JmVlpL2B+s543uzbKUQCdzvh324aqzPX5nsT3dldq
rgAszCU69P6xnJYDwMkt74wNHNaRhaaUCcbtxnPujWFKO4j9s0KJcQTC/U3YoJmrQegalqMczkTa
GUeDAPxQhvWiP0exCxf4XyUR05i+YtuG4fTC+/GcZ9v+DVdVR9MLBlFY1bs9jHatxEXz4IX6G+2w
Z5KtBwWhU/zYXsbPPetGvlJCyUXQuIQkPy59aX3P+JysKGJzZxia2mh9+5sBOMuEttQv9K3F80nD
wdVR4WMfUby+p7qZUig3WDoZ1OZaCRqMzAFMuuhqha3iTKvM8HdyYHy1Jn0fSSSivPLtvxPiPYu/
wuL5G1yrvN1ybDkT+LGlf+r94YLzw36v4zd8u2UE+nnvvVQym7TLWJ51/ykqZjv8s7UqkFc8jFAj
eNAjjkNIJpXLhQjt8+4LBEbRgPdJRWSrRMdIA0OT0lGr+F7vUx0v+P/XQxUf8eyBAJDsClmQDWSL
EYE9WLsdUqD/+XSHW1JKbIuWSoPRgVp+KrSutRJAbxFB5xfbYsqWH4L52J1Q/B0zpxjhudUt5ZfB
wCRYi4Di+IxEXfRhRJ10T48XRkeDqhIaHTXoHplldVu7UtoHeYrdDnS30RPq1hXpsPLsU/F7bWVv
5G7czZSpMRriPAFmjGax6p/+lOPXt75epQKmZHTN1KukeHXVwpV/4QhmJpqGI+dJlIV2/CYOWKxa
tZ3hyorpiPIHn/+eQ7tSAyb/jQTzpKopcEVFwgPAyu9GCCkmtJYQX3lV6iVP7kiDUBc6wyZ+ta/r
yULFSsX/FdyNdpRWPd9TKiPHoDTizWYvvRdyWe2ms+fdMJt3eSfWJGR9UhnhTRDVZRK5R8VcVCOk
nMkmAFma4ThV13mKxAxzd9nxmv8NVHhMov9CZWhVSgO1z2bfRcY/ylzyPNQgVM8iV0d87kUeEUBx
xAKH4acVmjK0R7CD8Ph6ujIjLNgao55m8q73QNq5wCg/t0ovI07Gl41YsT2dmD+2rEadkvSJk67h
Y83WFj4eh3viFRD+Okbu8x+Cgx/nLSH4+9IjG3otkR753hiTErjRaPuWAx6jeOzNLh/GWIXbayx8
r+HM+IKm78p04uiOc9ZataaTAoEPDZiiW9Gc7DnUcwcYdzoEnfOrvmNN9XF5aLWipAMMnf872kwt
ar6bwGka/6wi6IDCzwLwb/FLVbeJAWxGVQmsa2s6hvhtPFKzDM4RYb8oClyoQOHBvalidRxnQ1Vb
8D8XViinvMHY68J3JN4YPgqTT2MGOM+u2NhwPTx1T8ocQGVx7dyuNLOkQkKkADCHCvmQzzD3YTws
/s05W1FZLQSTHKPCVwhRhuNqAugw3Gifl/adzS/sIk/7ERPG9kwyowDkGXi0tCu4z68N9qfu6Hsx
2zM03JDknQkNjEhphjXxme9B/f0u1oQn8GbfZ/c3gvMNYinBepRBTtku5tQCCxwztajqN67qaaRi
XkZhc2p6ghVGdLGCBZI3LvHUr8fSpPk2znhm4oFV5RvX9R0CMXRXJsSOL3WRymL7ObQm3v4gMyPm
m2XRTX09HmpC4YtAUetASZ6Xbh4YpWuTkP9mJfuygkq71o2p7oVsN/WQgd269GtgtHVx72OtH/4H
eWCmirGyLfsaqig8ER77bvHS7Xv5ZIxBAYQ8Y8/pg5VaRdbA/8tKGeFnjOWyGc91+eMqsGNJTdjO
65CeFaaMkyOmBiJb2cPu1Z/wR1DLooVXX2skD8YGu3ycmJ1E+wWQCXdGmky0Jh1bgGwO37rSxg1Z
D7B/mr0d6u996poRFz+wR51ANZHnRi7f8s0/lul0cd2w3Cxl4c/SOWY4iTM0Zh9MvGQnkvio/2Zl
ODu9H5zBcChefNjh4fCmdkeWnmU1oSVsbiQc2w1yRoxL2Dna7zjd17XFnPWSujuCCF8C5bwVRu/o
zTi1LZIFSZ7x+Y31WRDuih9avYtg1Wq+WkKmc9MrHI2etss8h5w2GKQyQ8c084DbYlnSSMQD9CFL
WV8jfXrlEmAC8/GMXhqofwHp/A1niVEHkhcZhV+T2UtVi2V70MWeatqFixBgxrlC8u4CGPtEFFOL
kZCbnFsgktbPiKaQFlcia9dkEAfQO7+rLS9WnwypQp9NjnuH0m4WnlKhEUCukG8Ph8YLOudeTeTa
NqcKmE/Z19c1KCXTpHzoD5X5izLbsL9IQxEAXj52+JvIfG936Xd09eA8X/Km36R2SfHIROWkYaHW
nwxw46zkxj+dp2mc7c9Ap98hWKrAdPPgeAN8EHd6NG3pUn9p0Z3E2hLA0QAGCerz7HEYymeEn0VT
dtdt/oKp7dNEGR3Mq5+tYqe5f1Mf6c94zCohXsGUobr4QYZrxBf4ROPntWsmflPxYOhjrDaW3c9a
pIahhfuSsAIlSGvSlGQAmmfeth59ParQXxJnwDa92iev9dTUx7WC29mLIM6NpXtfpUH6VP0XldNr
6+HC9MOJfqlEk+sijwykwnFCzVAHXa3LsVoszwDm8x+Lji8/nxr7QJSk4UEacDgFYiGFojwdzxoc
3D+eRad7mBJ6IP6W9vanE4RiPzXQKEllIOZm2VKVdwVEKz0Yf/tncOt2ou8I8lGsfDhk8C9NS2zU
DZolQcv04/fzoE9aZUQ908AJhH8n6d5jKCclocz8u7/pI25nd88nTCxzFGcoQPnwjIIYsW/AezRl
PM4V8DivhaTMzdYjO9v4pdzwVwC76l+bpWsNazDo7kw1syjOFeXEUMJ+Fh8oUByj55a5J1HY5xK7
XImuAjmUvfe23IYnkTIZKTwwloUuxU2EVOr3s+M1ReIkxgYVuaEmAY0AgH+fzIzv8DKmB/98c8qA
rCElI1dxoaYMIO9HX0/nnA6YRqnZwrXGrgkTDtV25lbm6/jK08MkngnOJUQ+f3292i+m5+IyvuO2
kyq/9TmCOjeBLiwQo8WZMRH5T97O4hS2UZ3dF5RSUCFt+h7pnuyigAeqmRC2E15v8V3aSdtISH72
eBrwJPex63Aig3NZz96jYphrQZOUiEFvPoQvp7espUz9QHRkpx8qOvqfBRMzlwadzH03lDBRMgX4
Vld07OoIKzIYMEZ/dsXXFHdAsZZW4L0d8SBufSfs8N06YwM8t52xUiSzs4UZN9FwNgO6rfV+BlXZ
ll7ehQY5A72ioeLnaPOXKISwA03Z/FqN2gTT/Czbf37jEtMVfWPBpq/OqYM1HG6qlNZJP8BMcmY7
8NryVnFJotRnNoEPvKsXwv4BRrix0cNfaHUMrfq1p5Z9KfpC8QlSlovNlLWza2RiwBjgBgfONHCN
mKznamGgZLpJdUAO2h0jcUL9/Q5Bq4oNAM5UBZZWUlWTkZu0fex5x8z1SUWhdKIIR35rJYMTkfTM
zkOd0pBb+OczDZUd9OE/kl2K1JEdlrrmmtYXBUacA2erBgXkFU0ITUipc6sypSwyStj1vljzqTIn
eG0jG8BS2yQyMbR3GhDQsCWjQoCkPWHu1rcRqz8nuCl2tq6GaMR0oesTLN+UuUMk15GglEkLWVhG
xnPzy1P+hHOER3QhHJNR/5dNiBZd2uPYVD9fYkQNa8RByBJORvUU4WoQOiGqfXW7mOKljk4QI/Ni
DZ9MfR4U85rDL0HIqz/DjfQNMphmDIggMKqSXoNe9vF1GbRFWTtcHf0hH0v9JPZBiiqzEIzcAWWT
31bbl6qYc7wTVwBV09u6qvbmQeOeIap65DB8iTblBqaoV0lnbvHfjHTf8CpXvBIWPGhXAMujZyHF
sRmf0o8MfinA6/V7DzMmYOp/NKix5NbqDQWymF13T4RP6HwDI/aTVcHTVyOpOShBdQy1yNZHiJ6u
gv7kP8Cw2/Bpfx51OyC806fcirqYEADq/pLVEOnymd8DZdJl0Gc9yg1EndcdkjDlTu9AVxSBdQmr
S57wfpN5EZHtpZllJIk+sys2kqslu3Vh9K5uToztkvYdKzCAog08+bK0F02ji1YwfenQWzpjFhfG
ZWCNHYkkYYq+rpHPtiEE2/4OV/wA8wKq35rQxOcwigIIC6JeIVJpFCGH2+c5SBVK3ytMNZuN6In2
JfFffiDbxNFGUTrFYLuF6qEZ5pret7W9j9zZBc26/GM+JJaUcttIuMgXX8ihiZ5CmDpMiHNA3TJu
6GwRXMCCT+i3ZqqPhU+eYeX4XW6CYwP5vM0WpX/GY9zyVi/rKofjJfG0rnXT4qCeM+qlE3Hrv7mG
19GavXEYHN3is35mBDq5gj9w0QkZl3cAPEpapsRWpNYhnPnbJB2ozUcZtzp+Y5nALCtIwVUB8j51
Z5DbYOpxKjc7+w6VdG5u0o7a0AVSewZEbegp+Xi3T1eLMIsnYyNXoYbKzqmt+hhhRK7qSuT5DWSt
7RtjX6ffdR0nOJluoclNvdJVucip/Zgqn0a2kXb3PF6bFNzgcixOJjwe+7vGckEghXqXz+rhHjdz
84eDdJaGjWMhYSBcbRACD2KeWXpsOTB5dyCs1MObtZ8GL+SLNEFtW4hcBghQ6kyzeihdY129Pcnv
qBdjSG17ETIgWm+fA9PgjsMfCVw4CLxgn9rnFAzfBTtQzE2zy4cTlNhk1zCxxKyiw4D/9yofKbRQ
DMQpul2s3WhAVtkJu/O3Zc8VMXwkMzRm9OA6h5nmrfZEi2Oy959pzg3jA+N9VAvNhYaG0CCWDItv
ifBxFlCYY2xjBq69ckVtz/ZTylHBP/5NHxrSB40A9f06Jqq0jT37Nobtzim3vyghp8DG5cPz0eRF
7DUisnu4NttHNeyAm99sj6N1N504HambswQFEHWCI4VdY7f7ZggSzZ/wBeKvKJuQbEbwncL/XHxB
QQmfoAPXk1wcQNHXZIh1QNd1x/ErVw+/919nHV35DdNmFSFwpG85QotgkS+GO8Jb73zculbugvZK
H4OIJGmGKS/zjEYYipkWbx4MuzgOhwLP82uBTSV5ZBSzwfMN+rktBRh56ND0XQfy99E1ZbkGhKv7
EIAZQ8LC1QHw0XNPtiRNk3Zk7kjiSAgeTw0YC8dG1QTcGSYr/HkZcRdEXO4RekUo2jULLxONesEp
IDahF6jvB6WC3JneREpmdL1Z8Rc6k/0JkicGbmMRWxyyn2NURNYS+6cB3pSeg+HdPTru3aPIBa6n
fBNska/vzQd80OROQhU7t6gDnqvRc5hgbLaGrQ1NGDR8O++bM7V3BgF3wuHCB50isEyd0jc5LnYZ
ZmnP93I8GuzfJseodCPj1KkN6HvKFDP8p+A4NjyNUjEh+uHqPqBvS3/93Lr2EFze/tO8UJ3PJXCJ
dUutEt9NKwKky+JGKQyOtOHNHBVDzuB6wQiU0aQj0tBDPaJ+n2OwKRfD+iQMndogzkj2DSZquldP
9lizhJ16zY/LZOs1PrHkUc2bTJlasVt11m6AgubhQEoFLdvzsmsq/Y9DiSDaMBW9qESVrTqKa1Bq
TWHTvwx8a6rkMIzBEwm90BQlZenpX6sFp7uc+7XKtcxhDJiQD2xCOgEHvOxh7QIyeRtfquuSHFH8
rE72ZqaIi/fI8HrIvOdveYqbaX0x8hj1oYpQIJKDjdGDcWoG3jvPV5Q/OJjayXNzqMoTnN9Zs3Co
ROuMpe8iZuDu3UKQYKAwIwlfB4UFWm480CImF4ZjXbSRTt+DkOSCxmHzbT375FJ20nSMn2k0FUM+
aDHoYEE+ifmQQdUtCAhhIFQzetnlAqYZISAXnXrJFp/OzkFSYw98F/I4WP9HYVBiABnDfnHtKLHz
SJbJd+9LGnO0/RQFs5tWePqQMFpoGYxY4Mg0qoGf9X9rrDCPHc0+UdAle35RGMYvTESs4Cf2InbN
IqTspjypk95PBv7cYZopvSCG5VFHb7b4JvStcKIlMBgx9ZHhOJX7SwY4PdMaJi+7Lzsx3J8cXiSa
kH7ukEBvVQ3e/VzwrsAJqNIpcZz4fCWvg690g2cjKrkaEHDlxSJ5wKRH0UkfLaKNpb/eVe+nijOz
Y4ru+X2Iaw1v7n8mAgwQKJx2pChBigv5aN76xUoxcJBhxZ+ASQpQCu6cLksDQJH1q1rROE+7s2i7
v3YUMefwuiMA8aHr5eNFkVu1ZxGxZQCdLMdw+O50k10/uT5gvKXA7C9crMuy7I99EfDip7L3AwZO
IYSvdijSmVTsPkMIwDy5ZswES18xcEb01PjXTZ07XLwgty5mUdyWAnYJboX5MqoN6EGvKpnMtJBi
9TJ6NenII0ZAhSsAmtGrQAV+LAlotv6Vz74WKdOOYyiwF1DgeI+l02jIoBM+GV89D+/mnrWPQCg5
Px2rztX8e8D1dJowGZoS9S5TUGsEX8IFIWVTvS/M35F/58WK2h8ZAwhAlp/vjR8oG9o+7pOixaIF
jgT5yaSGgp9Bs5ICPa27Loz/FOuI8VxD8uJNRBOLqG5pIsR2oDe4E5PjvURADUT+1q6CrIMzKurj
Zo7msttGqMiW7KUd5nSsZxM2Qo5gJRTpI9fAs439NRDitbHCwRxiXqIRG3iZ9BwVGyz2FL/TZiBY
AZZyANjHSFmmniZMkPDco+/3ea5EmTrewkCAeTgxudcHiUXmJS9K2zkytHQhRaKdLpUxKfq1ERdh
kG481+ZaZ06x7uiaythfORcmeYFmEvZxu8+jw25YxNXnAQ2lU6JuWQ4K0gQiIJsEQ4mUci282Cjf
9ZfS/C/G40Zjpe3YGOqEOxbvxssXcRNHvkqgYBB7geVTNlm29Pr7tfCCwftwTrHK+u+X7jiNEItb
tR/Z8EuYFSeqCz5xcjQBJtSb14jSnfrYMtVOmZ8YutYrnDWIy32UIL+8xm8qI+x2lXSutSq2GBV6
mdZHyJAlJzQCYbXkMfCDzsM3ffzPnNpYyI+gQilkiWA8Yna73HtY0mqHcm1Ud2oOLxC3CN6W9eIN
nEPNksKt9BHNb8mnq6UoKCPS1Ys0EZARAv18UqH3SVd65S0HIr6n4N0EcKiBORl/MUL/oJMfAMQ/
09wrfLPg6X3pkk6+DhHWXkcbe6//JSV0OLhgHOafL+GnUKhABURoRp+VZ09O2j/CwILXwhco6afT
phvH0a2l/AWU1a/HWHRF/oer9c7XulxcTjfZ7bu3YHMIzjbqDa2C7qW7f3f+VirM6OkhTWuiB64z
/oJUySzd8TlTqFZYZJ2OhaJzXLjthc+jn9UdZb4hl4S2VuzhEcK8XPstdoaJ/BJTKz8m1WMgS3nw
AvlqiODFYptsN4ZqyPodAWkAhCJLm+pSoF/PV1gPbGCoS7U2H8hOUGYV7Non1EXxIs2HSTS1qvYa
SI06lw58CaiRY+4lKF2eIl7K0VYPeDqb3L8jSvUpaZtnPweD3Ah171dvajjgTQJJ0FClUXOzrrAJ
6sAeZr1LLquwSsXW4jYEdS1T/0jW7xr9VC8f/wjxuAadzBBIHvLDTdObF8xDA4lUq4Vz8uJiOPnY
24n+nWibYTnRYZqUZa6O1rYD59sZYSeka7bXD0RklVmEnAHEDqOfF5kxRJEyuxZ/tRutO4+8optA
3Oy/eGKEv8hUr9t1oEBTgn2Pw7uVPiNWcQnIG/gCW2cweZ5JJWtv4YDAD8k5DWq1B1RgUJsFj89a
ZEmiuaf5Q+4wclMSxZPzWdVNsNG6FFwFCxn4Dp13UGhpktlPNncQpXCzZ+ivlDjobJacvBSeuXd8
fG/e7t500E9z9e5G5FK/JdUJt6OnvXc4IjUQLYPXSxFqUxlYaB9EP6OJ5+fbXjxPTpfrzAHMFoSi
VyTwXrV0dZlobPKFJLXe+1OpCP/LZkb1rCKzM2FXuNkfwMWACnCvkpTiSgcQleUNnmwvX4bdcTBr
tQo8KJcdYJp0Ft0Y/L1yvztL6U1FDpZZNtSdNBuffu9GWdaMPJhvVPk7npUwQR3sq4rS+nAnABJ0
+NrEFCumL6AEhlpjdO5YcL5jl5sQKRpklULuNHEhYaIausTOuxdWegjiMvwZFDzmjnznABNN/Jmd
BoQ7G/ZH/CHUgP7nYv+C8KStnHZOIxDQvzZqq3zVIFRcHLkD4XaCqk5Y0oACHuyuEGcDVdLVPt1J
4af0PjoeXW4O6oZAvp48joN6adrapDwf1jrLM6fcdT+8jKkI1+wwGRx8NDb+If+6Gp5IXPBkMcfl
ESfc7ztJQaY4dGwS9vcZ/sPjjCCYgZzMOXyL+qgfV7xHdARy3f395CrxMFoeg7PLX3k0WF0n2Uff
siKDl8yWSd8ZZ4MxjKilqAgzUTMHx5SGFXgdgdx5FF7Fhpxh2T4kaHbFkKeu4N+PWWWo/nvmM46f
Bmw3PpD64ADDZNbenTpN6gk/CjhTYIJFZrFmjvtbEbe5Wbu+oCq4AoDi7d62GWJCibYKBhPvYWKL
TXOeTpkhGqiNueNSkn8nilBME/mAQATgcBc1w/HfGGzLjVyGDysw+yEm/38kY5GSSt0P+laoZLtW
veLJp2fiqZr+g2v3pagO5n63y5MASt6Vy/jl7PnWNNr2F9j4oXvPoSi6kPpfnqWUoR1hl4bGKPeO
7foxhtvrlkP6ZkI/7fwBQG+A7ZCo8n7VjbK/bgJLk/DCv2CdfrkYq9MQ/ySbrn8SiAQOnzrS6eEt
Ql5kGcbfSw0cukmDdzUwJyl+7JEA2nurjrrTC2wAkXz5E7zYKs1xG/UU1MhhAVS4RlvhyAZcNDz8
anNnd/Q+lLb3QcruupsgAncCxvOQtQKtEsRaTk6wbRYCJpfcNJXuzbwfDbzhinOSiXzxA6ZcRdSa
YOBy7e1E4WbxVsR9zzPLBP/ahMyV2lfN3MPE/rQqNmAhGl9OLOEcYazcmGQllgmKp9ajJoJowWSB
MUAu4gy0PXk5tofvVGm0iE4LjLJpAGwKmvEnam57LYjs4bfr6yR6JQITBQLc1J8s0EI1m7AWuuHb
9kHI6wwL+NIamKD5EYCyBhrTBspiZbrl71OQW61WYUlL4wDc7dmhsP413yWBHeA7WUPTdExLcXMe
uuUketnrVEvgOjfMn3Kptcr9+sZyiVpUb3mcb4VBc9pj2C4UG6gaTqxlzawt5Ae2j1pRagRTDJBa
qzVQCahm4QhlX5X3RoMlm2XYlkys9FJzj8fam184iM6jlAQrLwOHVnZReN/zsyhrFwFWizoOpnKT
sbNElHmtDVh9WhaRqJVqFVrkKtE9Kxsm/P8AFMapbVo8hZd0YuQwzX/5D91CN6WB/tHtNxYaGt2M
SWZz8FRLzWnXeU0xkL2oAFwTFQkzszLMWvfGBoPciPU6G6T1Lc2oPOBPTAw5EJTqbHpN0IgDAEfh
phQ1iX2LUSFtouK5lStn59Tgt5SXDC9mnCS8Vx5VBlEMXn8maw+2uuq8cS8rxpt9kqslA4JXyep6
LgI62O/fwb3jOGxwZy5gi6A6LliTS55beCzUDpO6t0D+BuwkIwQf7b3QytxKSQxjUF5W5JGGrzib
9NxXgTr+CgDgTBuFBs6vB3TefbBu5kqgjCyTIwL56TDJ2uuehz8JDC+/hlABklLW5g+WB7gjWkw3
wz+sBmCE1OtT43qb3WLORH/wam89vjf/yU9J3hvMu7ceQHNNDwQrVOt+dkDHCnTpPZNSmkHKjMV0
9w4H3syI3nbAgumxXfuhjV5peQwpX6qtpMb0gHK1tCSq66jJuYl5s29BXNDYRFcObGxlXNQ3OIV2
E22hBu7zXNpyKEyxDxiCkhDgt2JZMnsrscGkE6Sj/fUKYX6xotk49ItQIoyOc8KsEb6caF2U38Xj
sr2OddmCzvE6yrn4GW6t6KmcnFqRL3UDGwyIWYws59X+AIu+iuRUrBUWNbDS6C2IRgVQylnt/ldG
wRDQ8vm0Jx9bsdt2iV3UCqelmywpKbTpVJh7jH0bTP66LSZ3G2wMznOHYQuERW2WDUk7N9Ncwsb6
8t4rGhVRo5JG3kjDnSac8/Hmdzh9oODPpmXoOV6jsvtfdEHZ5hBL2PMomjr1m2oNWeh/kohH3PW6
SGUyYkDXsuCxJjHvr0kKLSw2Otb7uH7aT17rTtdizLrfP3R4b5pdTRymJtyasaLjZLeMf7yMFSue
++32Zbpud1aJQTgNmpf2vqR+xNN0TSaeQQurabqhVfwC1Ae4gpD2EHcDsL8Bd7xD+V1g5w5xx6iB
fFs3b2iPq3FNbz5eLF9zffaZYMKrbLtiae+pkzSswoanHi0Zi1HJjtf5L1fF+BOq4RcEG9LOqC7B
tBAHV0Gc/NdyFiarMy4A2qGovkDLjm/EbCafnG2bbf5xbpbXnBbEXdv9QeUrk02lEFAZgSms7j0Z
Wod0TL47ByEWI90MMgxPUD78b8aaAKpeLyNz3h570hdytPEYGXmEngh4THLJg5famOmWEVmGrqh2
3955dGsITzunc+MYr3xFQgzrFfDuhJJuAQNNnt4h3cB1BhuXi3jW+TH2de8lW3ackf4VfkRPlEw6
jFqaHeUswKyNjUonoOtUTfxCdwHhnKCy9F59eysREcFhWPYeLLKR0ijXCTioAr28Ony8z9tLXnF8
mALhnEbXKuFKDVb5aOACeFrgvAFR77Gg9/gSNUdCp2JquCGV6YxHRPM1m6oOI7gLw2HgjEp0Ia2z
4R92qOEHQvHH8mvTXuh8Iyq4stAujsXRN4pHb49KByBR3Rv9ahJ5HF8Ty+A4p2zOpwJeNcszaUQz
oPXOHJ0nCkEmSwfFDlPPOO8107dnT4D13qZ57mwg1sOKx5fEvmZvMjQowum2D+qIbwf5+HBZ2pcP
Xngesb40d6prFmY12uQemBG04M4/mzMFJNN3fCpdCJXuWmSc+bUX/ZZZgISOW4M/nPyErNHp8qwe
2s+s7Puv+XmHxiW8s9gcmTvzd9XTJ73J2KxLXsZPP8dUdcUt/PGAw/YZcgSd/r/GBH/0u6c+WdsN
peUv6LQBWrZNJ3r4iWIzkRP0gtqFO4LjVv/3U/ykOTSasaliaV0P3deG+vQrLJBCfJE5ADMwrjzh
eTqBtQduAZgXnsyIxZkTrkKCzYfhk5S41C8E63ai2ZA8cbDjUROiR4o2KlTxp1hLdp2j+NWKl5/V
AY8nWgYFfw77MnigFeFp/1VjoI4VzplbPjJjijohKhGL4UWDXi1dD2fIDFvroD381Vkx92FSA30k
r4hDWmLHI82DmRjU7GudQ0VXnZvNXjeJjMfDLZavHjy7OJ5Yli0DSZ4j8JrZ8EWeZyMxe4/AVtwb
je2nvWrcaRNhrn0uzXaL09UEj/kJa0D0t+DoLy3AeXsSpjoblhl4AEBGH3x0c5SBqSzBuEii+30D
QOQ7X7g4NQZTpqGS/UdPD8FDsWV0ZPGy5CBoze1SQhAXJUx+G2ilEjnURoaHyR1gg21jc+ShvUjg
4s/wCQP0CdtMWLcIz9J+B94LHG9HHhdFlKlimoL3HbdMHt3FCsS4ErW2oh/Qk5lKlBDt6wwKq6wB
lBadJZsGWpXmduQVaV7b4IedZ0aYBdit96iQV50T1qghYOmdQQuSuRsR++Gl8ZuUusxaaqZFEE4p
51zyZGRWtgDxkb/fUu/SX6LO0/DEF+T+KoLEReOa8kHnNEbvrVRXfPhiz7iW1r8JRC7rl6792pyG
unSakgSQbrx3MM8dqs3ZRDMpwnh7llT+qctY29bqTkBB6yAtgz9YnpRECu1zNwG0h/sk7dZuucS2
/iqUHnb1rXfI1HmdCFg39pEON6f4Y82Mba7YicYZAIfB9paWtFIfTxOw/FPa1qpJOFR3ORVlJMp1
Afv87Lc68OjMdMQoGxs95DVWR9cBR3clKR+rj2dR5T8knaqKTseZCiZOL6f0urn3mdBbJmTbJDUb
5dfLxOxE/nYSfrrFrFgrp33W5KpDqU7mqMxJjw+mzO6hVIyPQeZAXPNMQntPfJpH2ZyDHC6lGWPu
PgDI7ktd7HknFMHEhefP4cOKlaW1Z5DgidzD9DH3Pm8aTz1MhNns6je0kCWtsyzhZlkPxuWkUvGH
VK76flV34GCntIambiJmtN4L5V877Hm+mCJh08zNtuDqh229XnyvmoAMoFOQoqRht2C8gHfyg1q+
rRcg2kZBiKwYH3W/A7VtCxpfbOKVhYWYYQq8BD5zSd3WrbVaseT54R2AzWisk4tPkKdnnJYo+n9U
M4P3Gxxi/IHcFCKqBQN2gNUZHTgede6+WpS5EC2cllWKJM5cVziIMwJQfCIwyX63lWrSuDO6yIHx
ut7gEv6A6MSCNKWIuZC3T0mv/bqd/z8fitTKVOk+ygZlmcOjJYY1de3NEcvMj3JDKgqnUn0Jgk9d
sChCjP6DP2ZIBu0Jpz9N6D++HvWZLSejI7epnRYjQg2fwkqgdk/fYkU8ex53MYuTIbywlgymf/B5
0EEgZatqldsz6eicY5ar7V3wCbws+WBvsbPT5IoVnszkwNEB56JYUL1TNFDXbsLWATmH0+0zaVLW
9iwrDcvUqKAwCmfoi4RD6ffxHq6yCGRmvd2Tno0g5bPp+jwhehXIqlMGW5LhCZ3c4uL/WFsT0NCp
ugvWB6rxSpDUyX0/T7XsXFRlgCAF6KFPIJ2Lsv2NGBHysz+k/IdLctlW4WVhv0vQ21IjLixeVu8b
D6+udobOXDjKCbNNn0cSA+HEY23rSjVoU95KdW9q3A8w1XYazb8Kt3UEMy+k0RxsJrbS44chlDwF
3UK1icmkCcq2vrVgZHG102AY1jgfIdfRtMOZZh70B0/LKZkTcOLDWWFoIOXV7Gntwe9hL61/J3qJ
XMeYJHr97AjehM2mVbCFXe8AaICZMzy+6kWpi4vSKu+7fsWJaY6rgIn94+7eDmpdi86onB9TrUKL
e3SCof7UhiJ7uEenrGE5GSDu9kLh3CscDO36AAqmoikbIbvKO/wo17qR1qLampZotNaG17hPQzyz
rXrpVlarqaJOl+NQwWV2yoq8xytSrdnHGDOZ/IiZekYdPgGE0YTZfRbG7BIsC4UdxSvdt0NanwSz
kZPgf/JXzUfs1VisSCk97V6IgHgKtLsCmVL/Vw/sBbeGqBFu7wmwShZYuVOZDQcfl6OUAi5SROyE
bVKN1eYyKla22RA2DqBdwvNj5jgGCJvuSkyBOJLqxYsyeZzcID7KzgPQkL7eSmcWf/kYIShCj2UJ
L9EB9eAydXuHv/q2wtrYglrmFHezgLRN+MJ5v9faH5o1Opv0IkVrOsFk/DRAg15+LL5/P9Q8Jd86
2N13OvPNwsNFTwesvg+7anQuxebW7JFTGpiLDXJ3vmho5Qeuh1AqqQRLz5t4ZiLpUbw8tmf9ugpF
5zknSEredqy+pdW/l/fgf+SSHpBOd5y01ccmNLMToW5iIyHvN9bPWR8FpB0oSmm/+U32EcP3l2IW
8B3QU7I6RSjzahmqoyoJ8ewLCqrok2UdvC84LdchWO7AxsexfuzrDzl4rb9Xabgv2TPjDFNA85yW
CFj/Ue8/zs2OuykbUhDJUJ+IxwO+jKcGjyqwRAJ32QZtUrH0PvXHz1UiVj7O6c0RCRLa+r4YEz5a
BrhGhRJX9xo/lL7KAu7ahH3DqAtU92zKxH16H+HEMrHZzCaW5NzZXq6vxVu4GTt4mw/kWA/F03M9
bMU30YA0oIu+74FnCVr+EmQSr/BbVjLrW0sF5F1EvbJUYFBiLQVLrKpJhfaDzvSYyiXhiGkeZxNo
001/vjTaqMua5BCGemC1xnnn+2rcfVcR5jkfIf+n5uw0K58BbEfvbqR8fkfk7/5y3s4RsrMRauGs
fG93Mkcq86Y4LR1vccioqllAFuPT6idPHBkU8cRZe1Xnc3C6JOS9zx2mEz8i2fDt8YPT9ZArUaaN
NdY++3O/3U/QvSCI8UbeYqqNkrECPLwSOTALkjH64pL7ZZeemXNUm+Z6ydCSL0SSf8cbpe6PoaZ8
vzy/YDqpXK9vQOWJ8tFZIQIJyfm6XT5pByxqpIwOzA1S1A+Egu0Errt+itn+4Nj2SSycY2pJs8KU
BLn6FexYEtoUkWzQfIqFtw96xhubUvWIC2VLPs9aqOvyjhKOF/ViXWE6OWC5zSyesC+fl5BWIPdH
MUJyOFhEFL03NaJ2qAE1pRemEorDduJwKCVVpuBU6ReoD67ziH9KSq94Clc3vmbLwoDGQtdSZtQa
ncE8HY5iKsg41h0+4C6QetT6wm5XgtqbU8iihS053jj72nmggfx32YsrJQ9MQ3/1ALDdcEWVzj71
ZyHuT0wghaseWi0Zj/CQtX4NckzRrLZdSm9ouDhpCEO7g3hJXmNsl2X5OUCpU6gQ6wMB1QU9XxB2
/wLZOf6q9y+V1VPfN3IhO43usqb4U2WCFwplRch+IQwBWUxcoNV2G4AovAnQh24ydxWFu7GutzPf
p5VTre15eFUzLf+QgG7nkeLR4MWMGd0cc7TXtODDhVh/N2z33AnrVMTiT4Opi4Df+6FVLLPDmvJn
NshpdsD23L2GHQ+l46qdYlndVX+m4Jw7KLOQfx5sSPYSOLqAFeqlZaR19NqHQdITAB2eg6P0seLO
sWdis8t6zFHcMhaPwe/kBccgM2EVltZY5BK+WcsEq6uDT5k+0b0y3ejy924sQwxIDMDYcemieB21
kBtwqLmdijarKL6vQzrxuQK4o4hLNTWk2XG/XtY4gnVHAULOMmcLDZ+y+3MMLVYlIIy8L0Z/k6Yi
py+iE3GEwvQjrVdHVnBwij8WBRgmB/fke+nGaahTzhTuDEpSzkFyoe8u5BYo/29EaaDO0/yRjB9w
B31zgKbzM7Yyp1OtZcNJO/CRQTU54HZ/M/pjNvzeVVHFEadE2R2Jph+vu5epveJK8wnGueRCkdZA
oASdIGH3yfyUx+HtMG339nsOOqEufF+uhIuiN5uTa3HG8eMSSRAF0fcrX4vemx1RVrbh3i3gWaOP
KOAoutIZCbl5gQPxWsK46jjtCmN5UgA4OyUyVYFu6sZS/rL4KvPVh7gi7zcGJWM/w8cR4fGDO4tI
6PAuMzV4Kk4SRrkJXr+ye2L+ufXrX1iwmoakql4oRWSDzCiB8cyynnarlonBuH49pn5RN5Phj2W+
yctB1lYvQF4e6K0s+yAgfuJwOMm1DPpzM4DMxqEVtooau/oej6WtIr6zMU2k1LpeolyzU4kqv/7x
Fb/GWhW/IPJqJx4/b+HdCU+rYSWifLMrl0BuFN23AiO7drtDtBqbrUPfpZLlWEGQc75wJd5EfBof
neFh4fOBadtDBVGvd2PCQHM4jXFI1cdacNClPAQvX3EtJM0xkoIQR1+gl1kjnuHBEyxfh7P8ci3u
LUcqYv8hS85asmEm/1/81AMpB8j4HMH1TMruQneOFnfPjQp3rWNBM8jUA2YlaCYJJzoPEm8g1W6K
XWEN20ePZM+tC6yZHpS2/SEoUCbZQeDxMFHEFdOsxMsWzvbd35f5DfOv6QlkoZ+jMrLiWNe9cQw9
LL8WDzbxnD8+LZSGWMA0QZYy4eSoNPJDZdlxvBv/Nso8KjmtfgHzCWGXwSzOKmt6W4VeQKF3ikI/
asbvshyei313wC+4irlIl00L3MksVw0QIBiRzNZJ18B5IKTWRQptbPobCmyDkwGRAlATEJJSmHxx
ngvo5OXnGrn5bNrZaavs9QGvt2uPvzObRf/rUc5o1DfYmxEyWbXiMdKtnfXHrgOnFzmEyk6mHvQQ
S76vlfXS1mAis4MkLuP/LSE+ENnjjeuWw88KGX/9H/OMYDhK9YK0boCp3wqqqG7Dg2QovlusOtIQ
/xEJv8+laJos8Na4ABPSe+4jDlc6nS4gklVjPl9Y91wHZt98YgjLYliTKBiTQuyQPpkY3JTdO6se
QITA7ordB9ae8c8JKOu6XnMxH/OI+ICyNJ2zWi4TxlwGfiPMCRmOK9ph4zyHgTtL1x5E6tlNGEgC
RxOoyNDrz1PNmTQRq6T6e3A5m2iWY+3ku1h1zRuKrXLzEqb9X7uD3DnHBJv9LO6fxUyLV6syY9yA
Yi6OFVr0Av1G4kypVfpUdByQyqeVxUqVOg8CBWZ25/MG6PEvSgIlpHxI2r3c8clXHGdUmAxe7SDl
uDfkFakc4Kp7Cs18K30N/X6Wrcq5bLWAXpQYuwOXhOekfnDZpjwQuzMBR/eErfIqB8M+ib0SykbJ
hr3F1gFlRn4A0gH+M7kSZD5Ec7+On0ZMIv2JBkS2YFzQekTqWuhzpyRam8V0ooevorGLPJnlzHit
PcfwLSslBa7tm/OiS5/NZkiAOAu9IaSSKM/1lZgU8aWjMBOmvVZAbw7oxm0YUGeADS4WRTgMN9qF
0DUkm8sCNj47t92+G8Y8JXgW0hZKEe83LRKy7q8k1jaIeB/bCFwrTb9FGuS01q7lpMJUCU1At2fQ
5uDdOM6n082FIVh3s5UJWqsxE7TIR/DyeLf/dZ33TBp0U3fRDhAqtwxNf7shbOZyt3hhJHysvbkg
Gfqy36o6ZhqybeyXFsEZusC89mfDuMC1FSOZHEWO7ZkOuvkqLk56IUStGuHVRb6ehKfEFQS/Jt/c
DrkKTxcu0zy9sK/KPoNjgGYxIb7vozFjyv/ua/TeVKmuW/jnkqIenoZ5CGDVfZ1RG2k/HtutDn2u
oFGYu5JY3ryhncloqjIjqlewiGK+5iqr9p8QjD6BaWkx+VPKoaKSS5+d+tNvQG/dhayQYFxP85LQ
erZYnw8jhQi1Btei5SjBhataLlGwGz9700e7M6LAL/W3MVnLQ6qVRDQEy8kTDpnrATzIIBhQ31kP
KiYnp9w+T6B0ytmjtTrqqXjzw10y81rMYJdLYt67iW/g8QvgFOEfHq4CD/xh3j1olOZteeZONtZm
FZ+Ab5tZi4J2DZqK9xhbhkwzHzZF8rSpaND6HcsLz3HaD6+DEKmXDY1DLHuOax+jL38TExD+dbo6
gEQKMlOLzgcIaU1zr7qDBA4zxn8C1iGVeHtXd9/oG2rU0odAFx8q4IbkiBFwmZmV6gQ98v0LrQA8
MDZHqdvrJpRefB9KE6+0R5Rfq2jSsVxVqX5HVWSOLOBrQQnzNvJLPvyZRJ8I6X8bZqDY9lEXTMHn
wmAe3+GGexLxDZtcyqevU2eHZl0L14XGLi5kAFNy5s/k3hxn309MUOBVxeER3lsOeZDiaQXJt8aL
u91V2eqAvo1W95DG+NGcdkhzGv5mj8WIfOHhXiK2j3yh/I3HI/lA41fD95ta4tzyMFGywn/Lm6uE
yqyK16m7ZlJKAxr3mUzest50ukiBRvSh+Jv3AYn/k/+bC71OCziml6avOVnvG7hoQ14g2XxwmN36
UwVS2UnWjxMYTmdS37Eb/YvXZ/yxUaWICL+7fN/fI8ygpDmOV2pKUGgX0qYKG3YayeeTCHecE2mI
BnpR0A3Y7dPJ+nHMYwxwDOkEOouUES33dgtGDG2N9TOgRkVn+EseO8Ays/BJ2XvSS0KXjHrS59kS
H4WbI+jwOegXU2l9cfi4b/kdpUXOcUxcUAsffkuEE57gzcEGXD2L4Xd5qzWaO/rqjD+6N/eYHHhp
qycz0ii0AbHsR0mrJjQFbgfTrlglusX74+7ZFE+U+H+IiCyhvoM3jxEurnGykUa1rdX2ID7lLmYT
6oe7LvKkTAKvQuJiCkCeotPK3D+t8zQzfasAf5J0v3V6pCUc2V+9yNhiKutcoJhKOu7ApDdZYSqg
srxl6JclopI3WB0mjbvRWRXZ85mUuCpFA2C/m9jESfQEE8Kd4Gm9juZui3NQpQWlGFvaw2ZUtrr8
mY8MCA65r3uvYP7QaUkSKRM2z1+AquoNaKzBpCs7G/NHU8KAY2f0i5LFYDc5TNuKR7G7VcHRWouD
4sf+iKKFb0vf41/i0nwudxtzQ2L3sG0/CBkaPfK/Xe7qmY6lvA/c8H7BIF3hpdZxWB/zwfLogd3P
OdBuQUtUai/x8R1fLMhzikWDxsg+KVPTMsJ84w1tBXcX3N4I1GxxRiBhJRj225Gekbj6udohs8uF
k/bN6x/v0P3CNpyRnGnfb2PvowGd34An+r1qOubezaVotOoEzQ2ea+qT8DDsiC083P4hCgkmEOe1
QMkwAOoSm9aBC0wAREz2iv103FDl+e2vssgZNFhCshHHLf24bl5FDDZc1nU+86J7LRvulA+zfHuX
ZOEreVqSOenxu7q4bDnjMTRSicR5LLUbJEjYThd6YtND+H5zS5R4KByhN54NMK/KPSypDtQy3OE3
fnms/wGt/uZsiXMhvHDKXa5BTQY+sT5lniw+zsAmHqTu0K/ku7TQ3NdHuEy6HOGzskfQA8Mw4Woq
EBzRq5Yo/9jkvbPeyPGVf/CyrymuO+Y9RW8X8iFfwOziPtkhqga9GjGHr0yPi8CuP9yEt7q8ZZNt
93oF5qjtXhR3o7x+ip+1i58wUauKHifEeeLfto47woJzs7ZirbqGu88meAFaHiyUmxWGMpdXKh7E
9H8TH/HloqfiXTiMjPgSF9BxMeS4ZR+YhuJ5gFDguLGp6/BdWSbAzC5O2OlboLgm+KHLjwaNpgiy
gsui9JhKrplIp/zPHCA+KWJnTfZEa8zU9F06vMJw7kwsF2v0GJp15QoBw/Fk4gNgyAkXzD8xVTs+
33fzBmGqHEUJdJ9d/5ggPLp6caZ6N6VtrMjYXOYkvwBS8E+lUp2BZhjsaj/YFjuFnIkYpnPsPUHM
WMWZYp4s41YXD+yZcsKazbVepbTguu2sTCPYB6AyUVb7YKNtMjre+Eom/hXW+oK+/eHZ8okSXeXE
qkH0tV0EIQRJTKGsxRevRLks16E91pQghWSDuiBNgnf/gIszrPyV3XAE8AV4PssBwZpMsQZ8CSoU
KL9KeHoe3EfNHerE3rbXFJg+iP8sn9zE45EJ32Bjf/ET5Fk7Ub670P1CqnDRhPzdQdTjGeWE8O+Z
mtM8vxH4SLyLN28/Dyn5GfMlYsqGsh27WPqAbZJrY68/G8z7ZmyBo2YtYVL4/WCFuX6dPhBomBVd
XdkfUVfXrLAQDyDLYJQPOqejogljGQ7fU2E3uLKwZ6cZaLDMeYqKGQUoVJsweosAWW6fF8/65Rl7
r6VF/NLCJD6tPQsVxlR1ZoGUmyKjciR26/LO4l3vLu4/kPR5Co5apqR8TDuaPbjEUfXkpWYgXziv
GAiuHWmFaHvUt349+n92GaH8uR24WDIh+fVpvG7EGJqIKlCY/XQ6tgpQU8P33BUKZg/8NN0SfukJ
UChjZD1QnExTs5Nvs0syYPRMzcAWRDoQyfpzX3MED4mMLvqIelMLg2QdkOI50TOEQ3wcQQgf29wZ
1D7KRZWF+k2jjceFMKTdbHXjdCXTp2pwXNqhQQf3FjztvxS6j6z+D5yWrtzvy5r/poVt8VOOLb4A
ewyFKI39wLH3TVFxYNU1V0pkKqe7fN3P7I4uv4e1SSJuZIkcvwR69QXAdPq8P7ZICX4miK6pbJ9B
wB95EFtnD9FPLL95L8XHOTGKPIuO+6yFFtLt8ZSZDTDvzd3dWqvc15oIrkI3fUpBVZCGOD2/V3/1
R7jM+CA0/zYEcGsI8iXnEsa5v6VSenSjraWXkZ7AH3CjgvJwYakrBnNOey5XNpLYfeeKrcoA8ypw
i6mDTuLFQ2AQlYi5XQgJy4i/DN2W8dfopUQEyPxfLruAbp9H07Nm+wGei2LTlgDl08PqX2txQ5Gl
EyJpmIWc2euiOjYib2N5S+NYxG0mdaIS5vlzzXHfsRKmQUWmsuD43QwSJ3XWrLgQUcgjR0VeK0Dn
0x5IiBa6JZiiYYWcpWg67NMvtjgklvWpaiVwwVzKdtogUun4xYohrGcfQHwtUWMwwxzB7+ChAR4y
ZsOTUTN/fbZdk7vSGv1QUZhy31rB0TD03JZX8Wkw4Pq7CfxpL/3XskOTEd63/1HfL5XfSJcKmC8G
iQ4H2xCXfUsdgpFVNGbP9/5OJYxb/t7cO9OLXfGsYiBROCgUHLT0GmSsOEuEFdrm5SVxxP2Fj+iY
KWZMk8DQMNIe712VUC5eX7NECHoXINLZ4KXIWPViljEmQ45Pn6fcOGVhflgQypdB9IJApO95T6WJ
F2vHTEfddJeGyhvlWLiWzZCivA4qDvVYh05Ds0V7rBrUUma8yUNaE+VNQQHkPBPHHLqBNx/zPr9W
cLXH8HM672l91S/fKklfdemA9oOuYgTCFmB2JdfDxpF8JHmf8lH4+qpVNW6hU06+jYjg6xFzJMJl
Liml5B9UOVh5M25PxlEBvSC4eBvU2u8OrJEJJ67ns1vifxBtxoPB7zmR1nWKVBEwNj8ojQsSdO05
RerPQF8IY7ktPGzTKCGe1RUuni/wvwOcgVQ+o6iC/OxRnjxiWKE/DNCyerp/FCL3SnZ1lltdq9XJ
jxNzLeAeMXWmSyN4ZX9MRt5JU3phxAUWAIARAEoIqIyAn/jGVzkvd0OpiU4dMcRVBX51hMDFRC2B
TC12ebd+PtLc2447Kz20/0w0GEvM1c73JmUgZd30elqTdK5k+l4Il2iDcAYoA9/q/+JTnZOLfhZW
eyXUiSvVufITUa3G+oLPin2CvDszq3cVvbAqdjCEVG7obG9iIV6kj0OjvaovzmTjQlCvW5X7S5Ax
4j876YxaesZ7+7YaUTDALZ2S23ROMXp2HS8DGEWk3dSxgehfLmtGYdOl2N9y0pRzMtzslB03tQTB
6jHQors1U6zRH9MZ9v00wLa23TGUztgdsAPJNRaifNlQV1DHpqZUxjQKiQUcGU2nC5Ml9XPLfQkJ
a40297eDc54SUXxeBzhf3I5xXcFVIUBj5vhtU9ysBHK4BRT0hOA6Jf3As5KowV9XvTkMvEumIroR
SIblAlt1KbGb3kH+DPoqrM1DUmMz6kfXxxt3DJVrttCnY0cRbgk0ffWLD83aDPFqEeBLzXrsuRkM
m+aLfSW5whWDFc4nTphXWlrq0xnSoDjwsie4w7hOJY72RpAEopUPsN+S+lLM16fZjUfe1/hkyL3H
szu/BBKGMuxYI7eixga3WhnU52CRPXXtMnhqYecgqLhgQ/nTWrro7GLs6QfTBXO2BV5z8hECS7mO
1ydbrvJwwQZVU071yEO+dMU48zaBFzqI0SMMEPdCIfjKzbYQ3jc3u2owPy1VN25GZptUmLUuaavr
L7Em8Y7NYIyhs0BUCWw0jKhkusQFbZCucSlm7JM7tuTP0k/oALyQZV9NWqINHOpaR2gA50fzcSQ2
0g8vS8ZBtKPWXHnUTIqMOvXmEMIkmBlOCnYjZLjb2uDD4Lqs6C4GrqBarWRny0/eWa818L9JtCxV
uMTQMkpejbVc3ibrZnMlm+KmlOSodZSg1snssKN72gTQ4eCKj3aboSET9Nm/DjNvv8CW/syX8QWE
dhur8tkcnUrOwDf6t6XOMqIhje3Mav6284PNbGkKeZ36HfzBCcgHy9qXeeD4gbCq8pFhq6/kyOOs
D3VygC0tkduCyP2gwoul3FurkfKgQSHF6mmwjb7KMO07+y8wjw7GTiWUGcso/2UoTAPDPK+UnsjT
ZpazXgSloZTMHwEP2h/osc2ThtZCFsTG4Y0ypfRycXvCdIFW0TALtD9f8tnkJOKkW1h6FIQOULE6
QALQvxPPKkLLsv2JzyyVYE+QI5L5hPqrD2st3zp6OhI6D4qXE3jDyrDVrrkP+jXUw751N4X5KbGP
kGYWGGEjW1x9BWDGIuzAlK05n/OjwBV+kdDnhR6qS8GyPbEmnhtkyurcTjoKXRZBPS+8CKLgAjZX
2p49BLxPR6SYPBsUom85/L1gifNs9py+xQNp+tk0AI5NjAc+9LX8oQX6ZqWeIYJduHSMQmtZ0nSX
+fB3qOVbVaspz5XM39htLO4oXj/qiWWab1NraVxulFgmwgzbMBo8XGzyytyvxmisKbdQA/AB7cyF
FPR+SO3NtMn25tbXWT5mVbawLUjK717nm1TJXBKjxHXkrqcqgNTzjt96/uFs4h7LzOkaXBEBA5Cu
iNPN387OxIsuJ8LMbgMONXRpBci+fJlO1iT5vIcxw5orgvgpFiK2RybAkWIQA1zq1JE4vaqeflXQ
lc2HE8r6eGTSfe0fGdaU6F73oahX1nqfpSN5rDjA7HGUtUb4ACO//BJIgFQXuNtzD2y8DRR1G5Lx
UsONjDcXa85ilFppEcvmZnZnhWCcKwmFhosKGfI/WaYm9ZrGI7z5lMYdY24AsEJ+5RZ2VrTLLJ1G
2QanSiP+v6mFe2JjFs7sl4c2tRnGiV7lGohJ9ODnTIHGOUvgP8wyEc+oGzmahnPb1QA4sBWfKRAS
E/JE2X+vcPiygniqNhe06CmPqM9p5y13+j9huNfxG4vQmyEXDQObmPAK2y0lpeWpTBhflZuU2FM5
jfYG4pDiLJHMQbe7cAEutPJarWHWkf3bsGDwIx9zjClCftIvscndyXHHl6K5gs2LfeKCrAZtfxjJ
KwUQh3q9NEX9A5IfnZRuT1Focej0UNRhLLmVlXfFpTdiJO6gzBnSGoweE9Ft8gbeLjMYbLHzzLKa
2J7DZaPDvUuvV+Hq4E3A7fQkLleSPUXJVuuPB9BHFmBuS/d31HhGFlil6WkZTI21XPveRcy8iIpk
nLLbyHV2/k8ZNPTb8VkTGM1RsesK1Xcy5DTRzHHXOpnnPrfJNy/GE3VqPBUS3jYQdsMZxMARdY7w
jy4png3GU7z25HutMP+cq7Q7UdxBsM/mN+zpEcJEjOD4fzRXLOsUTP6FDKdCtuN/kbpJaN7D19lN
Ap7eS97Ngqy33QyjimvS14gBbBbQipYk/tsa+UE897HswWCKCjbHYSRX8V7QGycVodzOitrcWZB8
AAj7Kg8mhgHV0ToGd359dHIHgq2+Bdp9ai1oyjBhioYQsXiSIXO/bXgyHTuwhv2m2q/2SBesDHfM
Pp+TpBOK2BxQp80O+md0cwsbHZz8lxkyPC0l8QUFalondUuczySe9sRMBTIc9+C4AoLMRGIyx5aB
klYqNtQDLNOdmh+TV2CFV3MAMtmQDnxYEfEAQ6tRjJsgF6vaZ2QOcBR47qT6RaMuL8CnP9k3+IoN
Z3I6+9klkbMzswTXEllsMhGlTN2bZJmAL17ZWPKluvqwbOEq+pMixvQHuE0benIhXAcPnsCoIBIr
8oL3C7gFgfjfNzmpV+JrGC59HB/lrIQWAq1a/me49UfL0WbhNRDyR+ewhctyeMx9RG/KyPG3BFDJ
JHxEx5QrIbB0qvdv1BT9Hcanl8mkinfbkWxdGFovTEQA2nUpI0C4qZZFOwzqBERlNcRguxIV5euQ
PbiuRIPZ2VmWWZ7ZD08mqkkHs2ELfx7MZzvt5/nY1Zt/V/DBFDAnzcs7bMM8PuVoniV8jltEEdIB
7SdJa1RejHyPhfk7RfGSxFoXlQ1jl5WHgLvPqjQY9WtvEXqLb1NS4vBadAzJNr363qIZHyBIILRM
mg7DIgF1S8w0RpUuGZUgKa7y1FugTG65XwZvtKWiAcx+9GaaIt2H4v1lrjbIlGSZNr8oAe4Xf9FB
EjcLoKMWsWrkYsVHhr7utK979G2SFsQx91RLjAbT31Z6FfCJ7VgKJATqvzlSF8SplR91FmR/q6RU
WmE2llwGp3WUtfFt+i9oMZ++oQSmsKOk1MUZT/8fN/51lLHMV0u8bUBIPEbstx9B8hksDYmuX+/A
wOGQu7dftkMP4U6EnibzxvTyT2Np6XezIKrPvgrsl4QnZLGDD26beveqt97fek9nT5nPKfaw5/u5
h/D7TF2isWD21jzit9uhYecqQ4GxFjDMNHLncite8Hle983Lfx0d8l8YO5zAhUh7EIfmQa/9AlXe
Jq50lwwXR8BvzviX2iYAVVxcUabTniOdhIBn2y/oVenOWBXMMDTj31UFQYYodYdY06DVBye9m+e3
tCvvVlEyBARthIxQqcjUmTqKs2gammAiVl99Z2yELjsFIJchitoC+FpVCq293EX0cxl6DGAALqnN
v/b6WvUMlrOvCRh7e6euywTqY4XTE/wGVZtduCqgWz0gymD9/QNhpeAWdGvORh010ZOzdDNto/0I
jkwda7i2FsVUSbeWup7fQK/BQ/hev/De2iWd1ldB/oLWgDw+48rrtJ796ukpATpPGFPoIijDPK+E
o/dsyYWWQMGvDh7YlW9neH57f9F//kZS7/oV9XUXBUB5uXcHfuEvw2cvbKUBFRtCWR6eTYiuP1Fi
fhvAoyl44bQapwJXDNvy+dsSgN8o+g+rYLaMLDR9pLGdaSnDkV6JeAIX1GA9bcKQi+luCiPmMVDB
q06Cv4mXePN+sAM3gm5ee1edA4uu6PYCqm9qgrO9m31610ziDTr2AXRc12a+CzAgeY5bC4d+sCPB
pb+vPo6KAjr3oeMrEQNdcelT1Wm0j4pJmPTrGTf+sGG/Hzhq8sFwdyx+r5rXOTIiZozC9yUtS/bi
biFS3vfMkhaiE8lKMPxxG3g9MlMPJMeB+WopzxfJEo3Y+D3aUj8Ni3AxoJBP5r8VnT8nAGXFFC7m
76e5sgjZ3iEGuXVMxm0OaJF+Nxnn4WZ2VGMytIqKUS5wyhBlPdh4xaFcMDpiCuMheXSD2NsG0QbD
LzXglIQOppJWnJB/FxEFinLqBvqgNzFPU/G4dY4Go5eKGCBVpOTsJbhNo/k8OPTbGnO701LnOz6P
3X6DWweQTB5HOmo44zgQcBmFlaNd3995d04Rb8UkWEJmubkWBd+Rw9yOgzXB++C0+TP2wiPtvOkU
63Ir6I26ua54riNMqVaPM8MyKwykvsXjL4FOEJs11rLlIqoZOQtw0kOSa8ggMsxITm0Ho1TG4wEx
KGCAlv4QdfSCM+AjruIzCew9NKfoTT+gpYnqSgiuhHeWQtrZETksi5mLK3gaJ4AocOuLPysKlI0c
MLdtxUv1zCuEbcExwiEyMRD7DML1PzgJF4GW7QLXdJIbc2P9GyZtvZOYOH27ZBe0a4sX4TZTms7F
tQWM6usp4T54Ho83tk4B6kDagGhW+8kXQfH+PXn/6ZHjzdwR47Dhr73eia1YovdiJUb/DoJWqdcL
0jtTAypzxJggM2/Js0LgJFGrXMUPkrGEyP1TME3S/j1D0Gq8p1ntyUkA4prprFt5cWK/qzI8fUmD
Dfo583YX88pFrIE7TLzzmDCMuylyFMvbcRuzF6zWYHVCi6xe5B9n/PIOKYau847+IkzAkVJTmrK9
aXJMwx0FRdJkiev3FkVt5awT8sKRszQKnPFur9mjm+zKsmk3LSHqcNRHerY01TPe2JPPRVRnh/dX
oTGe1DbAGtotlabgdNUElNXilBk0yllE7Q9JlHWUsoshEh7FOCo/t5bqW27SBt/hfI95VISscRK9
Zze2UyAthU9T1bWQg6Mu4+GPiHQYe8wSkNZoVuj5GVAwOHf7p09JSd4/Vudnbck5eoOiIEWStFv3
WtWRTWE6uNMSPpV0mkFomKlpIpVaOCMUAghm+VJ44ePLQek7uueXugUhNmBqzK90nSBqZeHpqxgA
QlTD9ObNne59aAqBGeCublg7R/k2jxu2d3Ofm7hZHJVKB1zdbctdobjENXsRX/GGkxZJ8SXxPZMn
/ZvUYsVGMflLp/IPf2jD63PfCHETCMz/tUC38ju0BM477c3hRfp9mep2HI0LQxz9lgooVDzcDW6n
Cm+ILZghuUGIfH9JvBeKTSlW4kzauSBAEaNR4bV1Jt96R91auUH8gei73y5vVk9H5RANJ1q/ao17
CWO5ZG5q9fLn0WSzKNfCcL6guZVNf9YenTZp8kZapy/2pXFQROCngHvYGyF/YCe5rrzm1boZtvUa
SGf+V5tPvLU1fzjByuL34k4ntHvVKLcKu3b3f8a9PgH940wrswlpJDDVkntEaUudPsdKQ/2XO7KX
9NwCrkZp2M6WUb2vSo0r9hiQVmq0i9+BHWFJ8QNMr9l0Zt3iKbt5nE3Fh+6jUVB0+2omJW1nsjnq
oojjWjdE49oRD87I6TxKQxPW3fycL8bnT1MXBl56Az+d8i9Jf05m7LQx9pKq3PEdg2tl+MLuNsqe
na+gRxCOBMI8Tio/XfGoNfmckGIldPWQvpbZSSECmc/WgDSolp09vPDL5OSNpsY5DrKnG+cjFT+G
HgolYPXI8qBnn6YYoQGA0kBwIPF8ZOW20vDU+ep02LkkLB/ywKs3LeB6uBayui6nCm8wBRqAJ65A
uwBtz9m8XV55VV6pzEHF+x/JcxGyEQZjdr5WrhpGXnTPRMED1ob72LnniEGQNFUtHgYzbGgxobsN
et/i3pvNkul50HJ5VWsNJCi7rK/PyDbqK3zJoXALfFe3Dfenr8YrjOTmzIATMC8Sdw7SkEgVgTTW
7z8oVo0ngj9ij/68Q0d7Qgui2o9ysUlS8m5PhsMsmOyhDduAB8FocJtUY9g+QMJxKfHF+ALgioJk
NhP8zK94bmj75Yv5AvWZwLwzdiUAtrgjhRxbQcNKekZEqPSYyrO9yv9oGfoXhE9inUd3rFmx5OrI
HKGxiMCZ2GAlAoNcCO435YFmqLLMlxcbKiQrbuBmyRtQu6h+/Y8jOL6rR0/dKYiMYQKmWsGRfZkD
5kp8JF4Lj8amUJis/or/SqqA5of18JO0XO/b+3C6hQeJGTQkLnSeKw3hHtnB4r26p+qUIAUuCjnf
T7qJLMJN0yX0rwYsYmsUStzj0PDK1y0GX5eAkGbufY/g9w2mKkTtOU4YwcBzMHjvuS90vUFUpAjZ
o6yoiSuNxOrP4jaLnyLZ8pcfdagHNUCmaGG5tSe1bOav2k/DbKocxWRbUwDohn7nHptVnpn5qIB8
3bcfT6OmtV/bTMYeWSE5YPvo7oCqlnQ/i7q9AYhEdGDkxwF2LqLksl2MFeTsyVOmQFoLybi7Fuxj
1Kax21PRJxGkn1ziyn1atM4t1S8YhAV0ldKXO5iopv/8h2tWog6WikmBN+/MqlqwdzDLVvgdyJHx
J9KF5UmWfwr5DNTJvwJPwUdfPGi/AOuijBnUj9k4iJFexJS6GMU8OJxPSiNVki5Ipqh2A0u0fI+u
RwkCBoUsb2RKs1Lmp6L/OJg5wAa8RkZZ7HybB8sjxRW1H71YR1tgvGyWhkEg4v3tUZycdcgs6FPz
pye010oLLDXCv1U/cXXF1AzwzwglLpyW6CzWs7/BXsffKbYSiviE94hPir3ugmr1oVMMkn++SJEl
PjRB6QzMzuWpIOCiVq8iKqKYKM/PuQCHPgEHBbb+6LQaIkzgl2R5Is0iWe0s3LIxgXsJhTT2GSO+
1yLf8a59lCau2mvFNsUAfJPtE0gwhjs0hhtpfoZKP3Ru0zPaxQ2knu/oUiLUp3+8Z95vtwzWhXGS
WT0Nyb/oCYhIcaP5E/xCfEAVMKCydWj5Ftg/amBJFQYIo5FRmjx0UtvMnpDmg1FfWssefYK/idyZ
bzPQ/sjV8MSNLxdgWFm8qamDn9rB6+1Kp3wjLuf/vXREGBczBUnDX5ztTO6CAr6k00xrHNN1Mz4W
NTVyOBRRPnhhDgRoB/DgmOPw56+5xFJiIKBECH9KxE8cEyB5WzPH2tlMhiSxqXb9R++vH3w7MEA2
s5C0s+kLbx2GipRg1rsBITImaxd9N1ouKwZq6noGOhdf+ybSeXyL6EBeZvF9FSeh/1+2vJgkLsL5
6gTT+qFtbS5ZWSwk3cqA0lcbKQlaHXpMaf8wHW2RooYt+8/uJz7H7cOoCODZWVLTWtjfvOfHY0EE
pdib+DQkAnc3wU2g7lJrVn9YHBgPMLk4JvF9NwVpEomf9iUdHC1vKeYXAoBecXDddwjaofH46OWH
FKHzUtdJcP+Bp0bC9WYZ2pTuUY6QYkSnXG0QY2/tIsTODKZRU+dQNnuUxEuY86e1ZQcwaPI42z8v
50mXuXe1CXebPdwVQOpa/UI9/LpUTFWcP1Ck0pQsdV9xnwQ1HwWEAIX8mmzK/7z4U6e6LTsMLqzs
Yrapbc2eZkH/KDc3dClHN/mx+6KWl5PvfGW0YIF2/DMuEc4l9HYjhehwIQwLh+X0fxMauqDcXAC7
nMCJBd9ylVEARCjz+znh8s8g24OVpwVz4ySxct3PPYBGp1IUoTfbQP7z76p6fepQhP7COJF190Tk
LS5Flj9bPm4dLQbei538rP8zEIrngoAxXPpWwyC4T0hNE1waaZXebaen1jzFAXqQDzKRtk05oWrh
/MZCbdJLVt+NTUq6J9tp3sHLP3HnjLyOnq8LfPyWj/vKcXJgUGI/9nsOOoVpRDXCADEnsG2dGa4n
r1t5tlhUoFX1WHAsjxxcnBAjrAQMiwwAiUwVhymbtXzwMnjyKH1/yoZsDb08IL7wksafOkCMLswq
Og0vV654wxkd5Vgnd0mt+YkhXvTnoTZumPBycKAgL+Ob29zHI/kOHqEVO0roV9wrxt3oOEWWjuPb
mfi3OIlr6UljJwcpvBmDHlFSQ6SeUS3BFLEi8BCJ60tdihEGsWRmuEsYa3nS8MGgk366ZGcH/TOF
XSKnok+/SdoMQcyNZyh2OFd7oc3FNCxvVOVyS7P7ggUgwT1OCMjeWhduPpaYsK2LCWKiQXIgV6q1
pqf52OiYwgLeVY8I1/o10nE6HhIFHysKUxFUW+0V4va/kwQthoSLWsx3I351zraavfWilzydLFfK
HB/1R+PEzsbYSC6VaWgM2qTDoyuGqKxEb5BK8biXYjrednOIRxWthDd0vLoULNM9hWbgqrq6lNom
JSCNFpoQ6SHatYzuWWO8Km9YeNhkrkTqZR5te31iWkgVINLKPpFTWJUb4dvG1W3QYz5nx6mF/TwX
nwF0VtucVLmkY6XBY2BAh2eCibPHutv8wEYEURYnTCrtlqpmdUwO/BN8Z8p6FIv6WyiJyNsu/bHZ
wBCy4G5hHGIqXD9del26EyYtMenncBrGjx2p5Pp58mwZQaMR4CduAnAQJdORaNfWKrAzgRLRaAaD
9eGjXo2FHTyeh93DthC43WZrr4rvWbj9qgXxJ9rej89/x0p6b3W5iooPZMyImgv3FdFUOKtU/JVh
ypIeeGRfQG+Sf+uEJuGBtd9M+1gYV2OMOfnhoENIJtSq1LWdMgcVTDQnh0dsNT7GDllsYK7kzAE0
UHYXFcbDJ8u9AEjnKRZqYEHbLH1mhHbQpfHDo9j+SiBhCtJ37zawdVP+jYg7SkWywOomwKk3J8ru
zOhMmLuwPahG7DasZYKul5KuP5VXEm7PSW79bLuRa1So6rkOCDeala+66PapdXCmY/JDh1evokzG
55Y99DhUKbb1B6FZQhfAIqUjbSc9NELfW/Kn3QsNGVkC5d2XOWaBYK8/2wi0jHwY/F9KugNYrZZi
YTzVXmscs8zBAlk4yL01bULIH0ryXckSrW1ovov9XAZUoCsxMjnatg1QzYe8s98xl1BS2AyLuhmT
vd6boeqpKQJs8OrYEDLDzvYLGg6oDwKJU4SamOyAXxgwtSBL5mrE5Gh+AX1Fbbtb3TRutOiRX92p
ySVtsxMwB20HGTIrs+4O8JNs9AqIdQ+fxneYjvRPvIKWsL1RmTAyOuPSymAhO/hCP0435Js1DC68
Ljv7ALUQNC7qNOy3Hu7BWLBf7c0LHhf+6Rab5vSorIFVyOGaFzs6i+JJm96V4VHoxq2V9Hojon9n
r6ofqZfipLhquK4on0eUS8s6yCXz2rtKmOtNfyJsAMlH3mKlTrJM3lRZTD5KYVtQyrL/XiN6sPRb
5KT1yFbB2wCdOJYfG/AJ+LNdiYjsi56NPDQVgejAxoU0FlVqgR8yCwfj6YZTbIeIaI3iF9ojSYC6
7Uw7Ue8vfpAccUnbgDUVp+cxFZ7yyfU7MJsMXrM2+6mE0vT54e4IzUWpWoFBmGeU3fpiZh12jPJu
Y66KZhIgvyuD1Na6/G/QVHk/f6oCzMLWYDr/gJmKlNeQWuuUGR66L20PMMjL67wn/IPRo/i3yRbB
79oaRd6AbMaM8kTI7zPKUT/dOKouE7Cter1J762NordXfVND58r+LyWDnvQrHgzWXt34ewbZ0ulM
M8NZpOXgUse/N5rBdADcWyWuAfHdF3l2wFLLrfLzYYao5ChoGgvd5uGZSNGlRfVJZWHojVdNrFEA
6B+hMqLh65+H/xioNdK+Ax/K2XmiCPuVzKwO0QXySJwzxAjU41SRsidbFmlQ8ovtbp07d/jJKIWp
Wci0YUS4aEs3Zlo/RBWWNaysEWLWBAoZoGkVNSOfFaHGoSCpfj9tFmyghvPwtg0MQ8tusPT1A9fH
gvNW7/vSbnabTs9Xoc//9ueNdC5t1PuGEw2L0Dhn+BqcKpDi3qyFUFSDy+1ApH7MaSbuXfj/5Xmw
rS7MVIoW1anZSaMbNbxSOxtwVof9yd9ohgIghvH81L1sOicYPsCW8SqMs6SuLLjaNLdhHaHoFq3R
nbpQqG8kTQNMwsDJ9CTvLa4BJQ/+U/1SMY8FQNW7oO6myX6mhFDR+P9P+MXyhgMdWo6gPbUhzeEn
+J4+Rfi1fXIbYLniSIvI2xjDbMjQ/K7DIhNkBOHWzCBxGaC6Q4Z/7SaLiKjT207ArIyQby1/Spp3
TSxLMLB1i8XSks4irKyOEjloe8SSEHNIfVL1Bq5zgxi+VVshlx4+9xDOPk6I4kcZkNuOD9ODilXm
mIgpD6xxYIjndd2KYQZmAhO1hekanQFGyHXewvGI6gasjVweJkAQ8RgtGTdQdXuURYrJv2vYMp6b
Mx2gIFm/nbB6nOFacIsN81xDWyrIztDGrM8TzDNWUQvOtWEqcbs9C1ljn5+S1MfZrX0NvMSjs7HQ
SCCseOhFvUd9tY0ohBRm5+TloTfTDxvffIxO1pYpC4+v3OAeCSUWM8ryCWmvCBYkgkSSD/NHQ4Ej
/IYDZDm1mH2jEAiWFyOEcQlxzzx0W8ycawTfzPg7tQ8Y238kGT0VlPe8T9gUtydap6Cf1R0+UsI2
JLsXw97ne2oniDKVTMOm8wo5zyPTGmmQ7cLi8QD7M+2RuPVf6x1bOgfEBe5STKjCM2e9yfxMH++0
CPJCspDUtJgZNkX4tuR67WzTZpyCwS+eG5xIWlfW2QqvqoznRYawNqoYjzqNxejZWwvtMKhXLoIR
dD/rdekm7iCMuJNW+F443egnuBNqwQvVTZgiJB93AskApS3CgWuh0bYWfuiU5KpLaxVz5If/09WI
XVWUJDIUKA+JaUyxFjUwT74FLTUy2KD33pY5F9YgGJWeiXiB3IRzcFlgmcHHrFwpmWhPl65dL2Qn
5dFTub8g5YeJuBUcmWexKA5VIkbT0nXLBz985Ab0E1vQn2GE3zBEUxTSFhWyMShiOGPUVVwCQ7Uu
x+2vd29wl+XhHh2BdXkMedUGOmitF+D2RGAS2Y2BJz4n0zRDmLKPQBPiHq+m4Fa6/AFrCdkr+UDF
Nxm6axAB5T68yYsg3Zly5tA35FnPVmdnWeS7m0BPdV5c7sgaM7YjsAwTpphn+CJWV3BSY8EGM+GE
XkMqWPNayTuYtuSMQx+9hk2Al6q4jrOu93u7RvVm++QIINQe4Ni6mUg2HdaQlOE1nC6DPXk+x0cf
ueJKmFmfVjv6hy++14OUVpWWEyA0zvggmL+hz6vqJ5XbClZpe+df6w74LyeenC5CXS4h5HJo4gQs
ikJRnb1wCe0dqsy8Pj5kkLqybI+XEqQDrzFFYY/f8dqyZrXcpC1U2W2AwOtXmEuAZhgpiw08s50D
zOMdSPE/IyVph0OAUQGqCGhhizfmDIJWasmzL92huGuXHlFEu0a2o8nW/AXGv1LqNlo1ORwk/YX8
9/X5zrye9OnCbKYzMnR+pSMwirkDG1yHO5mapOnSbjLtmitVCYDCjUrVtnJX1eA8xhHLj751IJSv
E7nC21CU4wHB0bLYJveos+8+/Z7XmvBAbURZTL/JWR/ugFEz61WXtJ7hi8p1hXymlXv2OQoI4lxS
PNrVBdwSy7elMr5L3kaJJiY0qm8k/qG0a7UQ2AXjJiV0lCSoTqu+HErUKtsi9zzmxUG6mYKZhZXF
Wk3/m9t3LGjZZBvtjn0MEBjGc7+RSEGfDFl4Jd4QRyGnJfDZ/w79RpQUHegRwA09N53+E4ugV5fK
FsD6n1yaMDzzjcTiSnEKqojepvFDL3cwD64Im/NYBXkX0PXt9ULX2qdL9prbTmZN69TwGCEeDufT
FDtOZDoDtQYEkB5vzsjDoR71nHnNpgqtmpw64XJBWkRoIwYaqWIY+bmqfe4rBQwZZwmoTcNOPP3e
G/NrdFsrPvk6vJah/hDKu/bOMV2hGLV/o1c3PqMtyJ3lYeMPxbOFXCgKU5UcQ8OwyHPeTYbqcXEg
67YC8NvnsfLHoNxlWxwf3/zvR1s6Yd51rmMLN8Kxgm/twrzgyMuOko8xZJ8+LdeCGecg86iqhU2V
EaSex5kpponw2y8cT7yEZ6Gbs3tJeR21t7pccQ/TxeS64KCHIhcXI4XpST15uFpFGYR8DwRIp0gK
iHJsfnFyvUIw/WHj7vPczytOoaf1DrI+k1d8H/a1FZj2j4MYn3gl30GXtPqbN3HgtDmm10AtGhuO
Z88CGAh1wggG5U9NpzPbsn3BdgDIw07qPR5FJzcR9TBmsVqONK86XdDHbL3uNcxNXkqXD8vOmTcN
3Rdm4RD+abkBMhK1IncCjOhJQaMexwMDHIW4e3SObW1yVKL4ihIAUJjeZOIUpnEGqshsC5NdPRoe
EBfaP4C/ZW2YP8MrTBIVjxW8zxwrNsgDe+Fo64exDTUonXVl2CgivLa2rzcjXLT1lJy1t8cGeG3+
3ZMzgDlCcXDlDpa8njRCBdvc/vLQDqNs9IXdA9O2nrrdoHt3FLsCYjTMxkqt9+svOy1YtMaQ0Cb2
U8h7jc5gg+560lsbrIW8OkZJOMbc+ZnT4NCZdlxiJtPMX7DIrHaA6J2l8pNsdJW/b4rN8WSYY6yt
z6VveP0e8NXQ+RZYd/duPfPxadopK+ZlTWE98DSdJWV56gz6jtp442XnAWmCT3ax0Xdw4M4uIQHm
Og1q/1tnpCm+YQpiFp+i2AV6pbtN4j9FakJmPnoxJKlkNx5yXdZETMTN1CyBnbagwlqEFJLyQFrz
p7Dvn/L7me3sKjTE7E9l970P91eKDfEs5WDh0AyU73s3z+ry1mW6zwzGF8uVamFcDnqeLNBJX63Z
nN8gnOElnqxaMycYCUvMpowgvWcAH1xMrrNT7ztrY3xZMvYFdl/Y6bUuaex+3KOJh26mDyL1e300
oxLRw+e0W31DjxEomE4ZrJ4g+pTBoxOAmL1SY7FT5E9hzryp56gcToDQ6yhemH+AvkF/cHMUiQ8t
fhzybPU9eHoiwR2m7XsWh4WDsFOXIVUTHZ6b+W1O9Cs+81AH1XM7Z3vHdcEGrXPoocRRKm2CbQ0B
vjo7u8cJZnecDlMKSdoW0EO1fYtQl9wzawZRkd0HijIb4rgM8wBmKim/gqJi6fi+40aK/XUko7h0
lABsGzMj1dtJtxbN1fqmf2OStdYMo9EWeFnts/Dtymi2DgHYrdvoI6dBcAzFqK5EhldrCODoBfY5
KNcJn83xLrBxZIbo8I8sgrhxCME9c83ZyC9MgygWoSR64lxjwZRfly1ti6H1KxCBlP4v4nwfX1lM
1Go9p6wtdudcj7KHcZ9GVL1MAWOsJYfJD6CBBWF1khvJ9pL2WZZKoIsUgIP4PMgsIMl75e+yhwwB
MMI9MXTyQBQH996Yzx4V94Qrciud8CgKASL6fbs2rig45emZ7n1CaQ/FXuLHSkL8UVl6V6lRpE6b
k3Uosr9PAE3iqZS+72cgvSS8I+2/a/pQsbOXmjoSHnzDO4lGvelI30RkRUk7yK9jAnzprZovw7cp
7sRPlKrK9EDYRK47BtbjpC5eDuWewHnIvnOCcEGqyLfGogfMFiBtM8YFFm4IMTc/GGgRkfNF6PzW
4Bjee+24URzQTRB0khGN25QH1SojgqJTTtuAw5uqSaHFhzInF/i3MUq8OKhS/M9kQYNsMoboRoaB
HX3nX9cleomAlj+5wJRqEXr9NJ+PB2J4Uo7Y/kXdVErox7OGTaFgN9hYYOByB3wN5sKsylENsKX6
0yaLp8HVnRY9d+oQNrGicD5Z7COxO0fM87xgtFaQw8+sOyA5WL6aHwaBJxCBj8R/IGoT0TayL8kH
72dC3OXdk2/jzKkjiJcIsQjYIT6ubMRYWoL4V+ydmCycYFWqSq8tvmXyvXfYCtByhQtzVTujGHn2
AGP/T6Bx9yNwbkCSupICbcGl6ecD+hRYNS9MCjOXEoRrpFduO8r/+o6a8ms4FSggTY9EFP/y5q5A
/1AyTldlDUq9ATf04ZlYwThfiDWs4pj1b1Qnl0Az+uwclagvAJ4vJdV5jF0186dPCvusK5b/ZEao
BjgqAZLNh7P8phvppcV/mtVurFHyowhoBQlvWcDOgrsR4ruqMXI5XHLWdxcEb043FrzrTRLFh6De
cAeM2UvcD5vX9MsNiTqUvPwAtXZWL7SXSnuB3CdtAiVe8D/seDRDUAftzD6wCd8QFktQKCZwUBbF
m2RZieECvVD51WrUWxSu67Pe7H+vDfRacHPrknCoxebbrMJOg5Cr8FOo49Zx8OLLHtidEdWUV/zr
7EC5Hk9uNq2gYpMMTtHSwJY6N53nG+RFucUTUjYvhi7r/Y8M1HojA8JUW4mUB/nANR+sVtUgYW+o
yWvBUddG5k1RmO8LetwVOlnp7Aq7KW7sdWQXuTCyh/0BLWl+GwzwM/DFe7ti3J2a4Vwhfr6jdelI
LZNHzfSvKHMGRMBkJOvBOMRfki87L899dHEOMd4ci3J7KzkhspG9GlUM/EauY8gSh3lYmcDYNp2L
c5FxYXHNxlbLn0BFRqYTrZt4708jrje3X1Go6m/0orVtel/4F5Qk59PQ9BOwZLDWSoZz6AAgRW1T
KHI+hXmaDvSD8YyuhuXxnruh2wTJ+n2ceARILY50HRwcDQxxtM2pUNZmeDa/ddRSIH/RWXu2lelA
7aOfqpeXN9v4f5JhwpTDgYxBJWIt+ZtCaP7i0qsQMqrIsVwao0ZO0O0VeJRgoT4i33xjt+Zvn9ks
B9fbYtv2DY5e1DZnTkCjhU0AYldr4kWJCVgy8v8MfJqL4+As7D2gQ4pPHDvQHcR9NHQOWF4VETDu
u2guXeSnyVBicEsxoshyjtrezXIfzc0m17EWuoHFclbvwzCr2CWCPlKDKu0iu363Zu19t4y2URWe
8d1s/H0LkDP5VY7xOzNQwmppvQYWNNV2bjqxIrTpEW8276Pch3kP/UxcQJANK/ULCV2/37FGXjPs
So0aEHWPjFZTxJD3y/OTEmvF4AS56zDTUJYnU5h1xBrd5DLCK80L/wiRiPL1xzsNTTGHjN6iz7SF
0dNdY0onhV9I6UWYDdfLUEbOFNwzAJ+snV9DqVLzd4Nomwhz9cPEcRBZCN2iLvG0UwZzeQYXYREC
YloJCBsy5sXIBFWKxawptdVhJLxiDYnbr7nmncIQE0kfePiXtC00SGNUz+jFLfEUUC4oF12AWrmH
EZsYlchbP/QEUApA5323LyaKn4cdrDb3K3nEMDX94z0BDH0ZWUDf28OVD5dXYwbr4yPhUH+J4vbZ
Hkal3+2GlEHnx4dp9DBGQs4l43NDWYfqsWp/CNEDSHGwMIp3w/j8DaJBB3AAE1tEaBz63qqN+Awg
29rwtCl2yoxZfDvwUNOJcO/080qo/KOjGppKEQyxVg1gOKob6s83jEYF1C4GdeAmPeO+davugGef
cHeXrAtFf1MBeK7bOWDniNpjQJj2Oc9JdlO0QlyC1HZomLKeTIkGE/Xy1yRs41x7kmeT43lUoqH5
lCTT9/jfbnAT7TAwHn0kIblAz0iW7hSyk659F1aOfQmPezqL1XetbrLBvDP350AWMFmK4sn5h1W6
02K7NLjPmI2NuH7IAhdFZtQLOhKocDpq6OZf4BY1xd41EjlJLDS0PzpBG3ha4ImMGSSBejWiqspC
aCMYdt1vjHBxzzQSHjOFG+Nl0eB7imulC3MEkKoBhHLd2K9rasNfkGLUmrwang3x7nShTh+mEF+W
X7FTT10sD/+uxZrXAik4ZD23/eENR6A2rq7MqpOqIgTUggpi9SLYkRetcdcGHf6bmtE/9Ho0fuZm
bjuVs7Efw8Fp98XGrVehFVt7gG7ULMtoEyclMHRcs6Z8Q6V3WWbEu7XuAyhgVxlE3ImHQTEyN5j8
Z2pUboLAVLkjaljug5+nLDH8fJvXt1v9TMSpzX7IuCaqmJTWfMoEulgO80IGvVs0ue+GlM0wlnAk
/4dNscsZD4QMKR79geKSUTAyKEx+sRgwPbQk3C4DHB83yZiAmNPK0VEjfIHWU6a1Ye+SKoxlxgQB
B/LBtjc6PEIe06iMmj19If8Q+6GdaF0pjy3xv+6UG3AQXSvw9qlGEJxsRGzen/2T+r2ODoVq832U
I8icDw6KAEjBMEXP8NWtEYx2e13gOb1Stmep3OOD39t3lJOvdHSTNOk44cSXkytBvLzv9QTOpJwy
TNiSadPkrkIuAcPd+U+Weyc1qq6UDLm3ECfZqVhHMUJ+uQY+dACrng9r9pBcC0qLfIsUDYN29r09
umNFTRe9nDkRQHrCdJDHhdBYca6LgFj8BP/3iXvCC1lPuULKK/1PhlcA5tPeTI7BZPyF01w6Rski
FvLVszw2ncwnjojAZFvuqZyaQWwZYa7puapqeKfyZGd3zZlxVv2kLnnFCrmVUfJXXDaq1CaH9AE6
Zfjs71xoHLjsuaxCDiuRJNASDg/n3U+bkQ4oT6x4bgx8MIrXBTJroCn7Gi7tillcPnTdeFiQaJuS
cxJgyUke94Fk2C5fjQc27ppbIGOlwT+qisYMl7uQ0W1rmXBlb3IGMU+lvHLRU4Ahve+bVT4tTEjR
O2GqAaQw3UwNodD00jl57v089yX/efxvPElkSXB5xjwinkIOGEDj1KmHUYkHvg8Q96N6c2XOgK/i
SiM/cBecJNSEDZKp/r3cmDeQW7ck5LvX1+CHWITV0hMiYqFmVhGWttzvQarJgOOuM9i1vHPCWX6E
aXRWoEc1c/w7WuJUG0QenWzF9S7p9cibYxp2O8IiHBnlsWFMArF1Wf+gzFMSFnXxXqfy/54fMtCd
6SKranibtwOhLalbf/65IptII7R67EFJdvjRYum80EJA4YI7NJJiogZgsHWqoEzpV+onl+WouNXo
GUbVAdXII1kvUftGpwBz9LZxS+V6DCmnevT9bIAuAQq+pXfIX552n7XZcAhpfYw6BQnxTXXoCYh8
CmrBrjwcTXTxg9b/OcPCEq3qS7y5ZRncfc0slyvpNYSmg+MrRDYB3rEUizL4Sw9fWiot/AMKsqxC
QhS4apAwfNYl6raZq9cX1URZ/AXzJsIuSFx6FtRFBL7WhnR8IkpXFWyCQDgCZ6Vw6/g+l6PZPCDH
VJcR9G9fwtaXNDhQuIBqbWZrRCUZM1r7LNEfDEijKla6WJh7yVS027qrnEAavyykMAsOpPmZnKdU
ZPNkNX0Jic6ssPE47J/13k4XWEyG39PxXCUZ5eFZ5tWVkIsnhkfN/hrtMZ857+uX2+gpLHpBu69M
LJUPf5i3QG9uuahAN8SQORfjM9oKZghaVyhn8xh2b7Zcr76GvY5iYNIhn80Igmi8bgkDrMiHawzJ
L7bryYy24PjAPMGSK8n+f429D58+lMNSMi/VtPzqiVc72GZvEGGGxUsHZt4pYYrQR0mwEPf6sqgT
B850p/m4aq7ZyzODZGLqX6TxJ2lnKAV5NJIPS4Y6rkxjfE2nCgTFBnMBGL4pQ1HpgbCVy3IFGRFx
c2NchCipq4b5Mes1asRvttKTqFT3ZyJuG2svL4iIo39XK+ASbRF5wMOJCQAPU8eRyONfKAovnYK/
uKwwTFoNeRabj/uKFxeduxhcB1D976EVN5Dkm07zNdCAHvvPDlLe1tli+mq6gsxSFes8B7LfO7Ki
cv1dYW3WZt9uPPLuSxKoOmgA0TTKy5ptk+b7JYcDN2SP0WjMZtm3OnP3ClgAk4XMJzXNBDcBturN
tSY5mB6PKJXtxbv76lCcOz1NxxdQFA0mqB3gp7ORa5UHtm2f41lJ6/EgvHJMByKgfqNQW0QI3xrc
JrM19ojqfb/XoAzlXziWtFKmmv957b0WJxAP92nfKvpNEWoetwUygoLRDphUYozOgVfNtN960yTk
WrKdd5igHV9AAv/nWP7Nhlj265sVhn9yvGjbB2uW0JqML+AHGHQBtan5YvvIsu/cuUK/pW9MNfAP
9bzxNK7aqCGQrwt0x35VZraRQovCgQl9Jlz0p7H1M5K0TW3KeTIxyKRtFIIYwCK59HOPeUIj/ztF
pySoj57w8vou8bNUyupkILEEr6Weh8qkUenSra+3PK1dxnM8LebvzXNekJCYDaU4gFrgNMBQj9l4
Wz901vR7mwoCDZ7Z1KRyqgPh6xtfohphsWHzoHHAxRmGl57eDrjifnmDiOq/eZ7b46ncqBKsRtyA
m0wqA8rAq5lXo3UgcsyvKPGgWDMUy9s7DTUAgsZtocVDwQtLPd2y6L1Dqe9G0wCzhFZQUQ/ixgF8
wFy1HdbyQ2BbMa/gS7MeL+7d8kfcmUbtYXWFkFHq/tBMfL3S6VslW5/jTcK6pwUJmxRIlgXRPH+O
Qx4VnV/4Fj7rkhuTMz0y3W1kQscxZgWuJLN2hMJeGDUlZr1KF1Oe76CeuNoOY23UQF0ZDg8mGxb+
/oG2usD10bLuHiRTgoJVq8q4qB0oLWiU5zZZ1I188DC2dk4DvZXSPui4oWCIKRfgPJdB5wR+YxHL
a5WHQvyHaCrLoDc4hrEP8bMsCb+kGx9eXOgroGJK26HAnS8TFWAnySc2IpavBoKxNOub6A/PPbsf
RZpgKiZ7Y0x8GbWLZRIPUp5r3xXAc9UXtFH5uq6l9kJ69mOlgccEPLySo7AA0JIISV9zcYgRutJi
TsgcZH0suIGxW9TJ1knw4svOfI3Uc4gNJzseRECHDzwI960QnCEEEMRd7MMRtZ+zIYinCb1xhd7T
RSNSFiChTk1cJlyxW5AN9ouNCNZmQi1lSn9Ysd6f3jxdQW2ePbfJKtJQIsLQIY2/7yIR6cFcB3/w
RsOBSliyhKTmvJgDU96F8v70FoETL+8Le/n9vnPw8b19hS+tSFAzR2H+PWLQur30nX7WhjP7BR1l
6YiyUMOFLrgvWhf7rdwhugi+sUZitnjg/2cTNDkuzta9+KaBQcJg2PsJmvN/iRZBGqYqU9OFSQOO
+e5ucqU44Ejjw8soNubJJVcLeOQpfgq8r0vA3HV/2mOMzFTURYBcxi0kRH8ljaA8MPyIgMAui9SD
WB7Ep86UfoGsmucN22vHBzuh6L+inOp6ZR1Mx17E8w27tB1VgTCPvLv1czL9ZdAfJAHvLhmqRyju
11OZdDp8es2FATpUuBdGufI61ddELWlj8OIQCmoLT/d57TFjq41pfXfzwJJv9fkAF8RWOlbUIfvU
K4S0cIrCYsZXcdTSdEyJ+Bs+xXFLoRFI5BCbkVA9i8yCfY2rHE63f9PWaBOAc4G1W8dJtjUxojWH
pdsBaj+3dd1HsBcY3FYKFthAbzoUKNITf3AMs5Zc9OnB89qGI8A9xQUm577U+axFKWl/MJoDMhjW
vysD8b4HQUlrKkGCYENDoPO8NdqFYOiaTwXTp5vSmoXA9JnJlM7sxPVcNa7dE36dAWYeG3+UV2Fw
YGzCW2yx/nBrZt3Pp2X9xBF+FtrfiKZ2St+UYPLtJscHmI2qIKHkN+251VuRutjQr17yI13rO0Nx
S0cz70SOm8U/aazgfFll6FLoICsgl7PFl+5UfDeeWA7ojUoW96oShNYXVG8MI1UbhRSN7ucI33mA
EnAqoxrm8BTEn86bX/fLW/vZ1Ahu9XxsWqRGKzmVxHNAaQ749CdbFtIYFI2nQ0WUeRYYfznH299z
++ytDhfZvuhMeYrnf4faCD1zarMvT7yW4woO9R+vHX3wvt7Odq3Uqk9K1dKF7frbIIvIaSpO28Vn
HEaeRTesI85eE+oFMl9bdFd4FUWQ8QQA8NGf1WG0BabxzT8Q95Ys0ZQLkaPleDNXtYZX3mPVjR6b
x4gnEC+7eiSx46hiMDfbvCJGMmkeZAI42DM9wlSqyxCAnCTeMXkhlBraubsyjbeS9y2zxgNPxDwl
PeL4C+cW+1tdPFcJJ1upsnunHjfKe8PNUU4R8IsN9dSyfRJ8+hd+oCOvC2c5a5cJTox/WdPkmOZm
Rn4tRwBD7cPsRzsQecAYJJPFUc+eo+netEDy4PwzCVJk6+Mo0uTIilkGSZUpqUPPFvbGj89Hbt3w
22fjaBO4E/Z1ehmRG9wZb7qwNVcJUXrt9u/NiF0xZoGDBdnzZCotR1O9VGk6ibkfJaQTqsidHXgm
DIcph4lDrOanYK+I34a+ZyAFm99eDnJb1oVGC9KOFbIC2qq5Q9TJU6EkXPhsiYYVGCShWwMZV7h5
kXuRNUKnfmSUUQ8DxMmGr8zeOAHqC4nP5ur5TDYbvl/uWfgkL4f0hbEEmiab45eOtfBmgfCECcWh
Ic/CQvVOGaQKOCWJC+SkC5ncUDuAQIHj/b3k7rpVy0EKnzWt/7STfKM9RlLLrojt4pFimq7TT3ZX
fMx6EWeT0qAA7jCsx0naxQoMAzpUvIhonjHAZHRSJZxOj14iV2kqqQ2F9H/2dgM30+/4x40HNnxB
yoNT0uR7zxmE1161pIWl2hb+3JFTMiEJlnIvucGw2g9MXIPl6QMVZktCtLPCEoYg4rNYbTKuBLzQ
1fikQ0iKGCKkS3XvdJQVcN/69hewB3vVCkgPTiAYrn+x4hCSjXM6FFlDFJYrF3+HurpRQMuN1pCx
XcMLp3wdETdq1zX5ORPRwCfs7eMQgMQIi6JM/0EuqmjdjyWamcEy4cDXJHOOBnwS527Q1H+Uhwpf
rXGo4NLQehtWGhSAGU1e0afZTc93WEz3C+X9Us22Ee5BtUkIw7HKnYwLqCETULG+OW2+CSpHjPc1
szUTWgr4vBkHkna3nA6oNhSzQAozMjVW9TWaA1hlZ/on/Y2FxW/tEyGSltpdHFUU21upmR1kzTKO
3eEu7GxFiDtDYR0NJmgtq0ZDIFkLNPcBk/uvWxzLkvCl2ryfHdLdrVJcGZu3MKSUe/kqxCCs6V5b
kaAwEANCq0DN1LE+Gy7C5DmodNn3/Yb8elM2Rr85KufMDdIpbB5JknMI7cj8dry1Jcxq4qSoi6j1
FJ3ijzjsnpQr7ho7htIlAMSJRav8i9QbQlm8cgYa3ap+Njdsp9T/0MK54As5mUJthi1jZ9TIKRD+
8C6VS8wW4wGQA4iWswlpj5akHn9Cb076XJ5xFb/1qYXRl8kFDrMRCQjHwtnxorDnWHuq6hjrFTh6
YKFkiZFGZJdVAxW0iu0C8kdjXnuDPczJ+gz5YeL905qLVJGG7a3qo09zYWJYw3t8gsFlw248O1nh
opfuBH7WJuf+jSyCY4S9owp0geSWSM1eUhcjauIDeXpdQJNfvHB5xR5SGCoj/ifoRwqRsZjE7Mxj
vgxsFQZh+V3oAxNqHRfDvWQVwGAhVOYYZBOpjJRDlIs/OExpClAj1C+2RprIcKqztoMd9K6KSgAE
pWf8TDXgaMZ0wM/uRETM9/DbOGJcSNzHRnsJhz+hUu9xerPlAWJ7FXVYsp7MOsPYdyqfdrdj0BHL
+bPeuen7mK9yG3ZLrnG0W4cTFS5N2eBGFLwGG9effGMNiDWw0+Vv4+OFfb3e5iN5KOHRf/4V7BgK
oV5ZpuCBPRFTxGO7rx5kmRTBpMzWPt4/ovwJC25uwqo9iHCoJ1FvwOi0N7x1K2+DWbX1i2j4T7L+
4Ctg8UGqeB8LWKpMDh7dJIzYP/OLH2b5J6h9KSzZS+HT2GifcHEkIridxyegzQ9I5LoDsAKQxJ3T
eKp5OAeIMIwg2uLubc8x83EB3GAC8Q6tQ3tpPjGF/NLIYaIHVvIT7X9XnK3er49qUCmF9BLg7256
mJHxt78aRYos60jN04nUeqAp7kZ07xFKrTZdFE6VTnwJMZQtbQ6eHjNKrCwSslewEfEwqToNXf1D
2ybphuP2PfSX9/b9NaoGwmRD40xDhvGA7qm1j+x27DIOBFL3wGkLLcJUE836Nsyp38OY2qj/bW6W
9RQ5EOgU6v87fxlCbd0n9Cip787hqG6ERTatcT9cdxBCcCKFNFu8lG4RN1LG54PK1fxaAyoQWfxE
8j1BMmjOZDRcgYjUkpKD+1x5L5f5vEin+QPQPncyU1NBJJrrAJI58qayaVw+jvfS8mwodZmT0v4H
3gGsPseK15KbBGfRNSw2lJ8xzG6jmFRToXYtBfERg6rBAX/yuhARSLIBJy1JB0ULJnllZ4wRzR53
i1bqhIb5nzCyY/yp0qhReSOQ2r4BZ0tiom187Q0ZE9MgbFYth3m8FC9lTErffPMt18TecBQ7Xy2q
82N6Zojk8WGBAUrUpEBnsiXOSxDwm72/5mluM/3UYMwAnwSLftBL4ORG5wzto8vy6XkX7asOfBXA
nQC5wUYFrCB4P685pXpniBur8iKtUiqND913ghjFJDxcJOzCdXqwdRVwJBpIR2ZCju2X4mnmH38G
WN1pwjVFYkfkCY0oM3qcGJW3YySKowO7LlHcAy4y7ifz2/KSBdhnK8qJHbH8FWp3G2zx+xBiJfjK
QHA2srUsZSUYo4Le3TAVD9jXz+V2RG4Njf+wyiU1H7FhaYIHJyJbaX597rmrOzsHK8veu1+kk6zN
cglOJFN+Ol9waGLcZZi6BcoTUoufOQON/hZtBzYTZt5x8YB6UqLcphuoKTCgQen2y5ok7FyKkg/Q
R0xeu86vH90CkgYWwYoY43hcnZ0zr/ZKDv17i7ZI5dH1dG+uALnFSSjKt9hf+QlaXh5I+ihuENfE
LBrgKcLELIUKna4/CwgDAb2CV/zbHFe92puWBqOGEjq/iA9/sXS4zObaLGw9Wg0/ocM2auXf7IYU
aBzXQsCrH729FSo7CJDoQJnPFKIoAgR9k0tkPZaF6XWnnakpOm2w5ikK6jsGvRqpifEQzZpGaWqf
OIWtd4MZcy/FjejK8YPVL513ZRMwRUMG/Sf+1dWwOed92gcmoAuZJ46rJufyWetupo8Wy/2FnGvJ
H0jtL+M0GZHqklFIWtZS8h5eksolwNXb7ggwVXNeZRmeOghoRKINUb4Hg/A4voKezmvoyns4npxF
zlOy13M3yHVuYNTGdIPjTX7+sECbTGS8jimaFIZBUIpXa7FKhxUA8rXoFbB7RQiko1hdZfjSYN7N
0yugSikTwhWbIMg0lUVXy3QuL9Mmm5dp6fMOkMVXXJtIakpsBMQEyUu1ujcCxHIS7gtbEY/4to/w
ArdzKTWSzj8oi3PufHEOqaOkd7k7rotxqhoESevFLg3XszveasiC42FL2pKPXZdE1Q+6Ktu0IfS4
xFS6OpnY6GOnM1Nn+LYzfbkcfqvhkDqrAroyYkDCb5AG1d5ff5aSAyS3ZMPj1r9pR2aZs/52wdiQ
a3K/ooaSSRDMLUzJ6Hn/XLOel0Lib9qUeYAQ142jAuQujtDMyxTL6Dgn74sD0Qb4qveYeS9vMSK5
PUhR7mUyRncGf2LLKcbIe5mMNcosOuPosF+97FlzXS1mtgVnuXaUUS6AmD/+Z8jOC1ELMRolYdf6
fZZTkV35nuYWMZJ8wur7DpIH2PYVioJTrP4xqKftzU3dRQHBT7tfQMtNK7+FMIEEWvxwP9QXqX7a
XX6yU7aX5U4J3zMunWPaJ3W4hDi7BIC1YN+XQnGiEAcowJgfn1NmOTRPZxGPUavPtVK5+pnBG9fk
Y2HXgA+NVmsBbVY0cvYSKxrEafohO9NinV7o+YumvvV9DaxH9H2l/0DL4Gc3V0f3e7yYmgvy1FQN
kSo5S0yeRFhIlzDhlzvYGsBbGAcTYV8RIpNQbVz7ECHEzK5CD5hYya9dImGdBYKzxPclyF5NQqe7
/pbjSZCVdIAkOYNGtxlTjJUdubjz3fvI3CAEv0hW2JJ3YBHqAgEwtjMdzCsUs7LU5lJqkvQnC493
p+LStV4k6WUTg8ct9JX39R1eNwLRKwicr78ZnvwSgQCZRRKUCIidWVaQmM7ywLEufGZgLtweirro
/Oj90zEt6gm6R8HvF5MTY/COLikofK9nZ4vvijsX8mIcJonLjbdNntVYwTFnmz9r+fXOP7PUryfW
VlZnC6LVZHYiDJNj8r0dpVtz8+b6kWwqiiu5q6+w22wAgelJOLXQniSfBMR+TpBbuo2W+zaUwi5T
Ros5E45T1CpkjbqYF0DL4MJkEOhYSgFJiBBC32afi5ofV0j0Iv18qNjiJJjuUrnOdwMbozn5krUD
Hm4jO/OR3a+mgvIq49IPMoPhO0Z0tBjs7uxLZVa2tQDUlXYdc6tKzjO8xny3sQCpV7+VKIheoD1C
2OIlYDpXbnTalu4yxFtAoNg7uxXqPTUcuW0QUjIurx/0Y7o5Q6nzmIItl/kVSjky1G1+BeLB3ts2
zfBgCLjnHIiWcS3Tr3v05DK9Lxpo56Ldh7pdXdzTDESP9QPMjVafCfTNfLoJaEkfhIB2oHs6p+N0
Gh0R/LaB01UHXyBs+NtOCT+cE6P6WW27ReFAGlEGwH2nv20YaLast5Uu1vCpRzTyvNdxdaI5nuuu
lbollD6l9clIAe7bnAIOMasGppUIKxiI1H5FzqMgmwSvbC/MRINt9ofWV+7Vb9auGwX8W2bomnzw
zoVi5tn/UehZRm9bGVlR7YiHG/ZGMwV69TJFUyL3ZOD9kPJHxHdMuvy0bsJ1B2RcHTgPuXomuB4b
VEtNUp2SSiDULO4vUX9h8R/GaDGchbDlkiVREAGrO2D9+eN71wyMrbddpaHTxs2UzWpbYxPGUEF4
cgalxyKzhmMvYMamTAZsJcIyPS79G1n05Y275QUbgvXOXzj+6EKPIl2ue6UeYPp4t/8Qu0+nTv3p
K4kdYhtqX/w8Ufv5I/la8CDuhww3cM15FsX/5SIzRBiLnFVltVS9tDUcZDMJpnjmK6pvopNSjbMm
IYn42k6iRR1H/XU3kmk2cihatf3z+i6jq30ZKmlIqb+iu1HByo7Aah8MTfq+Hy5vFxYZO5mNcpSd
nqEKp6M32nkpnepAUWAx6vyvbfknr1dES6Q0QXSHFfWZFGM3i5jlYJ7CVF2kCVuX7sU0O6W98gEr
6YVDJFzxV7ZP78VyhP2PNxnR7R57tg0iC205PXBh3NFC8S4A3tEzl5y3+XXywMprNHaAeUFoTNAM
X/jb2cw7K5h2vNR7hkymseKAagxNdfqBEr1p1aqV4MIgC50om3PiBcbmWYl2DljGRpVAWrZw7TTr
EGw4uHFhAF9wz+hUrCCasgYD4PUVVL9tHix8nJPLxIVOPFchcNony8aPTV2IEt8FLjHn+ZJelM8y
n6qCjwVgfjzxzKn9Rnb3IyRCr905jnczESr4uByUFP422DC/tJmAzRv8S83vgebQBGJorA52+6oR
XvtYoEB8ZNun5cO2NX71+tWm6W9w94WqmZ7uyLfSLwXUAVsAJUIsj3StyAy44MhLrWWlUKh0Xi91
psEyC9E4TQDXfTq/TIO/Uk3l05YU/yetr1nqMkpFC/jMOrSl5o1uy/AcwAoJ/2959LxLK+2rzCLN
2ljrrgKoMOSVp1igeiYnOpCCI5dMXmZDW0pbYWZArHx+k4TUa+buhRHnm53yBxtuLAv6b5uO+qg2
fRyv9oG6mwUSOUR5ssSbIVUSGjpK1j8vg6D0d3qdUL6+2NVbtyAIsuru9EWoDft/u4PuQChqDBLx
0SKkHLsH/jsVUVz+pYDlkx1L93bLGlqc4FIzdNxQuVsH9flSSNJec1jhZ74XbWw5SO8RQnMdvMlZ
6xz6nrT9H3swlSeKd9OhPxB2ubdn0PZufu0dYJMzQgUwz9w4W72wv74CYMAMtoxJfGHzlaPG3UWc
H+UDbDjhzyZNys4tuMUbDutUETboOKCc59pEt+g3H3kjMjepkwz7X1O8jRfvwrSkSTndjHsDJtwW
0TQQlih1aawl6LR4sWeu8ujs9CI6BtNa1mS5SCbHyPH9tM6AZHRhClq6/qzTzTDGxAO4X9ZBKRnE
xI8nhQAQfFboi46G/KnYhOyFwmKULcpdhShDC5j2rzr7+mK340gZsdSGe+MtCDdZOBegF6j8N+Od
SQz/BbrqWIHEm5pq7qP/uHxOr55VVEngmdoEiB0+z7khEiWFOJoYW178i6kYACCv+IdHXfjZPS7L
aJXZ6XSGeFSzfZm3KI81bLf/Iz2vV7BTH5pbf9IH0QogaGHQtUVwZQAufZ1ufZm5SBiwp6bKdLLV
mTZbQ+jTf4mjXnnmpq2Ph6X0tATCRczd2g2eeR3m9LkZzAwmedJQnFwVTWZwfAdnxatfgHvQJBEn
MvPF8z2SQQTn1HiIIEAQVj77Lb50YUgNF1jx+v6Y2MV3Wpxw5t5hIxd/Fzq/nUGLOsUk4/dQj2Wp
tm3/FullMzfhDeAgjbegjWuDViJP9SM3lLURaxnlT4kvk+M/duSTIKnSFJLXDqz+6bJv333UtROd
ItLaIg8yxbWlJreb5PXWLl8kbnyQyAYuystGZ8PxN78XDrx8PlRtBSnfZi4lvTTRgV0QOuxbYTzg
1WWyC6ks1q0KzXdDGrWW7Bo4eIbNZTzXxDBdnTJCPuHrYpUH5xtkXSN+TO2t1EpnhItQH8eQq3dl
YVewzxfJumUQeCrg72u1I2LXx+PV5Z7JS0VukfNpVoVYq9y1Kdc8Mm6FUyP8ZtsUW6/cJdlwNr77
iXqy/w7FnUp/aot/uJOyLP4DGnHR4qw7rbs+YjTyXKHhVfbwBuPLyJNUboBN7pSNNnVABQXCsBVH
d1LsZPdrt7sB/YrY3WjyIhq+LS8WzpskdvkumNhwLJukIVCu3GtRrCjaKDutdITPjoYDEu3rww2t
Qr6hkiIF66i0qpKUDWJ/fDDexTiUM4HrrD4heJnqvB7CYrWvQdU7GtQ4JzyYkbtEV9g2H5RwjEvm
VfcpGnElMe5EPBekkvmxfgShNswjE7Tkzp4D7REMu2Q0alMkmYY8PjiExMS0/frJFVLcL/uubRFg
tia24UWdHLhRexfIfVwdDhcSNlLiLtAj0Bc5Rx06d3T6rdeCWXK9JzKbsPDuaMsnL6vcVXACl4/o
fU1tlque5VO0oWEQnStI0HQ3mcoeCO6rBMwnvK1i/cHCm0UQ0Wdn4RJKuwfleOV9TK24Y1PQzxwN
TyWZa3O/lRjO7XoduP31LlLx+TqgmeS7PggVkKW0L1uuDZV2zq0r5Ew1F25LEY0QJZfGrArupREX
Yj48wui6QR70ZgYXTOwKkQyR25G+QWGu45KgRqiVspn5RPEzkfru0lUL10zCy36O8dETFD7oLYQ2
CDlxZusLlNdRyAisOw6gZB1AC0oKPcjjgjKQjJX4S77mNbzhJSoZxWLQTA+bH82uf35FsCdd3zsm
/zbzNAz5xzE7W5tX+rzJzGDFwNCMYrVPOgWN5IFPu0STrBWgmb1SK1QmaGFGS0g/JXkFDlSSfN4G
JP2/9YksclNO8X5xMWxmPE5yp4V0pke5Waf5rYoBuzH7HInSpLhsbkzIiZgZeJ6wXMvP6qFVWt5F
M3ycOslAHtJ3MJ4BIc5tKcMBxgNbVzq+Qyt2xoWyHs2hTJ5t3e+zTNDP/A1xyi58i4DLpv+j0CkV
MXHFbzGP6RenjOpi3N/jEknhBiHqDEvBoZZWdC166d4eCqlAzaGa9mKByO7VnwfISolc5q6Vfppm
sM26h4XZviyhxu8/ntM1mJLgfGw+OJAnhOM21PEb0wzYAVLXzsP0mqj+oUqOQbRtu8zypDhgYTX5
ufOggxh29hPY0Hh6ex7ySCZ6jMlS6TwfFEsNLiTWCUA7jklc8V3UH4jk4Qm93B2/gRvFLJemEY1g
FRnqvEd6Q/kNyIp2UOxCJo15lLzq/4xnTcwLIuhNsNT42B6bZDGwv7A/9jR3dxDZSBZ6tqGHyeFD
geEK/ySWIgBBGAp88AYzf9fqyItn6S8kRB/uHFbKxqbFUxNN9vflFRu6GwjAqtiI4Cq7b4yLDsoW
A2xum8wJSujYU1hg4vjs9j6Uat6mpnwsbHNtiQ6qMgHl1ysg8B4EgKoqU8A0OopUeMAKzm/1+Xv1
F7kmE0VmqgWye8uKRzS8QqJyggvogSlK8sBZY1Wf93NOs4DFI5yX0/ICQxgOtE7DQFWvvmw1Nqeh
LJhbojttgyMC3Zp76ai8DNUzidHGicX1mYKLUo3B1C0mIRv0OEhzLkGDzc+1llY6wiaRA4w4DWzd
aP62WG+swSpKtrZaTMRpCA49ET4Hq72focwkDiqLDHvsPpKd1Y8SxBw2hxo+l0vGZEK32RRORbIQ
IB+u8i5oC4dZSwIrs/Oe95q6ew4X7c+R2/col1p9k/72sJKmroXIAZ146E791saSIJ2Ts/51NuMC
a4tf/LXgCUqdYNjD2LlpihA4Fl2jvRkH+Vt7uZXRAzkIadrYKD97Dxq6YKu9pwlbaRB1TPiQR+d/
uUXfd6VHlmYyBRjBS43oLJxYoI6TxFnUUrwWo1j6wHPiNbTVAPec3sFpzxKiVDA+Gqbm/tN4h0Kf
S1NBwUJfDSOe6RIPNSSyplbXBHLUCJY2X++sQ6y8Q8YR8kq2df+ztoln/T/TbLdIuD0dQW/UUTtD
PjMYKPIdDgcxaYBOPzfcUO7XJZVPCNFyQM7YW7R3txsvKp7lWrvQwY1Z+KTCSKe3rZWBemX8AgHe
rK9wFR/B9iO0jcLb+6/9L5bntTQU2j/EUFt0/rO6ePtzjTOCkXooN7eVa2/riQ71gZARS0enFHhy
EccbUqVtSNKFsFSim4p1sJDKjnlHiBRYKJSHQVfEDPBXEPXNob/iZH0dLPgp41eTfHeerEVFXPEt
q2ZHauK5njy//boxM8P6OUQNsAUqvk9TyqO94Y8+PyNj0o5ioLmGDsmD9HAwyOih+tV0TQSYIg9Z
ty/GM0aHGgbO0YbGSuO7g46ZNZ0/so2/aaYDNN/ryyyhLYWyf/VsdlxOKOWB1xAO7GOQfB07I9UA
rhcXIfLskp6SKJ4Wk/QaSRvgPuGYt6/QrmJC2/1IhZiSsZXouXb8QQto84lAxoOO01YX+v+zQEQU
ggjgJFcOkwyDa7EZWPMTW5YLJfwsE2Li4CnoZWYd45UWcxQKhvzowUW/J7FdWfGU4eDEz7z3VZlg
0Oeq5+pWXDuXUkqsQT2Yq8C+1SoI927SrShD1m+iwGIbWqegIeMJzjTpLV+RoPhBE1zJ3ZrfmPs+
mib6Xzrx34gOy+cVmulwnM1gqd1qMfYF9mmHqv2odLTD4r5j4rvGUottT30nQqpmlcxY24BhMbPY
UPXeUwjAoIsaUcQZmO8lbcs4fbaGznSt0+6U5lI+RzpsEaPYYsquppUSimXY/E/OyV+qfMAisolT
J/4aJy5hhB/88UWk9lnYz2XRuEu+DVQz5g+ObWiiA3iZAHISN7xg7sNDrTg7+o0Ayjvb1pS3uBW7
i/DMQSsP3ctNY/YIiLgTfRiMSY1As7qjhF8ELWpt2AVdNHYtGlXtl1WZb1KrTE57/1lsmT2IDEZY
YLFRzQxHe84S0XXRRbA6yjzJ5wcZaltqMnr+RkDZx6McO++6lc+sPqV8LelYNqLo/IlJvwXRB0rz
5AAjo0C27YE8Mp8jG7uC48uvNNGUbt3wgvCv3qZ9HB0yo3r8sIdwi5tPbJ9r277Oy+poCF7HE1I4
qXAMkYXBArkPWfHhIYmSP69XBpZjejzWVFtcoqUcGWQkoccT5lQ0ezxRir6ckWsZwgZqh72DrPVt
6guLBzuvMfkaVEsWkxU2n8FePylKI6YAFh1C3Jcdep+z1dnRKF6Yn87swM0wKS+em98EC7EVtpZF
+1CRGV3Ded8EIt55OsPOMJyWq7zc+7EPoBg2qRKINQHqNqRl5jlR6DRrWadBI0JdZ9c+Zyo36JtY
HpPIoPd9I9qKiXtETU3SpoOI7dAqVfQG0Gy81llVvWtlIJWhHxv2s3h5FBv5rzqDOHOBIPCONxgS
iSGk7r/FfXCNh7BQ3aVn/gT/PU0dMY05RjQDILjhIH9rYl7e3PGFS6bxaShLtu4N5ggOegTOmh0c
xdwwjyQmZ5VlF23vdk7emalVWBa4d8RCkA6Y1oVJb+GmxHoBCsoQgUHtP4YYA9VimelWEQyTup0t
qX187XMF4Nj43cv85ie2IqL9X964ou8OsrXyRKsrm26hdzcB3UzkPW2eCM2j0y/mKzEISPTiJZgZ
DTtite/bGif+BMNttsTj9R8uAgOEAn5w+b+bm14nc7WZc9Y0ZeeAeLcYWtl4Ro4cNv5Ub78Gr5P7
ip2GYRzekjPJQs1zIaVfayd/c4NrLsXq6IyOWhnbqa3XJPbDeOzaWB4V5T6GpHKcRXFQCicW7U3M
8a+KrxnZv05Jj6lsKNPS3P9a4F31AU3x1nE98mgXI+1aJnXI5Ro6iYL1c5aFobKYBcNDhQ2VH+n5
vGj0CVIKV+VsC0AXG0ApjzkNbGPIlgf6QKDvUCyQDbl84h/Y3w9Yeccy3Ncb4tTwmr2A8hTJRzRn
Wr+aNerrvCHcIWHfmrJPzmmHpgf8hRI4CI4v0fuGaQ3Mqnr34r4v6psO/Zm3XA/1/pzdv5vk12dM
+llydJR5DQ+bwKrA7yJYCX8XHz87O603HT475KMR2WYKL16oPxPSTeVFd9kT3jOs2ArkcQe95p3l
5I8PdRzz5mNCcbsh5CEEYiFoJWui2gygyleIjoWP205fcosD4PFfcXjo2EWMomUk7RMqoBqjDIQR
8gCfXXfpFNmCwNkXd0796t9dL8xI/EvgCkYoZ7XdysQJLAwVTN791TQxWVu/f3zr7OEJVIvQQsb9
SHx9C60lyrkcQwPwIW01gGp0rkj2gpDnnn0e9eQ4koTMAFv/R+idpnglHVlVvdqKfTxFW7Gcl8Ex
TLpr0qxnCZBXEjvLtC3D4ZvigEKIBtq8FTtHHva/u9fAi0P+Q5TsHCgvKoa0T381ES/XHvpTEnb7
Q05u8lCHqzux3wMbuglku86kKtwTmSH5KgGP9isgn30j9H9SlMmwkpW8muatAykkfZaRocf6hTfE
SYj0qbbi7W1N3wM9DBI2FuXc6xUYSVOhqfdIh0f8liQqARj2fuga80PB37iIScPZ9BTsJ2rRl2d4
l9YDV69YJvc/q79VG57SnwgFL7n9yntFajUhANG51/iTyt3pYKerK2jWivy0atQ80kDjh/Jl5mNG
PwATMhx1MnOyLTsQtcIqKtzBajJAjQoS4mAGGXZkvlFR8mZBorMwTQoKdf39faYHkTBcazu1U6mP
zhJ+hKdP2CL56+6aQ1+HJaib9+shI97Nf/qooQAtrnXtaPiDoSlJA8L4aCVltBqFi9uL94OzelvS
jHpQJvLMA0QPbucaBpseyjg7azxinqvIdKj37EESQjMIXJMNZmOS9pMj3dxjutXXSsZPJHrBxszf
uQ0GBMGkv3cjfjbC3GFTWQWrDdYtn/meJCk6dXsiCit9P29bowgQe1tfISi4Yiyw0WA2STuHOSro
1G/doRZThb0dX6uKMNML0TvR2b+Aga4F4vsu1qtUkhgX+RRmCXwgZBo7B5bu+u69b3QoCpNKl9EL
9ZDgGZ2TJUaX3EwvKPMJMNK2BAKdFbNvModDXXNx7QW1xwIUroQtGKloJpi2fWavWRhS3UkgqhJi
O+uWlSdnME0Y9aGVkEkgQsMVKcJXWzuuP7xmL5bekFTvnYc2q1FMbGNL/mGSyhKdXNq+9MLOeFjr
LIWYwmIXU8L21Aq1agBp3uaCaajkpOJv04+L1mknWX0LVDM+kcmssMLUK6B0j9brMQOGmYBqyeBQ
AbKxKaqHGIaF89fDtHdac/w5eGkL+LzTdjPSNZ9gBmEqACerMxUDiR9dvbLhFWnPYd6+Enpyjd0h
4PMx6KZUZLTnpKtuWPC+vlH0qx4fYeuhGMcjjvkXwpMSFP44P2UEu59Gn8W/EA534H2/vIW5nCAm
TPUFE1IKLcbNgSrJ2a8NaduQGC7QXC9/ZkmNb0hTNQ29STrxFBBdaISPAED3DkkhDVgBy3w+vMVw
gOlRV3VFdCAcDeAF5y7CIOKVAx6OIYXMyJ8aR9PqsRGmjZhqImKv8fXz4TzgT+LJx+9QUjhKpfUx
3zPoJlS8cU1OBA+EDNMFkZnfr4qjsJsZMeMsfFuwHnSOUggl63F4kODL7lV+hU2kJ4SsJQmMbPLZ
Zd47B9vqHMc7jpkPRRxn4WIqwvttgrk5vJqCU7vRh9jr73ZvZmB9BL8JU+qQfPvbyuDFGsAgwM22
vMYM2uOy2Ub+L5ArawJ10YIFDAgUSEtYiH6Vd65YBP7qDmKrCG6Qey0qoBvk3F4RnjzJLRifpoDM
VsSUxhyryro6zWX44sKYQpOJR3VHhv9a4HEvVSn8hIKPN66goLQNK/i4cDcys0nyWULMhaY8yFGn
k0SF7LdEza71um89ryU7tsSDJ9cx8TkRUzIX5thQxUN7pXzt9MjIC1ywOEKmUorRZ6luGCxTvjYe
ZclHI5R53xhlnJQofMCZfMkLDGKUuDFYbQQ1nfdwJmFhWxRK8hxVpDwNNxNMaG0/jbVulHepJete
gmYdoW65ofvw5/sRyBLJHDaH4RDm6dVtfwUurNk7m1q7y+85VT3wG3oghUv7s5/gKBPtOX9nNAw0
kqMMRujntnajvWx/RhnqNESqlyR/tyXs3NMGLe6cdIGaN2wgzUnnB24+5t++8kUWvbOFEnHtLm51
9dRXYrFS/QTXMgK/6m/FKzJtpMVR1mhyAgGfjo+gD2L+2qxgbRh+upI16mBpjFpn3jS6feaWq+mf
q3REGv5COFJb7o3K0PmKSvvpm6ekTFLYt9eFz/e4/0PBJhpW1Uud0bWhi1p17sCN6OBnMsMCa+w+
WMvTjrSWE8+OsOhua15/JlOPLsl3aiZ/Gb8O0Na7PAErL3LW+kSHictLWJVro2bZ62gDiDc8wZjQ
YENZhwbKcvn7vqO7isOOEV5Q6JbV4Samu12hiBk71VMC8MplciDG/4oSjTSVAuKIxe7yE8lU6foQ
/LZPbhhajSpNoapBntVLa9T77vkEECMZLtqVVFTRSR5eSycZl5Og8xLHJejdYhVBRz0Xo9r8FNup
FlSH2MVx3EbcynSWNG7BXAx5RlqUfgtdDr4paaXDzVydPTKUMSG+IU2SQwt4UI48bHRPnxTaSZma
YLH5dzZF0ciFfSK8ki6UHquxCeWrjIK56de5jdtYmo+SKE8EjN4FN+D3LCoPF46zqZAI3KFSybN0
7DA8gdOp96bEwcKJ+By6RmaoreI2SADQxAp1RONaQ7LNqD65SBjZepHS8/NHHNH+lzaYHYktXC3p
zLzMm10TEI0FT8xXaSK5uGUt2EM2t9avM1MHF8AG46UKZEoNp4tbfCZ5ScIwbAKQ9qbX98ofrMZt
sX3muAAEpssHWihWExE6DgeeIB2peeZnaPl+erTcEtk1YCsqmHh6ZI4j0oKJX0HDUrrtaDfH0NUi
WeQ6slw4YIh9nD+GuAJtpM23mAiZAtkqWnnaW+fvqhtTxrOAMoFMOOHtAsw+w6BbOqLTmXtU8cvS
IHVtnn+sjj+yQzgvAmxf91ADrukwsSaDxLqO1sIxsNh9ugRg20N6m1x3GgxxUKSKmx4s93jQwdEJ
QHcBZLtnHkIvRgGfZAVU8BMlnrT1GyeAWwhxS9gxRJnbCBBXULNOlj1wCP1NwiCUWP/Bie5FRL6Q
QU5WeA70w3rraAEbm60diedel6mwrRHrsSMS7mUdzXHu8AyqBQm2QZbzUVWUp8WYKJoaiBfFnzS+
OJzdtjz25gg6bla6Oe/yPit+q/gbCYCKwUqUi3Yvt9IzMrxTP9axuEcKESiEDjIAql1S2B5OZdVn
6DTuWg22Bpqbi0kF31Y7XeqQX/QeGmbYmWYpjxI9vhcCtFzoSwt4M7WN0kbX/9ZaR3XmneFDcI+M
bWibXM7Gvdis9ciKrzn9fVg4LyIfgQ3VAnuOX4gyhUyBn30IgGz7B9bsHRU41xYGf32amY6/HiNX
zeI1k7MmT92ajgwkSlsVtgSeswnu7218v2AIunZfuK0mwDb7jzOQYNisYJeyoNCHIst/Ngmg+zWe
ui997dBTvGXDEoWNsiGqRDnpEtRfYwBcg3TDvZE9fgCIZYpZ9T86me4w2SCEIxvcpnakvUcG1tWo
rNimxMrA2xG8m7ZY0VsEyVbyXYpHJdnG0bmwoU70YB459d6ga5Slt6zQzn83fvrniKwnS8BTBIes
JHwJcx7hmwZ9OA7nm73VKLB57POBaBIgrsXJNehM6c1p63EGOy14IaMck6LkjLIWejS7cfc3RCgl
pKPfg2xK+0byyPHeHI4J8spdSCeTk5bsU79PSUfHaAYMa8HZ2YdRJVjF98puqJG69O3PqzV5L8D8
zdiiczAtPOjW6NqTrXVNf54UkJGaBzvq+em33B00gyVROoG/pAQt/0hCpY5FySPOTBcKRMfVdvMN
n2D/NRkgQPV5kUbaowHbwcWyzYWm9E2RHikNdj2pKlWlnMa4sRDdohZutMKa5CZNl1Wx/pjo1+rf
qy45wI+c5karpTuCmhs9wK7zlF2fzFcZcsxJmiuXQ/ok16o4qI4mnI7thF9CbjkMQUeC5Mr4jhdo
ky1oLWT6XPhvd7TVtjlOeLollss81Wy/W1eW2etcNbVwGU56qylHZbHsNu4tCwFCBDAlwe1Q6k+0
aku/3+g/oHKXz9AdxxY3d7eBxskuYJjSk0QEDIJyTLLE3iAy9G6aSRinCrXcCqkT/I9FcuaLrBHV
VvlGwNXKeV0fsuL1qMuin7bwdUVKt3GQxA15zkpYp0XTGhFum4qqW/Hlb1EdxhLwiYjGZ4PeTfeH
K4j98Bp/X5/o1w8lpu2V44QIlNxYVEugkh60dK+87Fp3pCsgZBgb+i5OXF3kx4Cy2hkIKiYonO71
gBEUQf1v/vZIy2rr2fhrIqLmDg18FcRika7SFZLPtuFGsa7NBkutJRtlHpWSHzeq2lFJ7LN62aIu
oU5mItReM0FE7GqTBoq0T7C9CVJAkPx34ds+7vfuq8aLM13C05YcAtvWA7vycS8GPXGN4LJDHwud
nipyJPUJI4kkEJkOpSdmbUgMkARrao9k1AdMckiK6VqEMDMc6cmvwYdfDLiz5xMwUKDOzQ+BDOVL
BHKiNwuTpX8V3isHOQm7IIfMyrNXQ7zI9aqFA5N4PCFR4Czipk+CPvITiQh7xTIBkn0e3wQWozjC
oXiCOsdet3Z1WO5NK1xFHBiI7hGTGr7tq4u6/pMiwm5arLO4OE06gDJrS+cZDDcwWKeGg8UMNRfD
bg8+ylwoB1maAWNO3ba/7/VrJ7CoVUzfYTs4S/6URj0QCKWHvQ8iNkTI4HlPkFa1UGq1eymoomrA
FTxKqOv0gGdTDWqlxK6rjnwVMXhwS49bFcrM9mE9C3SDrPazr1cyegpb2kkiv6nPxjzK7PldI6hf
KfcT8OCi7aUCkH/0ie6mA3nLvN9WfcM9DruMkZo+AqTt2zPqyMcY8Ij95Jg46o1n7xINiJzzOy8A
qvw5GR6zd78GBCeBiOJQ2dVp1rXYjSuc7sx55vr5neZRnTRmCxkwllXG1OHXhPJqYgB6w0r2aNA5
jDbEEoQJGPejqrGlrN+tbtvz1C58s/+vmiLaCVU+R0zK8/5QtSGVwAfViw9CzD/fiFz3dAwSB+ue
EmZJcqfz+d1Yokk15U9+JLQXPUrulnIAnu7iFJEMPu6bwDIiW49VnUWDyf8IEmr4Z0hOUIxOOMWa
zYEcdmwfqxMnYmuBuD+DaDbYpqgSZ3eIKOZZJsNKWsWnlRrzRuqQsVLPGHvsY5UINe3Tc0XIlJWM
tjWGv0MWHWK/huQpk36HXZkJ2mnbR7eJHKiQFN4IiLARo8bJUhpt5792t/kIsQ5yt76of6EfZXw3
2GBnmQ2BQC2d9pm1Katgw19G/H4uXvzK3KKVZJcJujo/fRzftNuYqNuR64ZQsJBiTDaVE1Jn55Xz
lkmCERQt8DrICFMbu7O+m1ETS+X1ZHJLTlT9PhXRPJrczmMatyVIICr6YJtCT6EfdicLbnEJbEYg
kn1rJW1Go4YPJeF6OI3uAQXVQj1Aop3VRBkDcpWmrJKR9JfO2vYGrBATqCqY7xdrNStJKqY6sRad
/kUc+3LXr3t1yrK32CE34hUfHfinBmbnQMRCOhdbLDWbw/vSn+cm4JLxBc2wuXutPfVbCEn76PGf
rJWtPXnKU3DNpIIl43FNPJedNCobDm7iSrafhjKTKtI95UO3qtk9tgyZuW42UavMgA2mOaONfpAu
SX5B3HskqLl0UgiF3zVV3RJ1cE/QW9dtibFTzFD9ctLd22/OLnQwXRpDjqT+rtMbiL8PZT2m9/Jv
Ev3eBwap3e9LAstEuyZD08RuM3ojQ5hLzWOd3mZ8MYJFZsP8wr+tiOX9kr/wwgNRqFAQgTmLuNNi
lxDUyEunzl5adGn+2KBqhGW6phVdpiXgL+kASHEc/6L+Fw1K7SLaz+B19k31GiXtwLsTsS/5Yq68
K4dtWDRZa5IVx/bOa66Fg15Ji099kaMj0PtonUyD+bYdCimKBeuk9l3L86iBiGHVXfFupwfsJVtV
XQxABhEQChNj8NMq7M2d7r4KK9mBNo3SFAJezF844yQkZu6zfFZDXHbtCmumLyCC/0NqSV0WQBrx
rvWSvVTgbnDtHqC8yRNsn/F9s5Uvhc9I4TgTuwwFVl0PlClMXEWv23JMH88g0mfZH4++yjllNPxq
tGGszH6ZfQXOdU+2yOj9OfGlon2wCAicjduQqI8ONJOq8x9FB6IKJLnIbfPiUo3EjUrfjCBKnjlz
SvCt/LuYddod4XUjr4OSFfkSGWuPBqn4MaL8KSlAK10fHIZAbVDKzboxlaepuo4UJQe9ds3AX/io
BuUpiArTQFZdQoaI9DjKIWRltNbS+GxeEg3BMNcCTOBocowb7Ibpa4DGKjjByFx12Ue4gBZ/vIlW
FDADQusbrJxXBV6B81Z2V9Lxj7XdkiV3MMoa2EM6oxH6N8i6hxzYXP4ge19FWvm4pEzHae4yElyA
+MDKVvpkO2olg3K/8oV82BlCtGYLJsxuL7epxvBnYYMsQei1GEFSyHWOMnRsN8+kra2EXq6e8J9Q
KD5/DyJARJ6++0b6xR6AtV4v2Gm/CGUul3qlWG1/8gwCGMrKFzluPEHsD+SzbsP/qdQLSlAP/Lil
wKAKlmN26kG0SD8qBAVUyQ+Tctqsrm1zAM42ZrphJGNGZiUseMR5PnfKjnTG/nlc8MQDjCH/czs4
rzkMRt1XYKiGY3Sg3IKIGzH6WyKS13ElUAWYVZywEvCtfa2V5ERe8qSOpaBrvz/grjqqxJd9DP9z
2ronsErp4dTSLBs9lbpz68VfPPP9tzKx/jtgfV7jSUt+RO4gJ6/eUH+k2B+V7N9ghZIGrhpldU7x
aP6ksnpJBl074Jx0+hXtlm3mnzTJQEvHArJ32V6mSSKBit0S/OYJp6LYyOzwVTdikVUkqnVarVzi
Yb19suHoIfeAytEhLA74r/NIhzqQ8VTR0o99a0r30j56a/iaepV3k72vLREiUjyGdzqk/IyRp/TN
AvJ67KTUqAAmXElKEZd1Kx12nBCTToSoEZHL0hLSMfq6JwlvibsBDIUN2s6YAUkXjVydAjm39S+O
C9WcZWyd5pDV3EVkFqMKzR0STpobO/ods81rPC0hyJE28VbFuF4yl2tv5FnHxcFfNmJtmsvII4Xz
UvgjK4LfSdzIo1zFBMsKZikRxoYKPIqOsX4oyJ6Bv6bn8X/YVJ3aaHnMkzwp05lxTL1mWwS0SGEa
KIODQlQiQKw0uFVD+zP0UIRouFyh6bhgtnXQcUMlh3vz3cbTfAESADu0u+6p93eTdHmqRlQ20ydA
soDEhEgsdNbnMmd86wPAFGyKXCs5waA/DK0N7vA2eV3DqaiSreYDbl5dCzL/fzRdz759Asi3nmT2
/zt8H2/fnzwHSmA6JQj7oabAv6bKHFaTCdkhDy5Cc02ItnStCwI5ZUhaLhfjZ68O9gcw5bUJfCFn
P8NP909y3ktfqq1zbmm4tQiuMUdEElbWZ4wm2k2TpfeCJ9J80ygW3sdKfxDM7oRaMjqzzctcA6hq
41bPpJTK1j+xDEsNIGGSHxUp9SpMNqO4frFM2cwN9ACriZRitKKnarG0Dt4GUj+W8mzMVmF3fL0T
kbNrDZvuzRxN6wVy5AEWkydFXDl/dW8L4sbd/0RN+DvYP9AWeC2InY+lf7ARdQqMrK9HuvHXUpYZ
6g36S2d00vLj3D4AbuefUCCzN0+9WWdDqMb7HCfJTQQKKAnuJN68+FMznahvqdRVU7lRMBcj37Tl
ermjRgTETErgylJEin3kiQc0bGg1P4wen+oTzJ4vGs8BxuGnc763ROc6uJCBCWvE+C/hZj43T9ak
VjPJ6UrxoU357A/E8PorlFGo9ZvFW9Mp1+VSkGT/SXlCmfQI6Wr1Xs5Qc1ziBF5ruA9rpzZx8ifI
WZonWEhSEUSQUwW40y/Ldkco5p4w2VPWSwoIDQppkD/d676fAurL/sYpERPyBIYlF8Kre2P3Ly9G
nYhowiA20SfG5JU2Timw0Xgj8ojgXFXERffBW+JpfZw3A1KmXu/Y/ECIMkn5Sy5NxddGbgdZgAFJ
hSeC6iqvYPmflq04jsQWxJ9aFOUNQaQnPjXL5vb4FoCvkRzX4ye+YhmN/EIN09gUgP5FymSpeMR/
wjsl+aOhUkqDpFujzgFyaHEKoLDrx1L/gearV2+JjuQEKUJsJqcdKmlCasCMDNFclpREJU1+CkhV
BAoDg1LZ60rkOHfQq0ICzxHXbhQ/SegKyUqDibXzNVqgixEjP22xaOC4uK4OxbMIrKZya/I8FBfb
9/c2oJfyHZTChIaC3WUQFrsAvTsGd9WPRb5zTc9OPtb+yzvsw8bXVkA6m3E39iSMAPYrNnX1jzcr
LEkGcngeTxeTvq9cMSjwOoOdjmzQDgqU0JMMQIapaMuYO6a8r82sjz4rpyKOzSsfmUAZzcTCmevk
rJovR9pO1CnCw41+ElhtRlS8N0s8cVlerYCMFFH3K3wieUokULxDUSGIYm6drKIvanx+NGyLv7hW
FWLnG57bzJMcAIX5M3gby+3fx55btyvk9BEQgbOCsR0mgYb6Y2rkeITOQ5m981sJTHS1xGUJXuOb
NpDEMkgluZdpm0W3w0aStHTQs93hhv4+XNoWpzMZVCJmL3fa9aHLzB9+DTOfiiffiVxHC0QZrnQu
GKUMcExju1TTkMjYAkTlPZtw64c3SGvKnTBqgmD6o4jqTuL5P+Xmlrywg1kHijQz9TuSsj2Lhuzw
Pz6WulNbdg7/Tfd6vUvM4oK5t58l2JSvk684GODuXO66+Qcdy9zF8JxpN+GbDpoXbhzU8tcSfh+m
KWyFHfcVwpgieQCteisSacfw1Fi2IkcXzQ6PjKFTwBb0e6j2CPndUAjc9gNl70qYmRiyh84OWdag
ALucD59Py0SOjTarKRKL8kAY4quQcvWK4sc5UyeIy7duY8lXlZwey+uzGPPPDfOD48T6X9bHdj/h
VZm4x/XG0hGBmJ9Atzr2sJM4Qe2ZYI4Mi+30M92oGSLBi5dsfLw0qi6jn0PBGYo8GAg+WZKBvUEL
2m6EuvNzyAaY78IhKStnYyDcZLer7wyevnP1EbxEQoWuyjz1///hzp33oTdS1RJjT2K0j8mIkZD7
qL475dTT9Bd0fj/68XevPTGDRGNf1B2xE7ITQ9jvqIPVi05NGx5JPmC6eOEqZivJDO/ApwwgSJCy
9j/HjwxBYZ1DiOIXAmtUpkZ65kqo7Zc64vT52xtnmMYorMyITRzkgIbMuZAYcW716rUxI7S5SSQ4
fl8bIfQ3NzuwWv8NEQdgfEFWAZoMHWegYxn4sWuVpnHjMVkedLYNdH0Oynnq0zJPtc9pIR31yyjU
AaIvtX7tJqES0fF0muVW00RI5aSgsuFsB+J9O3p16Vg1YdMZOTcF3mZNITlA9R0zjfIn0Rl0GRcN
87+IYHvPg4ECwC/xLG099Z2UoedmsGLp7o7kUmu8l9hUKz5JIjZhSbdRaCPUjaZDG9T8aI1Yf4OW
arQ3xaPTcZXR/0jRFD4nkVbgxPHRgONfKzF7Roapl5Gz4EKFV4WJk4eyMvXKOPok14ljcBwzmXn+
YiErIyKlWqkDgXiRR5Bl6AtckU0Ztxxh3PrKAHRs2w6qkfHYyOoesY0S2Ys2wKpDwuorquodcPPS
L7DIVJvPw0o9QCefmkAQMzCFKKSttX74daTCeopmZOUVwXIzmqF/oBWqewvW0O/+8AOympZfoFjH
COSgUtwLPOkXm80b30rO6JNvcJSlRGROJblMgspzMxOlrvCunUUkjRfdDOtedB9Ffqi1QUoWXAIR
KIMds3W1AmBNKfraxzHAtE4uYXVa+628l+pRGjUBWPeI+7UAQcYk1gPmu+YKY3POhVrc061XKXKM
co8gcEmlvOFotgMlSA7LsLN5lQF7vCgRet2O8B7nZ1csy6VhWYeHKnC/Oye8vmb+sd0ityaCPfmR
x45w1KCctjRSR2SwNoAt0XkIj6/cy7lpi1w3oAFOSV7JhM8cX1rB8ywbfYby0zKSYV0IxL3YiEyd
6oeXv49d6E8QApZ0j9K7jGd853zoxKu4quKxE7uPMHtQoleiHIC43ba6/nCMSa7ok5uytgoj1TJr
eGOJLYwdlfr0O5JytAFq685IlKChAJ6qOi7OTRasvnP4pTzXGwk/eTPjOYA+dhbRzrm/XUL/V7jQ
pzpVEsm1tnUeiFHhdcIR+E3SCAwDcDyVBqeLeY4gm8ohQ0hfW0JYTBs3gnu5MvgPiITGVAl9kyqF
Owl+HdGd7rXyUd7NN6MxTS2uQUVe9NS9OCTl4MRejnH/rMSZJhie+FBdZVEJj27Nh6UJP+1QbHTe
xmSEKZCTVxvQ+BrgPRcI6KYK5iDrZakyN44Halh2vbiYgyJEAq8wmqogRXYXqMitnGkFah1UKFT1
Y3N9X4lzTeP6YOfrE0KnymMv7E6BLVUfzdPGnmg/kHCBYHvxCPFPuLH0jgplDNLYKsCCm0T63W0H
b5Cz22h3nRvfFKRRxTU7CnidSpFqpi39Qox1Qv1rM62Z3MAJjxdHh/qw4VVwaXVrciHhWnvsILD2
E+kbAn11YGZc/tFSnYoBBuhKGWZqHkBgSX7dTbdV3bVmUXUtjUk3y96TN3Jayw8DVqQ7DbvTzGA8
fm7lNbS2djXPwPzQGuky6e2TuRw/rWjTDoYDHRFLSBW0nVxkszA5h19K16ZMShfHYrhHAHCgXvch
9KtDIgcgwe0o7Ij9WAigkkw5+/jNYlsq2MvfTw1sQEXfAfDM9v2iFnq1v3zoEevV/xBHj4tijaia
yea8ggPYaSRFp1n4hThQhUUXvzd6W7ET+zS4eH+iw2CMc/5sBGMaB0O/O1ZLfsIZBOT/bLtcj2z0
jeUwsXrL1w/upELImIRbq4j1Uk134FDEnxozF1eopsIoEtusUPr7reT3aFEzcH1Bv3O566UxtaN0
e18ao35QuSsYRZGyj/j26VMHdljjNu3jF6dCS5SMWxia+ZXCfp+kx/cxaukLuAfRlOnKTqTWBaiz
/ZTnbQDIvpWDoW8ijn2ZUNVr6bhvTKxn0QS2/Do1EI/HIOA2OcRfoGdhoRBGR0tgPpx3+y2G7DlS
Ru+UwD+h872aO9GbVSa8QImtOf1GjfflE23pWR/MpjfGO3a0GOm1QCbB/ivgaNf1hH7YsUAyX/gp
wPzD0Rt69/DxYLnsAQ98sxui0z6bCRae7v9iVD+ffIU4ecEPim5mWzJ5L9Ozo1gQe+Ma+LJ2vL+f
hlljyH8XURhCtIqZALtKe25PK0P1Ye3iSwyv5kGjSl/cM9HMBTDNWEY0oLwALHLedjUnubD7RZox
wAYjDQIlDH4u1nj9xOIICuQozOsOtaiDGbg5fWQcmr7StShj1Wu+3qlU6Lpujg16zOtZnufZS0bK
RJx8ZDi5svx1CgCHUbHr60bz98x80fYVQtV3kRlzinlkIOWW3yHT1UmzWBwQUCxuxewaEHmafzcL
ElH+BITZ62JwovyzQt5Ru6tYWKIDumcIhYaMvYoNnPA135aM0IOtxwpF/iEZB6IfxXBbHA0pfjTn
1id51VmntxVaRe+AzbqxWFgHCDoGnDij2bh0gCEQ8DN0VCit5JXzUofIkMmvJIV5UqSP/Vk9Z6fe
Ke4tKZyhKtT7yqF6C2ZZ56Rbsz9n0Q6wBdZ7Akb2Dt4JBXZZ4C3YKZk/lRWRlI10hGwjcC7TGa0I
YbJQ8n/tGDZgSgDH8AoAvEbnNDj7JsXbhHFi/rfSWf+8TwPKtGI3NHCOHSNDWpWsyr1712UxhK10
xiB5+m35aq0TeNeiNw7mTJ4Y0LbelIqh5BZzCrG/X52Jp8x0MBtVPuhMp+MZAq7GjusHjdmZJoLT
64zAyGBCD7LcGzzYSk52ZX9D3mNP6c+GXFaMlvcORnHmhAHHxEnsK7/tKLSyNm9WhUqCeyYoX+61
XDymAkfBpjVGEMZLADmzMCUJUb617QlbfeKJsxrPiNzwLWgXj0Ln20SPzH7tZjx2oJfJPSPSwR0t
59zBOOW3+/0KI3NEIvRFBF2CiQbe1J/5NFDtxgTN3jczOvZnSNJamaEd381mVQ4qfjs5gxxOaJ8y
phGMYiZIlqO+vNNBCgM1Gf+JCiukkYfyZ7JeieLfbV6Oq9crfT9JzTIiEA9tTvBn1qfwgBeUNBHS
g32a6SQcgNqh36JRDPmn1N8ykXrY2blp1CR5gE/PczItRs92tJ6CFab7DE2Yxs2trtk+W6glZylc
WE4+Fo7crc08xsL2Jb84wk3FQgQ4pjl658MeLIymBjibbG3VVCHbk+46Zy2p/9Y0eykRpmhjg7XM
bvkbWCMntuGhehO/fFtk14+1dOrmc7ytC3WXk1VhuYyxcTz9VhnNRC5boq3K7WAxHvHglRRE08b8
h5zCVpOP5ArqCslZ7TB2tb6s7U20Xl8zRQyF0dXOl3fWUic0JQo9YQBQxdKsdTHpw8n81ELkiPiI
nH6Y56cQH0bYvkxiRtu8KMVyzMggLblG6VIGmv+FMdRsIjnIA8SQMsnL5aCYm0pr9O49GhlP+9gp
muhk1Hete0IYLv4VIoaZ54RnIW33AnK8vF8EvLmVu3CPM7knbqP9F58pG8xbEPfXhIgRwDJPbNyO
DR0tNmcNgd/6SElLk36LyI5CopCxpnVIxjTRhdoluqkyS2TQQqAzHjNxhu8J1WqqOinV7Glpv5rn
w26GAiOs8Kl3AsM31bA69tXZumC/LeQ4Xyf9irrpECvk8oRKr5BaanrxAoK4fhw++hloBc853LY+
J9x7l1Etxsr3uJzhtuSx3fyUO32fJkhNPT/Elj/uCfvKtpsjPpxs14MGnJGypf4v5Bmp7NkxIVza
jIbS/Depc4wuSbRZXOenR+wf0o4URjv2zsts/LX+DdMk0LWE26eZFfpQ9S7DrEDP2IOu6hk2zqSS
BgGjd1j6oaZ67KmM/cbn+BjchdaiAdh4R+k5wxNxCTzNKUSFvEiykgWd3l8ixtukPMDIvej4p7hl
5XVOwjlT/W/DVLiZwCLMaSxBr+e7O/ZbI8uqFOoIHG/INygMVBlIaHNE//MBd/jOPD8cpXQIgXQU
B0UUB+LOsc4y5CN0Yo6tqOaH4gVfwv7cyGMx4oC66S+DAW58Y+HOMwsjHRzzhUITiGLWbDUeLxMi
viCfKnk4fssCQEDP8ivX84hNLrY2pIv6YY4dezKg6cGFi0GWL8iC59K64r/o4WmGittKonBOQxdN
CdwkV9GSQ3QRg4fyHK1pFWyINQ+kIe3jH5nmiGJc+CfIaphsMiuj7Jcnmj9lVs/yaCEGcx/R8MW9
ZvPZ6/ClcmLkoJwfglRVuvvlXfu4MyYUTBEOkU+bocE9pZqV4lpcXEiqe158rY8EYJXBbo6PDo3V
TOIPim1gTik5tUc2aN2zKakD1Y7TetalmaXL3LQyWEjk6UHuvQgWbIngV85Q8ufeMyaG4P1TDNCX
q7V4lEGwIoM7dt6FTV2H7GAXShtUZwiA0TxspX5p2JN4SW5pPowJa+7iD6rG25vPnHU/uzwsXJQT
2HnnQdppILkER88Sv3d7Ym6H2S2XqpXA2quPydHDGxjIrdjdg/vi0FLqeBSUe7udqbrFdZLjAhu2
JaV7CnUdHVkRMTDk/PL8CufY2xPCzViZZdzEZlpbANDgElgQ/pxVM+TwvpBUSxqO+hJjQX8sKVyv
KbU6R8KXAYISF5i2lTvf+E24ERjTM6Wx8nbkehy+Jgsdz7e9iREYJizSvqylf//IVx586InLZ6EN
+1pEX5/SJnVG0zQrzE1YEwE5BrtXazTJimrTOjhKoRwjr4y89ZPgQpvzdidDTiuCWOKxVQd3Gk/4
xmUvWPKTrsDNCSeFVvv9Qf7quOuebVWOb6Csx1KnLRdt7XN7DJOniT4hxV0sC+FO6jIGdK3qQFGS
IM4B3xZ6VJFniKXnZi7XPSP2c38WjN4gJPjbcfsT/2NAHNHMd4ocaiFGPHzd4gxSjPjTy5lETxtA
JaC3P9wXVGXo7Uhx3yubGIb7Zs/MzKPQKv3lqNWwJoNnepQQEcHjNrR0qEvYrOKpG7bKUTPqYvGi
z89RJW8O5GEdm3WqQnyYoiO1L9bHTjfd0C4p8H0/t4ReMlTXHDOTd8ftp5e5wl8d8O1eCX0d/JNU
HpQ/x0PMRLD5lHlomZTyqVqc4JS7VS27936swSMtDbQ10R8h+WmUCg4dmuytOVQrRF0sYGEEpjFc
r0GgyGcRIi8VMRGIXHUXA5XDsWdC8h0HP3bQyhuUaBcJyLkFtZLBOY5YchnVuBejhy9HQLbH3MV3
qC7ZG6Mrd2c7VvzkzlkHlenifb90z3eGxjlqzKGniWeYq70PTTg2O2RJDuL3YddAfjEKRZXUmjwv
UCrVHPl4R91+Tu1Yd8nyYmqA8BDfm6/tEddLshGzAsKgirYSzM56lsFG+n/+cwmEko8xxliqOEcu
M+Ybgqa/tbtQcYCM5o9y3SbMGGet9uQj2n3K3SXaOKg/EypvBj9X/PvrO8YDBOlwWcSdmg7pbWUJ
QfG4L9N27/W1imriGGhF4o1DcL2GLffOjGLZ92p5DPkQclM6SIkO9K07TixMMK9Wjw3E4XY3NGu1
TZZIp1/Hq3dczcfRvi0+0hIHUxvgBYtOk2GJWw53FzpxAh5bW1EzfXDg10G5RDpi3lUerGGSa9Yd
es5SPgSyTEiy0BdqfUPiSGjso/YHySlXhrEpqOHnckuorvBG1l9hxKUQ9CfQz26QPAkXUlKC4qPB
9Au7/ZrL31Jz1RjE9lJq8Mb1hvJTaU5phzKeELp2u0JukhbBLMCVUXcHscBApyko2wjr667iT8qx
6eNwOuy8t0kbyPIDbR3vs3+p6+RftxWNNZ8n2RAPKlzzqfuPYjbdpVntedt1SdfK0OHPmDIx11iO
CitC6HVfmZEhaDOgkv+pntIgbEvieeUsOz3ZG/URMks8iIwlTbs/ggZpcOAXYgmr39IBuRYaI237
1mH2N5Apq8uh4WNyqMoGD3fecOol5c6kMJW8SXJsslnmvf39FDnElYBzLexGdJfhYc8za/ygUVZa
TliFcunix5M3EzH0KFjql5wmBAgvcqRcgiK4qdxflw0FLEcs9LoasBs6sldtJ0cM7AI5ARuq4mjy
7KfrtFVT6fteCFl7VZZX4zA8qLiTpmdENOCOZBbSAKJhKTkKEoYtQp4wPqFdBuD+uHJfU/9nV5sP
7+ZnzyCB6pRmDjvVfXvrLTuZRkSK4BkCM1KvVVFiwDYkPoDaII30AvWoTEp0CxQUqFSKef1aN6Gr
E+Kc1S7FAhfTwEck6Oa0wRIg1VzMm4schuVSp+GgOyQ7T2BaXIGnXkQxkpe//gleJ4Cv8Y7Z6UU9
33n/g9XC85fvlh8N9RhaPpmQCCObU+845O1GxXqUL7YvEalLcPzma8f4YnLjp408fFJkpMDB4ovu
wrNe3DyOv//7ivvHnbmkVJ0FYUoMoG/6GFQMhCeKL5kNihxhcazeR/4VCbOMavUn28Bb+n6c5qiH
0rHxRimnD6goQzGr046uCfGdWWOCmssbdm0aqUhWy3JEzuagPz598ujCgtpBMpFNBu5Qab7Oovrv
tt9FQdj0g1kiryV5MaiTjGBdbx6xZutEGBqJk5aNmlMvR1JeDwjnuDU/n/8FqbIx/qddID5T3Ref
r140usK/HA/doFs1cd3a2gRwB0M6B2EhvyYjWS7SKf7BZ0fwXrGLeBAPDhoR/BBkeJW78V1c/PQb
dRLOgIgSrztq6FTyFuJkAeNo4nKlxToYJoBUWDvKpJsDzZ3kZvaiHjqM2JHggBnkr6XHfzbfOnks
jFBT/pSKajwvu9gnCw1Me2yDAK15ft97ESyficwDBwe4OaPJKTjJJXFGXxrKOj3/EzQccOZ6VTBt
g3gOnj9MRic9CwQ8x09aOUnxGrMIlD6234Rm6ByxUr2NwC4/38A8Ip1sxEBxqvSPqlReIf4KEWwk
qJ1Y6B2NDOjP16Rfft0OVCrgcdWXKw3YDpjExD+crqXcdu+hULv6sPjcp+ZEEmsEXH4bLgAeREu+
2DlgnvYteH06oySXLgr4OHKrHSiRa8nibDLYMOnG4vZvs+ksrU4obsHlfhIgXKWv0K4M4nXgF108
SQmqqKO0OsSMfdn9AhI4HxcLtBTE2HD0qVTxmQq8uATAb7pp7yu/hAHM0JOmFbQ9O5LNLoU1bF/5
rqdUS+X2Ty1ja3BwdlDeeX9HvxzHsnjreHa/QkKsbTpd6yi6VDj8L1CZg+YYZIwwGgZl27w1Dr8j
aoCNF7U4Avu/UNq2k+E40U3gfxfZ65p0smBlg8fLEN2xVa52/vr/JKVI9BbX2jspvpH7Nx9Fje5H
Nl1rnXgqhJP0sdXJGfHrC/VI0vxAs3EBWo2YxYpVffovzbmxCkI1ZqfgiGmXC6LuEd3wG4cZ/DoQ
qT1Oih7piCFty8wTWry9FPnzukVSRckfRIrT/tybN0oty38SFOS2mn4ah382183D5gzlkpEcU7ur
IKGgNEmtrhLyEsIsRP3dNO4AiO1VEWArUJo71L1v+0fzgj8Lp5QhyVd/sUnPRrUm2LfVUUAFplEB
mfDsaXCqu0x0Q6FAAKw5BWUUbKU6qSY08Ag8tcbfKQkv9YkdT8hz97Tn5TvVuUS0oFrrSqjlh3+w
gT6cedFUGzOifA1hSGrrP0rQT7Tkf5PmFThAAucVCYH5G8KhYobUiFZXCsAP69NI8Ux/yVg2M4TC
0LpKUhLTc9hOeDEglQIv2BFH22X9vsSzNfPq89ZFfP8x7yJK9W0q6qi8GFHrfyArabGPdtAAlpBY
WrcYW9ON4NGXRCjFlub65Vn5pOPRJQ/NhcdJ0qUxrtNzHRax5fkruLiByd8Odjwnv+OzObd5GN1J
haSxet/VGfH+g+YWHOXcCW1g/smZmk7hZSv0Fm8fGd9cdNjSDptEutu5QXRSn/gH2UKa9GiLZL8N
ji9TylOeC7SR2a/aTaEKX4eq9se3iynqrD1/7N/VPIosIr0p3XauTclO27EbfxDvDIGmIjIrqFyL
K8MiP4NVvxfZ/hgd0QuBPhFgCsy2Z3MzqcdKle3TPl6KjFkteDFaB7TrDg+h2x1B4KU0JDoOnXiK
hKCsdxnsc5GwAb23EIafBo2/5W8S2PB7Zy64vQa6fp/XlGlA3J6k4TfUUUzS6CXa+7bxmKeguWRB
A4m210SBi4B8XaqNT0CxddVcpf7q5SomNPIEN+pstT2JFl13Rw8LPPtvybdLmLeenXtkCpmRnL5J
CZ0l+k4e4r18KPJC2ClBGtbsk20IEvPGKKyeLzaMTeBdnI8lmS5douc62stfYn21omimgC/U7yJV
ZGAAhA22QFbEFKvHrVJDCsHqu3FoHD0PX3TsybcmmXoMdUwGjK8f+UvnJjNuis6AiYgzPxhxGeOC
sDUP9e6SNqpJOkBPluC9Y1pwtebt8ZI5XEpyr8G62j4EqJuG7q4Rize6kl4yeXyNqsHNHaK8Zzyj
WUlK7KbuVFPmoENV8lxLz8KvvCif/Rf6qQcxcfxpkgf+wwEx7MObeoXMVeLn9tXIY3SJEn/M63OT
HFn2wllVcePKJNt4nmpoYWgGbkQII9tfMgYa8qXur4+hCuOdWcVx5RxGKpi9yL8L37aC469cizH3
bqnbg++9sthwxacKOVNTIyUneGdqfLloVscYnRLzyfQdSRd2/Xx8yqEJ7O5a3GV+k7O7nNShhEFZ
I84JyjRjhOZzpYb/M9vl6G9QqgvLIrQXZ1nD3o25MJA9l7Ez6AKYUYgSOFr5qbyqaWcfJIEI3dF8
rZMWa4SZ84qQQBEDJeuGgYAlOazzqPriD7ybDIY+lzXOxPnA5Il6S78cznBWOZQ790oUqJCTrdZG
WXEKRteCTpO/iRq3JHvWX9JpEgjms1GQ0O9AGOoJaWxjmf33a3BRE5hI3grkF1bJSVLjtzDDU745
aDaKeVrxknVzOUVrbMQ4lR25WhKXUt57Iw4jzCc/c0nTPemwSPd5u15gQ2cER/jn56V15mRbodUj
vfVeXpdwtZu10ydl3HRf7hylLHvtyrMWILkMfLEDwGWhP9lHUV3iIA17WpgZ2+GzsD39jzXrVqC8
jEbD/K/k4uUY751T4iscxbsrr3H443pf3hfB1EphbUcWHAkTYBWIeO9RuP6OHPhCenkoxJhuWnG3
6s6VRDAWUtHIrS1OJz9aaeu+tRh53z5kCETu6WrOd01Fy7UQl9ylUWXga270ikdqWyeISklRYz+2
Zuk4zIkJhVuv/69e2J+jJduoquQjoFgSOX/9WWm2zapiiRvpIGeg/TmUkglwt8NVvZ58kfxwWAOM
0K3Z53kvCbriALaX3T5J2agwPsykykGZLS071svhPuv+yARdnYwqtUR5LeA9AvfRfudD7KUFNDBK
k84w4FSgXDzZLvPhoX74F3kLqYCSWVqYO/zSK5DE2UBZGMmGUEdwCKiLqLrjj2YJ1SduLvxhwWgL
fjhdjfBe1HGSd8Qkux7B91tpqJQWL4WbJRSVV+5DubdXYpMPUbg+ojD3HH4+BZdx3lsgd/E4dzdb
1vND/gUXi/KRTpABLPDG9Dst749JYa8pZTuJ91ysal/nkWXys8nwcEl57yeyRu195NheabZI9zBU
LnqxuhJhIDBpdl6Ve/Jrf0cniRgxFDQX45OdvIijpGU1RTxASbPYlPgW7eIDQoaQdqnQSLNdpvft
o7c532z4Hlm9GulrpZtKiiz6EUHEqzxRrZTq0iQRyJMJWAsLPNVNeUVw6SLADqOUkLoFKSjodU5j
WVWmPaEcPSAN9GBMEd9rvgE3+qoW+4CEQ/QYD/LMNJzqzs7ockSfrWyE9anf/zdqoF6IbX7BF2dc
28OMu1m8KWr8Dxc2IsKiLfFZrv0XIcJftvZs4iIbMUaSEHuOJfkYwm49xRlDZhgFgqYsglpXOZMz
oWIZeKPu+6NrWzS1Rji4cZR8qeCV+O8wGWnQE+aEpR2e9aUAvKwQanMPCIuHYX1zgy+H0Wjt7WI2
u6axfgvZoP8FR9jG0oBKtzZ9wOjvodwRZmrelKKcIsFIydkDYHyIOOqqFKSsywPY+z6GZg9iLFp0
ajJeItJXcWyaWyPHov8IIVSD7di0c2yWNHwi4wBzdp/ScsbwyG1pMe7yX0izGvrLyOQSmKlWVu95
/eNb2Pul5Lml+HsosuS6kLenUutyesgsvGfAIezq/0uAfxnVQ5geN5CHchfehP7PhQTwenNPh+qj
aP0md8+1YFUYjYSMsS67UfBEzO+RpA2WhmqTyvjSXA2DOUeHbwpPbCyueY51B1JoW29V1+AkqbT0
kO3MMzTJAQhjaT4fxLNCVFDXu1zwEmGmFt0mI+Xmao9CihJW34ZHIypJucPdDoakXxikoDsYjSA8
SBQrkJxkjU1cSlMTnKUW+QQRUI9Efj3Q48CaF6b6kChIH7kIT8aCQwGPySnNUK/FFh74vpekMdTm
Qejhz3WdYK//6GwZUm/7dmM9thfrNuvWQlHZSCtjq9znp9u/ldKUUo+DatgFu+RxqZs8v2ckKwk1
MQS4OXdlUZ6Dt+hyYJvCm4IaqXaayemqSVnikNiLgOForgXZhgxeQzuQ9cqhG/rSv4v3VLZYxKQ9
iQFtkdsenPMkLrsGDUrClt6hNvzoVTucFTJp4yWEfV9TduuIWegGgOgAoWqe433Qohlz9Fzq7lfm
lOPCUojdkSxzYJNiEAMPi8OjrZ6qvbnpGP3zOMNqgQLZtrck4tdI8fXzhVCyjWxBPDdcvgTARqd6
CFsQzN6eVrUOn6RKYjtH6ktrTfBZ5n87FzPDi335NvQIiR0HBuyywBfYeR3kriT6UHdy1WkZpfB3
1OBDNc6BMFjOr8F6zAc+sj8jWj/gUA+uiLDagUoMRMBfhYTzC5ZY1t+afaO9qUvosCsWai12dHUj
05BSGx7S54NUjBRYoP39Zx77T14je9OJdtHqDEVuesePSDxDnVuLbt9kqp+z6UlzVQoKG7IUMxbq
2eizz1UY80+LcPczB6FrJkBhOnnG3L+yVl21SMwoWkB5clMLLDsAlI+39ucTc9bsc+G+jJQTDP8d
03ZraMB1vhVe14yEwS4Q1aac9ZMsjpBbCvvhsguOXlbUhbfs7V3mGN3gcD5JsmZYYvxl5xV5EUbb
nH0q2vyyQumKTO4hc12BYqViCeEHF0wZoi4OQDEQtTIrnF9hpdHjoGX7Ro/pWZdtCnvfhNMzEb1U
D9QrsbNTDIBOaR++f8aY7L6ZBX5X468nBFIaUYjyR8W84xSB6lfMo+XvP/0BsT+Ui9sK950lOna6
d2Gmf9BQf3+PDdSki4jVwuqG+Dy4OOn4L2oMutdHxLFVRwFMQ9pKGx5IYD552/URxl1BaJYVpztD
yRHr8bBFhD5jidq+qrK43C6MqtGLUkWpTLykcJsoSFXuNU2mt0Jk+8GlUhuieBkP/wTF5BYyu7ZZ
6MHJDbtZJsp8f2n1SYDGuKnPJb0U3cKk1sD6BdB07KrsChisLXXmi3wySqh8fz+YM917cUxgOaLJ
nm9cb1icD2LclTaGBejPXzXxWq0eSjFiWGvwouKOVsVpkCPhVneO4R4HDcLiHe6O15Msh0MnSFxA
/+DFUS6U1GZnnzZ+tJLjSCHj0x/uwaRwg12z06UK9EJ/iyH7df5V39WKd7zcSIaf2xlmD80pL+57
XXjpeeQ8SCfZgsWIvyJyQMF5YRPg71ZSHpxFczVX2Tw0TJHW1OUwxYG1iGq6Qqo2hUB2apDALDIt
Mp0Ae/VQN/2CBuP4H2d92oIfEUvtrZ/CJbs8np1PZurGpOqGc/M8PZMJbqwRYpCksgZhgY4q43q7
xKGPL7erkL76RF1KZP8IztZU2WNbqtn8HuJqpt/bVgZw1nJLuPczChgMSo7LdnB+7OQlGz9tKXce
COO7bnkMvWijvGnnPRlTuzsbJLnIzy2WUIp7ZA6VKZdQop0FvWwyXgT3hSKJIZHhxTnzaS4yV4cM
/gPkAmR70Re+MDR6sbMk7S8pOYhJOF549dCrOsdnvb5tmvi28D+tf0JkiN0KYo6E2eXhhY5BC0t5
DLnG2qPDU1nUFqy5mK88E/8VHlXqCT0y0kWbDCAIkG/J8QjeNg1giiwaDL9vtMSg5N6fAnL5CH4q
jycLWFN1fPxTd4iQ2nLjF0uH/KDGrd4Bma4FTdpBoRvvy5MjtYJYfYWqOiPnU4nECEIOSnFPRDH8
3QuR0BwUf/WQfpuzKlKAkVAAYloSPFkeCRZDbiS66KeSoBdcygQtZ+MPqhbgIzjFI8equmAWivMT
PNPkY8So0fW0fRMdnJTpwIo+ETsmUXVjdT0YG3dU6ajMadhIa2XYfeEWNcRxIPWio5n7vplZi0Y+
3Ny6hiZ69IL8jg1RtWlpUZCxR/SF1Xz5zXxZpy+EeRFgfH/toaT4zjkrE86PUl2zsyNzdDP10apr
9zuldhD5YChVf+HDKFZIShfTUIHlyezrCapQ+h96oLy1rRdkUvRKj/KtPfDs6IdsctFG9nusUxVN
x+cGqy6M/Gf+1mgF6Xmx9DIKOKQiDZENvhm18J95mr1LxGK91PVo3jgxOZEzlOcXZTFUWhkk4GU0
f96GMMdeWkBoU3btQBURcKHPG/+HuwTX8PqBTZ60bSvhPJXeEiXSSkgUrvVW9rKXaherECMtupYb
mlaoIDHjrbdja/i6CqcL3IJ63U8nURk3nVGfiFu1IfDL9QqV2p98DUo1oNbql9M8HRArNf0vgnCy
8dI7nphULcvO+XBIdXnpn46UiZGnEnr3FYapuNbllEbit5C8OeTUZirqCQ5AtXOSCMHRZigUvATc
l+f50yhktyjbAGE+nAQ9DQFJIRKNVPWdi/Ve9GWDfjm53YnPAv1RPQcvh1uxnsRCAlHmFeP7vEo7
Axv5QIxD3fowKIhEOc3SUrRcFjJfbpZd2dB3ErrIuta4x7cU4aOE9bKLu8qrDF/gfUmpOsAfNNbV
jkzQSzdKXGEJTqvsQKHqMf5LYVR1Stofc1vsqqTl8k9lcYF1RZHYW1+HfaZYTQx7R/g+wG15fAOi
9NU6e/TTzljQoINu5Kw1jzmJ2eLuPdLc6lwMB8xH07tWzfOLShLKu1RA8kPact4MJ/WhgXBg0kLA
M5AkicpgIzM61xMb95zfQV7CWnOtafSaMIWe02CR0nWsucJUR3EeRICBfXvlPYMbjrTkj3hd7C7V
Mt4iP0/mpQoj5BiKqe4JoKFD9A58vP+hIVHSzcFJnDi/eOnlBe9kxo6h5tZL/hwLPytbpN0fSoMT
oB+zphvsD3MEMl2GSwVlq6AVQCUbO6Fdeje0iSrNqL15THg8j2lFcFscGOPJdP14/lKNXzoBbGPW
zq54UlvjD2A7D3eSbKyIICk9ruL8ATJfPL/4TOJvHl71DIA82XWdZWl1lTQxYsnYdf27mQgTuJSv
KNAbIVXciZDKDIpZ1Ff1DwyEYMwY3rs9DeAiVTY6cn1mgD5Gpt2xZ6aT6fVXJzQHww/1cjH6Rtcx
CA2VSM/lCRxeLfYlHIKLvHWrh18h8btE7K3v7Q12Mw8AOv6j/M1/Y10a+K06gK3SCrRkWcZU5jtH
orIQh8ZZsbOJFnRDjxDwTkmTt77Cz3jFujrxwrJhYuagIssTzHtKv+R9FaDSXUGfsBv2Q1w5R4vm
PdQ8hgnR1kQ8aKFAnC72PZfGxA8ZhRsFgoBmXvnSStqtjnfkeHRzlVClZRShOM0bAJuRFB79xUaq
D+NmjyQz5Byg6p/UCYr3IiZaq94X995D4+6cyQAEfYVmhsRDh3UYF4Z+pubfnQEayy6FLRe9N344
HfZX8ltwywolNsTkjm5xSyfGKFCDUXrkEe4fQwAf0fDWKcKasYij6KqrfFkhKGb5u2B1UWJg9UJE
bkH8V9s8GBivE8DdEmNjb3F6Udt6PRcU2qBzblVfnnYNT0s6tHi6ZMdO+aP7e1FP3ldxzxiTbueQ
PsTPuaPy1EqfC9MiCrk2dlFOKnhoCA7QeJO29WZWZ0kQwCrI0SBgid7kCuMSRcY7/7r3+PiBP59S
6uodLY8Tkukz8Ix8FCOorCKKTlPea9HIY4vzjDFOieLaEjp6eGq5tA3/rngyVfAMuUnd/6E7hQKe
aSB44lJ0qFEHuUQXvZVZKKc4c0qkReZq/GEfvKK8/4OVUZBaLhmsxluEa6MAG/sNwsQTfteqnkv4
tFgCIOnmUqx0ian5O567p6G06Ket828KzgRRL8UdCrrPF1/KyuUnaCOW2Sgt0TL97tOn21rQfJkC
6Chk7Y4MKvZhc50Ut5Dx/dMBm2/Sezdr1rfjYQOQomPSNGwV1hpd3mraKTNoUZrJnqiD4szF1Ss7
nNy4i7Lp4ku4IJ92Zcr/uySFYBGl3czGAISfbB9FVnEMAMPzkeLRPLxkoHF693b47KtEy781DNC0
VbchIm4oFU4NO1IvcL2T2QKmAytzX7ZVrYHbdVjOssE4nxhIxFDPSzYnPrVtHA3AaMHRnOoqrG1B
hlIqQ/szdcPN5DkEiR1y8AwSMakiDhGNsF4DiaoGxBIMthFVHeZSg3VILioX3yLr8RFFMR9U9egm
cexn26Ir5oh8Mq+rNzclW2DQnNT5YvvHdypweh6E4IlFptt5iRDTSVaHnb3hh80PUJ/HffAMxop2
MlyL74LVzKBKVQnaEdt7Enbg5qmekY6K+FFYifF8Hp895YbcC7/9ivGO6eViukm2pziBiE1i8G2q
d48RwPr5xep2iOtJhmDcJAAq1a31PxiGJlxNl3wij5TK2AprtVjIFI7pTdHWWH3wyDlsxzwxWR++
lUlbRof6qqryabnvOv/98QWnRALl9NCsG/hw0UX1o5TvFYIQOSXp2zfMWdklH6NmUAtq/Ds7U/v7
thuJQPcxcvzKRx6Z9t2hzqHU8OX2vP+oPTrC3Z8uiuPjQJpkoDqALU2NiH4GP/X6QxKBBltksu9h
6nXdV6QQQuqPhEtq673TCGSdO4/QCgDumEZjMgFkPrY36TeFl3MAJaEByadbrXrmGPeLU0Ate3TE
LniR6JZ4c4N1Z2EmUpC0p7swKaAmUZrlbqfprFisurjLSYdNHZF1vSSXmXJ860VrrzalhzQDoCsl
4Bgf+nfYjajLI4SnuT31/JWzxzKrgrAa9ySJqR8u26pGWVip7IjZmfy5GHg34ftVDlA2RgRSaxhW
7TF+46Am6cYyWgcoKK5uPdiyEc03S/r/N3S6o6mWTCw8XI7CI4CXeK6rMixnP8Oo+5/9fHAGXY2z
id0LOeL/iGpFB6fM3UmTuU5lSRlzWD0Jm2wW08JkvIrtJb56G71rBQLDVufSjhU3OycLhRaSVfLx
Ku0lLEkanRFohFJ0eq5CTEfe82BDWX2UklDs77UKhI5HxCelxUO68xi7ESZhybxyDfVs2+QzD4wS
81MtjtcQpUqv49xenlRSiP1xcD+29McrTydn2m2izH1FHVIa94juphAiwo1m8GO7WU/dmwP4Rrlk
CgiwH1/JC3wFopWxxX2izGmmHLX/hecEFWu45Gdl3d9F+Vnb8Oy059YGz9Y50unqcTMvOfY/4Fri
/xS8BdaEs7covCh8O6iTEXA03zsTzt4DciQQkjiup8h5rEbX0spW/J8JcMhh7gTwwLxIrqGVjs6i
HRWwbnmYX/Lvj2XJliGkF8kzMhxtVTuoZxaJd/wWsRSrCdjbHGnDxkK0ax/ntzj2pUoODPDM8w25
TH8misBCdXjSDojn9c3MaJNKnTTTYzMeafN6GYoGRJ9jm3RoDyMbk8q9uPjD3Gqllv3Brmlw/Rc3
WOxXNDBOp69l33yYI/ojduZjvjquzx9biUbe1do1HVEOI28CH+3qJCCVDDzqsSC//KDTyTiZSRnf
aK0jMkMmRRaaEd7FOzUDvuvTBYJLmyXeWW76e3UpqQWrKdwSR41fAcY+jKqzMGiHfWCRxYSM/kU5
i56bNa2IQoWgwv1RMTObEj9fhgUAbTFLbtTTtdEzji8dZk3DzMvRJuT1vkAg8gZdLVAx5AXAd4bY
AeDrdCUJP9Dt5BvV0G5Z45MYe8qqrxPqME/UivIEukJLkD1sLnqfl38iwI4lZZX0KybR7mYqF5E4
o9kTi5yBqny3WwewjYmVfHanBveyOiujr5K7fGpCnDRyjQXYt8e0ilgbX74ViAuYgNHaelRdpWA3
pFXGFBZn5NrG6QeKmyJW1igCzpJS8evSwlMkNrMQ8ZKCFTWaiGKVKAyHyDaFZV4CaDAEytPchfCu
Q9QaIVImqPaNEYba7LhiSKFxLf4FBDukV9od52wBv8KQIv/mBgdzcSYd8jCJBLWlYdCTiiURRHfr
w+VI2Zlbf43wpeidOdY2v6rWqxcBlrpRoGnJjvyVd2H8oxZX25q+E4p7NUKrwZHEFN471NJa0FZ+
n31FGLZl9Lx6lgyUu5E1dgu7Y35p4QU9645st4zwamvBOk0Y1cRMpzNJpWaZD7IVDX6up+RU6zjR
zh91ltuclYcujJ6docrLWUqHJvRSD/xsJClpDuveQS+pHsn7in6NaBMPKa6tudjGBZRQAxagSaa4
Q8CcpFnclvUueKVvBGEfL16lvUF6VOswuExKgIylN7hHUDThLxym6jck6C6frgGof4/vwQorW566
q2dIAIUSLDbWdI9kvxPW3sexU2aQDa5ap/Pqfjil8P91Lan4dmxHQT1HHg2A0UNN1SrNmOWioCwS
qIhjMzw2zCSBjgkEHNanoYOhxdSlfbj7o2wwzEStjO/gaH/G1DMBATbUG3YMHec/tT95DS7y3qs6
tIjOw5H/sLrIyd/XnrsUm0mh1XPwZfAyUHxItbG6W+WhKE/69hU+AbbP0Q0DCw7p38kDUDrDOS9x
EJokGotTzoxeGgqbPnBtGSTMx+q42kPZ69M0j5uEcio+WFh3KZ1RiYrlbODH0uANBiSKVRKrnggD
6GDvWhu5eS4CrxMMbLJ+o5/vRqLIBgyUva7kd1OfYkAC/gfD/J9hVVrK6n5529tKCmdeRcHeFhX8
fWDMbfJFbMcxhN6oTsUpUVZKdwb0aF2VPeNdJEg+wrVPLy2ADvACONKwp0DRcufUXHSqFgILzOIO
o0ol7xe32b4KVm1thS4qNEvsCV5nXEEaS1gBtG7BXaGJZ3/GEVIaEtepXnaiCZi/B7DgMoL0ktS2
AIAPjHd+g9Ou4PNUPqYU7pePETHultpbBmPsM3PyD1mEpEkAMymkXkT3HMdxy2DuCX86IkSSYozf
XGOJUxp7c2M4+246gqa7DOM3OBow5Sjkwo9kb7RVsU1wqVnAWSaK9pyELBdh3M0HZiW7JJF/Dhbo
4Q0PG55/dxNcOGdMJGGvwpyTOOxngeA3M0m4dEN67SDW7LqFitJurnxNEJA1LVZ8gATAqjFuajFP
MkqjdnX6rP+srIxD3t495GZTsXTPRNHNdp8gnVOgsgto3cBi57n9ah3NBPmCI7TO/12sUTQJhJrv
WVNVnUWrBK5PyV68IFtfvxkHf6gZJ4BgMI2oJETmo8fUzstMrv9jGQFRwQIaRbKi3QcpYi8CnS6Z
By7cUPo4bLgyteU3ZNYs8GdHxqhgdJeUQLbNZ8JVVmm/jMJR+Yu5fIemaizsPeB4ytl3SyadLig2
VTE8f2Fg5YZahd9eZWSA2/itpV8qdwTCD9JiboAuyWrP5D/90Qc4jNYonWCTjXU5y1bOX9ry3H61
KrtbfJOx2hOSEqImLrIfSYr2YXQmq1Qzx/OYvBNAwz/O+pQuehkb//EVXfDU/LUiife0KvuJ0SUm
MXEacWpD4IcoXcjsdzK/9icVIA7tHN3zaf6l/+gYm8tAroolMaGbPFfzA/WbTxFX9BClrxlTa7uu
0CaWPx24GxwI6+ZJdx4DFnHY8ufxkqoHBfFuZH5/vdImS2rVs4652BIsBs0gMyfrnM1MX2N0+vRJ
0sx6T4jVLzT8brNRmVr7ztYRcK+eOICmm6xenGobJypWHUEUp6xS6SSSMwKIqqIiTifNzpgBNgu/
0C2Z0T01/F1eniD5sFkyG9+ptJmEUg7DSB+ab8Mu3q6KNDziAoBH6sMPnuwQSM+ydluiQpBKR2Ke
apIE4529YJtmhOvJINuOxiuFlk0T5L+N/DBtqb4gDCxUZt+eSasOXd8ZA/VGGt4Svuh9QDwyxmS7
IzS2jLrN8yb6bSeONUvkcCCI9djY/VHQqPoe+/Dh7t1AF0JNU3h79P0uoVhwl2fwwBEgzKK3her2
TDIC6EtaMOlet6uMHax86cWwER7pcEi9k3WycSOizcqr0PRAfF+qRx9D5Lv4dT80/1W7xw/4xF7N
TSuNTw2G7fD2ri6lt0gkxw3KRqD92V8vcs+0nphu6YMAtkijUPT/3wpggJ7GCqqr6yYgiazGe6Ji
D6+VGeFWosGodUVu4LoW3td2OyCFTU10Zcxd4cnIG7cwN2lVBTlUj6dZpG+XnZMBgjBCSH4Mpvyd
JxaTiIEQ8Q+RhfXmKL2wSr4UOy1YE7QzpSZtADMmzw2xHXWkEnnqqhUAua3MaFUyD0bQwFsqDvwd
nimem4N1RS1RPnDdXlWn7psRPSYemlA9zNjpL/cgcJFARLbAtb+OYl9fpCn2coHxU+M+Yt3G5IK6
+vIc2BUbCbAxHbb+Sb+vSICUGkwouU0NXywrDtDGSvBgF4Ted4iatTqXQAi6ikEitBT48efYxh8j
yYOxCwHS+VfAILDVYICfZQH6gGHAlePPiarA3pf061T5HEDfMcSBq/lLsTe/temEZO9GV7pLMwlc
Oq6Xee6k+rww2yVp8jBvJvQKanZqTKyXigoQOChEnOMbg1N49bmMp+L2FDlExloRuyhpgC+yrR5e
J3hqJzT+I01I2k9wekPanmm+Esn5beL89ka7yoF0KE4GlFSUKFno2VfmKv2Em3J8Fjvkmp5PM7Um
6wSqfJsWgSZPT6g8gYyzmFzllsND7L8NQFxSV+PkEUikml4vKMVXs1vJs7V+bfHcj7DEcjeU6MGo
Btp0dapaU2uJw3/j6jNB5plBz2e/0MxUzQJl+P/nlHACa2eDbF4L1TfIO7lEIpkYVrtN9bNVHoIY
/PzVHIIWxgmGazCdyppn920zf/vei4fQYi53BxtH8qweVszv2AA6YTfDd2E+2VA5pewLiEKQC+hw
vz+oN0/rmgqdsjHXBqQSRNXyp7Jnit0I4Ia5s1XZUBFWVaX1CXNBVVN31kbaTcCo5zsAvOLjQiCY
JEWOIieft0yWBOOVk1K0A0ihId7zJT0p6r9fNC2RZjA6XiBHpv5XTkBkqjUQh2Dk3dfE1hb4+I5f
gAlLZuc89kzN3N+XDfw7Bakb4UEZi+W3olbh5WWJKI6RRAvJSW+TnRrhFo80nu/1TGEUKzKccnjX
Z6c+FsfxYWHBqAPg8IKQt5NVDNCqdr/Xw/hrE+oIqrAsBZgHCCq9jGlxJZnDP5xzVNExYqUFUuqc
9jrLlIthkkvsQ2oJUsGpaVlOI9joUEuqnzSvumRdtmOHZFoghgA4e+vNVVHEkkVSB1g8F1wzkWLb
CtYt+dFetycRNxAenxM8QqLf+M7aufGS+uLWPTEZoap4AFXnLiE/cosuaOQUpKExoiBurVbe8q8H
KKl+naLvWdMnJnOPZnXOhDpSdee9pwx+8bU0aKlMboePbGOFNCIs0ys9xS9qSUR5tc57syBexuQu
sp3KEr9K6TXrka17BWYZUGoC90byiF8NKEGMt/sZRZrJEYWDqc9ksDbzdvxJnrk9pcnvyCP6pJku
bu0+TAFdDkqftdQSWJbPfpjkM94LW++CqoOymckT8B0Vza9uwbK7bq5Gr9cXmMnf0NFfPpAp5q49
u2gwkO5sbILQ5CK3BWodat8fuUgKzmQCOGCYaq0I1FZdpPmwOAntsl7jiLhZWD4+B9LrWCTHUggu
+HJPihb7V+HmVXnXrOcmbAJIySSYZOWLkIGXNbaIaMg7FZ0zgQ21mChXcVC8VwSroj925uwLBs42
lsDdyCGEUWTRvEf+fNam5ARywcIDig7KmZ85XcKm3Zg0OI+t6Id5c6vhy1zurYRpr0uGllhBu9rL
3imXJTynD3WT7L9UnqYcJg/IUKXpz1DSSa4VwTw/AqwNwJ1f7isewv6WjbwkvsIiYO28h3URvP79
YIbjxSsyPVgxzoLBC8VsYlHpYpp2vRwAqw8t0B9kkrU9ekFDqasAxyMM7Gi1bsM7o4XCfos7pCZh
lDHroWVcDKDA0cK1OTJfQkDoFKh98qAnsmOm8GbsjcO2BmAEPViPDwy2/mjpScVIqC+Bs2sWyv0j
O/ZAjCJEupqcc/LKJGt9Vile6kEVSweRt8R96sLAT/t4FGZQo2l6YPXbS3QXxzf+C04t7NToWcZm
whDRBsAabk2kv4QomAIgoYTa56PvbywlFoLgHcQoj3snqEzgJVkvNYaEmvPmMn9FcdwVxULE83WP
+MUvqbH5D8r352oPaSyJJxRFBMUEEX2X5KqSkgXMcL8jMhmWYXNlNYmk1ioe//CjEfnC65SiBONw
wTJ4AR+U+OsXoqwbii5PVLv4oUz1066emXgS0jsZAo64FdMxUFzhKCXi8Yk/f5v3ero2kNuLBLeS
3KfkokA7NKx+WQcr/59BRexYJ0clvsPT4ZSGdK2k4m9Rr5ekkzMemlEHPsB/POknemYHmVXH6eaK
10E5cZgDZxyAbksxlsdcXlHoAEaHyx307Hl4S40d8rrd0yjWflDykKYuDj73L3aH0kjHsdIyji4l
KdZvMuOWWhAxPR4yCbniQ09urqAR6WqMRhXLLcegwmFZDAtW48jyWvUlWJZLkPWvX9JxfkiUamsv
BulpTG/VyzgmFq8LrjzOXd2Ay6jyiJ6RoRVFiKi9EAEcIk353tnTjmnaxLMlDHIZYXQEJt2i9tTS
ypIxB2ksZ4iWZRA5eIu+tGOTArt30N3ybjRf52C/IzYElByoJhbkoy7sAoei8Vl1f8+MeJpAjWLX
rD3mwzLVM5Of1dBseQAWeLAjludf3sZTCCu94mAV6z83mcda5Eij00xYa3d3vL/HcToiXsrzflha
OXaHEaa3N8yQ/kJoZSQgy6zJf+PckPXN2zWmgEiyl+mT7J17/fNHlKJ3grE6gN432FNZ/4m0M4qC
3UahRX+od/Ni2grgPYMxrSvWsWZC6OU6OnU0YhVVPb68csHMf0p7AMmerLzICekUZ9obdAb7iCsC
Egl6oueDAofFYYO4U2a79JKNuFCZSFcJCevrqY/FwPyxrTZfEiEx79tlRRn9kA2w0uJzz+vv+le1
m2nXL8X35ogIhRFLoh69IJloSBEw4aaeZCtVaizVKnNdaoUpIGRYvi/mVgYBxVlZcgtG/dlwiuX1
fVuGoSGmT0GmD7bCzG/oR8ThAua4VfTvEfz0yPGJWt/D7FKzpQcdHq35kfuiGHs/AvgDZpkUjqd9
SXClKZ6Z+cmCx43+nTxfTLQqzWtkJ9ecVkinaudCoYLsXi0Vq6MCcw5An2G2wlyPJOYRpNPTUDbh
Haia9AKZI+I19598MfNJtrtaIhLLXKIGtMed9lmQNEV9F6RXoELSDSipJ5OS6NlIkbv11T/+H+Ud
hMU4vpsHFr9v1BLdLhqIShvJsCKVLXYsKaM6YNoASWmXFKNpAB7vyaBXOLUNwrRWp7RgOv3JKx8G
bsNGHsvyZp/Y7FytVBRgYPkwyHP4aEMCfCbkiMZ02d9GOccdcJuJlJxt13hSD8KUMO00WezcPoU9
S+6rNsjlXtSAwO6J3gdsDIp0mpThIo74vu3q3rbM/fWVl16UJFoYDUD667w4tK5JKwM8GTXGYjgt
f6XRnEuu2mVzKpGxB2PBA4uOb7WgjQEXTCWns5+5HrwKxytj80atU/CuLeRYyqc+VaIr9iDojypQ
9JmtmCtMA9T8vL88rQuz0ptS7j/WT6pE6onaRo17GKAY2wMOntz4IVYQt4/IpfoewAdRrLgO0Kz6
aZbgXZbtVVbvp75SCns3GsowJfZ6ZwRg5vZQQNtLJ9c3BI9N1EK7eOvgpRwGuID+omqYaCHhRdYa
ZS4o8EVqqYs/qASZVcgVcexOz4TvmZbc2ZHh9ZynDwl4zBd9VxjuddMdLL0ssWMOcVrstUJVpFwn
D/PZaGmvndeBIGIKoy01+lLSusvr+gEYIkaB61vi+saNrs2klP+Q7G9dBym/NhPEN8xV0EX2NJTW
MaKF00YOdoNJa1a51fkoXucbGgU/6lQl+l7+VkS2t3DCVIJK52EiHOFm5tCGEYsO/1oVla4lIvJj
XT77DAIiLWgRWpgsH04pGoRLDopu2+of4UZBpy8M08Fh8itPdtywM67Tc6ZW5i91ViR9PNHnYJJT
uWPtHXBwiXf6pNs5bRElEpmei8tLcH+406ZG4IHnzaQsjbkK9NiFguyZD7THN24ugsaCvkx4PGUU
Y+PjYavHFbJwMQdpqqoshag2P+EFPlm0rHuUCm2r+h36fo7YKdRJ3q/rZRDerjViJuqjrkcJi1Df
sehMG8ngRtObIsuwNWLNcUq32wqf+zC17//mlOPG5LmP6XKkaYVgU4pRJPm7NsOHsj6rKCkSM4un
9E6a8Ft0S5M/fkh8HYV7O4j2RMORt6WbasZEY6CrGUlV2Qn8E7zmNGXrO5XHCwgM7C8sd3cgI6zb
RxQgOq/EdRtb3yT8/j7pZCvD2NmoCw2QNp+xjhoYc5bcqCQ9WHSaCRC/WxmuZ1N4TfZNrg347uHt
vsPBBGSVuGsDKkcCB9b8OWVA3PlbPOn3y5+GzPdMwqUIrwFm1odJNrvcxHBCJSFbAP2Exr0lvMnA
i887fv5X5+O+YBbx1e2PXOd2RGhkYc/rPGKNoLpjydAEiqjniSlvUHXjCLWGuqmcrV95DEWfbEYU
vd09uhp5rUTyvY6a4hkqGFl/4FVs+DybvwPMorx7zBMy01ZR2gdn/SazL5wQdAudDEyz48HoOFnN
rdpBA8+fMpl+SpQjghjV/9j8kOFLVSRdJYje26O22Jl3QP+9SV+hu5UZBkwVrpscZDQb2KuYYhhw
/z6S5W6WEKrDwwE8qlSxSVarkAHOdvorrKsv4n/PolTRtROsvBtbR3ccqmVrDUtvPB4I2ugDakEh
3/smm+8Ns4ta108RU+w6Rixy9GRCVBaJY27+9Skps0fAN961ANMogUXhbNArjspsb5kAd4ko7pwR
84TrrdyIQdV4744mB6ZDdcGNVpS60PKG3JdWnwXK0rHpJmnAnNlsE/8nZgqvMKmyzfObELe/csRt
gAK/4/8n1yRnBUcLBMP9LVnrVhcQcv9t6uAsj1gbjNO+5e+RbB87yHY7sJxPC/aSbl8cPlvSc9K/
y/+iRF1joad7R6SWNPUxSjJenwdj5W6baaUy7ssGPlXk/MF9wYkDykKm9uOj+rcyKq4nb2qbT3tp
rc6uhYQyeLuAIAsLrgDE87of7Yp5hgyi6b5HdstqPwBZvrSzR/wWD9hxUghhCu8NIw9sc7FgtAAi
p9Cd+Tn92KHdxOivERqcXcurj+FAL57MhcBAIIc5CC1mpcibmP2zM+cuEJix5xIXujhd4AuoYkmi
t3nOagB1zviVtazFxOxWQkBguZh/CJSfuWyISL+IBHU5AKly2S0sFghg20B3RgqkIDfGuYx7nQMZ
jnZlmlBH68YWTPhEtY33huF6ID3B95H7FEdrMmD9pF5DHfs8yq7D27WZAVFRfMtlTcbpOz+4GVwI
fZf1o/9pJtMwrPKjVWDf5VOHoxBtvieyx4uwZUShaO2BBp+QDekiewxMtlwWKVi0ASO6snWqV8or
9RDq84cQ+ry/zNg/P31iStIK2HHSIdhMIubCIrD/dvoURa6vTVnBK3p35TcxTzxwbJeswvYMQ0MH
F6x53TlL5Riw3UBJJ2ngxW0EBQfcEp0Y3lSls3HUerp2nsIer8JSDK4IUgTqtIDJOIJcXSExh3PR
Q8cfH7QS6Szl3VquXeTf9h6ZhS4+AhvbQp6GRFGRS7M3m8eJqotdIz2hj5/qhe9v+fEWhRRbk6KF
5fey/0pSZpUrXD9/4YWUQho/B/hpOUb+9OL/uW9ZZAkymsuulEcoXB2+NDH+gABijcRah08zwlTH
wopT2Db+G44mLYkJEZ3qUdrJPhlxDr9ffddX7yZegemKZfEyJRL2+QRqGl5lTkgaab7zJDj7v2J+
ICdozj6VgBJi8aUo8bXrRDTxVk4VT6/+thk1F7JElgzoXvOVJ0Q6l57Eg+jHh3UnHXSbF97R5vtq
hTBPaZC9Gf318v7Tz1L+otAENBHXBMcvaPUgcxLFUaVTRjmGZ/LCNF6PTCdbi5RhN1yVyJJrlMOZ
lUoVF3W6ER2cfEWsIvc6W8KwpS33Mx6bCirOvUAkMmLxvPns43GJ1hzMS+brBmdwEPNnPO5NETDA
rNFFQSmQyIJ3SJp95FF4qQSyQ7RS15urBzCRnyzhkMUTX1/evdxn23ROMMk64cKoIr2eIPWBkPDC
aCt0m+l6WkZZ2tc/dIeNHjsiQmjNHQEWzRW/OM0jWEEQYh6ageVIF6E3rR83DPikVYvlnzyc6Kn9
AyWtra7DZj1BPKj5Pc281XOICMtU11hCRq3ZG2+LXk/ACkiVNqUoIAQSzExN6/mb+6HrvANRyCKX
WVKfr0aFbVi2RYJfmvbYBQgHhCSA1QWcLWTwZXH/1BcLJ50KOqwbM8qeHJQoIl1DEg+sLgIz5jfT
5BCUjOPC/rCggLFrfZnFGwILqpCkyTjdwMpXN03nLxalog+TDXk7pSHqDS0GjJhJOFcG6DjG/x2l
aI5Jt+1uJ6MvQwktofaaekv8IggtMNW38iAKk8H5gN+kQMpFprwoXsPdYlP0Hc8GLlvSLUu4w8Q3
tNr14z52LHQKCqouQAwYkFP73ZKKHI4QhFcaFPkAnXS3qYCo9SCVxaGFafTKUYewUKSHjmiP0n14
Y3RpdPybeL1/ykElHXihjZr3V1YX0eXGuc226OL8pfZOczCc/2DSRDIzNtFqda/Kcw99Kbxu4f5f
RaHCxLUjPvcl/u18LbN9pgxkMCBf3gcjUG23Buk+oLTA2Z7KCiOKOcDq2pAR6WUjcCoFjwZMTr4y
EViY3pN0uBf2oxhodzH6a1oNUMJWB1RF9smvBGNZlj+i81TyrYN8geN9uBVkvjnZUnxsxU+cxdrL
rCkllJ3EvIrIgXGaOt0sGk+zeCYQDCTVYv0njeM5mQXF64gjRy9IRUNv0ayDXdYyhc+y5Bc87qwv
AegRbANVbjaiTQQMyOlwwYWnGkWwHNOUSv3VlCCI2vukuze3DM89qyQPhYTCPmBmPSjIKN0QFlKx
5nZJjCmtUwSnvxgavJ4syn0gaalYKK7eq8Fj6j4hmzDIub/qY2wJInLtW31fP8ZmBe3CJ3l4sLmN
fE3pq7vAhBSVS3ULMtgPgMITf4f0aQNpSwpICIXWCrU4lfUcGYoWDmLWUiLgawvUuWoMQMdGbtl4
LMCtWXccxVwkGe4JOYLJKK+yMkOyAPfWIZmeGZk3bMuNmkFLLbF29aXmCDAn5FkoDN3pdDmmKWoK
VKtZ8ivvfrmIpTXKb/KK6r0tvOxeJ5Mfefvx4ax8X348nh6gdKN49kbbHePKQMl+K7V/h4vOhZk5
Ko9YAyZv3R0DUFEg+uG4317/H5DzKPJ7JrO2tI5ne43fkYODFyL1cCA23pvVUyjPh2DVXD2EHo91
L1kisfST7Nh9GsHDBYR2XWURcqy4H3hUWHC3AITI2VjaBFXWAZUgcbCPXvldP/JXG9cX6OvFCpOD
7yMx8yB/OxWG3Sz5PTCw3TrkmJCGB4Nj/QDMpUozV0wA4CDvuo1wwO91Z5qZaJPmglyIUgEeFZr+
/hOEJBlfTuYmlzTSHJE7EQd6jv67z+w53jr6tBSUkS0RRbUP8wJxWF9ciAs8AIyYEBV0DqPUJsVB
Da53bg18nzRyDH68L/yy0EeqvACmj1VgKMqBbNpoo/gHs90oMx5CbryQhFecFdhj1gyjGTE+rlUb
EnWR/07m3ECL/tZCyIevmcw8tDcaY+2xxtKC6FZJETanHSQTqruSV03SwYirsN/VKJvhTB4Jr6Iv
dTKh9dYTBkWgIge2R7Vqw9LsoPssOFMjkYf5xyAvunX1xfjASpS5IWMyopMU65WLb/bxlt9gkS/j
usSQPY+k0BaSNp+2kR2lDEgv/1K0wx4XEoJJ6TN28thSyWQLI7IcPTu9DRXRJHBwlX0oBMcg84GN
u/+8T3SooZaPjJg6pmQKax6YotQ1krFHlsTBwCcxo2lOPM/deeGGArGpK5GCradbFY1q54TcbDes
0f1C5XBngiMHBgC7zexLCMWctvbwppdGtDzQ1B6JQonpOGgh9wTosK3IU9E1zmXpoiyk+P7AwRNI
OJvuomIoPNTktd8WK82ICzFHQehNpN3WqTn8H7EchLaQx0N7XtR0/Y080U9ARwTmmvkdddCC1KsU
gXRV13brJ5i1YBh3JkidLyu/1id8enPXjuSUbXhyFu8Q0lIcytz+nFMVqGs0hyoCKU54jhxBnx/a
Q63V5fHG1PZDSQZN10CCwQqZ3HKLta5LiSNy5OKKa5sOQjsAAP20i+biKjuh4pTtYv7dRaC4dzOv
OmVu8f+4yDKqRhMeETxLJX80OXcbjQJNX5d3Hgl1UDbIAo0ppirNp8ZM4TbznN0zXUO6yse73/2m
HiUhRGRg4OSl0bJi/IH9qO9GpRGQy3ZWHuLETG8lYH8uaVx8W+5EFMYvUdN+irf6Id6ktnrQ8qEH
bsxfehlp4X011cmG6mz8UqD1h9Ih/xXVEw2LNGL+fROg/tbDxDIMletc8QQs00v+1XXsfqfQnFA5
PAUy3Bl1j2A3IK/qYTlTnAudsy36TXVYYjOP+opKxHKSdJ203/Om3iQUf6w/3N4jXVrZdmfqxRm+
FyBeCYNFLGgPoioRkW3/vgQ7+PWny8GSkFlv50qrXyzpQeHdCm2xAFpqC66g5QJIUKXPyNBOBX+H
D4LG8w6TBLGhVReDRLaZmPatefZfkvJHLOYKnxzr1h4jfxdrI/rYNFelELZ9hCYzsKtetRNSD8D0
aaHPkNMCj1tsl8qE9+t2aNfTYEs5nAdhjBOxAKOvqmLoYl1loc4Se3q4WDKDQFQr2zYzKz/M7Omu
kRlpOhxsxV/lBZl1xy/uTYY4h5BLaYPk99hUdypMpV5EzjvZ7c1UUyMP/DfNXfB1G4QSTa0aCQqq
aWprcenvBljdpXVxD6jTcXNaEaNeDqtwv0A4Bri/niKGK6mIqLcz2xeKm50Lb6FI0obulI527b1a
gYGBVUy2exVovj661StPrS1J+ECfc5JM+Ux/WChES7SbU9om0KJrMdi8kavTtOORv+Hb11LF+3/9
BrceXyw3A4Hr5isutF/UZNW9wLmTvhbPhx73ya1VVQ8Rt9zf4dGTaErSQf7iuBoFKjNSyByF4WVa
HwVaivIv2gJ4VHmZ/G4ODbOwOG9yKbdmXokIU+Bi2r4Zyi8MTZ/q4TiX0sp9CTallnUnEF9CLpov
FNpBBKAl8DXV4zc/H2GrldGbHuFkZ9sA/bkUb6imxR8b8425NbujaHTxLTKLLe1tsUiNo5D1N/u2
Z0zk/ixadNHLkuoGrgHXWWw7rZLk/hSunOnLBSZXyiXqbQszaK6npegzbKMB2DcmnlF2aEVVGydn
HHqKFDXN/iuljoql8+Z2PdFRWBrQVIMnjSNvl2wLuFOhpFCkW9ag63FE+fpWE03P9YuGjriH+Dm7
0dVTdvv80mvXTgss4xLmg8cjuxs8xx4180JRHdJ8qbCZb0rRfgCclZvlgm5S7JA0sdyWzG94fEkE
VeI+aZ+xWX4YIpICm+xRAMkNEywBwrki/sHdqsXKW4lMpEx+obe/9kJTfm5UT/y6I3tnlqABeiuP
BVo+bEN+s/3L6GDK7tz3nZSh0I/zaOSvUH79+Xehiv5W5u9gib1aE2CpXcbywmqUtX6G3PZDWunS
sLDAwgdGxSOM2jRS8G3iOdM5f8i7MnLVgCFXZ64Or+0QBotfBOLRUMGwDkL7qN/bP3ZCZ7u8X+e0
oT3dA9ijYWHESaq9xpvgQYsDYPFx2snxFxxSb2Ra1IRqjg4sIllmUPcsyf8tWlLX04TAeRMEjETc
WedlcVEGHKY3cWGol0z9Lbd10l/KHPnoIa/fIQEQF5KCAzj14YHSmecPsNQ0Cajhwj787iVy5YWa
Cq2CKxdLlL+SqcYJ1Z8yjWo5cCJp2znoNcyUK8pWVMW66oKpyBY7KqzoXdFUbswfwudnQG8KEHIL
uAkTH/6QBWUU/qOw7LAJPOiz4Tp44Sl5tyEVQs3Fu2eR/kRyADn9M2TxvVJ7eWVheCtFB7YMFX+7
aKaWdp4InKcRVQwA7rGxAyNzwxfgDeRglQmcTRC+8vVT/SAOGJex5ItzTHKIG8gYlYhIrB8L5n2I
ii64NB9SsFpkCp9qtKuYOOVI33dLZ4b0BuPfW3t6yHmvmPTwhjXhshUIPCw0+WL8NI2pMDUPx+nQ
EFqmfwFf/sokKs5LGp2DnFLznhRBDLSXMkAD0ATQujBOMKrHEoFtd3pn8/CWTyd8T+3t7+SkuBBY
672TxNgRGhkIUba2u01b076SmSeQY2Y23fYsQskM2KAHAHv1hIaXZwzVix/0N2CV4lcEKKr6DXzP
pUVhWiVfcCuIRRjMHzZGVEGaabwQBqJTw7V83NB8K4sYFqvjS+pf5fmWh8iUsUfJq9in5EyqDw4h
D/iPbzleRMYFZ4dQpW5O2rrQPbXAsDVQ/QWYgCX2H2UmfMwV7L4hNJl+sbjT27xQ3lJCQUcU9fhy
otn3cVnosGg4RrWY9SdJSPr9fl/UagvQ/wonU7EQ/fn+UtnLVOqh6SlYcBafu9/zWHQJN/YtIrEm
JjvvBRbhpJ5ahdHTbulvV4vvnkrZ3xekTspAsplu1aR9Lg45ezc4mZf0aGplm+pEqVQYncgbTPS8
zqScIzOuFTsq8ytgSp58EeZls3ysz3yv+3Qc6jFQrzLWyq48qEFvJsg2kfhhYe0yxC4Gy/kAqu9G
F3xlKmy1SvBs6qWzilBZiqGN98Qiw0zJgOlC6W59VXTs8swU4w1D//Dxk6YgfbU/EFP+TNoudHd2
UEcbDF3IQCnron9L5hlkNBaZMkVvhRR6EvXeLBZ71Hdu/XgcKJKCbxcD5Xs9XozsOLA4453Ak04u
nrjhUSYNsC8neFOy40FRM0pTv+0bNhKF3wKyKh23j8Q4IBu7zgC2O6FZ6/0V1rHzur+vBiRxR90k
vLPPWCNEaDyDdi4lpCQGpRIMciS0t77g3PVJBy+4CKOG65Dv7h0KThtgWh9ZoaagLE44wEXZrldH
efmNI5rK8/2CH/9oLiJfFyvFMs2/MNkzXwpLjiVewW5GePkUqDGXSXvFvTiX164eHn8UZlOCH00O
pRggAD50iDHv8b7xR4nVXtXTP/wGp8DSfbpC5eUG+7YNhAeDRtBHshtWIJuHAufcUtA6Wcb4CSUI
BRFlQljX+j2hLbo4xVw2cuHlJzCcfj+2y6OtVyw+EL/pI/MU8Djcf2UabzyxvX/7bHo5aQg8M3Xf
uZp8Uix1LntaWNwIrjR3MUtL8c/kAK1hJFcdO9wGcXzkrN9xEeoUM1RLYtzKzy/oaZcqXHaZ8twK
Ckiq8bdkTzVwmvz+ZmocuzKZ8YSj+y+yd8fDoGC/yqfkJbi4HnOgrT8XcN7hyz8LEWtFsbY479DA
rz4kNJX9bPKK9xnaw+i4sPuEOwH6Jg8MLJS/w6qe5QAybiWrLFgTn+KBG9oey/Mci/43s5T0qiVF
dwrGIoZYFrjrHLrB01Lwjc7uWbUWtIGIvZKwJH3F6L+5eKQlKpoR74H9XHaCra+O9HSrBdzj8e6Q
FvBvSUvxj1fIBON97TbxC6aez8qDdDiHr6ciDYYasVoRAMi7Vq6We9T4Kc3APgTveiwJ8CZCAeLb
sNMj0dlwBUjlxZS8bbXOn9RvTOz8G7+Hsy306fHGt0Tw2Rrc6rxgzxPVFI7jQScyTOvxbiZzKkYn
lS9PkVwuDl55R9oLjRb591Lw0TpOdi31syjD9GSGyhUHllNl8MQnaO7+E4T9GEXFEShSFNCZpBB6
Kb86Qji8c1dXMW1m5fRpxdJVnPdeG/jwKHEraA4IKvGN8vOEtrOYNrXu4blwuYWNWU2PVhPpDGi4
cg6kiBCleND9HEj21dVpwCLIOKV9zVPV+Zuz35gUiEnoFPfLt5oj2rpVNRfNkLcpGGX82OIdgiP6
zJm1juFZJPAk8NH4PnoSYzgC5Jo1RDzzzpPrgCs49rOiN8C1+FPsSo6RfJG15zNWsWYt2OuV2yXV
jX+T18atBjYgZOUzaTjtT3v9KUTbxayGU+XrqGqT9LJFeg+QmybTQKmlFGJkMkoX6e3rq+J35F5p
zdLPIy1rRhHzaRifuGdJcYBwgneqmvQCJuOY0EeNlpT57etaKHoYnfH70uX5O1GYbH5rJlYF9CsB
D0zpqv71ObodP/dc/Kn0H4QCCbBsoBbRvZssggnipf+ZSgf7B+3hGHUL8U7X1MvZc90s6dYE1hxu
wYQ4spI9eHb/ccajpA7X37SdCskD5KJBo4L7Q6MnEIcpMVLiHAmQi4A5w2GmEDYqpllH0hCfSbjm
p29+kHoZ2of7MWjTuDN6VaktU+qKEydxCtKNIod1vEC5JXHrgE5YxboMzr6CujBSJUyh0/YslNcy
wM4gltFRO8kow8hS54rPigAJKfGQ7y5BHDQhjBHlMZZjg5LcTkmL8J5TIo4rtQTeiT/LByTt9pKv
bsU2rK80jYk6nU4yiPmYgr4Pz5wSyYcR6kDJ7sqjSA0mNcpwScwuKyWzW47RL09vPOpv0+4O+XRB
HB+95g7UsKf4zuI6z8hTJX+ZK+o/2OiMzfkM+AtddZB7Cjd8di0JkZvCWtuBSnXnKGV8/zlBNhNE
B6rp1buRgBedsjFWgjq1IvqxRsvwKngXAgO7ge1kLa76w387tB+rfwVH7sAeXBj8nhS9BQjarpij
e14T6tA8R4vMO71k4/DWSOcYrEAuBU4jLtDugVGQvHIaMxpiGzl6BOsIbgEg5GqcGULxzaeMQ4Ty
V31qhxsDJ1k1yR1nWNL4fjQPuauFXTnxwvcAy4taInjN72D/ZI6kZJht6snwqw/JaSaBNjq6Y5Bu
+0zz0Yd9zeWIz5aIZbT/SgbzWuuLUrrP467y+YN2CuvkEcGMhQFGUAmPgI1aWyVXPBNbIV62ofF3
uu2JQ16ikyr8xzSLkjXu8Zrg7ad5rLMkQ9VqkjKluqTWMGkE9k9thmB+Z5HwHV0vfg9DdFNj9dEf
XOJH37MLJohG9H0uUzUMB++8b9lNehhW56lJclw+tyThdl4aPD3yJGK5otQsjYy0ksVj37/YeVL3
DZsINjI9OpEnN4kOwc/P+HextqA8qJvS/SigXiObOBZ7w7lrmJQWzWprvaP592znTRydpba4zGNs
zdobqocaXNk8H+TBQX+MnI0aAZNPisF+EAN5HkSbQSeOuAiarnQG/TeWxWgFJp/TzxwyNqJ6vBUE
JWzvaqVYJu+PU8xSi+v5kK1Ybjmpqx8G5AH4VpVDCwxVztRzqydLm3VmkYbK3XqfpkVvxn32WTPI
CaOYP/UMgNeSgdMkFoshLEOvnCwpl6B8QYxIJ+tjbkQOUk47yuYsyhlkcLBcXOb20lfbMZULagGA
oqaUvsbjzqT+8uXP/8lWc9AVBHBM24WM+LVjG+Epytz0fESje+1tMG8H8o9mT65Sr4cSnMuXimem
7fyL9Aj8kz3YQsmFml9ditSjoVuv1crorjDprmxn00m0NEAJa9xx8bAIq0a8R5lW+6wyiMtiVAzP
AxnbmaS215K9tlNKhRrchjgqpbQFEXfi0t47cQCRR0gTdmOdg8hlb1wNFtEbrcW0+CfMTAjizEtu
s97Jm6AQzbA/Yz4+fM5STIfN3LKl1a0W5NPLpV8u5JshRRiPjQusjbzP7qrk8wBM2muKi0nBiZ2Q
pABMLNLWJz7jlTLicegcDZA3YLTSS8ayQlac6FeFpzSRpP7x5HuyV/RYZxalY9tVpkW7DT+Qtto5
UoT6CTLsP5A7uqQSyYQngYUZdlQ67fPpXhjtxmPGbG7UYdMyCZ7GLrvKtx/erQZjg4UORRYJG6v2
BobDVsNCQeSU2C/oGLiJRaHLaDbVNrUMGtoFuR5ehYU2XUMDev7a7/FgBU0nAF9UyvLhlzAU3Yai
jAS11RIAvfmKGiJIZ9zH6EToCNyEA7pGWDO0CwwQ/vjzgg1NHy8lSaPnQ65hvfHzA/kmsiXnJfhi
+LO1SBkUbd6D6vqmTTUZaNQh373UXN6jaTuHdyAXOsoDRhncRtj+2ZgiNTOHVuL//hSguZ41bSIR
l8iK6XCeGR1hXoJHOJtnPH26EKBrRIbH+qiOgTAEpqlgGT36aE0DisJgY6CwXYhKG8MOU/MRjAiG
KHmSZFplnJE2jIJzPa0rfSIJKhaW2T6ZAjkgA2+vx7ZNh31/71+b4kO9UGT8eyxl3nmBkK9NmTnl
gg81oOj9sBcNWD4FqS079S2uIaff0hjCqkerlcgcpHDYtiOZ4YGsKvce6//kF7haR6io97pEeKjP
JyWsaLUfjjTl+NhH12kGneCGdL1TrH7l85lQJSO3GCc1ggjwPb3au6ysYWp784khVDHIbmJlLCWY
7GgL+YgI2t+O1mkQu261kjRQS/f/AqPoCg9rIXg9MfX5tgLL51XTvHMD90Q6u+Db2ePHWl/mgCJa
cx/Uyh+AwuiB/DDjAPsvy6dB/+vLwMpJLwOqnpxe9CblDOCMCNX5sWmzAJcYURpEd+rIiKu8ex47
UvjxgrdCcz2IcKg3cOIpEqXWDdUIAbY/Yk8yfTVx0ydmN7fO40Q+PKvZbpsPk3PNxesdZ5xg3HqW
4EV0jzSQAsGTGSsqfafEu4j9t+XMYgSq8rwiovtYW+KNKQ3TQEWuIxI/6B1JKwOxaRHC8vNZtXng
yUji7/6GrolSqUAHWU+jpG+lEGJIyA==
`protect end_protected
