`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10832)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/Y3
LeD+qw2K3LM++tksXDWlRgF/znF+Jw9c2JQAPXKM9TKRvOl/czmCOhE3aNSoCh1FUwlKG7QK7XW5
1i+Y/6fuS/CW01hotPrez34/+2hYr87se6GBDorysLqVAXMsLY/YV9B7HhDUSw8jyNyknIEmI3U7
WudHo8vhLWlCkMQkDcMf+Ivoy8TEGZRjbwDtOXoE24Tpyh0y7Szqp8vQqEDariMqKoVn6oTmJYLq
2DpWhIEswln6tRI/+zBSleCqwfAdmXyYA/Icw782kOJqC1rm3rVrW/fPVK8K9QJVLjxlLtCOUsdW
MXHfW8zBcf+OJ6M5Ps5WfxcGaSo9F93JhZJwtp16qQc943Z5uL5S7F6uhx2/2/JNEiZKR4nwO6YF
9lApKneiqiV4lMknv2GfPf3Z0yt/epCJ1D6rwzHUxOS1WE+QGHCe4rtK8iJJPU8gdqWBAV0E38zX
DrRSC8OcTDpaHRsM4h45UtUZ7QHuncOnjyjfle45UXlGJHuJmqtQtKoBHlkWLaWs8IxPTRJdashu
kUk0S37b7qinz8QPzVNDizIo7tt1mrqBCLYTAlFjqwSpg+Q2GoQNpEbhhjJSmvYKPuGddRJZO7Wl
OSphxyLgZzVvmxDSH/t87kHgGHsFgjp9dviohojl/U/zWNmgRey6ALjcz02ZkQE6vzh/zBsU36oI
1XLzZdPOsmsFTW+hi0YtW4QXrws+XJn0lDvqAm7a/4zSUan/YXPqgWJAp0UJnu6AAEQbDjLTTbka
rmLtzTc+KBM7Qh/MrR0nLXOt+vB6+4vpyFW6VF57FxmXcsdwTMv34b7IGNAHXV19xTd61xcwO0FS
hYiDkPuuZYyI4HEIp4JXLUgW5zvyHVNvmOFASRRNUBRiTkDYHnHp7Z/O4tBKX1n17fF6v/fg3mwS
2JeiK4If3PXvktkxXJaPGyiZmPmt5A4Bthy7HLbet//JHNLV38xyJ74gKq7QU9oEASiPXGEAhbM/
x9I7SkQ7MIJFc8uqyxac3MnFNurIiDEeYdHyaMERPao3PN6xhb/2oFOdOfTFP1ukLGNEUsk0hPd1
LgkUtfW5A20Gbm2UqEhuCsZlhhN713pRuj/0GuH8RmIBQvAjd/LXyOWfuP01wImCTKOjz7332xEc
vYTB2ZLyx0dZNiESt3YthzquQ30BRv2JZ/yMS2L3RICN8EY6volLZIQ9J/ZWNZnto43SN9PZ1A4d
KcVhHcitoNxEjWlorIlUHZeWcgjrKzRKTms/5Qvq+XK9VFq4xnGh7Oac9iup4UOYCOq/mhqKA4j2
JlpoYNdiV2q/qk1GYiR9lF2o5Ecimhm4F6Qr/f/9tQ8wUUD6qfkiHSEpOGq0Z+43W/6hQ3pmdtRH
CP6CKYahbYpyAC5P664kR3KSyU3BSn/mcTnKBa/6NWGyfV/dwudwQZYVTSGWPphViyNhg4NXBZdW
VpNjfiNyjHV/WD/NL12VW2Cc1vUJznM7Ohc7WOPoxL3rTVqMbdkgPi1PL7rVXfy3t8gZU9LEOkRW
PzJtI3ekd0GtH6hpTLnCd4KmXpUwUPsqehrqFsbkKH7YNuki4EFBpsExEHrPqDWOzpH/kcA6Kdrc
YH3a3yqe7rPGOTbbq8kMXtkWN+YItZVlgy9BxRaEYkXkPwPE5k9IeceOrVP1c98Iv+echFZLGGt9
j0QBJm/V8zqFl/WSHqF+eE2suXsp689eqNMH9JYhg2llYDoxhhS7WHFNPfDyoEWMj1/FlOG8ECsl
8hbPn81Rxh9ZGPDmnWU1rLYxp70uYzLoDW9knjjlU7YCZd0swAJvYRhXsXf3VpO1kz3iv6W+nZMX
Brg1+/LfOSXBphl/YIzzMLzLBGrPVYuVX6U60QduJlfeyJj/jsupLa0YCq10Y7+A2WSQXESFHfnp
Oo1bNau5NhQE2DlB0tGBKT9+EPIslfIrUiX61m6Dkfx7lrqNHGsqror8LWJv4D6YsANdMsKop3y8
ywyUOABWxCDeC4c0Mvj7ZXbQ7mSXzmcBcrunwbWP74A7PloqWvI7iteJV7lKc7ctjR9u2w96DihV
W/DwvdUVHlOVlxCx01PJRop9W1LKbTZpY/0ZzTe7UocPsy/89bc9AcwM4aV8BP8oa3Tq0MJrZOMO
mP8yNtdJbBItrltMSYPKOFrGF8h5Z9v2p0WPw/sstYnkE2z48Rw+6hSemnVMd0wzek9T/E1AS1oE
ZrA3f8QL4jIonmJyBqQNSc2KVR9ezwV6djyk6MGEmqbDiHCADFai9EZ365ggEep82nSHyOwH7e7k
WAk5TUhv+Z/kHNdp52dLfVakxOtEHSbneCdm8hkeGJ7HytHDkfG0EsgZqwM5A1W/2scrmPjhfeMq
Z5gZil+FLHuqDgpnlqk6GwlHJoOLR6TnOa32UQ4VybJP9TMmBagp/su2C8/eaMBKHBuRVk39v7FX
8dhO0ZLg26Y43Dp/r3gPiA1p/bUv+HokNtQflnLHrnfgcNwAFuo4ChGQr1suF+/6MEZ39+YYcLQX
aZIHry63MB6k2POVKN1jUp6i5HvsZkxmE+SYqfeSDdTzqzoy3kdlF3NsS9UON2EiPWysa2Qu1opo
tMApEFghS37Yp1yaPg80jFeZRC2laiYChE9ZVjVUsteBxyUf277ypkGtcghPr72TPqQ1zQtbODEV
01nBZ4KzeBhaYwC0n8+Xh271Ug+NcvgaVLmitcZexDBHRfooei8SXKptlrX0Oj+5f74mAi29Jmga
Yl+J4Ze7y68N+bzIJgr5GmTFfbhcQWOQtM+BOeiDagj3eW0qeSPaLziyW5Otu/hbEIob2UQETk1p
onrFt1MwZK1hw3fcZGOjClWT219Jhfuyy3lsb9z/1Y0t7kkhyoXH0NKDKRuDurkJ0bKhY+0GCyGQ
H38L1GYASu7gN5ku/Zk7VkFeHIldz1l6oisOIKm7UGg0hicb5B93f2Pf12QemWqxMQgJ63mSrLMV
boU5NveNGoLsYDtDnaV2YNF+CNcyA/sJMBZrLAgN/9Y9uAUXs3U4HPLd5x0+voXUhAbX4JvYJBIt
lCVF1LiQZRVoZ0CoPFcTPy0oqZf5t/B0waoz6o3QOXzVHLjS+SJmInj4IqzXOmBxM6t77U7imk18
bLYCgkajPq5Q2BsG42RmIsu+QPpn0N4hg+BdsyTRZhPEP6EAVaqRoVBNIdfJ8gn+tTTv+OCdZ0fP
wJmNdiPolTNcs6vK9TbANpZeWuI7a6qtgKNBsOCOdc0zhjb/RF52S1BKEBqc42VuGhh6X5yU2mGb
ruL1Fd0poo8hfojdBetT9uzutJqvFkx+1xuUUrZIfuYOY3VMlY5n6iS6tCuK8VerRYRMRQ1w3ZNW
TjZmBq0MOs3B64bLdjcA+Cb5wKYCtVDrfS1jPXCYnY11vEYxa0lbOLvnd2vLtQkTwluYDygDt8eR
Vy7ZGhDBf2KaHmfrIu3ziboSQ5DFEaJ/98YCNZiiNFKkMhf7LI4MzhlYsZmfTO1rnyW2+tHTEJNb
Vm1wWgpcmdwKzr0Rhxk2Uwp4Zs1oWRzaqP4vwoV5uNojWi7ExhmzYYWzIveKtpRYPtLHtGkExIHu
Qz+oMGppLj467koDLAp+7/pEV2YTdWBgRVZ5iYmLY3GJh2kJ2Juu+zZSQNHTkft3UKzR68NQ1zLM
n7jcGITc7aluViR5H6+//SM/bGsG4Kvy+2V8oyxGP2E3x/nFEXbTCAxAgLNHL61UaSx0ds+Ez5ys
i6/XJM0O9VvqCv7JSMnSO10V8NHMcurN3FMnRYAg+lWXYyw0oxuj1yPd6PBQbWkbilgoKahUtsGf
6EOJgVwqxprcGaVbDnvF1JRFyOCKl43mX3qrXy8zJKDu411YmcxHi3Bk8y2aKoHDRL3W5UlIZgNT
CMCQ5BRuLSUR26i3PRMpgJKRkKQxUmProV8N2At+xoa//NDwolylAs8vvDaZPdc09NwR8KIuPY+i
IXcXws1G7j+ILMONmJDFTJue/N5eaoFUAr/wOclOdmgc/rtrmF4Ty79+4+psIMaaWMFgQpnky0M5
KzhfxG2y7rGbtb8p1pXn8EU1BPZ8mkW7DEob30CYyRZUFaYbOO/r5Hy3+b+PyyCTyktwYpAFnSZc
HYHmYnlWiD81t7b/W/1UopwVzpOchGItDRFfubFBl8vtkZHcAzS6DPnply6Q9MziLsweBzycLBVo
GI/OJpsCMtI1pzRDihZ9BAjXT+G/gLks9pRWEXOLI3n2Pz7N0WIZeA40ad+WAsq4LMk5x+l4iqtP
HK4oN/x6a5ava+CFXTRPIMD/kSNu4Eu8nqwP6Xio+DvOqie83kPnyG22o/Tc8uCNLF9aAcpQob+B
25b+QcWTQsINxzFVXuEE5CMn9r8laPVjGpwu3fCSfUVLvE3YP4cVmxsdg6+Ken3i3jJbniLSUOg1
07A+m+TUgVNYEhTMzS3NBVIBK/zRYEqh3C0bAlffm8a2Zg2NdUVxEkt06LmK6+5FVEpIpruyiJox
QmHl9G+aiJP+WQKsJsZPLjo087QDRIpBP+eRKs/51DwzVc/Z3llXxakQVx/3FFOuJP9aozd/0JRN
4thG2HGr9IvTj52/RO+PiDCDV4CY+OCWdUxYSIVRdka3pCYV1SLF+P3MtQlto7TjDtFUIeGBHr4X
eeVzIfwrcmPqIRv7h5nKfi39Bn7LzZmOyMw9qJ8h2mfu9QFvacSjY7A+y8yMEWu/gps35aeppoC5
k7AVTmKrVeN+zvSv4pOlot3IWu+XC5G1ondOW65X5107ehRsWMbUf+f1ZqaeXT5Df3u+HP/YDD6K
1zVdTW72P1jBFDYCx/R8JRfVk/M1GrFaM30Gd7WAb6N6tlW8lx0r+OMsoJnFtCL5LEGPZw1IC/ND
TelVI6YHOQU/hAa+rb5+08bg78IUvlNNJVlZEpSujUMH/G7Dve5dPC9wkP6fy/gc+LjgZTh9nZGO
tb1jw5/bEYPXFTk3L3dIS0NYRYkQd/1vkyyUTa31CJHVI1rcOrgGfYRr4hZjdjppwLRLtzlSzzJK
JplGO9CMimZeHRo5jbxvBT7Lz5H64ZJMOaEz8Tl3Ic3rFecWLgVns+A+NiO7P9YkGCRQLQ3moyZk
voCSbKJSPm4Kx1XO2e0VjYy5ZKCkT4oLlg5wcQb9BCxOzBN3GPL8aMsxqGz5ne4TEEMnlpOL15vB
WAfwaJecivPYKiDv3BAhmQpzyRSPjxLKtfyQjCmZvDCdDgJEgf82evIrZmLF1iS6EpHQb+qmdd8b
MzvjiDXCcd25+/ClS4UIFi3We50726hVvHz205fw7ypSCfycy8KwgPKe0vddYzFEez2h/qCn7xVx
Wx7/YBPH96PKaiD35ZTEWaExvpDDHuaAApHMzl5OSDvQwgwW3wE0J1bBy6vCsEWJqduIP5fCx2BJ
yRpqLoUMpmP7ge2wNVw6lX8fN6Bakejbx6puGrrA9j3jLhWzw2hXWSTRsIlDznTWG4T3xTudfhQX
E8BqBrB7ZF5uzietyzkwwkOP3HSavcU5NpaBnL45QqtQ9wW+YRfBli9J72QwS16YguL6CW76dHvi
pbR3h3QHQnEoULDl0M5ulNSgQAgu/Fr7Tz0xOz/Zs/rjClCqTpK/GMJG35uBZdTmYx7vusJGU0Lb
9+/tZcsW23zVJN0kh9qL0MQlcf6LrK410CHAGVagZ6PMp3XnWNBUOwta/2moXBG8qnv2ZBMAgsH3
s62ZGKf1D/6tggwiPpveaVxHebP4Mou1Wh6f1tu53YjPwDflJoGYn/f07MIeafix7Lxgxagr/FIc
eBTX1yq7EDq/y4ymEW+0BWzEyRpGpYDQIAH0d+oKAghBjVD9SApT0pYXY8jtusfeRFXQrtgNAv/w
fpErcHnLUyMhIUZi+oC07tAEMzyS4FddDNYNSEgipEGUFWxBTZMEH3J2HtBgPKxDUJMUZYYAL55F
P+8iba0ZCvLqlrWdjx46cCrhEn/11/DOHiQWe5Z0Ywo0+6IjGM8q8ecYbdVbXnKowfrsKwHvx35f
Fs24cJqAHlPaUZ4kvOLl1nynYOkHOIbDgczW9Y8g1nKs9/gsWDSGEZTuL4g3oz40XnpS97A2Kydc
fuy3FlPBh4/dJbKnFuzP4C3M7URSJj12uDvfMjV5wjwnWbWWELNjHGsnQsvJTLcZHYjyHJJh5ObW
w9hLQFYsePGyzSahCw73IIrczkA6WAwLxNxFQIwp3fFwRzQ+vTxZKdWZvTW6sqy/e/bbcBXMS+F1
KSFDAjU7sLUHaLDzDQoF6AEafv7HsRhSH4XynnXupuzp2mUP2FoSJOxoUVJqyDEq8D+IpTtLlOc/
ukKUsrZSEiJmm4CFecdwy8uodSSSlk8W2wN3RMNSY294+g1rYCfXpt2Paf6M2EBnOP1TV+vLGVpJ
jKnPZdg/RX+NFalEMS22Z5p/LDpmRrA4WwYAQUrZHsLGih82Pch+vzuaDM/iBDzV4GhesxuCJl+D
ak/xy92aU/v5zGonqKVBtm4bGERUnvHXWzy6Vv+F7xhA2b5KYjh/h1Fhc2G4+f2/ZMQ2MqwMJlda
dNzgK5UA5jYklaVFb0ShTJtaAFFp6wv1ZsinDxoD+X5Tx62+CGiE7Kq5jIc5caKJji1KlGfY+6mE
iDce6Jk60WhP9hkhw5gPQqXsvH5LDqjSiWXywcJjayGNUzAAHcGyas0U+aCrLILpxumNU8ZXZWVo
rBMICw+z/zXTKbzlSL74Ct4jKvq0QUUn2Glq4P5HKrcU4SIIMPHfrQGHkeKOPlyeQbprjmA8PoGx
zV+tvL5CGkKfjihWvzSqz+j8BKCTAm0ki9vGa2oHt1Nj9x4J2soUJzZM8/W4qDcvnAFDikCrVaDY
76RXxPP/AfcVtHXKZgRmZeIZcuaiGqfpU+4rJ4ZEPLJJ+qLDnBImvHq+913EKaEo/+FTHID/Ia7q
hK17QUETUoM+IMdbRHLA1Tk1jI4ZQjkATQYE7UjFlOSNVpWjESP6NoaSB69+3ZezgjJZkBTc41pL
KY/EbBvA9mp/eYcEa3tbu3ukiUhwqNrYfpsufinQNhWcQuU5l0580L4HzQwwlnfTEzK0ajT1Fliu
4oT0KVQVGPbmSoGVVWNTr2gOoXelYey8KM2/y8RIbBQdLKbDffUHW4sFGTl/wFbIB9FAqhX0xqnz
b1W8IZjBo9DA8mg9ZiVhZAr5Fd93hrCKG+aunKRUdwf1MBgl/02TFGI7XaXPeQ9HvxNtzVkIsD2w
Y8+12sDBYH+USqK+AM0DAXWgyZHQoc8EytHTeGHU7/JWByZ1meyTK88SPerIMtl5aD1dN1OD7Tu+
ZnXiVwU5QRuGGdTxwUvk4i+DA3F8OHa+Xyix4lhr+964U3K1juJZ0oIYu/snDOtRXXVvjoZeU3gz
LZaY2AnViQZPhl4WXftxIY69qxKE3t3M7OlvLZWHm3b+yGIgrDniM4AAEpxRNGvZVUUqUuz2ubta
7BwjzIuPXCwAPw9qaptLzF1n+1IlTK7baH3x7KXzo86jZDbwm/3AB4bxK9XrO+/TGhh9hKRRxzlF
aVEALyD1AYww/jLfyOMYpVV2nMjzh4lAdzkiVYX2FxrVcWffALEG9liCdAtVZsaaZth1wnRQdNNt
NldF6LHnoCRkjx1vK5M0vFPNTDhIDvE5fhFeT4ddYBQtJ1fouWkewpjxkMaqM3q0hsYz+AOdEG+q
a7C2snPOuWLfD/W2DEOyaSpKAf0CiGP5/Pgg9V3P5xRySYp9N324emjwI0rEn1LaNGZg37//Z9sp
Lnn7aIRGQwsmylukVf5XSx5WSzQOC+JoUAYf4ieSgEWCPKaLQ6PQ/RUHQt3TW2DywcsF+9KH4fOP
24XfnfYfwQA3YzNdl+BmYI1/xZZ/5BGWb+AXIaqA0T1kCajytZ/Xh4NDer1y/f3xiO0ySux/WgeR
MoF5S7nXhplMZPAMOKhPLkXjEgN6hj3QEJ3rxl2vvednibOrmiuER1IivdT0R8b9yYfzqZEKDtsZ
4dSZH0kWp+cXsLxm+PQMQN7//ZoObT1HTMYM80bvriju2tEIN+IebmKDnsjF2nGbf30DZreNX3ct
aliJW8h5fEaxDJUeB5+PdjKyBOwFw3ZfyXqW4eV8C5b/nVqyD5dAoO9qgIwGA60idAeACuIpybpR
PB5XBBv6An7IsKr4WdpE49U/Lbht64wGmRER6Dc5v9+BMTImxY+SlFdEgFRvev32Dn/NTXf1TXtX
YYowfLAq6LafhEjAxT2KDez3yNiextXOSuTUbdJX4VlgLupqtfYZ5ZAt+Mc/+5YAxK17BUu1EU8J
BHjPCQHfxn0NRhRrI7exP9EFr94ZGyCmSYAAJ6r9qsCBNJ/uyg6USGyz9ntKYk7AxdEIk48PbawO
fjQ/I/P8ZT4hSnvt6uAyYszLuEpNH1OA+q/khWkPj9Ccy5BwglpVurD041ScuaWf91bTC9OOyBXP
S6LV0I6/8APlwm6U2G3f/OfE6L3DMeqQgMNHTym7wVhZZZXMwcs/fThR695ejFRbrK7ngfdgkMX4
D6uz3Exuel7/w/rmmnww2LI0TKJjPzxXjpIgqvb2hACxk2IGT+rjMSMYVUqIDEweMe2BONgsWq6F
XZTDq9kyMOvRY0vthtTVqARi6JXFIrs0QubaNAr0HjZ3UxJu2vBQTUomKZ8g+y9VzJaI1DUxeaXV
WhPR3mrVQsVFLPRjHyBQG9S9Gc5llS9BZpPVDSoHKmbVr2QaEHevMggHPDLO17d61cPN/wIBP9Qm
/e21kri1z/2YjZgfQe81i/MUXqMMwDnn9rohk35J8DbmsMSxJ5R3djVeA1yZSdlZt0sG4j5j0xo9
CjzMxUbUe/R7U/dwAoMbc2WJ1Q9dI7NEe1wuhko0yVIIBUdcg1BxqY6kWNv2RG3bBes/huQ5sM7p
imtuTfoR2XlBVASXHoFxzd7wrqVw2ZwPQoP/BPJMJ6UQan3a87oJCKEvO33q4jlz1kmxsc3/vfvd
ExqEqlPjto9aa4HftZSr3Eiif1R6cGY+3G4mRYKDrYWbRo1XJML9hK8lg6NQbyZfXubUidc4a9RL
sVN47fdA/IBJYQAjA5XA+rKoBIhB0vrQlxqSUsHfQv/jAhhs0iQgEWmknjkCxCfCiUkvn74NPseJ
pMyvdyEmKxKLADXY9Us54vyHcLoorRQu2CPgv3G82EJrgRZL14ulDfNIz2FAOARENNbH8u6Fch85
412T2DjmxSEWN340RO3eoXiKlXd7ErUYg8WxULK3HhN4bU0US94CxnkPhX+tcVC+K4lLlO8AAy91
iT4MzQzrFDZWZvWeF5MvBJut3LCleR9zFyBfWoVgM1i6Ux+iaApWBvUKJKhtPmu3s8egwDOg/chQ
7azwoDxbB3kQhJovJAsmHuWscz27Ss61BtHG6sFxiqWsdl4rumJDnE9EY3r5T//KanH0S29BDvgR
BWVLCVrEKSlGKs1ZOEYfaYt/j0OqI9CleuU2lpFT0dRFyCbnLWYPX5Fyu59EOEDwqHWXrXZ3zMhU
FRPZZjnmDDPPXuQQw1bWiU7aZAtl0Ca4mV68RwvOPK3dQAkAf31/H5UF74N4CrZ2oqw+15kKp2Zw
bTPtcQjtfDVBQhxxw3aixHFNqhtj2Ig01+vuzlk1zWniwFJTup8Dmx39u9Kn/+ZJNIWFo40rAVqX
Fn8yksKs6zpTB7GJLjAXyc+1zg7msDWRZzXpcE3t7jpMUaRKx/z5DuuGwOL0Co6Svkk2SVwNDWWh
h875oxd7KRK8/BthEyiXLmjcG08J6nqKNliOvxSEs43FucfgjzDsLPVJYJFTSEENeEyp5WBAHZmt
wJ2DUAhUO24sMNoce2X/RR7zyAud14sG/63mmZrVw5GxDxIh5+9sC8hCxDt7NkUgEoJ8X8VHCUxr
N+piGkBhGGelE1t8PZ9eG9+lgKNWLe1qc1WRbe+qMyoG1MIoDbtGxqoL/cT67neyDsdWGDio732n
40I8/x2TSycZyLWCeK+EvzmvFh2C3AKJUCtzJWCSww4idejrN8gRcSD3KVNpdS6XgFmRwzQUrPNm
zOX4My1DeplrLc8cMsmtVysuVda5nq6uB1ofwxPuhO91gzsgup5U4/bUgUEQjmgS5VpmapMuM451
gQBjhfr85MlqUN6EH0R9Zh+qB8+hemXY5BaoSoNgO9VkCjQ2wDBUwUYr0SO+XQOM06iVvNDLUJ1d
WLDUjsv7lRB3pnaT2RD88IfZQ3LeQTUtt8HdBVVDHxirprz0ynlLaJCQfkMf8vDcc2qmPTrTJXI9
GQT5p/xXAW7uIQfE0Uj1PnAN2GFuMIyJlHhy0vk5n1gcqNMSMkmNqUWbvZ0d6H+sFPaEk9zeK6+a
z3ClCZY908j4m+/8Y/cIrEWbMTI7q0dCuIurKKKgOTFChTEGjt6QtJ6xyo9ECsHfXikgVxFdiE2M
oBW+wH0yDaewDvfTd6vNJrZ99ju8d10Wv/2IeEj9fdWCQg/0wAwaNmTzDKzY3it6iYje9Wuz/1ny
LyzfS8XQTmE2RXPlNiq73KdgwAlk70p0IB1c/NvZhfHyynjvsxw9Bi7OVqb+OiIFJCApnmN7ILHd
5RLwEOrWWs68TyefaET/RrNCR5h6m0fkEIIoOdKC2o3fKipo98n+UuPnmlmyIyp6e7ZzrlGeVz9/
cTrzG5RRVPOTNQffG1Xr4PYj+wX59dYh4azyMmdf7gFDDKGPET4jzjOUF84sD2X2M2aFNbJKJpSE
nYaGlDtpc3k0fI1a+sJ3/UtlXgvAQH//k95S+aay2LT9HWj08cg0uR6AMhalCcT3CRj5AKU8GITy
U3p69kbf3y/Zn5pZxExI65XUznm3RaEi0Lz/MX4J8Dr89s1lCbm4G7JmC+7/MX8+kTzQfVwMlQGr
EpKYwQn0u0Cs1eAp+PoRbC0qciIvzjHyJFFKk1X5X37vMnhQ1SdNBk+44H0DHkg6yubXqkclGfOG
SUyyBLAiaHJhIPNbHNA0ZqQCAZ7iNV6gTu/1n96AsjoWwF75HA589Olnjkq6qzECV5gBVPR6vCh7
IHgfc+xY1uLcPwH3Pt+JLwnp2hfeIapgZJ0uyoEQf/ThWGTo8/LCiaiCqwr+lHtGUbaldxd6dNhW
j5TSJuhPpuuE8CUJxiyr0JJE31oeQLunDtkuogIp/8JwhPGq/r39osvamLo9SVDnDUG4QUdOnsfg
Mal8BwfmqH/4ZX25+oJRAFlgpw7hvhyncxX9iiwfF/H/uS4dVCXL9iFLSij/FllQFmSEy0OpFSuO
7KNoeWagHVmnRy6Sb1FbYM7+6FekMMsKPGypAVx/fEqxc7eXz0RdPorRbwLMwnQE1NYeXcjjnPlz
NZ8+hdMfwxAuILx8qs+jkO4/CJkt/2MLgsAB/RXcjBxyT2GioD4CuABZnv27zAinMvKD5V7+JtxG
klXlvJ3hA/hOumCtOCXpEq98HKTQPnb6JgqCQ8ibo526afGrz9zJ8igrQOHSIF7jGvSh1Ja2ZToi
C8OwujliUTaRjwQBsCB8oIKyXM/bvj/39PZxFecbtCRbOIJTx1KInpPUWAQjv3daNvcIrE6S5Dpl
PEJZvKGxTBsFASaH1qwBx7SF4U5XXF53TwpHC9CJ9zsN6UTWiJ5Sy2jbQBQe230R2De5ZdgL0jps
S1wOrKd0dmqWxxn/cWGfok7RHv6Rv872buib7twozaY1/wS9yqf50Ue7HgFOoxfaoy/+RshQ0hRO
Yoketcsevyqj1RgDNw2DfQxhajZyBWmlgdM1YDE7M+swIn/kJBqm/RqEJGbTMNZhVNcRmYZkolFn
DzGxcE+E+KACsy81CrKZNu9mo76WPOihfxmwoRuf6hXfIL2zoNNbpwvECpocoAmaBSPMy+0Ym0rV
LZ2eAfS7j9BgXAmLzPwnu5NWait8tPzLs20qUHB1zrwHh620HyFtIkHF4+3aBSFawqD/BjeWAST3
0DIgMPqMiaGsCWl9ocdsZDq/AztHN8CE572z/Q0CZFg2h3neDelTnHkHCHtXlluu8wvMBVQ18t3p
VGvvgo6ViO8EKL+zxvR22st3yZdthfapCNhSMvQQYv5NlpruPncBOoZTxrUrp1VGRZuIbfLpZMV/
kPQr5FsUFL1Sc+9Jt+Lyc3iW95kWYWDsuv5n4bQNxJGjfo/bxzef2UwKTDte83icW5Ut/PlB4VZL
M2FpOxVeFQoqJ/wMFZvTir0oxxo/bbm1bpe7gYZcovI7zVQjj+lDS/bxn+E5vLbq3F3umw8N2btD
f+BlwjpNRH2yceeIfCHHfGTYvRKOfG469rDSlWVWs4HKoSpSJldJcqA9Z5dLvWuSRWHXNtQ5EwsI
5dzkYGGqvBOv+sFoNHUYNP4YsiCcPsAZgLRNB9FDwGnNNvGZuO/0Z9VcuSZScX8aOe4ITwrhJT33
UdkgPbIzUundulA8WpqKH4q4UULh+gbMMFgFCSUJbeaugercpIL8ZJOJNnPGqx/gbwZLTzBV3XlM
hXD/cgGxIjZmt2icNTIRTc3cDCc3HAwvFdp0CEX7M10UsrKHvKyLuDgilPNZGUbsAn0sPs1av0nu
5nP761Ckl5ziQxlkSAYk+/I9eW4ak5d4B7LZs8UiZ/5mpa+1DglZleMbFyB9wQwIQV7/Uu3KITPV
gFvcfaYg2qeXCEvACjgj+am3h7rLdn6HzFcYnbBdRO8FANba4nPNWdlYI/j6ifVkqOV0yZzOn+79
GwrfC+vjMp1ZTGkn2BD8eCvyAq+62Ig2eYwD6Rm+cZ63sC9mYiQvIQzyCwMQJxxjbZ8Xl84R7lyE
pz+3FevWbwd2PIoX+ZtU/57I4OOslCRS3CDTKXEEbehuQs3jkI0Bp1YlfO++EdrcVZUBu/wdMlDz
p0BGnJJVREt5o31Rt1nDWouOEfiCJ4NeAoAXAkzh7eFMPTTiuLKzspLqfXHAPX6fh6Xv3ANs+8dv
L7kW7JjlaF+vorLXDRNWj3yn5qbXCf/1TBGeQiStN2JQU3WP3/zrPjR6gkOct6qEd67OMc4n9ZCb
t0pr1TNVYCnOE+huJGRmi2NY7Fm0+I7DPy8s6ZwnfUvYRpBincXYPprU3wC8jjntyuBWCQHnt8/6
HbGbEfnGTbpeKCikZM1qWrB6ciTsf6gyNdcIWuzOzB4CSv5Qnt0pkh7x6BUoyStdOecnrI6yX9Ef
f5KNLA6NvKhhmHN+gWTkuk/9rpdg1S9HNm4xsuPpSdzE++IBbgucdpV6HxqGtnpBxrqNQhHaz1BJ
9v+BfS42ojtYVvE9FePQV5Yfgp902RILMAVmZEoFx1gg825hnt7VrLgmbVv3YnIZYIMtfYLLkMdv
8ScjcpSZVD1LhDihatQzKbY4EdEVnqLQgYzBe3QjarP7r+eiRytN1TLkK5yqcQVIIKEV7BHOl7LO
I0LgSkiHhCtIFYoMoT2/m0+hbKbzX07jGBFFVuBq+ykjxk3/7DO28M/opfhCdcQLQrcZMVNxweXT
tI7KDSbp2tSaQqq0A3HEIo9Gw1SW6NqAbxPs/WjR0qVQfAjI0zRohM4MDtmogR55zpOKjH8YfSna
tOTqKzKttI8nLr9dfh4om0XF6nnXgGW27OKXDV5aUTI1tTgK+sGmFuo4Ex0QwMNK7dZJeVlaP8/0
K/vs6HYB++v1NTt1lBikmkj3ENefa3tIWGJeh9LvJFsM40UlMBEFpHG1wEiYD3MyrUN4q1m8a9Rt
9f9orYQtwdwT1FFmuRNvQiR84KfXikHvxVfL8nIZi2bzEni5WTFHXIO4h7YuQPXs6XgZjKCxVXnY
0s/NTDZohoVa68HSSrDSoCFtSCF+0gMekcjHT/TGkqQL1WyDrRONkpTbS40U8V2cu2Ha8bzW0JIV
ofJBiFBgRMQOAppAok99M/F0kHZ7VrNbu+bzY0efG8SBwucH4GdRgNfjaUOZS6dchSmaKDMWR6bC
nc6q+hQ/vwWyyOEfqW6aXzQKwwxcle+5bxDgaK1/ccjWl/05uByOp9u2XUaobaZSdW5ISuwyGHFH
I0vDcZrJ2HtXG6aHel+IBecvUaqxVkTv3SWaYM7SEBAVyu6rFQEjgZT2CBXAervWqje335Qx4VmN
+wNrptoEgYvTyCW6Cnfjs7asslVLI7mjp2fohmEDDcVkqE/ZTtOgGoEFYQ5BrsJlWZaDYAPf0Rz/
nFIn5E9l9b2WI/60dBfLe02J16XYnjSrLFXf3rD3PuWkQfHnyvxlVsdKci4gpHsK1fao+Zzs09Dd
hXQvt2MMiSa0lszTt/YvHxw2tDFfBCqFKPHCkVLF0EdrXoB6QOT9YmqCzDUmpwWtPA47OUmKqlQt
5aY=
`protect end_protected
