`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d5VJXu82JfSwswDjhvbEU9He9tQ5/1Rw+4/2nB84LUuT0wfekcnbAADJNd0/JtXdeaCUlOw7Zwks
Bp1VvQeB3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T1a12gH9+o/WCd/uq6lAozrIbwFwnflilDyEA/rZKRAxvRmKOSqBXtjVpxVSoEgX9El2BLPK+36k
Vd8y/iFx5HcwlteYeuYuGTvgQerRA9ycH4Qwt9s5DC83MaSGod9ecMMI8PPrmdJ+hCOX8sXwEsN9
IHAKBa7h08XDRsgW0os=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZE3CBd8eugZohbo93EvXvQkUxCnosHfYT2eG0uuvFgW4E1aUdxFin2hcHpeAodvxBTyPhYz4Lsqw
3nsUxnz9hTb8Lhj5XnlqKx2mVFP8Z35n8lJk21C09QHBGoSukklDPI8dbQUv/KxN+k1qsLBHfCBA
FWz2UAwKlgCaoOPe87s5MUwwDM1/P/D4+XgEQCRDz/7JDN7p8ZFVtltMEx51xjJOCvfGoEeTzG2k
908lkYgt+B4pvwsuFOHwC28xicC9lqwuIR+OiqTI+hvqIl3tijnK9dhEHXmlIo9PqdVp3p9K5niF
C0wKwI1gK4zk+Z+Qv31AV2g5KDXjXxSpUgHlpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1K/c2Exmx3hO4tktdfNX/hsUCqBDw6bH/vDRPja11f/SX2mhefMgy+yYp/XXIVeJlyTPI7AwLQ+m
jPsm9qUsxInkPzY00BDkxz+XjPmDvPZhWK1LaTfp3S2KuDInJ2AYP1AwgClVQtpRFpipBFYqQeNS
QrfV5V8iPYsCh6rtCZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z2R2Fz5uoP9gCKKJ4H8ByaZdL0II83JUVbmmEiqboGhJOssYqqghHZS4Xla1DO6PE/W7lUbFZBMN
taobe7WZ5vLL3z9KT5znQ5u/8vqZfQZBnNTCM9ij+NRl3PRmkUPrtcd6xURukGspBspXFvJDNTq6
HoC8rJF2dAK3E2hXtQ2qzFXYx2JspRBZw2ARE4ENjzYZSYK5AhF3nV89pEvyjDlChnkSNr7Ec2sz
zSK49rQXLtbokqxvvzCHRCEs+NoMqKlklN93OyjJFAIzYffS6GiGtNeycU755Cv+/fAQynybNWn5
4vdHnb+JcudvHzAJFK7/azTzKOJrOSm9uJYTZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18928)
`protect data_block
mvi3i3MBI7n8zvuunOT1BL4eDGhQlMnzDOzVrYI8XHOS3ZoKFTTDP4UmKkCCDyXvukS63/BOGJv3
NoJdfMFYhDx7pjz50AatTRm5dOIAKktHZJVnSGt5h4GNaEO2RZrMb78Xxh3U1zVrxlZ3qI2EnJOc
mfKzDD/4p92cen0KIbw0o/47imUtaRrkguS2FWGYh9siVclH1kL5cuw48mIsnse+TDhuRB/CPf2+
aE7uqWPkucaGk7k69/AftSp5jcZSdiE8ReN83EeqSKUNwluOxTwdBW1DXFnFKJzGQbzmIiEAvIZu
8SqEGCQm9xpPTizV0/XzQH3z68ahiPYL/hjiXOl4N6OFp9WziYF89PwlT5z+Z2UmRzAzlZhM6lgP
O7uzHXVzH72i19K0AEAZmWjYDL8f+0uuWysD9VWEhlqTSnh7KxunY6fNGQ0RoWvSbROnlmj/fqnD
qn2qN/FqZWwNTvpweJuWzcXG+aK3p4u56bLy2+dmnjK13Q2gd73/AfJ/GXKUzdAzLl7VHSDFuWLA
e0fj2G53uwPCJ3ppVO04wnNmI4HecmJDK01ZFmTndzEmw9lEGPRpIXdcaQFtGkfGDk1qLGZDirg6
fzxLz/aH6u3IjYG2YxW4zI7fKUXnmkv7XClVZuzGFzG2Y6CEr14WaidNRlSB3AVEJ71+mj5/afEJ
dz8Xg01940kAqcOPkXUbam+vSDziHWQ9ii+ID3W3hANdZdMW6XJQERbHL94TrU3XMo3s9YdGLSsK
ewMMtC9Xl9U/8Wc0ZD/yBsF/EyPvpGWPDIv18EAFwGtVAOqj7qAiDJpAQWtl9kLJB9Hx0Y/EU2Hk
U8ndm8vP4hulKylPyW5y7bHnhC6Xx0U4hcuzhjTbQSacH3MG2No67E66R3KpSF5G9cENvSv4Z9j/
v7k1Md/i32zsHKjW/4qNxsq6eCxyb8Kt7pgEKSITPdfiGjM4Yxb3vNPuPaCEqY417v75S/xNr3Cv
MU39w1KksVAdwfUB7Pf1Y37PHCuFg1JXk30sgGeLwGPt+GNYKSKmL9RlRnliYv40g/okCNKIHUHB
Zu5OSd/ZofovAFjXC0POoVSCKyhe6ibDYad+5ISI1BOWyojVBHUAKvNJRN2z4SI3S/vUpA5PoX55
TwRgMC01tuJQ2Ac+tGE0q8HLVZFVkTmOUwQ95z6YrZZ4JEOPHiVv31fKAXPJiBvMrqgNGeVM51wi
WD1bhHPDB4VN4kKcaiNI9yDmzwdy6jbSdxw3YNaq1Euomm5m4TiBjTaD6Crv24FCmJ466HdHWpcR
V89JdqCcT19lXOaf0xBJbsZyXXGuNduWejoxZuUM4ruurRUKqOqNTOLNdoDifFOw3r2eR+R7PWUt
7d4waFwj8UKZP9C2BXUtNZGcJDMD/2AL/U1UMeGEajOzeBzawZRE+k1FMgl0nfdAuNd1HF0hqW9l
F2kNASq4dLnMvXhg2XWLBzXCqE2ADLEzKnHh8T0xc/jmfGIGNJovj7+Gr9NjkOUqjdwH/uFgZAxz
04p5px7rIUsNVVzOsDNi+oyVFlNkE60BbIMS7/Qec3jTH5tHQd4uIf4MegSKB3+5eukwHjZVwd5V
lNWyW0/Ufn9mL8EeFKYwwpdUjnRN0T6T3MHhqJTs20+lkrc+2LtUvFhpIeNNz9qNgNoGlSfYSBFZ
43vL8PGOkFSN1AKlKzJFB6IzqqVmQXIhcdVKrhvGC6yuSkyk0wc5Ze6514A1iPzuQjYFQdnpr4Lf
5a6651gbCupHEToGGrFuoTXaHUMiDeQeuYWVdDWZaZlnYiW9RkC3O9Qt3yHF2uib+JNvtb0txC/k
kHu58LCZNRw7R0ROTf107lxJvIeef1BJ14UMXz25T66UIZt7I0bReX/+O977MkK7nxu0/KRoly5h
8Z2DqfQWKjAyy3R5bBqeF2Zl/dSdeQgqPFe2/2yPXepxJIXFTzBPNSnAn/2X2V/mS91lrjOCreJH
yWWkG1C+Hn8PQiqx/0JNB6HvxxNG5VYJEvUfCXHsJSj0gNBaWsSRBmv2I1O31ApZbjRS51wBThFv
G5RogfL3iq3AqsJbIxOxzIBOoe1LDOA786eef7zosTh3GbwUJprc/WkH15gQ3NxbQoXF0qKiO8UF
HFodQ+F/pHQhLl15w52SDMzGWludzO9/ZkG0n/LKWJ06zRxJQRev0lRRrfX7J3GlrjzYbVinOE0Q
bLRXYhhUf1NrAtYzglWu1zg16CNnX+1dTH0eWBhwccLM9yW4g3X/SyO8ne+wY0ixv7oNY8k6vU6R
nKe/SY0/2Z5FYVXWA2WV62MxngLreWIcZfgPsfN9GSwMmF/Ht2hgTGJbOOJZ0hXXc476/PzDDAUL
+8O9M1c/cMZgLbg1iVYYC2f8OyhpAcgvvyOYikxyrxElZLcEQE9PsONidcwIVMNlLukKSPsRtY33
3n/fSXsDDisZB5k8QJYXvx1HqSk+QQFLM9vH7JCFh9k/lT5m2nnyEDJ+FgEaqGoGHgaL8XgpSm4g
mpRdy/oSoOKcoSzIC5EvraZ14TDfUF259oLi85cUqhx1hNxY4rmgPt/GD5n9w9dDwSUv9AGOzrSB
24t1NnmDkp08EekUewAe6T2F96+S5JPkHr1C79wQ8RcczVDV9RdXuAdUykoK5lffCpjQvwfE9Voh
+agreKxt9oTZ1lUF+DZ/5FlJi3eZQwuY2xHaiCAuPDvpcuAOiBZxGdDRDm0BvXkv3aw/zMn3dcQO
d8glhI2C5Ggt+RE7laU8rly6mAU9CaQWnoZ3G/cdxJMj+cv9ElmW19LVzwjhYK08dVK9Xqo+i6+N
cqtWnnE3LnRf+29LrQqirm8XGrX2lxgqXAQuB5uNq2HjW/QHunbIq3Gu4O8ytc7ELHb4XP04fcor
5bm9YsfqGQINM7knC9fGQyOb5hDnx/ouHBdP8JsMwZP193nuPEMwJGX5iTHmpfPiyxrTt4xHZFEz
QaphTlfXAAN39Dk60BABdXq0KE0aSmEvWrsuOJN7wibh9ZaB5IWGewpRc2hVH6CuLpueZjpdv9Cv
vxBNmjLKfM0YC2PXhGUW26enLa1zlZbLjgpln6UkjLdZWhZPijFiALXpiep0GMLhEBCcuHe1e+rx
jz0l4g9o2XLx/VVS9Awr4fADCHSfpfeaoSaxsxDQGSIazdGtVbI1Xq8SiMhSPbEpSz4vFLUFBD8R
2juxZwcA8/qS0k7FhOsaO5jTUIqL8cz9Fn0/8bVFMWF949odlVr4xPdncOA6A9vI8dQTHXDGMDSA
vk5hjmzND0HwC4UpzPEK/v+V7UldrDz8CQLmlJCrIM7ONz0pSwG7dPhHkamDhzU3Y8JPL15P7UCx
75mW4U2baR3AaAUyuFsHiB4Qze1oGhYAY59kjvweiPjZLdMiz+3OKe0BXmYY4vD1yhI8iWdZ0kLK
3Ey5SQhux3IbfpjgegzsbHhscfLV25eOujWFwilVrohd+9vfi02q5DC2d64ZfHcC4Wg+JQwk3GBz
Fs5vATsoKaLLzduFNUqI0ZR4cpu9lUmxdnQjGWukI2XLVLj7VQcrxm5c+jW41o11GtDnUxFKGOA+
afU3QwjsKkZdnMC7EesoYV3BoH13ozgkyOpNqRUd4GMIWCv9nXx/2SpHhKmBIPm4fMzJvY7nUAbe
g9iue96m5XDz1NXGYVe/V5W4wA30/uLQ9uQ0L9hlLkysrNXX1gWOe9Ohvr/fSdpY0OjFxx9SAmnk
Z88GB8eq5//wzpbYu8TryhZi+S5qXLa/RRRdfwlVulAAPh8x1xDcZGqaZHPU755e/zD5SfjUxdmK
E3JGWN8LcsGrGbPUbHxhq4TAcHIt/OD6oYBIVO1bVSTxwCR3DNHSY19OVOeJMpfN8DtlrUYatL0E
h0+XvwubJkFywRMslUucl9X993Vhstg79gV25+En6SfBCu8Q2PMhuX3cBDk2lS2IqjRnayZzWd0r
w+uRlgiIHisM7fwSC+74YYJgLtmat4+9lxFUTxRxZjuL7Ck0UP+dybktFQfrtySowryWORumyD7a
ffUsIGmo+ZJBLGlDdarfOOGmWVxWgHMIaz0VvrjCox5f5IcNtSTgWtylv1UQJICMbCZXa/Iv6Bfj
QX9MjuLooX5TSQdquAh2VawQO0Bh7M47ZTVQGBsK5j7UcaY2PzZBcFfuTO3aep/RIQiB0jhuh0Ah
4jTtqK9bN1WukbAPZkKG+EK6nGRk4r5Ft/iiFHqyARZEobRMGHqAcmY0i0M7gKu+khuA2IRTcqve
GsK43EAgcd9z6EOgjEwBUfogxIV4tNWCPps20QXnu7X11CYPoeBqhk/D0Kk5rxwjAoSAB1GHtID3
ENnWu4EkRRFk5gSj7TpXKEB00d4uJdaN1vAZT/tiqAIcBxw+elseam0nv9VOkRcsWYCVJqDLSk6E
/CN3+yErdc1hmWrTudYMFgALq84pNwajDMSQuNf2kSMZP9wOqsk/nAPFptVlEZI3K4kISHsFEc8U
VmRHEsQdAjUy7/fmzhx5Z+VSEoEwtC5svWISZAOjW/WuOfe7fg06r3ceye6d+xZkqNL6xpHnqRfV
CZhrZ766vmyMGvrqW79yufnh7WVJ3cQwSAyNIGLv4frxfOYxqJkPA+LDEr4D3oKvz7rMTigTR4A+
sEWrwpsaNylHjn6/rzUFkJcCqOD11Imkr3wruYIJbHdGq+dHIUzNBSdo4QR2daheIDY9a5rDBOKP
mD7XZdk1hTHKgnUExZJWwcyKVM7+DrN0scGXgI8TJhFIf0wOddX0zoRrqkmzzLcjpk1AnMK1/fRx
0NoQoHe3zwX7QZ1ZmV/QESu3FP8v03LCWtT0Hk8zy3uOgk5w/Iq51VVD9SDqFcy4AUdsC7HessaT
sKLtITKHH6NQ2J7Ssz+NGyDXyojO5gVo5PrLTuFXjoZflfWliMl7Oh4aKCGeE1GB7ngBw6y4loCE
Fetsh6d1rdvsX8JPiM0HC1FrxNASZ+OAua0EIGJWsso2rvBu3LQuwfuDRmwxWXWNxmM/ESNkX31b
7ZWg9+1MB6/9j+TG6/hR4frMt/4aNVrfV+vg2/DVx9tqC3C663lRcg3A32qNr0LR8mt+LiTbWNwm
4XLPBVhiW4RqChTSgXQFMFAV77+E5tEnCqZAD/Qp+a6gQoWjEoCHDo02jdKfat+LXNhP3RrJnPS2
kbwIArEteRfDFbDSwi5aDBU8iZG75CWT05IzDMYgAG/I9k0tYmEUkgXutGtxslvy63lbONxUFXbk
pBkyUrtNd4PRXyy3BVbeHIdD2S9Mbn4HNy7e5TlCRf7vegJ7JIdf3HGxpXhydVaSbMaBRJwA1Kqa
IsezNfhM2fr+XXTM94Ak3cFOpzvK8AmsxWSLPCH2PdxGbHbpbTPN8GH0XUtclzamkntwoUfH8peL
zB+qQzyHWkMPglNdoHXHc3gzaQvJeztGfcyGsyZ5h7F0b4yG3PeR711rlAxCY+sZVa2ys1QAS2qx
zkGetjxcC+DF8Rrc4XyMzUy7kBUw9t/Bb08gH6IVthngkkA8U2o5YiEKgY8tGqybl3kp7sq7z99O
dU2kGS0nhv9ZUU9rpqbogbBvv6x4oJjYV2HKnbaKPRYvHJ7pJ/FT423wCWkkgJqPEh2K/zNHLkVv
Y5UyQV4hKA1ca+lHLBpGmvchuEyMaTH9Da1xeRB/gRgrGRxK7941m8M3B9XyVXbqb2NRnOjZc7Qk
bORJZH8Cr5BF4zUoyKZU3lXZnJyxVBHPcsmfRYDTvl85qHaIeOnJnwKHwDQ4CqdrTJXcHdyu17v+
BFl6Zuv043XzkxfU3W+adfO1W8rhDxawz5uhjk2fjvAOafiy3tN+9zqNsEQhqeXCkHEfGXLxtIA7
MRnwBJXdZqgrmfzkDwa65zB3wQGc0KWi3QJfxLMzgzoxk6lbreQJ2TjrRoZu3LHh5AP+ZD0GWrzZ
OlItrK8cRWf1L0Ul4C10r76Tnh7r22MmDKHHrIpDT8Cy5/GZ0VgfxeYxHiWAF8mX+KTHJoaeYXJc
TP0KB3SnKZNsbLdrKyCi9DaQLxt47lSx1AYJtu2M9CuKzYySj2THbWi6gIDdtWm1UMz/Wk86nreo
PQsFXFGaocXFc7HPykIHpwqGv6LcmP+M5pMPasHu+7WKVa9WZZHGovdtElkt2AuMkKUjs7D7t/fD
l9UqrLJ6e0p/HSJ+OXslBVKB/Fg+agtqWmVYzcK4xpX3ObPsLREokd/JmMzhL5naheFWLVfaT/zs
nDw5DGXwbqdz2IDNeqOUK6gM4umMK8hRrM/HJIWQzTyDopv3FGz2YOe1zVktGi6v0o1lbfjYNdCO
lM/TjMA9Y4XXHMmf9urV/4QsDphEoF7q4LisSID0GX+BZiTtvPRUNUNhE62ogEQ3SczB9Gtutuap
GZAlL7FFDhrllVG78VZ9fzofMc4V0LchPYSHRvwJWBWmrveX8n4jNZCutLI/1a6yAEJ9pB7CcHjG
XM5mJAovpMM07ElSd1KXxLRkN1vqDwcuEu7o9mSUlbVjl+0pC86FD1LiquN89LVAHoN2LPfdmKbi
MdQUFZE86+M/VD/cygyIfGGPG+396Diu7YPvG3cZ+QNxNoQM+fAvQM7CaWfTrOwvhkqRY24tV8rJ
SVrGbZ7Ru+s25UwOxuiLLdgoqS68JOV0MHVgNByINN/kppDcIjiOw6cbFakaG61zLVFySyc4iESc
cbLNkQ7CDdqjgKMVyQdriHA9BIBSM7N5jk9ipTDWuxfhicuRx8bkXWrGszQXyL/6/y+O3UHakId6
L/vqO1fPNGrGGDu7v4fy3X37hGM4MR3OZN/zonShmcX1qXlVT7fgVUDWLLhBPgzFg4mh7yss9Ypz
kXQ2AyDnpmYtKMotesvYInk2GeHyD7K4ZLcKO9LPqRfrMfupuO3F22yRFked0uodrpJwuNOcKl8g
vbiI7Z/LMlh3bOfJYhhwhj4mEiukpU++np8g6mPVFsywOzbviyQWeuoXuUQvKIi/p8A18yrAhaeN
a6DPZMhw0xOby/nUZHY+82xZ/5qKexKaAX94MnqHObqQW8U3V8Nkm5lxJrRJFbM0AdzQQxc1SKyL
1gI65koY1FSL2VCEC9QypEAOYA7aIhhO+Z7aXchY3B+wr3QJWbCO0jo6ltShbt3xaunb32LrOIIv
Qwz/nTMQGophmVIurTMHpdlrBqswrLV5P1RC/b3hUOsXlL72FJCH7y9xkPamZIKpFNBn+mWOXJN4
U9i0rb8U8/A/S4MT7tLMFK8LQs+0s5eEONC8dLjw7ppW/jDvP/UOamtEDufMR2W0FPmK18xJK60x
5hvdiTt30/S6+kIWlaWdx1BwSmHgBwTEMaaLwI36pt2rJYx1dgFUJeXwi0nTvHCNsuNC11ZkqSSF
i/oxNxnt/Loy6Bg96gk/lAzZvDCB3TzeX70tL3cUlW/LOI4O5fsw/jWcsOV3CTExfWCrD35lYpP2
ZCZPgMao0su2/zEQdfdPT6M8NWTIUoqNMug0UooS46qr4aideiHKVN9SKxA8S9f2XrqEJwDqmxdB
smEaCskeBxUv/mP7wkS1tqIVy38RBpScr+qysEvKZjHhWsB0FXZTvM/NdAelHYqRr3Kimrp2EQT7
CduPUYHZLu/GxjSR88zZ16fkIIezt0WcO8+hZZHtEx5y1vv6X4R1Rvu7bCLBX4Ds6ijXPmoa9qVZ
02GZBaBLaUqxIFlZEeIwrN+UNlPXLplUAiGoeKf8mwmb7Ygzo7dr5erj3uZTc3nr6dWTQmI4cnnv
fz3WFmGVZM1nBJy1l7KaQ9Czp+2q1+HOCFdzd27HM+OiBRyx0HRAEXzN0OzQuM9eF85ELk9cBS8r
/+nlfsUOQ4w/z8b6rEiIdHdXVqLRalIEodAv78Fpx14mYl+9ul7yYSzQ+iClgMWtPyb6Z+IHyXMh
1brrcfA5NkgKzODiDTMMSIJHTc7G47UYBC3aF21/w2v9mfEw9kbDLMeLoLRla5dNZA9fdcowwVU8
Y9GvipWROq0Wo05nbC/3Z5C+ZfWkcDnMQTfDLXllR66OKBwa+u+0maQu/0OGd452HkngdtGY4jgL
jUmLhQsfdBt9wMuLHTtiHmyG2pOr9VjXApB/Tdxm73LpuOjjzA9p0mGhKW5VPIB6hxbjE19jjNe4
4p5Vfl3mwqS25gRQ9KNU8xbXGScZbvFrnvDW29PqjUhk20YtXN65vTbSWkCFaMooD9Oui5P8tb88
LxlBJWXE0Z2dEiSWrad7qK7DvoOhD4a6idB7d6XtEYwPPE5c0GUzkwLW+dvLxDSyb5It6/wt/X0r
eO7kd00C9FB9BCSs2qryQdMPMT0nslgMEbRGbs6IMDsotYQUFTT+sPaIS4Kuwd9OavtUOsikMTGr
eEsLo+LWTcoBmweTQn/eMFgKxkXio6Ugaf6+FeDt8MwrgLEZ+dn51gbxK0sFn1dStZ65oBhJo+xA
5I2sFsxf26D69T6NqJEMzI5vR8peWUa25dIL948wSK/XbBfEhzK5cWJ0+QumseBfstLVoPHti5XU
zWg0V1SR8/6XIWQdS/HvFfZvdae9QRBS9OEMsGXqh1vyGHHtWpolzW/rHwZNV9bS1jdOx0nnZnHC
cJzIFqeIsPTV4+k3WhHou+qW7pzAq6ZuxagkBKXvjdxq69C9pEe51yTr9gYcJqv7zI2fPugqaGQW
k74F/PuO5yof97IE6I6095o2q6x36ZwsZaaHMODcWkthGa/r4UP3YRMc/g5l9YQ2JXCMkVDVBCli
5FBaJJ7IhiLX38kw0bIXJx23R2SqarrBfNwUhYqPiO+JayXY2Qr2d14mh2vVuvNMJJsMKinSP0cD
T2Dmaznvnfz8SZsEmusG05ZmP58fk1+qi3ZO7t4R8iYibB7UTXAoHm2/JGspskDpJQCCcBFGUYQT
O0yETgezJ1SKD0nVeOu5vYGOqXTpknhG21BxeOYqhS5DpYU+TyOwUwPZ0C+bAvqep5yqJ6EABvuu
m3oIvoQFXOh2BGJHdWeOVQRc7q0laET13CfZZeA4MK2VG0PFt2f0CiGkppczDFi/05LFcTFHA59f
yu5jFIRm16sbDWU44GYbCL0+LXiOR+pO0/SCFF0Hxo6Jg2ZVNhD8KbP+O1HQ+V62IgIBsVzIw3IF
9PgP17uwxCoBenbDhgUfwXUjv4tqRRP9MVwQjvT4sSjKnG9W2QAPLzweqrb6kZzDRRnrscrogXr8
8bCe0mixfT6eeSnrnc2NXg5UQXPwRUW3fbtzPyTw13Pn38rC2ydkZvNLwBn+rxuk6IoaehhU0zXx
TcWMoUlYjNyoHfaj0t35YW3HE8lTYZE9TER39//RSdKpItjhCQkT+BCN9JTl/yzlqRAmtgQceuNR
r+M5V4B591xl6sIc5WCh4DLhWQjC0YcqomXFdUe94NHpPrr1A2BdnE5iAi9B5bWKYIZ2mq0gw/EG
nZYWJhyacu3ZbieMy9w9jEGDESWZ8iBAhrQRgMY8VzE6nfdpq9/vl0zDU34vqyh7bn3cFdhlP6sH
ShudYO5aEbCwiNQH3DP9jjOi0pHSlda6/aTgiJ/Ewk3iGjvP65mrPjSBXnTGVfWeWKns8DUYcJjE
PtlpbunQ+kSeaLEZWyZq8Z6LFEhpvXJbU0iFxT/srg4yWRqiXeLwsRJE4ewwuUGY+n0/V8/QzJ3e
1TBkM24x0DqZJmqHwsnKSro2xIJQ7Q23wZ6lQ/aBcNgveRVmzCkfRdvdxfVIfmbrhw/60jYPTcdI
pA1qEWQmXmICl7+0x9Ka9I/d4I387xosbOkHQQPWfRCNUhEgiG56/pYGnCOSXwlfNYQ5heYwTV14
Dlm7U7TgKeO5WlyDJZxQO2iSZhLbqOHD+nAXljNlTuNacubIXcWkhYvPp5nb6MXpL+Pj7FxlgQpV
8yWsEbaEzO95fDRMK5j+o3s7p048YXJeVJoOd2QW5momyvAsBwzJ5YqMdRlStjyDcAriJ5T5C51Z
sq7jdK/4U5hinIZ4u6lOC8EUL1/BBRO8CtUHaYCEKKoZ3Zg5cZVtcw6cI15f7+CZgWg+/TpN1hbT
yvelV39f8N2D/Ig23yVLcOnOoEa+irACbrfE6dX4NO0S1P4eF2BxTlvbp54T+dM4rSviHRfGsCi4
9evyZtyASigfEKfKSaPsjaw0zxP8PA6LmNDuua2GnaXtafjQUUdh9R80peaJ9Uuot8HOwRg2BdN8
gEresgwgESoWTiaGLeABoQJCK21tpQizs5s+bUCQv+9F+PeifdPGU5JCxsc1LITtbr048dRmEvPr
dzjxS49jN56f1HI+dKdVnpwbmMlzYAWFIAObgzq0Ie6/MRnBeQr0M1hJjxnWGu1fxdMgmysgukP5
jC6mtkDYx3Ep6rQuAQwttxcZ5PdZbCozT6Ste/RgeRBp4NJaaTKggclCbdSnDUBMAAJEtdYMExq9
ikgwsIT0Z7M6tsgU5q564NVC2B+Max+fpHLxdeNjB5AAwLTKSPW616Z+i/37wwrSiq2UZHXrYNa+
is97jst0CdLF7AiTM1V7x9F92ACPA1KPm81h60V0RK6H/GsqVwfH80cV7W2lw4SJGjSQoTMjw7CJ
nBnnwuDLCxzMuOSdoQN8eW+VzX29P415Qb1VhF15MynvwTcq95sKdJzyQa57XIET7tEiegkZsP3t
GZ1Oz80DzhDCXeHI7Bv82D+X/ewupUWPsWNNt9KyKV3UmoYz21rt+GkPR2MCq4vuRQ3wJn8o7r4Y
tFvQ8lHnFAf1KHHUtdTZKtVDcd//i7ZU9QN3Aq5EKYKREJrleUstP2LEiUmNhwf/3oJ5PVGGzhGp
y0qfj5d3CAkA5B+xlsOZJZ4Czr11g0oWgNvlA+ydu9bHMtKq161TGXRQ2U3Q3ShMtHCkw3+8znIf
TMK1shFuC1aHX+6MwiazsonbiDGobRemw7zlJu71kQZ0s8XZn1nt4JI2o85nfeurmlE5xZwqWjKM
/1GIgrWoxPu5bpIsQknqrA71jDX1CeyS3XxPcueyrQcmuVi9cHfVn5jwzQb5eYTb0gTKB+Z1TZiY
PWMvQGUZdfiOJOmXqLpkt4Jwji5pVDICOKqsAyv9nGxWuFXyy2xPgdQJ5jLVnX1NjhLDP0wdP3LI
LQhr0b+b4pEumo1flawoagTCP6KR7m+W8Tme2us1o2jaFiqNujI2He872GG0vr6qfLmL2XmIXkzp
5m+jt6IDdWdd5XlOwF3TnU1qjWu53yEHtXYihbmwpXtG1pQBlw4hx2I2GruwCQphKuktJaWzF34Z
5w3D+8TopGenlPhXsVvGAwkmspWvv4WePy4C/BMo3hR8XS6igPs/EHXhfhU6B+5b26/0mo7gGZ7n
U2jhW7OzT7T69e3bzAcJ43imrsnZfeqx/UWdwQPxD5MXs0vnyLx1afvomWxkOJXxIUxtFeRiHhv6
nazGarBKdi9+o4m8zyjQnYnQQoNVuqALQMv4xZhYiyQSfWL3NlNMhrucOquJeCRqKvlGEfi/fpwC
Qo7FsmSM8UpVxjhpvsFn7Ef28yLTkdvp8iV4X9xNar1S+81bRNlzumh6U2hgYcCJkYHtvlRcroyG
bG9FLeHKnMZ5Qh+m/BirbynPREr4O5gXXMfC6Z9xh+NP6WQ/JVX63MByU8Dcs/5qPGT0JaZMbAFE
wtWyGFwj2BRfGzbfLCZyrSHKos8YCCGm1txhYR2s5pgtQwytfZi2BNBhC1m/D13y/l3rhs29LF20
j3OI1z3gLBQNNMTzw1hMCdKUa7UNeopm0p4o5/NfJsfjpTYdeE3W8L3R1+NniWcl5MbOrch5Xo8N
qRhf1fvZjTzeXSB1phSCo8jXHu0CnX27C05hsJ1byGww/uUx4bK7QDZrjhRX1x5r18d00JY4xJ9N
fyZCHev7ju6ojUT6TDY5vnnggLCz4qwFOIlw1Who9dWSWrIeBGsNi1L2r6KsvFGYB5u2J3wyuplv
Dmsg3XU0EiKTnSUWCDzl8X6HWiXjyF2uV3v+CA/EXJqPF5NQtuNCATl3S1QZee3xb3SBfF0UeoHw
G2iLhSFkT2eIYuEKqE5lEmVTJiu/jFA+FuHousOIx5gQIsrGF8K12mH0qbK5gx9xgd47vMIdNsI3
AGwJXNJ5QcnrgeLbb1YftgwKbTcpO8N+3A6Le0Vk0vojZunbciffW2zzWi6+Rl2ut9aGX/Ry7ahL
h8tvhftcJbYgw2K0WVh8v4QN7uNtOIf0a/lsx2O+3voHXwVJHcLvWhemiDmqIu6bO0aoxkRq/Fnb
4CPXZDMjqvH70PcC2EF/HnE+rdHiY+TmcVFYboT5mSoBCLC0W7afhS6rbwTBOuPjfaPXi4XxbtZs
zImFYhwG+kmMKz5el3QufL1t3jmqQ5ol0If46Ykt5z7VI4FKbuFa9asR30Ch91U6kQdVy1YRPrKu
jrSSZT4+KykaJPEuVj9M1Yiv9QeEG4Wf1rAsIKWrzgK7IUxSv4kmZmYFrteHx5V8ilPe3vw1gtIh
XyqeqjFr4kw2ZXtRbTeaLB7H8xwDL/Ixm3qg3gg7l1qjgtMEd2NAE3hUVGFVNq4EOUaNt4rhw5qT
88e2p8h7cWtau9PGNdkxJFpsqRPZwwap272Uvrk+QcKEWuUHO51953TtLrl0CezlrKOYR2CjocEu
dX2Ukno/UX1OO0bn39mlM6r25JOjDiPVU4TMSwzkBqHnpNsmAiIp4zxGLNDn+KkigzRQJL909IsN
7H/NgaGRDWpqunhT6eDu3ZoeEPJPT2p6gk0a2I2VFuL3WutIDgPSaQ9Z3Hus3MZRPp6v/WwtGbY/
GeHvMVfl0ocRcGs0lfXe30qEuqHJb0HQ0+0xpmJsIlj6q3msj8lOErK7iGOiASV416i2StFANLU/
CU1Np2mtE3AMEg3uUpb+LsRek/IHOqMqNz0RoaByKS8B5QmOKbK/MU+qqsW/6zjbthYEOtt5FIjw
JNJ7d2MQV2br/YzxjpbjtWXKg2gpUvqHmShenHa7zrTbKGolzkanzQpPbUUYwj2uiCcnEVHZei45
22QhZ3HXfj6B1pBsBQ4NcrBVoU3BtjkQFmbh8WFeXHlAWaJ0Qhz4c5CqDndLI4AcxxXogaAuJ3+q
UCgSPmogIFSQk4LEgZv2mKBACBYPBb+ATOqahlzZQmgStV5xVxmdLL+7VkoGPzBRO9Yia8i8B2Vd
jmXz1ekYOO/sJEIjKAjGzaoIT2vVJjmyl6+Q+O6NbqW9L4YLow13N6twxj+Ho8Mm4Qe1T4FufnI5
1fDkzIcshPeFleKYl8Ry/rxEIRrLvptrI659gSTJuqSAXJDnwv0uKFEBIBNIwHWgOilo1JAPsFEa
w836RjY+UV6MOGAErwNeNJZs0Gl59InoqNgwmlaJaM/Hshmio8oJFvCb9/RGmMcmj6VtObt9YQRW
6aMC3YbNW69N48uxc9pOI/V9KfGgtVBbVjq3NXlqo4gQQZFhdICKz7y2AmOpcDGY4TUH134uisuA
1aWYsvb1AqHQqyLG6KK48U4hqdIA0vnB5CoIRywI7hCurDRUn8wQt+4Pb98dLmNez0Wo90Ces9yU
1CbxUKMmN6MlhCbGsDItQ3+HdAHPRRp3J3BS//DUeba370DcJJdU110N/cumKCcIAQFcqfvMmUPT
OdkTzh34Z3rBp3uUKkTDjC1PesD0aVBEXAbVTyydj8X2Zf5GHyW8lmkn4oTO9895eHqpTxN+aOyN
RYzvE+kWNuvO0xO1tNDUZAyD3aNrDggKRDUjArdZjgvPYqGFjmjo5vUdkG/nKdXARKo+S7M/eZGM
jdyvZnsOD7AXkoARXp9Rf7tpCVc/U3jh9Q7WvM0e06LvgooqNJo0jlwYa9Yyc0yVErtPPCIMhyDL
xUGhtwGkskGc3ihspMwKjuaVTGvhZC6XwMTm/6fnuu9AwQMDoN6SrmvHYs5Cl4ZIJe3N6piPJibH
Hg05BKEm1PrvrRV+bt98LhLqx8vGUW/3qIeUlScpmzidQxmQ22ShXkshsVqgyvSts3sHXlNTn33y
DDRerw0EaPZ46GLuwksIs7quqNLGBgYiGWd4UzE/4qjdw0lHy6/Y0Xf/KS0hAiXKvwD2Cqwf+iZd
Jl7SvUaeK1zyoxxSvCRAxakfsK6531mwjn90q7kxrrqCORx94zPpdcvfa4BZmOM1lwiukbpryopn
XlhLvlP/uh408aIF8Dp6c5IZAf7Uspetn0Um66BkKhozHIyX4Pv+f8ArTDcKzkoo0x5ca63zXKJw
l7l81aW+b8RVeB49PYAycExB/oUY7NSPnHOq6KReqYjkozRNLUR6d0R9YbthBkj3dzwC4fSANmTg
l6jKXg/MEGxxqP2NCLTha/dtIu2TdFEM0UC8XMulE+4dKr/KjuQiEUHSzv8P8kMw9L/+Ul4vowhE
rqshFgFLuuBdzo6HRFM/Gqswl0Ye68tdBispRfd2fmy6rvhoH8fnq/2jNrfLNpiq8EZt/W3rRaIf
YGBFatVnrpNX36FFE7jon3JRJV78EUTbP3sSvhoi0TESUYJBhnt45VLK8q6UUi+gumWM+dK2oSSx
lx+5bzTk83LHj5v3e6JYyHEMk8SXEsThvCWD9b0tx2Ogw4U4aCUB1k1JGqRDXJ83wjOI6Fzd1f4K
Labm/NKbD63GFHp4tqk6ojYAQVBXd+Nbz/Ko8B17/VGAO4Gpwf7uqFNHpsdluRHt3XHXvBWT9juE
0dwml9KwmuvLlJzPEAXHtD3zx0F2FwDm/6TmcunMtz80HaKjpBKjc81iZAtfp2UfwI6xAsjGLBVp
Z4VrWu9W9MFKucguSWF5n4ey3OSyojASndv576TAdIas9vlhD86j+wcBInJ/pocnZXT2Meria72E
r6lEpSfmrODEOTkGJXVCAz5GWAYotpvaDIy75FSDADqY3wxpT+EdttP1qnjX/icTxUIkhRomUkof
eM12xw313d1kNq1l74kGO5suLlNFO0X+4DeRdnBbz3NCtj42S8HbYj9u805piyMSeQgOJa5Dxfbc
/wT1LXBGtbK5mlXt1TBWRffUIJbyiXZZl7E4uuwLeNNUKKU3LMEIduCWGJh7Jwzn6Tn46xOG04YG
E4VT7rvZP74ErfG3pFVnTmmVGUOP5XVXCRtYUwbeo13YEN61WIgW78r7bTMZ7N43hPSO+upMJPUZ
fAR+8OY0IAa16MqdTW9oAlWh3yLatIz1DctCrWe1EENqQVBaBjgey0xLUGFoV18sjkJag81iAGEB
Au1eJO5ju1VWs75fFyb7k53HKpoiqSrqqB+qc1+pAamN1L72BfpNpoJqkNxKy75m6fcms2+QIGzm
DqF0g+WaQoCaYMOn9Xc19Vw6r3bw5dRDB4GYx3tPJZXq/rHsHpqgMLUG40YqenrijMoHKmu7I1+i
krKay8ab/i1eFpnKYqNFuLEIVRM7YLnenylMHCaSKWLx7gqMXnMsMmHWGivgQ1UxXVpzWk+Nhk/7
A48TX/lylidxgnI6ctFs9ZjYrk925bI049Nh8RDB4xH3edytaaIrLUJjrZzNdFDXa0KQPNmIKu7I
S41j4mB3Tt5ekT+0t+YMToYegUSsLBVzx5qvMWShhZ1CYIKSX7QLYJjB/PczMgmVqQfMPd3gC77E
6lOgIKtmJAG4uQohMZJaYNnyjeHQvBc6g3qsPqmPCD4Z1xDvPRHXR1lHuOOBL1rWALcY9JRIpium
njFii4HhTzk6zA6oGWa6BbuaexNI5g7XtLSrCIS3xu/t2J+uwjng4icxr41sp2QqTIEXDnLIRlcL
MvDPyLf2CZy7Ry7CXWOZev10UQExqfkYDJiDVpA+zzjrl6v5ptXCdkd3I1tiPAayiuXut3vpe36p
UyxVtaZxKz3bk5nHVsT+GoyBGlh2iz7HnaLJic0BrMcvzzSAMKwB8Dcus4m5CT7Fw0g8x++gJ2TW
yU1T9LhpU7mr26YvwFL7DtHuCAGKhzMkLnLFESORbIVUtlx/p25z1+tR59tiJmn7U6UpNzB8Yra1
yjLzi2CRtmzVKetTd3dH9DkMb/3vKutajzjzs0QMthr57bzg1MIgPbE8Hchhg8KIetxpyB8UNr1s
zcFGYTyMCJJ3E1VlB03PLDF5gD8DiALCGJUWeF3qq7049N4nYM5MFXkMT/3JrnKTL+imKVsZ4vKR
daD/s/FZ7xGIkva1OSXesH+lpE9/PV7aMOcBuEt9pmHcIv5Nx7wXizqYzKR0rLsXRRJPZlMWfh3j
oOgZhUXsYja2RQmsFz3vnDNSBO//WJbOnH5KzB7ewinAGztA4YSy5CjTz2n7Fh4gN1C+z99pBjyB
vi+cs7nsLVTGC2oql+omn7h9zs6BRNM49fUFy53GWfdVwxLvv81qiKvyQajXG7I2nqoFrTmfqCqR
W9BzE86iKJPCM+y4wuzmNe4eZu1037oizjc0eet4RuLDQTd+d8VzCrbrSBbr/95dJ98LerxSPVh3
qMzSb5m2tj2Xv9rMqDnxkUiZrMYXEFWI5ObDh2u/DP79gUp2DO9U8/ha/+Dbq0BYfp2dxIG9B23R
zNAi12UctlzgtOa/2CtNfoaQiPrmRHPErwMrzgouAQYIDT05Fm3QG9tPCDS32QVuoOi/08vBH+Ae
7xBebQhhUuh55moy+slin1gJtSHWXj+HIQ2TvtUb7lxsy2lxtQKfBxVtEkr0twe3rcXPw7mdppQJ
97asS6Ej1qiJHuM/vZtxRh4NF+uBy/FHIfG2HE2AThiYrI0W1yCQ351GtL2xCHzNxfU+lR7rxedP
Tyr9+/WfxCampbw5P9Uen/qdKgTKWYrT4p66eU4hl0gb6YbHzmOR5jAMao7NHdcCJcxnkvBpGn/3
yuWo4POBqFzLu/zkH1aqFHgQsldeD26QQvVMAqxi+X0QsxDhY08FQ1G6DUV6p5u2132CW4cevEAk
ROXevhHN1tAqirBOwKraDCgFgyB82g+ghcX0Evm8AZQuwx2ejd4Ind7HyDGRebK/GbeM7pSsAgfd
GYQgE+NECrOKhILBXOXEHQJ+g0vYmEx427nom7OdFg1Huzbg74bTtBQjb+lsqgiI5WIkK6H0sdQ5
HhFFF9omndTF87eCGbC3Xfeqj4QRXJKLBNnl+sYvqIS87sXASSeYFsC/DYlTRxafpa8CJs+MZoeg
teOmZrfBb728fGu9AoqGkJTP2wNnDg/OSSv58AvsnGYHldafeM4T7Rux2VLFQE0+16ckUB9mtZ3L
iY+TAeL5xYlJJGo8PuTVTVMLQ+zPRpmwaZTNPBrUi1LMEflh6ThP5L9SPhQBHGyFSSSuiQ+EKbE/
NClPNBvmQJ91717zNgk4ItlaVJOlON9uJxhvm4HuMFgdR/SVYnYSIYidpk12/A1fEhV1NKLf6aq5
pFPrX7Z52uh5B1YZ0C+4x4fiFmgIdTEZFSWsIN+8aKhyF2osydxB548sCHnM90VgsUpOxp7cCuvO
uFXa3HocLiekRKPF504LcNRMx9XOr/wVYe8WxIeKrSFtzbC6iyWVaXGM+yZ1sziChvLvQcn4bBT6
OV57hmr+FtLTQOvV1KMsQNzIfIpGWIltS2VZdvy1z4XDIRcONRkkOj6KTzjfJRmXgWAHirpysBUm
ycxxzrDGneVDB08ByxApGzADjLF2VQRNVo6Gk6vpYhRJKFvPtfJHHD6fr4Vlx2cNR3eFGgboo7qQ
R6BZnekLXyxjmmVWNbCq13ZCfUGM5HAhJk+sYOskY6EmyHr1kygQwcbt2kjsNqeKFLqA5xhRAwxZ
yZp/XOeDDb26Dl6XM9RPDPkO+dGQyqimz5NXmK2FVQLs/8tXmoiPkjSbUuDyriRhQP/NHinOGZxx
zDU86hHObCauQFEQBwvkjmzby1hAxyZSDgp8Vjq+M24ZtLIgP82eNaChsS/4MKx1rzMKppQOI8J7
ZLgGQee81+TQ7k7B+SoQjwHtKS4/JV+G/sJz7VFeQoF7UMP7r751hMJrJ/vA8S25P8g6YIoS2xn9
na5aUs0YEQFHRmEdG2cddbGHEZ05BUUxEzp0HSiZm56FtCpHqhlb2KCXfc7eYvRpk3N7VE6ff36P
EtWB8o0gYxwHLWcuvGl6K9bADAmY5/MQNYAZYFYRMujRCcF8501qcMrqrY8/iGBtpgsgE0AaMxpX
3WeJhgj3K8vjreC1qWFOOAtS16nM9ih87THNbCCp8H0n8pIfscnHYgELLEut1kmDrBDY9xwQUq2V
jhJu4NoXxL9QZb2Df1gNkcH9PeZ+pSiuQuSIaLh9YzUYTl0LEnUdwuo4cp6JzxnMYrQIDW/c6b+2
kvVWEAfjz65u9HhUU1KALvQNxQH2Z3+/OTSbjkKXYVxyRJFz43LMsZLpBn0R3qQmWYHQMJatuTzF
yUOfqTFGVP9p6h1hUJ2ZU1z56muEm4/TH4zGey/f8pzwx1o8FwdtHZnQe3mKQPx7a4+a52G9S6nH
XSIMwDSp9J2G4b1hXO5n1eRk+1inOwnL3hxrhC0ZgTc7LYa2XfR5ITVn2YHgPLGE0b/r2LkHtpj+
FQjBw+r6uH4AVOw0NFV9L2nxyapMTbhN+mnQmP9oRxEbEUZaqujYm4mfyAVwRl6VxkwT4hMx+AZ0
BIYEkO0zhXFvIia5pKfcCbXASthWIupiaYOkNUiH7xceyVOIlXTbkgO1OAsyEfANmTZ7Y0zjCKyy
sz6jSZTVZw0hFAOaJZkw9oa5mAveDUMQEFPi9PFScb0le+0I0acn/UxRF+hmaR7Bglu4Fsb+MEL3
yQBRm699a6HwagYzXmt2mi+u6YR4C2C8Ui/WTTCts1SAD88v8u+sD4qKlGj2u95fGIx5HzkSUQsI
Q+TT0UGM92dTcKZBJ2Z1jBnQEyODHHVICi0j1NnLjTGlaiu/3Kl20pXqA7Xr70eqtdUD8PsUrHXN
xfLLJ/qnewtExfp4QNCs67ghy2mot8QovPA6Xa+mGK9H1/YDFnln0GtyBu7w6CR+8aQ1ufQzV/Bu
xirB5bQRkkjPDGHYWCOy+lvUWPgt15JV3+GlWHJPf9WSWkzcUy3RMj2E6xs+3YT4bCrufpfSJkzu
mGG0lZTn4OJyrC6bCR5fA9YKdSqXINbGeeX5XduCvOoKZcCTnl97HVjLYq5V/YVrn6FflqZ+T5fM
5HqinT56ikgopuzoGOJNqUqI9cq8Hm9M64SJOhjBx1gtLswwFuVHnAgfXOED33TK4jdhNnC+cJpu
/0fmmNd+qxezVjlLuGwUIiGMvsBBGam/LBLlK8TPkgg7FtCs+xalq9ef8YwbMLlwrgBi980ldLQm
h7qkeHG8m4v/P+OkjPpxD7ah2gEe9eibadwOLM/tpOTE5o3KNYjIuLAlz60v6NzdLwmUFjXjfooR
bV8UdFH55brQoD5ygVhZY312pT+Xha7OQm9TTM1uSTKgfWAxObjZ7HMLkP/skjS2uCdrJn6A/dqV
wGIOCVPBUrfHVSMOnyRuHJ6GlsKm/I7Fikw+2y3ogjuXpEpEarWKz2K3i99PKwtOt3GDVFh+Vsn2
JMDx84m7PXEbMCHgYHYwWfNleJ/4mXdSxEx1s3WcKX00Fojbb7HPuS076MI95LKqElGkn4NpY2/i
0tuD6dorErbdOAFpi+sHmRwjEvdYkGEch4UohwYBKM2XP014G+GYmCQ/lshGaZzZquBfSAVjtJMP
e1hkHNNxruCEQlc9+kwBBBPqrI9+Ze8E9ngoQf3nCP8nsRmmLwgwgTOQQTJUZtNx+kjAoXQ2+otH
mSD1M/RPxvLLlQ0kwEmfPexys4d9Kr3gHbyo7OPiqeELPnvFPn+vYiYn9U1sBeuWn0XzXJcHtnyU
WID2zLSFBI466mShtkLuCa7IN2y2clIbJAQWFkCcjQBbVd6HZ762K3RskGmC9omcMzk4IeSzhFsB
NOB22ls6RVW9OmY+Q9YMnrinp0y+x+wZq1WoTO9wJiw772QtRZgCcg+x7r7a52jsF+h51X5++IN5
2fExqBjZsvke9bawCEDqeR+f0HOXJSBK17vEYcV3PSfHdKwFRhRJ4uttr9l+boF7POkFuzcLyCu+
xJlkFPBNjv4WkeETRZTeLt0WaysGhpYY17r4mXFFWlXRiCO4orJCvPf6Cc7WwOLqiUadwR99W8Yk
KdE01YSfj9wxVxnSglqHNMXA4lKAS05cZVGBh8ZODI7oIjV7ZU2TdEjNq3yvP2flEN+oRLkZ8m+j
wgIQHgXXNRbBlqVcntxCTfmgsn3lMcjhIs07Q9U1pV+Kpy+qYfEcLsZN0s8EwJjfRCZB6e5d5cgY
tZ9ePiGF6bUdUmzoGcWa0xrgCwoolkMVockl2mvVH6YsgIJm/D6ieVpg89i5NKGWb8VsBaLY6Hy7
iamQX06qjdTlw6xIr1qezWd2CNNi/H+jGZqWKy1K3y4KbZtUzy7V8i1QJ1N/jR9nILmlZg6Ney6h
pqMCmt6QnK4lcx5fLQPaym52dRUCHntmjUeqeCUrKXrJKaitScwmtKZ/eCQz9tjTLJuevWRUUhMO
eLGmATTgnE5EA7bYLxOXgwyrsfsK7wzRJaq64y+6uKUFv5NYkP790BnPillIF9gACr3yEnZNYIcG
wffJKftHN7aF7BRJ/DVP1V84Y6f0cMqY/pheMZMUm61kPrE/Ao2fvysWTVZEtfHl3S9RQwPEjNn0
kR3T7dRtVeS0OztSLB0Al5YRC0h+FTTx4hO2PM4Rie2NI7qI71Rp1xZW2Y/HBlynmai1GaMUisD9
oYeAlQS3UZGzEZMkvSUdBnboiud4zH8YGSXzzO3ez596D6WsuZ0xa2mz47TPdK9jXrGIKntMPLTH
tPquUvJVOS8yCyKRp5KduCUQjmJXx7O4Gu6fgoeDVvS6IxkyRl0ZOSvdvVKw6L97XFdxarqFK/t9
0+T2+rim5W+9nqaLepnixtaGdwBWb4HHevG5s9sBdfSxWtQH4XRm6uiGLIBJtSOh7I2E8/cKSlQG
S0QxP2ijMCmjcrmGSK6xTgB7QsODoxwG7GJrgN00+L7HVSK7jYyPSTFWhH0vU1ijt6fuEqNW4ZIa
sjJwWpQgjYc65xjwYeTLWA3L/YsnBhuZ6NsIdwqvoC41QHJbs8kvcfzXIqfkX5vkzEdW09w/RUuK
gw3IgNsjl+ByVf60kCNiCCEwoD2z4Bz4aG2QWaZY/YNN9/rw+prAD4R2Dmg4HLvQOhskpjqsKZKH
0C4ZELETczTuNqf/EzLHKL9DIjIevKJop2PdddD5twrrpWccxreUfHtM0MYdNuKzUJbkLHBirws8
m1dnKQw2msQpv5S8NokabvzilcwqRrDWLOKeGzJLl+pl6godTeWUFT9xEd5DJm5cYc2a+iUTvj3J
/UFB/3KaVheA1Hp2hbTw1cdXFxS9pqNvcT+Doc6P4gszjywL1EV3myMvNKyedJo3fgZ+6MMQCAPy
NulImo3Cge6BBi/pcXhJOdSgJhF8X5DdkFh/AK2rotDMyFtHwlr7SbM1+C26r9emFPsw79dZ6I/+
9tSdLuzSiypZ/fZWKEaiLNAE71xq3toALv1y75HDzg5NhZMMiGycdlQQVk7pC3YRl834RX8WNMT/
srTKGjbK+fMh9JSOwVoerJBLoJ/BeGLCqx1POMgVwUPE7AjL//1VmiEeAF50HKOSUGgD+vboAEbG
bwziao+sdyAPniZl0lyCsiAEAYIrxU4y1wntR+sBV6Uz2g0krD6R4k4aQ8faOw44S+bIoEJag+Jp
gaAm7pNMEkuJf2/aKONd7aoVa3REfaKnjHO1NqWhFeRQAL32iqQ91PgnSBDtKM6RYzaATgKBbFRa
7r51GqIxPisjlb3rieaC2cLqJ5XF0m96QZ+0wS6VgtGe1EW9Ag7NvoXDnf/Y5vtLaeyf6PKdZHh1
Mpjy+hroy1Wy/t4Uo5o/79Ju0AYa28rOYkLNYnjVKtqdscEq3H5COGhKM7tZuubNNRBnsJav48Ki
jk6p0Bw9lOi9Z+Bmt6pLtTfcLyMYQgrNVVvbCYWFKzK8837DyEBcdlTuYy2s9eCOvTFYtgpBw5sJ
ohI8yC4MrG7l7iD6V9nj2ZBec7qM28HVJ+51gd/AxEztw4ezQcJkLDEtfB8cPqip9K0Inr2/aUWq
/xBNAFOrG4MdmZeq8q5QPDjJHmC22V4lPE4/1nfPJYTUH/Kpqka6udEoksIhMES2KKvD/NBlyvm6
TfVtcCJ+JOhXT5vAa4CoIVtDuuGuIrdlTHdi256ljSmG0D6/kTMhBj49+b2++Fh22Sv5l4656BHX
v6LpRsHlm1Lzd5FC2QiUNBFqfZB8Sqjd2CulsGhBxLlNSPjSxPqHhCrDApErlpsQUtHtOoaqWWKy
cmjTsxbqNtrL+ZNLcnqRgpiXc7hXvy+ZeMXWi4df+7ty3orT/StC7MQLinTYhCaREzz3YlLdaIsb
VnPlTaTFPsEAFCuwh8B0aC8rDoNlyQ+4mRvnvw7b0SsV84qA34IxirtLCq8TBiADDkMYxuRaRYyx
GzOXAAkzxKruZ9JhMiYCsM11rbhFD+zbTbS1W4OgCr90O8Qsg0v9+OgeRaphuR9umzO6gxKFxv69
Vein7HmfQCVUl91jYuNF+rMOFm61GfrohvTKRQw2p/Kc78smD6a1GOs9NQT36WXAbJdACgkmDtML
2MGMafpFQYLzJcVGv8YBHkgWRYX2t4nqAfZ8OUl+j2KQMEfve66C2xwOaAIk5FycFLr/OsVrjB8T
VDIMzLrcc7dPgLgXugZ4C01vOZunqV/42VqfG4fvHlnFLJKAHC0/BDSw+CS1IMn+oYGcVvIHdwg/
jyPBmeDVuSvYhUDjZcNFvg1RoB6B/gQ7Yhqsy10v6D9K/k+xYLpXPbIDT51oGcnrHSSzM1x2wee7
5dCB5xD7T7uAiiRArVhb/EZNTehR9W5grkH70UruGZmzFamS6cJumVKhCgaREv/GOpvRcOpq31++
N1nv2mN9JDNQewqYhQPfzmw3Ur0hXNwrWHzgUEjyx1lighxQ+1Ya2hiBiXInV+ytPxNd/VVq7OYu
AgULM5aWO2iB+L8/a8Hn9U3k3aYhVpVUfzUxhpBfeEoXOh0oRHRdyj2dB01yxepgTv4xfszDU/LE
xi1JmM/8xga9Nx2ajIGBclRbGTE8i5juZGa0/RnXWEGMbHg0BbqoHFVShdhaD/h8Zb0e+LVtRiDA
WyBxop/Fl0jhnQvo1hJG6FYAHqJL1lFBIKRIMofikat3sDQ365zXw8n31qiHgjNxPbY6Q10eAb5B
4QxshUXQT9W+//mbhNLWxXpViT0mWGfvD+ZUYyHf9i0CzjYwP5wEzalw85pB1LE0mzdvtsVgCzDd
vyQVu8AuS/clKePVqd+Lti1gezXm86DQKoAzfuh2VOiK8/IUK9v+AaiC0Svx3LRRimOcICuQi3d0
Eo+PaID+AJqETGuWXsfNJGZ6t7tOBkiRfoQWMxXlIMmTY6V+MkL1I0HfxSqmOoZN8VeUQ2C73imH
WxgWtQGPP3PmaEUUZSVZA/CMeztuXVaa4uLs0BX/K9DM2WC/I4vSLbAvWm518ixrY808PnsVa/k+
O9GQakk4iRBSTofkIaD02HDrdPnIKxAm6kC4NY1/49PK69BiOXO34IPbMbAzqSJFIsOveDHzp3sR
E0s/aizTevZvVJch6/JXIx1X7o2Es1GxTzojyTZ6bQSDRQVG2F02YQfDAOXdGrO+pZVDcd1lxMK6
EltnSeEhn4qwwZaCZsQZwoSWAwfJKDuNkcgalvxO9FCaEMLIeN1SOd7muybaelJdHndARvaRhEFZ
P279fAaVzYoZ7qRuXdAW006OhrAL8KpFkAo30yag9mfQLtV8SC8KKkC5Gx+wA4lE2ttlvusso3Hy
ktEkxEbJkMWIB27iLThlFYp/+jcKSu7FHxQJaBYkr6rzmQOSMkNaJKSsmxUmfSzIRtp2QuwmOWoH
+fFLPmJY/Bf+mGDQoG8v8j76hvxKc2hr0VJs1KyG1a/ZH3vwfpk6vMkxzGAIUVXW/AhtAtEC28W+
JXgiUdECdrFbqULwZ1uVwRuewHUWWOpe55ab3nywMtNsqF9hHpt/fH7RWe/Ub8DnBu5vbKl8pL4T
QbgwlKx9NFJvrHFYMKiWWjvQWph1cJG378WPSO5+5jt/YBe2HJMvpDL4WA1Z/jO8hPI45ozEAc4V
NASzCvWtvlqEEX/a4UqMe+AfVqA9qN/aFxcMgISAOIRh4Nx88BH8CG7wSqblbmTaJKVd3KQpK8Ld
kS5tw3OwrXTzI6g2ldpNjnBwKaufLhcRKsKJWtRQhm3/I8nsYJJ9cqRdgVZoEuGhnC9/HuCGt1sH
pUwT5TJVn0NiIr820CtONm2JTPmKE2Z4ccTEC178/GnvZ6vnexwE71wZWLn/To9x/020+LV96/fJ
0SU9IShF51vxmxszCdF0cmxltw61lf7yKzxKV/j+rniOkoFvslSP4AYlRDlBTyft4UwAUhC8XugH
/ibqZtElcJVEFR1Z98bGlAGJ0wwUIfqFq9pHAlcoApP1sfyj8jJDCoVV2lW42L5ldrhHd1q5BmPh
my2ft96JyA7fUTPzr1Xpowzdjcdb4wtSUMEmdIXW4PN5jAf1f0a6/F0NgOD+0aUPUbICyQ93QVBU
V3qqIkWbEGFEG9Sxi91Xhl40c/7bZGnGYDV5sVezyJfuLthG/6aEtw68KgbuznOi2ZH1cZ04gM1m
wqXTwKJgbw1A6LOlfPxPJQL8/EF5BtUHHgoNCmwYm9miviIw9dXiRzYyeB3tYJphL8Qv5JbtxfUV
aKETJIBWtufJaYHnrN8rz94GUlCCODDWgj9A+X/2nx/NuUfvhZwkUVQwAdqNR9QB3Z3i8DAPUY61
FnSYM9FQkn0sATqJDLl5MIv5B/woagzeWjT3Y3ilRUi0w2EvgH6RDom9G1FlTRqrMzG5VfRfqJ9K
HgJXEs1WaVrRHL+0n1cAUff6VQkoNoBu+9QahiP6fLdndf2j0YSshje2TygVm1TNH/BcKCgPHu5C
TY++L31Q7kw9/BS2XW2qPEupuhDM2cl+/naWJTtW8p9D+t5wJSGoVg+8tJ7BExvUl0KR95JWAmMB
exizEvj+uWkTQET1xrpgGYJQ8SRDBdV05pBLPjcwEifiDrJeBCzihzrVpbVO93rCLbNeb3PLCluB
uqcwS3P5+Oe6Jzi6ReMcHmwsaWPT07q6BJ6xtV0P2pUM+475V8uZirJc5eOT4kl3lttUNvEDkVOu
oxiQshOxjZ82KBEYEEoC8U1fvQx+cPnauKHWzhcqx07ue7uQ3KBVzbnEqvVTNJwqmKPKlWbsDrLH
2rHrhg==
`protect end_protected
