`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 27440)
`protect data_block
td5QFuuLITbKOtkE3oI0mGg81uxEpl4OzFN3dx3S1ftkr1FB28AsEjJ1JzlMER3jugQ0XxNHpZ6B
MQSg9LCC2ub5LNwlhvbYEAYYqCK6ZgIfuBIOXcuFFCv38YT5eHX9DfFv82XjsC1Pwn/wMP5pa47z
RkUFjUxny26VVLkcvVGgbXqytVTR0La1xotifeEjVydMrmZYXl4iOFvRKQR/0EgKCt57YTzbnIky
JLh6DJGnFSWystzWEN9m+rQ9crfQxmwyJpBFPQ1QII2LokmEvRvosXL5x6beIuBaCOKFsx0OiJz9
Fg4/beWAucsxlrFBfY/gzEkeEt5K/rjVYPngc4Ri0EFvyyEvbMTir4tc8QjEOnn9jRDkcf/RS36Y
ET0rvaIgmsWQK48R53jYh0rnb4crHhyLle/Ld6omDaWj/Xc5XOaz7Yz+sXCm0nrOX+sXMiBfcHEx
TEO1mvpCCwn5Ok+cna2VCI713hpjMb15nBwhM+WoRwyBnqoe5vDKSrQjaVTuWrY2fmHYY68kaTt4
xpCVojqKrWy7a+Wamu1mLLgiwdDsDUp6PYRObD8mJ8yNnRXCxYEDjTYwzNvwRyrh01T5LLpJqoAU
sbw/DUe18Jk8+2esJjmEp5zF9PntzGnMXA9+Fvu/mFahWHYm3bdAKTbe5ela8KxKQPqUHsgyQM15
EnhwMs8hnDjruyhXcCN2lHx3DukmuLXdqsrZICknWiaqWHUu99PPdhun03ATDEtu++uKQzw0sW09
64H6tdsC94v7nsQDL5JTFQqvsJCDcgqSS0n8mtSh0BeDXUI5mQe9umSEdBYNNA6BxUtHk9iTOOq5
nBkxTVY74Q6qr9lYZb94esrUFHy7pAYNw6r9uqSAWHq+oUwopvBh+pGHDI06L2Oj/Jtap+BUfHsU
GqdxBdAo1DfPL3XcZlxzJnc8uywtdTILhafZn/UwT8nK+LeSCbCmzTn0oRagUB7RgwZOmpOWvV6l
BwrNUBDfWk1f/ME8J5g+j4FPYi13d5gGlNil4ZE0mKQE1W5dHoe4+h/JYQxBwYHw4ovf3J6NwZYm
fpdzNj7YR7ClMGtgHhVngXMdbXuI2RTgvpJEUcazZzUaBmtq1o4HDItWBAZSHE0cVJ245qMiB4BW
/3BFsKtO324KIUVUgJiRDgMOI/4ZuqtQJRNrI5bPkv4u2Ot7nKBrYaXsZ83Zcyc2Ia+MZQfGNyCV
xeVhpStbJLmk/1gpRMqA0tJ1BDg+7KBCYdbqIT/g7PaIXk0x5eHwv86wdj4cMn0b5eGMF0whx57h
Ofkg1KV+Y8Z1GfYG0v668LTF9lOIRxP6w8+kfVBYM4vBL2b7cMiRYknhjD0x2PUx6iGZL7yL5d2D
PkIhLbsNMJV9eNZHNUjeUP7jEVQNLjfqdBhmivvB/lpv9bhgPvTfDyxXO8gsI93LHdC7QKaULDZg
IvbptKSnk+7ZZFBpRQR14KgoB8KtZZ1WYVDQaTOG/JNW1aKr76M6wgqTJjdsR4S5xu2fZoddBIge
xDLtAloZ2bLorOMs0WRXHe0/H+jER0cA+zouuV9x2PUF5VeDVeaCloQ4vpT9UOo4wwVmGoJD89VD
iPWQsLEjyWhiobmwvic+xZZu2HAwFDYhsbplu156fr/tvRbxOpaRHyUp7aGO2hT5o9ozgIH92AAx
ujHnIgCzONa1i5y6WmhDPjc5c74YRxJe1c6E2l1obKOXvrfdVpmnXazOiqiloEP6lU7VBEoSK7sg
1GBH8m4zZaLT3wrUOCZit9bA1gLJYRRC6GIOzJMlqsVEW37m9bGoEZI2yRjt26UJak74AmZvzNPG
lZinFl+r552cMJptP2oiVF+CYiR2Z06PNX/+ylaLN0Kdl3mylfcqSrKGhYn+w6HdoSLh7UmJH5Lx
z4FA2bZF1wjsKRYP+8j2MUPu4suN2OZ/idT7ORCiG0L8dyZVniCTeKioH7FN5NNk+R7infm5RUIv
+YPBkd5pxTYqrbWfBxG3AYDg8tzlrAUletO0pKL8sA8TA+Tg4GcOLI+u3NJ6vXoevXrVEdGIhwL0
nJZquKUPzHPSWaYlrOiTGHtp6bu4cvcfNJa5Gx82YDV3mHX1UIPsy68odnhhzHf+5AxVclQO2TDo
JON/knNhKALNy8aHdNJV1Pl5GwY4U49xY3+Z3AoAwxn9z3GwLJbGgSLUEFFFb9AKnE8QEGy76OSf
3YohxSpvLynF7FADJXIbXOjfR8NCqXHlmZ/FCLvUFRT8BG+QtGDAQR3Kv9XGECWw31lmhtE1ch96
gSoz2rnFpee3G7OslLRAQsfIHrzOJ9hqA4Nuih445q3DlQhEQ0EfbdYcmwTbMVR47lsjZHt6WzF/
M7DZD5Qo5kMAzrCgpfTfJHGIGXEOhjk9108zSckoDBgDSyFyzneHjxZvLD+g8i34s4muAMnexZKv
S3vb9sIfjhYCbVjHoF8eRwikZoYvtZl48DsPqnZ/Vc/q0EPFGUt5Pe4ZUJAe9BsPJRXWOFhceR4t
QauH4t/phDuuFzvexGNJ2DPcZmn9d/9tKk/H/JyfNiQwjg+rfXdknqzdkdyNCuMjTZ9esKiPTCQO
y73apM+iWRHHD4+FHaRuTZf9fiahWaz8O68wG+dqOOuLqbbQPux7c7ZR1iFR8Os9CiY1lPfkk3Ia
+CoZW0ThoXMJFowQrFHFdhOqSpJE+1hceQ18kQE6Gtu8OgL/iuArj+2ebqEwT8d0XRYUDr0Evi16
A9fzcb0WPmHHnNYzvB3X4aIlYVeNnej620gFYFsJKmzFK0oO7duGZjkQHisSzgQjcpzeApJEDD3M
TzzTMXG5X16IavxWzZ7N22nCPsnqXVOEhFrRPAJgEdqiiBd91M4ImsDMDdgzG07+syrbdkjyAKRH
sNBj6tBUMj61rbZl3J1ei0UaB58LcV7yywxqICg77PuSYOT4DoJNMjLX++dRVIZKOwwniIHBIj90
5MaZ/mxZiLECrHzZ1FmivVZ764O3/Xx0EKBfpnScjuUBnCmWoVTIesUp7BFhZ3du1I1wl9TTAyrc
khww4z0ZzsFigGvyXQuyusG614X7uAgq4BoqF+xhEm52GQx9yD9WCsYV8nmlgBKCSep+be4N8xfC
4y84hStLX2kC1p/DTOFpN+bcxJqCTwVpCQjYomp4JenTcXtqnV9DCex61yhQl9agW7NWcvS+0ccs
tdZN20eqMssptd51kMPs+80SiqSjQ2hM4WhZqQpWn0a7kekjGAihoJbwFSvbEFPuflI5tNiwIGge
PaV7R4WNn5Fg5+X2wEr2Lgyd7VSEhkw8shMZpoI/7oKYgoUYb7MbOefFl/B4+jdvOZqOp01umlSW
sQQcpXgn6Y7LeKtpI23kUqvbeo7vhFUN2id8CrZH648XPBS9hXGPjvnui9fQ/TKhnMqRAS9X2gYD
c9ZK/2lGPKM79qV8FE/DA+MnTz/UkfFGTnjquExm/y/P3jSv+n24BnKTId8pKcn6qCOyZC/HiVcY
ZaT4RLF9xDtQdDk1AFV8ChD+FWHKsCo2E6pgfi0LQPLnuvtjAUQ6tCNODDuNDinx+ot+f6qxbAyG
LCFfPycu0740EYE+u4Kz3KNxYQN1e5lR6QOCsPbwgE/0yx7ftOqnIkXoMpEhtk23lpk0Gyuc/cac
AK1wixid6Cz5++viAQAcb8FL3c2EMztcCxCawVyoA2eQjA9G+FyEt3G1e4T4Uknulcw4NSGCG0VW
ZBJRmbySLNyW30RBN3bU9+viJFeqAV7HZ6PzTN3kJiAw3fvX16NtZUo6ifDr5SKOQyxl0spODQLu
cD5nIi/tBfkAFfj6pIwUjR5CH3QGGVccJIeWF7l1W9xWjQH2raxnAsikG3V6bs+vYjDkTgDNYQW4
z4AWaF/DaZDJtYn4znHiCjmugLfXL3cMpsTupESLOu1J/aObvzFtBG5tzni1Yqj2utkOQTBavqM+
h06eCX35CXPZSkJt2w4h1jxsLlhvxp+PCRzfiTgWpdCPHSxDs73GMRHlhuBr7Cjdm+bo6RN/CL1e
oCmH44oryHUpFNwOVTHU+WxQJ2RThuhOeIoq+KkvGFEjMX9YGyYTOrvEX0f7x2ykdlGFIUNPUHtA
LaWsspfBdV3UIkPrVOrx3jYDVY1RHj3hX2N9e87ALUcUS0iD9Mm65kjghYxdw/MUjCNGlMdxF0JS
xyeqyXwAoI590ckShITsxfC+Gnu136+fgLR5NqL2GIfwPv4jF7cU1wbzXtUvHj7QJHa3X/EU7V4x
wQXK2pkAepF42tNXzfHf99X59uVRuG+n5uRqrocO0Mf+pPuURvFQVsOoCKGgIJlxVygZyjGtDkwg
AhqHd8E1/t4DgtxQPegOH++9qdZg5BIrjDBf2rqjkLc2vOeP3Auno68zw9ecUMnZ/D8K0rel0NJc
Beuaw6KuCmHJs/198aeJaqtMFwD6MhdJBZEiydjfoYGY/inA3HJuTIKyYGiN5gVPcEeIIq3gmcR+
Ix3VDjzWdzqyso64e9dRd2eH1qD0WOKB+yHmh86jqo0MR73U4l3bzgfT9tV1R54ClTv0ccFItVJS
QQTnobJIwoNfQ5/e4apBiViGYs9Q/QjcTRmONai0jIREdGLXlEGbszDQSvKANQ1KL1Uj9WfpUsTF
M2qqMiS1Vh9LhwNrcRb4KbNkKBLWMR4UaAVCt7YvFU/3JE149AzAHHHhOiweI9xlijbpmcVigI1h
NIYzpsmotwZvSr+zMp7sT6Ruh/3mosEEeaLAaYM2qa1urHn8cPnsREq8f3AVQFt2zhaCX1pjAs60
kvPTJEqXyqzrD3JnZmSFuPhg8SHqMUGmyDYeV2363VhgsWIyIQwgmseGSnocm77kdLRvUNXu4F3M
XDitgi+NF8mwv81MdtpHvJ7kWPNBdbcTBIUzF+8I2uuoJyZ/blG3GSaYoCTYT5V7IRQLH5+JwvId
7QBcMc+BmLsdPyAVRlEkeIv3kKs2GIJnGPxNFDUbi50Jl2ppi7vAJnrJV9KV3btEVher1ek8Z+O8
1rWaUdJMsNEB2f9SxZ1rgegU/wldXVmFNhxKkgjeK2U+pVSNvWQKH8X3pLLU2cR4CpUSdk0iv5Yv
3TPrKZewL/gYXocbMJJjc7p8cjFBEFMiEipD9qqPRyvGT42niI8aDtv3PnSRHx3dEUqrT/I03fqg
YADdL6OAhJBYfbqgfDHLbYbuf/Hxi1jgkqjgYWB+PqoS9jLrAcqbmH6IAVqi+HdrqjExx8JggUfT
4ukU120avzk2YuSOcqwwA7erJfxydynNBATtxyawET8MA2aeZUekgk31JQPmo3P4d3KoQsisQzKj
V32T4FTGEeWIz+6zy7QXa7lhP/6lliYMrX0FULWQ6FYoZtcPgS8fjs41v0tuBdOegKNm7mxeVAXA
DILfjLv59sCh1sje9/2/uMaSo+T69mFpLYQhu8cKVUSmVaal7qKDInKHdQSY7ZueKPjkzJh6ioWU
9FhZOyhj7W7PLUquPDI+ZzBr6gK55LBe/rWw2NZQqZ2cJz+oDkg0eGCrZ3zN8mHaicZRE9w63/lX
TeIq8MZNqVJ9MU5S59/RlKhh/8VBp405+p9lprX6D2FRibqC7x8WJsPoR3rT2kK7UqltcLjwClQq
oAOJUhW2zG7x1IFk4C//3qhXVxJF7PZbIaJCsigLVbRs8fFsx7VifZRXC+QYanm3jLSuW0tyHI0j
zjFIEcqnix/AP5Op7E76lQapUthEVPvB/lCIqD+f3wBGPPzGNh4Z4gmuZHdADiMhZT5IMQdxPM6L
f22R0fdBvf+9g1vTJ7KYL1fjtJuwz9AHuLmxdcR6DTxcjky499dl5UJgTKsA2UhvjpLEJFU72t7U
QREStRUjCteBTQ3aM1LLZ/izG0m80F8ZtpOHlP3rEHzlV8mbQiag/q+bjs0uZD+u1Z4PAObpKk15
ot5i21/8zOelcnzLd1Ysp05fSwb6JsN0ONjCHJSjfDGKUoPG+B17Zsp5vOLvZmYdzJkG+qe4AbEO
M2f+WxHY6M0KS8INZrxhI6aoR3om8SiNWR4nxviZdQ97/UMG9C2k6dIEd4rwGsp25dOXylD6oyp6
pUFDtNm8moadLmwFVZk3LGBIO2eq+yPBDZwrNEHg1IEHj4XyPJ/DYTdqaaRDPKXu+JjtrppK90ca
sga2SCWBV7BJ4tI+xi0pafz0TbGSXFsLNUt9J1omyBKXxQ0oez8UahtyAuw342MrsA779/ZI4tkm
ZVnErotbnOBPNy19Y51hyipfcQLeHcDgDGaQ78W6TySL41uA47p791bIFNy9mlgPD0h6XNnhz511
o0MMLANrjVtzJWceav1WQbnN6cgQFDBiVrxnuoByGIX33QV2REky9hpknBMefHRU36Cit1chT6W3
wrG1wvO0h7QiRkN3zG8cc3p+IWJaBGrvmkFXJ1YuCNKwJjbhge7csjnAh8YbpqMriknjagUv2PIM
+fh9kWT8OwaZ1GN+vyENb8nM7IzSEtQAm+vDtvf7touHEv4qgzNFTtfys9yS6UrieZfVUV/QH1SW
v5xq4Av9EBRkLGf/RTtpAXyXnyAnaVgm2tKJGYbB7l2Yt/eQP6YhjyvJp1T24fZ0C875Hq6OlkER
2vEFKdW6y0KrGRddLQQ1LBAg0gYvdthro34cha1pH9AH1PT2vHEub0d7kh5gJb9NMdjPuezLBHIm
9R1EVBNz57YN7VbK+y5bLnAagJG9HKQycfNbt4ev7dZjhHJpslKJnabt4EXWkf8tftwC1Lyf+880
/c9Qb0qEYTDKvUML1CNFusgX9EMAUZ5IEKDGZTdNTW2y7Un8V09FWVT0AlATb0AjYgJhUTSo8Xih
BI9TjOmis1ZXz9JAzVtWbzQSbXKcfDj5FwDl6CxpWzqQwczkb8cq9Bw/NvhoLBwPoUZ+tnYYt7xf
5LG2OXl+Y3prCVns/3Nivkeqnf4Vy6SLFklbzQXDq/2Wln1VNtP8shxORTbu1izyFUKX00eRbzdy
Xnut5lPCD9PD1eouNXC83wA3S3+XOBO01nFf3UWwun52Gb+cnwI7D3pQ8rWX9H6xFNdWlc5tLSn5
mwEGV6lQ5rjsoRbyDk6AhghMR3GIt3ReYqii08VjIFBIQTvcr7pEfiG6QXw2ht4W6Tc9JTYooz4u
MYz/d7lL4gPfuB+26I0rEWaJncsBP1R6RDZ/ijisUduL2x7JTS5Pijh4HyzO7icsHc75Fpqk4VZB
u2fgF92pcOkmX5P11XNs/wS1g5qkgeBG7OiLfgEoZyD/pTL+GKXJ/JR+3WgpS+3ioXr27n8w2QGG
Ps/ugoYDz1deuhqJ5vRMO+ZI/Kfa1Dm7ccr4wpNbN1RBBDCj+qabeUC5hoUzqo060p41XT7fOEy3
+UC+77OYLAAiIdW7bgMFF/ZowofEbgiS9VjdcCxR9ef7fK48G0LNI9igj37f2oleJIqJ2BJEwVXm
wV3Fgdjjxx8Hp8ZxnEK24dM7Ja7WS+Wxo9nlyxgJ6nlrOvhs36oBWNFIkmfUNC5fG+ixh4uwOZyH
CLh2hoLVUgAdBX5VSBj8Tb/uLC9wa6gst1W61ngrLxyWpdnjT+Bn5MByYk3m/bO7FFo9me1Sn5jj
LvCEEldleHn9nnkjD3umDCqflikIcrbkFV+q9mninzupOEn70pYRZXgHTJjeBriZUaSUT8/L95E6
yPEgZJoWfqJLYPchLEir8VSjSpbCQEClwaLVG1NIZdmWhhdOtsV8vsa2kAIJTCCZZQQGK/+jqetI
+zXWlZIztgIYTY39oGKhoULBONIyW/ks557Y3GK9RjeSZ/bGTz6fQs++GRebtuxbZ3kofknG35w9
2NTicGFoPzy2nRp/OgqZERPap6axAfchhET8IeVVlYtz+CLqPXVLe0/NhozzWFj6fJBgMb83lQdr
Ww35MiJKgIRoSZ2rV8oAJu5LAJW25Xt+oDx52yZKngeWovaqg2CcRjzQl/SIYM0J2GvViGCipgaJ
3ChDaZaQdCEvwBB6Yeps27KQyl2hnOMxc/XaGRRsy6951tNyXaeQpHA+jxblg/nQq+nv/pr6Bni+
GVGCF5MFMOATqwA6/Z7CmEXFoiujveRQ4i+2K7y+WvSKdlDOVqXf5qrY9Q+/17t3u7jgECtZhwq0
Q6KOGUcFZoVQ9zc6snKh94mKCDDQutXsIlVBCKSA1/v2FatOaFN4FnsWqQQG8D2KVyqAJ++wsZ4j
iSwT0hOE66KiAGqN19Kl6AXez1JkC3rjK9/RcvuAr54SGjpaAF4pcAwVO3OWd5AIA+FYL9eGHbbc
zGMDCXZPZA9ruFQBHDalPWRIPCF3XfkTtkp4XhEUJolX3Pcvt0oAtS6Jp5sPQ++6Td3PO7ermUJb
K+0EVsxTfMzzmKYGYu0dlo41hS4cQL6HW++XZqxLGoB6MM3wjOjFDzqbPtctUticoFCjvevXnZ82
43wDMTpkumAUwy8FcGjAaMlAulwyg4vzGuBvfuXR6jgzhYqpmXtkt97PXVxPJ1OkXimMcB5HF7Ad
DmhaoTv8Pub7PIaovp+yd4IAxfIFktDdElEi9M+eH+gwnelGPP0IzHbKy5B3z8PfrzWl1GHXGVfe
kFUrkjjfW8JNw/1yc+S0hr7Dh44nifX45e0mk6xWf3E3rVIu1QCuJx4hJFLrL+8zb+YOoflmGtnl
G3SHoSi3rj6bXE5HV/2rM5U3pQxIb52FhaMZIzrS9UPORqVp9FuxYe4SI1qvZk0hVF7Xs0QFRu4z
+sYsrowG+B24qnb7xHLUEsjITF2YEN06o037mQSJW7z3YnMH9ckOhM+wjq0ZpaMiK8fkNaGzcEOD
qHfL8XglMNQaHQpJJEGyu/AlEVMl2Y+qtKOhnStD7ZTTkXb553sCRNHREqN1SFm9uhoCRDJRSoFa
pFoPqB2bN4vndFErpD6LXaj6LTLgCsKWe7ZInj4pZc0Uwcr0DGk/h0fjsIRnYPFqKL80VEtoAVFI
pM5BQYd4XeEGd26PNW2DgeN7XJX9i7dCvhvybIDfPpaRGF3D5oMx2GuL/HOnWP+6wV3muKx3Y+Tm
pgbm9ZTkjnV3ZmlAcsB56zZ92kazI4vbDVE3MYcabsBOCWqit9vx+vM+VXFdAsgnrZWKStPwIdKZ
FFULI08Or5d9VRIM1rczOV5ypmwQSTesBJ1/iMsnCJ+KpmJHJAwivh3A3mZR28GOLJDzJW7aJKL1
5LC2p5hDmpw2QpKIeyFLOT4XRnhDXclCSx+KOM2vLJYg9bl2PXyAyg0XC/HKDSUF2Jto551N59G4
KSJPQd/n2JcXhkIBQNB8QEbrzmOqzycufVO5qG8D5F6/5nYPeZxUnXQ3exNjnzBIoAy92Izjj0aE
jcpfC2uDQj7QrBy1guo0TOdNzv25qSJJlwBmQZhN7UQHyYHH9Vu0EOqD3Qm5apZI2BJF244rriY6
qRQhjO1/Klk9RIthAYOJqLflcPBEejUYJV2R0mxsMjmBsmWzCdo0Q6VZbFAaswI0FwFPub6mfQlT
HBivlIs3U3LarhW4gGXcMC09khRaCkPsZvvUTQZX+2pywjblLfkjAFdSoI/JEA3/Jj0FYEc7mxuS
R4R+a4hOofyIm34oeT6GOu1jF80Iis87CqYQ/ZzvQ8Mj7FuI6d6c/WO/eJ+sRhLYSCc3ZR2HuREL
ngbEjncFRiyR0fqRzv8KkF1FV5sTQjF8vi8lCaEHiaT6XowuNLEP/jUhm9fyn4YAQzOPA6E61AqY
VXwcE8/1LLf312Q0w6lMX4RwqPjMlZRhh/aRnRiOiAWwsbj8pj6Fiukuqm8YfTIn5+MVxIkK4/Be
5eQzE6ZkRiIV69Pu/D9he2JzzpZ+18fDiN1OamFRw4Du3FOEodioQWIIcyEEZkv1NrmP0VDAm9Pg
D7ieFNRU4yJFpiUX/4HUT6JlKmO9yp/cjKBhzU1OWXrzzVgpldnlcSr63t/lqZ20MV2z0jc5zL3b
ihQSCvkkB4cVIfjUF2WmrDVvMesn0PB2hgOP4tN5t2L1RwgPcqey3U79Ijk+6J49hUL5O6EFrNGd
NnlFratFlps9ewW9u4ArrxZb3W2PZHICdm6fnb5AT+k0LoWbJUhB3FcGImCjo8lyAjMRU+G/J0vY
pV6ybb6oriezEwTXTMa/ynzkhBR0urVdYSzJX9QtsJfsR/EAc5ZcyBTHgmXvKZWOIvTMgNpEvRrR
YNttNQgMq+nX2zz0boWNigybzZ2mX0v9qzc+N3ZcZUzwJS895H2eyBtJKiMvYfbELNLBiLb9YSit
7+1JZTtQy13ukQkXmGRIWWozUEDrg7qG8P4swYu2SK11YvAyX8P9PXteDe0Yt4VbezheUEcm/rVP
lpkib9XoDIszRZsk0gjWP6XFdQOTKXIzKf3dlr/23lJL83T4o++yiDoPE5uEAMuZYNW0Fd0bvNrT
jWeSu99VQpFAPD+De711GuV2Gyzn5B1YJhD6O+93b+UQiThadgUZVHTZ4zDKCx11Vegr3RAICWxv
du7Cnzuqf5SmMyMmIf3+8pdJ+X/m8khacwgR7GVaUt8+LvmO66Nh93KzkEDbqekUKq1Uh25ziRH/
s1CiJh/YpKr9juY+H6ZHNgqIMY7HM9wpWF64auqJ/WfEITzORDnR038/YRxEYCisA/e+knsMKaZm
wFvYt4yrVinYI535Ejk9c13Bnhv+f31cXrC8zvYUhUArSl+aFD1k7BE3IQUMRif9zpH/0fRYq7OM
FvQ65PbLA0vlCU3LamTzEvi6yWezJpyjsqG9wIwQVLnsz034jGpojdVcuWQuBIc2x0TOnvgbQIR8
l3xRFBv3jV/eD20MWB9Usf0/VEn2ZwsQFDhlrW17KVRJ0oPuZ2W1KvwoFEDBb9JbpeBUfirMewpY
Pvlwj8J9ksRosIFgEPDsjg1mMwhlivE5l8AeoMsFykbqNVh3ZvDZt3mYKvX7jtBrKfh6Bf0z45wX
UWOPHgVZ2pqPjDd7c2Quz89qwnufcIoBL3oW6gIa1bzxdXl1lr8bKPX28KT+aInAmXxRqMu/V4eF
fdSuqiFrjNPKneW8uAHUQmPGb3CgF+NL9Pisu62x/TBSZAaLfYy4sxbYX4KjI1DfD1RDYLZm86uj
7JhqCi4nbLIRMMbSsERIKnq38+RQXIEZvSBIIOx58HZ0EJJz77DAQ1ZPwlZz0h62/ZUxklah5hKK
Jacj56NFHoau86Mk3Oz8kv5Wna9a4GmtS00FLbd4FOVwXaHvql0rvMOtSv6TFsxnLjCqXOHRHZ6t
KEnNBq4BW5WPvpGVggGjyHCTKhgfyS+hMskxs3LVATsCQa5AcSfMLsVXqCdQNAJGzvR854tR3jgH
S4lBmArT9CZEAMKAWBGfc1qKcH3snQU08hzf/gRTOEOg6EDupHR8Wo0qnMpEdb4EPwO1XCmrEM1m
PfBX7ubVwTsGdVmHgLW/BMlePX04tEc+63MUZ56fVOahu9pKNdsOhyCxWPSY59ZM4UycMPDlMvIN
asYdb7eFsDsD4RoVvW7+Aa9xDxHOu66YZoRVdnMGkFyAEe+wcpnmaxrwCYi0goomoBLZeP++ffMy
FN8vYP+OEZdr+CCd2EVdtw/6mkeN156XzC4sngFc5dIKz31IRiZtPVhBt+bSLAT6KRxhIbjUsQud
Ow5B8C3x13Dq42QtpBM2ii7Z88nafPa5F5Xl1lXRjT+xpLGB0S0sS+8ix1lTS0QCk05QtjHGtft8
PWafnQe5uFIgjfm17O9gIoxN1SB+KOia0Wid5J5wVzv8TvttUIzjXc1zUyU05zvTUbYeen+v94fJ
0m94bmEgtprQRoXy6zXCXVm0lEzkizdbHnTPo9Rj2ftlHCU7nqmReZkHScH0o2rvi5/muPLwVRxe
U71WNpln+P/lFPrO0nu1FOPkqGzQLAREsRX03k2HQPjCxjtVQoyQL2bw0uq89zwnfxrXavaErCdS
TrT4+d+3jQ5dhMveIB/tKZmvSBKydwdG2kBrtOSdbGDRBO+7BNPMPEqcqSxp6ebur5bEXfxFzqIG
r7qFrTM0hxqS0Z+jlVsGeFxA8gPWfHs+8ARrzv6nPrnd1A2UNJh2sUpJo0Ghr42nC3R+1S+KjJsh
FOH6WNXRODNx9xUCZow2LmhDqzc156Ou1IEEz69Jv4Nq3RmOfUD9xDYTha3fst0mDXsMe2cRS0X2
p3ETml5+0LubKhazV/5H5f72F/+mFUlOj4RQzfEMU7Yt+eYANSECEE2X2KNU2TcvmJkVTkc98Gid
vqYJs44xIDTcadd/zxyVzQDB2ZdwfF/cfxS/LVX8i7F+PCPhxBg7MBssSX3ah1jM6KxGh81bAa3K
F5UwDMKEW1q1d6xnKJzSkLCxB0nvjl/fN8Wi61J8JXBWlc4KAfNtUsK7SVRWqLBSyYk/NFMX55lb
0yrmR81iL0HiHMVGP8mThG6GMC16eWfn5soumQL16b51IHTWBio9Aiq+W6z2tuW6HCfMDs7JzHlg
1VnfvIDJEiISFIo/mbMSUBEPW/w7TYJ/u6y2RDQ1zjJHWRq6cP7hDtwOJnT7MFfOKSsJ9a1fuqng
dAg50BaPhwPdBaOoDE4qO6wJ9LC9qK/Xm+5g2b6VI1iHmeITv3wtcCnEyTGQG7rRzrgESC/u8nmi
iwH6K+rhBrIUKBW6aShp7It0ot5O6WC9v6pv9f4EcVgVd5kj4MYTedgm1mJF3FQgvR2Q6nFr2P/S
ZPE9cqB5rM/YGCl4DBHofwAJJAuDITTJdt87aotWH9vrAIhGz9I/yQpObf5tdBQxkvokfuwMh61x
NQSNePH8lwnctgRPgSxYB4iiw1HDNrz8Fu0TK3mBGcyWmzMIDiLFrbFfKsx+QNrM27bz3gHGCsfM
n1nCXBr0EnkqA1Z6GVo/e67tBOTbmSi2mA/9IO1sNNL1WeGNMsgWONfL8x6tO1PfWzlOzbrl5Zmz
8VuUd7ddowAoxrUYXAhaWJbbymKH16RjcEmiXWmA7lp7LykEQ4QiU76ZOuiJrhhOvhFLrAQF0eqe
spQSl0Pmos9HxToXANkrV8RIbExv+M0TYBJBFEruOmXFZoy7hro3neM6/OJ92TpCzR08kCmJMQNh
Cu2vPZxYcDrR7OQAwZINRiTZRti9mQkgGIuOUKSvlJIcJZ/hqcP7fOO+BqLF4hoQxfHz8zTbv9U9
ENKM4/S4q0fFaTdZJbIbMRZQ2ZLfM2Cg5BlvBZiNublF3UcoHHxrsWVEavB6/LD0X52Wiy+K+kXZ
Q/5fX1VAkkyeJrYVsLKq+hDRPlElmXcGZpdbF+15aZudr0qJgyijzRxqHe0XTldyQrbK8ON/ebz5
E7UwLiyUGVAd+p2Q+de+IhuqR/Xw5A79DpqFz+AOxWtMgfV/bM62XFdePxyGbyo0pe+9t5RN+TLe
lzrMN1dapzSSUFuTpOtB8sdJ4MfuaIzB+6iGbV8ciI2z1H8Ox0sGNqf8/fexmeI/uwsMJryp3Bhb
XJb2hfUx9IPWhs0Uq+B+MwmcGQC6XvDZZRyFQrM6yCDQYvbGKYyV7Hc5/cOWU/7kAIpmPxF9vUsj
N9tD4UGRXU0F/NWqcTU9Wo/FTDWzrKtnZAnUXR1kFlw+9f0SiPUwmQlz/a5e2CurwNF96e0XQbGf
iooRNmMuOGeqnQ8vvo5zdcDjwN8qfDbEPARUPYsB1s2JidiIcbtlARCM9xR0uOB5VLbWiEMUZ0UO
zEeEtgTxXxGAbRto7p2NBY5AmvkvhTH8oAX9UoNKFyCXzgZmnhNPPg8a9bMUSnbm+7rx4dSiSCCi
1JWtJntopKpIlRioarzUMb9p463JV4Xl8UtWd9c9MQFs8MZGYc27jQZXYektZtvBog5gjkZFiUOm
G5E5RKnIZ9lQv+bdfWTT+SiBSMnT20voXBryBu/RF5wHxmto6BPg/Wnxpy0Q4LjIJiJyc4JhBpwE
+CAnj8JM3b3SswCVext+Onk/d69HruwEsmlOMrAmlEa6Xxmpm6liOuVnuugj9miwgH4oVxykCTOc
Udru/ao91MeiFECWSXopr8Ixi+7J8vnw36zbqu1fniFRwdOfXpTP7EJ5AqtebGIK/m/nq3LCteQb
69aYkA+ov2jFIxZFqvITYrBG5CBroh4zlf/aX+HsxJn/5J4vOiMt0HRjpRRGbpAuC7HcJA70/jPy
AzEp6i2TjEF2mzSPMpxzkMlL6q9KbgzwDhhtjFZt8bqtAPQqK1m+1kXP/aPZ77PlPlLjUofedP7z
bBzIGislVsP62pEKSdI45ckpVRM9hrwYrZOwNK204TwgVvm0YsJF48hXBzbULHuGb9+9zuqKxdfv
YFdo08MmAAvTwTCSQUme1LIeWQiQ6XsvHkkyvPwv0PFRZHjLf+kVwN14V3HUNAz6lhq/93ncxBPq
NMtakdWmJyca6sNZJzbdA79nm7qJkYslOPRKOIhHN0xFvOpDZMdPxXqhvt6RTko/L8scaBZnnhty
4AgQXyQiJIML4JqAJS8XeiYnfMfWs0gMfpzREj5I933j920/RQpEMY0szVZ3Jfafj0tCtONgd4zz
/qB2yP4vXZg4rxsul14tr57qgLC0ap2Ik0dzdPCcPKPXcoeQiDiAV7BaQZCJEfOt8MTGrtFFGKUR
B4OM7rKfsDbM3Skg71TbWo4aVHJe3tSPoa+q69PEgiidx7KG3FgmXHFtvVqSX09ClFmP9BOxidzv
ZdYf8Elf/kXT+cCx8Iqj1A/55lb7ovJktNiMf7FJxh4ENvsTuzx4flH+hpaE07yt12wAThsbHCrr
GNAh88GtFzLtMTcmNTSOIU22MK3B/sDPCtcymuyumdua3BH7LRHMVO7y7ihV00o4AxtMgIjoM7W1
8CDRSBzsMK288R8BG0/w8xRLciUg0DZoxKB5hj9t0qJQ+GhxTKEVW3MGGOlWkYqHH8UKph5Iwqrv
S4p3P0vLPRbUschcjJ4vOx5ghnuMWMgCWMD4OAxy0aNogt83JoDEyLug3x+8S1qkdRva1M40l6pA
uS4XwZat2YajSVhIuroZkUUWIrfq8rV11pbKC41ax2rvgkWKs5ETKxwYMvmnvl1VKllT8TYnkSSZ
8E0SOjj+qX4x+rcRBiFd3hGPUcVORfXaZofkXd4CjoJFNOgtOuDtx9vBwf617FWUPjHCsga37zHY
oLP5cgF2+MrAxO4Fcw2bVvB5B4dW98Kv+4sANWrpzH/Xbql+uas926kwqyb0JPeDyzvXorharft7
sH1AQW4PajNNlbhgWYwK1XupX9ikLFLlXsh4M51bvqZGHuiIRT6Fp24pou6+8uGpdqtMbo/CWsAh
ubzDSbZJQ1EskqtM3rwjQRifKZpHsvx6AukFv+EIohjOBun8A9Q0RIHgVhfZ5vxmeqk2fijosacr
RiRNqiZMQAZNPxSLRQLU2nqiNDenopjkXUoFqr3VTJ6zejZAh/zDjcyupntuqLrSQrOp7i45CDPO
slQ/VBVn1OAdk7dXX/Oe/Le9Nf1JNZmmoIH8+2A3RPpkvKxRpN+jgzaktdMD/X6CzoOjvt3Y0K9Y
3fh2jt/u4yaCXjWr8LrWTx376gsCNJbimtSfqOiAoGoic49l5/L1PJuYycFPjr4mu7h8g8QLOTXY
lNwUSJAiW+lF1W362jypCl/2NhRN45jcc0I+vUsZZ7L99GFPefYal1HQII8bdBKLFOLibK8g3FYI
h1oMMwnKSguoPtYy+rq/ZVx1YKNoiM3U8iP9eNZltE8tRZceyZBqX9mTKZWBzEcG/8icnvduXbpk
EtmsOhNYouGDNEL7K1xdblecVUc/VW2krt3mOSgL0iDfMr7yox/S12W6NN1fCQihkBqyyWgjJcLU
vFbIxPhUV/1abor6ZlDLTX7YYZ79Ivo6EsRy8uamo4/bqtsHq2+uJ2eTSk9xdCI0mB17BahrZTbm
jaLJeuJ84uzQpaxoaUsmyK7AJOt0qPwJi418fq9R5ALh48AQRiDVHdj3BZBsZZI9dPs3PNv0AE+N
ZYXsgKUX6ga/fKFAqA1gdc70Kvjy271ZOvps9VBsTO9/+ywS8YwTQHJBtLCFjUyb/4FiCKmKacEL
kaxehaQIi65qWjKbHYXRiAq49lyAaIvdh9S3UPlq9B+aFdtYnDa7pNlSnzBvTOgTdIUwmlXErp+/
CmKuocuDdripd7q6j7OhKwwfniMq2UBbhUD7W0ipqTe/GTMT1v7ZyUdjDjqYalW3Ut5b1NDKwO3+
qNpNtHovu2zn+I9CV73DC6d/+0ChzCvqOb56RM8GwDvfXzuGOCTFgXQSnb97QVpgrfiYK0GMpmEf
yKCFE7kLcPXConZYGSNOUOnsv5XieAkRoZtUwsv0eiw9QV80CQjnwUwO5Va54dQ6F7WAndh0jto8
0wf+U0oKy5Cln9nLwovpw1IAEW9HQKBCb9ZV4tx/tS0yOsFrFszBFVIUxwqJJvWe00fOMj6UBLBn
1jvzCeTLWBd66c8JxQM70kxkFLlZXF6LKUjGtpZApuSj6PYLiQ40V6Tg7xgYbd99W72smbfoVG5n
FokCdD2pZZHNskLsf12E+z/K2bTqNCr/xZ/Jmop5J5sIVo+kP4AMQL+0MjCmkY0+dznm19g32Tom
Zc5Dx1bMeYX2HNV7zwKncXQ/BbDcB4hDl2I29DW8bHenZE/CVrZHzPB4P6Feh2hc2xO9Xql/Eb9Q
J1DJ+Jc2Ocrc1gcZjLL53WpTMyczSZtw7eWUggRAa8wyv2ZB20nFJy+0O8IYQqo7Nl8F/iWUQ/jh
fLdUGC1wf9lpXmRDht/V1YhgbMFfjYDglXzZyarJUF/6iFOuWxZGajKQUmjXDiyKjVR1JgKShLSJ
m+/WdVd3fNuwbMFl82ZP9I2dLp2kmjpZo/KXIsp6nfBnzXOZ8EmNXRKKchigb5rBt0o+3XLvf1jD
/qYeaX0Ppf9Hg7uPMQ7XRwVmwg/anOZbXYgYHNBmVYU2njPD0X2xXOH9S1Woh9BFjxPh/a4YzeNl
MWnsP0sSMxNikmzrdcaUHJApp9lPQMMo/XE2C7Mt3QGg9pE01ncJB5D1RP5zRA3CJqj/lgY7isEE
oPpNyLUh7XWekt6EUzzDOVBQAXDmEPNb/FTV4leEYKe3YMjdqU2n+5zaM4ei7Lqpc3wmft0CaIDV
cBMDBGRaSuJ3jWtdTyPiYeVhf77gdXPT5lUlvGQDhqtpLjDifACxcnhNDi2x5iY4L5Fp3Dme3C8/
FzLvlgHbO5qaOvSV8gw8bA3l/7MUvZwVujM4XUEpn8ft63FU2Q4FJYKP3ch8ReUG0lSDLPFB1FSG
L3gO2F4RhV6vA2iN60MzDbhvuXA9Y/rQ50MYtkk5HrKbL3uh7w0SJ145ag+8lHKdEUgLgMzyMc/x
RXivkkLHMWIqgAtDvzoktVl1MQvLzKGuK2bvkO1oH+l5U8y3RcSwVFyrcfjVK9UAfw4ukQliQUuR
Bwi/Vqylyv0GkPB80p1nW6IvQ42Imf4As5d7kej/5bia555KZcmYtMkX4njYTCK5t7J0k2EraVaK
ytcHwnSTBzER8EadMNiFAl6kOOGGnja/1sD4OlH6E9C0cbehlpUbOKVJknlgD2Pxj3du/wAA8hEU
EPa3QWe6EXWl0v06Q3xbXhEVx36t/M9UvTa6na9a9yrQGEQbYV0Qt15NSr3iSIp5OogfAWsSC1jo
q64Je7Az24iEpgmC511dw6Z7tCdQiW1TU3+LuPOzhQI5VqA4+OkzpLfincndP0Kbw8MLT/68Ruv/
CeCC7VjRebVW/FwDMPhTWSQfnH5UBnlrWBP2SH+Hmhbx1vY1aVT76kv7+s0nIhd+FoWnOkhPgRV8
cMGWuauuD8IMNynsXvXzsAHEtSF7Kqa9ECdDVXyS4OCoHk8iHQfbB4/Y7hGp09n3fFFOgpZHBODK
6BFnCz2cwIdJZnuUAFMuycQmc0xPWKwG7U2AMkpraQM0Eg6irkV4Xx0jCnXH8lEp7RdsxW9AXcv7
zgE9ltKMh5RBPjLloPL1dggh80Rp/MbbVJTChwpsF8gceUmgXd5JDm3Ieh/7zPqsUyTHbMGbja7G
KezCLg2yuoHyTo1xS9+r/CfX3clZS4e8r8De39cEPZmEggPQkq3VIRqQyXOspO4dkF9jMZ11n09m
Ddg5whzkYf7zgsZqaE0nADEMcaKhD58fsr8Sl4oTbU+nNBWBqvS3Dbf9I8giEYgXxuK30MdhDRI3
PjLpc8ewGfCJwnbVg+5ksI5rrzPKO/pR8lsbGdXIDYLyxzY9XSo7tb1pe3wHsGJoK/KimYX/dzq3
w4X3z7s839Q5OuqdGy4ixAcmy2aZEzbrGUQwnJ0nPwvyjUsq96PpSB+Q2gYymH/ye/OCgd4UqsMT
7ULUk2uPi5OOLfwfLL6gHfZN46Co/SvZ8wpzBQr9ZZf3ZwO6GA90yf8Sc635hufYqrXAeCawwPBy
y4v3Qq8GEOuIuXF4gx7ZKQ00lT5hVsJnUyUEhMtSMsnQTrXdupd4qRiR/+luNKLrMl4UUjjNqB39
kkmFwIOCTRITBtf0q+9EQ4cyxV9ujt1hxRZeuHdMdTuZDhRUibf0i739LoKRYp5d9JQdR8is7JKs
w0mLMknwxkIBSVLFm/u9rpWCzUlFFN39VEp86KxNzk9v0KAN6TJxt24fwCL77RWxp70cH8V7I9fP
vxdrXlwBJH1K5jLvV28scNnYrmcF2nU0UEDMfRN0YFxeKSQgkTUHLzZxfooBRrfhJM3MN1K4ry7q
B4nrPyrIvAWGL1vnGFBfPXxT38Qb5T9Ijs1wfr8cK/F5xD8ymDL4dS/39GLB8UrAXV3aqLMeOQ67
Vy3aH5kdcESFqlAw1u+jDaJKlg1WoYOROjpiXqXra2HVK7euuI9BGUhzn2O8CerpBkjIuXJOcszF
jooApBOdjN47k6PFNGU+7xhjzJn6b0zefCisjZPlVSQLuiAdV2Wtc5M/15UJJ2l+NaFIT1CjHxPv
l7m7xfLKwCWWB2OhKcAY0t8bZtIv+7aZF+/yIVYdR0830hHRR0EBOxkvD5XfIVtzXEQi8LxlR97a
WLMxyT6FFiEl8X56BFNWEwmjdvpYmrusP10edxjlsJEV9TbzfMHKaQUC65v9YYd4qu32eeVW8H6A
T8u9KIl8enfyavQp1K6rGZR5FjHYExjdm5JuwLZREG6e8YTynX5FOBwVddLpcw74LVmXnJOYW3a/
teiHdhjKDO9hVqSjCHhR50SZhu3bGkex2PsJdgnbg38Z+C3xCaruNBVj/IwFWldL4ju5OEnDz97j
3zOw+6KNDR4uLM7D9lop2bplqe68hYhUnsGNxX4WseBP9XWIrxeaWQb4iHoisaXwDL6L9ZMltXIt
6ZtVRaAr0H+ivgfnITI4RLng6cDuBmLVclQ3uLvcQ3FrdQGEzIEPV6V+PpDhCmAncNcA1EhjJwqJ
6dgBwtwBiLUeg6EILz8dYwUJyU3mgd7hTA2ooPEqY7F38GYEzRU3tZn0YlQUpPf19k8gu4hHP8K3
lWIPsbmZpkFTreXQmyF0ydN7JWGJXABW6jnEcciNIYBXFVkqob29Lv9RFsdZPDJDHDrFGRS442Kc
Me3qO9YELeCA/3KQtC3+Wf1dw8UHlqszzhAfNbofjteT0Zx716unHiejzGO8IZUQF77w/UyhMtHd
C3lap5+21nr3Uv3CFJDvFarIagYWKa4gUc0zYTwkXnC1YLeFjxDIT7CFIcUKygd8ana89kZfVDn9
i035L7x8//LHTlvpUXWzzzRiT2S3t+gfwe1p6nkznDvZHQ9s0KxhX4PFUrC8rm1jAJeLn6wft2sV
gFXJyMVLJl/F8HUenlBSm+5eNp6/3jalq66YPZiBkO0LOBKl9SCoYCfkW2WZ6qlhLCH9TddW5GLU
nGHyFT4jweZDdEvqleVzEaYvdUFA9dfcbjLtf2mrzrTA1CYIXvM5r2Q5hLK4KzZ/UEFi5IqhnwSe
4AE/qInU6SHYH0DDZ+QPnCac8gCJmWAW+cLLagL3Hw/f6gP2UIGGTWfYIsqiKt9S0MLd3gz7oXQ2
PpVAKNF7Qv3YBdoyr51s4CVmgCrrgD1BCOiqNuGpgDRujWon8ssq/Ajm3vTPDyWIOgNG+hzaDLh4
RzJKyAn1Uc75473sBAXLDdLedsNm2k8wFhcAwlef2Pcd3xxsGu9uIn4mq5uNGD9e+S4OKYtmoGZG
19SKrDZ2QpP+fvoHHSBcrI0r9WvkLkmvX+JHOx7njVOqXxwbxZ8ko8Ri89AhKI3vowI3eQWXOBHN
zyKhZuSgde/gvxMJH6+8qrhhNaVfVEFAFhHShcBhFuuNT5Xg/K1ayNgYzWdbW5K1qEZDVkHkVrQ9
/iY2gnJUn7eMKDPQWbsAKshvD4+6D3J6ux/Kjwp2u86LWaKXiqm1drlpo7WAiDJdGXhRNy1GLAAE
IjoRh04WMYF+3it/aG2ATfxYrvKhrGq9YqB3hh2+u6Iid5nUql8v0Q1pKib1vbEpCJ+1npAveQm1
rtZU7RyJNHgvXe97nbTJBpKbeWIsgdhnfmY16MLASJ4blLV6aer+nzqIPBHlsGdQG93SDFplVWdu
TNXYJGHXvOwoiYjIR7vSABetAdWAQGZINpa5FDYDE5ZV8rS50hwi0TDRcthFoVnpXPCBradMJeXg
WNiQI/XYMZjotjJxQm0uXoyUUmbc/CIof5zsw1/J8rj5wKz0xYnshcKb0uXQ2Za4peJWoD6CkDH6
oMZn9D7hV81lzE+1Q3nX0FBAAD5HOe3WObrPj2HFPMc/hkGFwVwwFfwqHD6nWNUHZQwOGWFhef+r
ha6n66p6VA5k/sQS8/JOhmmVGqIBrptTpo+nSOHNb/0ZBvxB4ZWkpanutYkKarU1U1VIN9+nUXpM
n9p9+3YoUaXFytW3m55+yaHb7gHCRmFG2rfE8myaTmSxKgkw8iJN3sdDucBF93JtCS9ULOftxu3G
n7QDD7kIVxGyAyMJotLfeU0im7xOugyqIXZj0t0wzIiuhPL+iibNO9y5WRmR31NZK8qgl1/Ki/VN
sB9Sj/nmGPaB6HCDlxZjsmbWU9RKjOPTnBbZxLOla4AwWp3zMYoBMCqWeZSnAdg/9P1hSpNzw1MM
fanBAsOuIou/EWyzS/SN7aw0T5rGULUnWz+qxNAwoNu9zfbQMxQKxb2eYnkbJI2xoG++T7iwbhuE
FGtDUJ/7Q1ghX2PbYkalG37diEdd1dun2r8Bih2VJQ2czJF+0sPuFwU90n2Nty+0Fzwlb3eatZJO
4TP7v1lZcwXjdhQ8fY7Vc3ltna0o5y+u34RC9N++iKcO18S2RuRRbcEGcjnvY87krkhKlTay1XAv
frax1xN4Vvsfxc/m82mmbFyJkUEjk7bsLBOa6nQ4r4iPmSgPfiC+mzDuc9TQch5IgkC02nyBnDVk
SV5d23uUYdcwo+UbbQ0YocMC1AcWxs6D5jEok1iEfHpicRVHelCSoIk1X2Gs0cBWOk+oWgPgtGPk
YSPmMdh3U+xOFC9lI2zohzHxSbga3F5SUiEfc6SOax4jPwePHX/ddylOcXLB9iELaZQV/Aef6EEi
T6wHQLe7GZoVCxRrWINlQZFQafKZA4wIKWsZxJpkK4h1rLr9rGHUFlQDZXe3h3IN0dTx1bi+fAHJ
ve9WiLLLA8pddXaJ60nc+0Qlx0Utx4OQVGAXsYAMz9+OsXmaK1oT/MVO/+s6tmrfz/CJOr1LbA5V
huTBZ04/FMm9E+X51GtNqStAxx9a9aujuECO7rcA7rFVKCX5+LtD/7Muui+LXx7EOTBnn7mQClE0
3vnGekc3Ene8y8mduTvTL7reEBDKn2NoRarjKjRxmJ/NBgg0f6TAZi+G1qy1ZGTpTlNVJU4yqkY3
++q/wmZI1COVF20uYzuK/3kig/WMdHVnbxLpuos1gpTuL4FhhHUZNN4KzgD57Nx8F65o9LeDLIiw
+WqbGNM3ww2YGyUpRPHuwziiJ8aeGyc9UYQ1OD2f19WmXlUdpwVT6kU3BuylPnr/zesJJcwyZ4Ud
pH7OevpqePPJ9GrhrPY1xv4D7CcdDCaQO9WT49VmV22o/VLAzkYjLiHdlbzNq/vX7BrWh9agAsx4
7BY2PTZS0iMX0ySWoht2n8FbBWEtIK/53h68lQSQ+kVPgQ+aWxpqAxGtGJ1/DsYH6AwvVG2mcooc
pftyeL0np2vUNBkpMV2mLW8c0xBk42KJwaJmRPkQqufaybnl4DqAzZtYPkURdHu5t7hKuQeKuPTp
m05vf+wuSbSFhBk2dC1otMig2zFO923R7o6+UW1NYSnkLIWhsatThqQZ68Gn7lxk1XbClslQb4sm
bSHahlcfcct9aY6JBEo93In5eZWy9zz72018O3bfX6cJriGszRryLV0qfgXmedCbvnm1IQU3JxcP
oq9Wxz9s+xmF8nfbdoKbUYeRVKRb85bNftLS3SR/4fGitxotd5jPlzzBpxwZ3ckhBGiBYQA/0Odv
BkPrcxNkFGOUBRxTCAsK+55+6G+/IPsf+PGHjgBLCV3J8cuI3mLgBmnOSjl4+Lt5x1LH+Sd8Gswh
ErCtKHH1tBgndKtKSl754mKWEBoUy1VTAY9SL4uq+a8d/5yIibIB3NRYkbKNlYqte1Frrr72oXPR
YmDdyOnBSTl5ES112bxNOkfJnXexGhe0SDt8ZymLnOgt1zl0R06iXqkkNzTREL+O6J2K5WAkjdi6
f8eQk1VX13tlmnGSoWC8iLBJbueh8TtJ5oUStfO1rSkfPu3Zn7U+Nm0Qc6fPuhBmn4K1ZAUtAIei
EGPLWazCRSD5PhQwymWxZ/RfruXzAguGEO5PEpxKOeAhvv/x7+tICabj/Fq0Wzmh0W38T/QA1sOs
5BXroukxMsf2C4iZQ219hnq4AH8Mq75bgIT56Q9RKHtipI11wfc2IwFyMkB6A8wZ2ChuUadaYMto
tESIKUXC3fki53SFfXEvvsPV2013jWuvr6gW/iJ7jIU0yJpGlzy1Ua30pqR7Ev89/HP73d+/s837
zANyPVEcS1yFvppNNX4nRKQLv0ULw0yypv6u2a4yEx7JKovn2YG6Vs8G/wC9G4Sk4GC4T7MSym+x
KGIESoo4q1lDEsRb/3BZ41yqwioniJsLLGUv7RCg/f3VMSz4lIIJ72S8qmcqRFsmW3nC0xQoVpSQ
tRBGjhLuBsEJsBj+jRlfROP2GyeyoQiGCG7c3k8au4SshAp/Hfxz6ZFKCxj4laJkd69d6wgjbAWr
085iCkP4PHlNgD3kk9LnAzXmYecEQ9PRphmifMJr+xVDAhbzItGj3C8nik6QzEjN76vAqLXGS+05
nFmNq4q9PB5EvCDzoM5bSiOnCYk7/RfK2AaWhgbVgWQH6JGVQxrhYcVqfZ0eeMJwIJr6dEk4KrPY
XelQL74w7SrGUxfySYaIEuAPVhZss3ZDlJ1reuFFGLpKvT2qaCNzXWYM0mhkJdau4eMkbXrRjdUP
Cy13YC2NnjZAJ4FSpICImKLn/bdhesQOaZoKUisahWdXfzJPq2+20kGZSnonTzijrX9zoKK00kQa
Wv7wgLzqQk2BeHukZNtkIOhq1bZJMQGNXKUXz2G2Vm1CJcSuDjoKwOk0b1uJ426b0G6IrRfNC97X
tG3Aa/XvC+tzZkjjsx2bfShesQb3lFo01Y5qjEH6uw32T8lsqzgf6p2Ji/eDvYmpBjURIm1Q8IXT
D/wIUaDGDmUtads7lD5I4jMJxKZGsBUl5qhBnU17muCwahQ+j/ZuQvD7ZbCjpcGw20smHuGQXM15
38YxmLQgdchQTZ2e05ZZ1ctV61hgQmMrEgzdhLrntQT2f1O8i8E7aQrKNY5RguIby/n/4W8dtsxy
rsOHYcWKviOPAr0xXCUWwsY0LdneKHKD8lHfPzgC4ZWRPNf4GO07OCEaOWUTImNmL3eLgabUlzIw
ig4ogZVU4KRdQVNMVKi+T/AOaQx04wBH79AmSAm1w6E/EzfViWOT6ZFTQdsYkOi7/9DaJsX7zSGY
Zt/7YxONdoQOzaC//hFRLyM1X+oKlQoZno393WpmUYJ0yZc0mYK9NRxq9ua+bMt5kMCDxk7wgCPc
sze3yNnZodz2K1aTReu6obQ1a6Uvnsjkh/YZHmMh2rqMPwptdnHsu0pkcpjJKulV7udTro/c5w/z
EDl+yC8jJDuISBteDYFNADSR1v9siLH59WU1JLK5Wf5Qb+JzjOoCdoF9byYggjPe01QABoC57nqt
nS++JaXdFuTqkxypJ18bCzVg3aORrukUHKQ3CYntsSz26uqPP6r5S6bihJw9asO0NzAggYVaPoBQ
7vFI02aQsaInjiI6Lp29NnZS4FWcm5hWo5TME3r/ifyLPgRV0uzi/t2YILIGc5gcBdPb1fKGAVh+
zbWKiLnQfTH70eCsWzm8mvjsqI40Vj9y1a1hhPa61ssLHaABX2a/eg3GoZmKWKCV9F7tpHZvI0yG
Dw9A2fW7ByJPWk1XYigYx2qlwG/hJ92j/7DVO08OjWHXZTwHhu1Sx9Lm0eAZj92CTGN1YTzlc97B
ZkcCu/6rdATqOZLTyo10zvlLKMXOmYdzr0B2rpPSHx/r61VCeV1dbat8KzSlQ2GdZwIGU6skqK27
YO3AAfsZ9QsHbQkBcA1zKOy8Kygnk8wi130fILRfnZJULDvaye6lXdSotJ1NCE2/Ds4RYP/7X+WI
pwVyqjv4PbTsIjPjN/IEDhDNYzh7mAIVQldZAkpu6zzm0NxxmtwZ7WHibpILPFFjBfLo4MTe7j37
TTmgACN3QtKFh4oLnHbqqJMRHRu2WYNwyZDCaQDW9Dmc49uOpZqGqONBBQ6v/nX6Enbim3aW6b6t
/NNkW+i7cKqqauWEYLWJwpsrcOf3scOYAyyc6fW1mVifEpHbrjRU3dnrxGcL1s2lWrGkHPhKklv2
mtEK5Ry4aMrHYzcLDxy8N+6sw5kkgRdZDlcipRJFWm2EPYFkkB/1jfzdAbuDHWLf2yrC3NH3d/5S
xCr0Uj7N02i/6BaAlzzrdCHeAgRDxE1SBcYZhgI0+bKlmnKcCANVPuGP2oo3Yf+9dRfMejYYbZoI
UlX7Nyl4WFoYCBu33hbN7ULX2VAvOdmq05ai9kxVNFb7qFlmhyfWrUGsv23A2/IX4OHEUi/9dTod
Snwu5LOoUsm3azfVOUOhkW33uWOL+Kb4CV7c1gmN5BFHfv/56uzdT64sakT6oV5dRDkcOLz3XwGv
z4/NBTevVKdY0MIgev2Atd4bSIUH/ueC+bM8vakT6CBDVi6wSNtPi/VyYfbjFkL+G7uBTWGVdYUj
mqUAzRNIUM3zHupOzmfRmPOVbl2doWadMWXIgRMmIRU+3U9C3b+lCFomciJLlvG9IfUoAFUSA3kz
e6wYgnMfWAtfHLp003v0B7RLqcExHsIFsxsTvrd8NiH2trc1wsasQ5bVoxq+tdNoIig1J+v0nNcF
2CxwDcgubFcZzFcDNE+vs+ZPlnkjfvQzfkFJM/ahzXWXp7AkDxqQyt5BBJFJWqEalEizDngvO2dY
zmG9UyMUWjhuCBtwr+aqo/mLiWda1I+ldMDxbSU+0IZRzVLxckJ3yOFZsiOeNkFGez1dHB7thKV4
LeqcLuQKz4SBXTttp/t2BmxfowCsWmqpIyP/DbVUPab/Mr67CI8SSk22dRr2uwfyHTeEUaRs8NwO
Ft+ePCwBuglcADVvs49cqAAwfrh7MdcPTfHk2GUji7GRw3nhWnZcRZmDlDOGN6znqyP/MW2M6Ac8
QIVlDeXGBx15Flw5mL/5J+1g9ZqvEpAlupzGLT/zEFGM1yIOnkDZ0fVL+9R4Ez74jfFVT6ieqjyH
nTk/vrYxRaSlNvQryGuM2d/gWYUF6A1CPDoVJO664S+5O/bC2M4sC7GhEpwIPonukjGS2OaTVZVc
nxoil+SzR0xixTbuC7p7XYZE83Yx+ZG3/Xzu/COOhdPP+PM/aVvcOZ7RNc+UDCwepmSeIdlMDLkg
sSHj+wM5k2Iyjcavv0VV5292J3/P3Oo8YDTZEf05M9L3pQp+eewD2250QVTgwCYQSw2BfYj5xFkt
JtGd0RcvP0t/tx+PG5aEG4GIwfU7/P8lKYtyhSgu/LYOCK/mjqL+//g7c59/zw8PRuA+9lk8/Zfq
hBCDTo3S8TRbik/8Xpq/qlmqBZEs5wK83w2svo2P0343EJZNeEY1LqTYUaM9BzlpZpk25wQf+RRf
SdRiS+trMJx70laMmgy1TlufXy3cXBmJdgTc+Th1VC4eOrUsEw4rTumEt16A8sKmOC4RKfOfh/Kp
i/z4FFR9Wj9vhGRVSPkxNCiOzZePLhOzy+V6wFy5gL1ONqUlpzvs3PT5AqYAChTqU4sxK4mksL1P
XvuBSzW6QGtxaYtxYJpldHJhcDPjYOWwnPTe1up40wp9cpRS6G4YkVApUcswRzOL74YKgL6y1lE2
bEihA0awnFpGYJrB9EG58sNHcpRLPI5XeHwfT5Iu0hv230AKlMVqTEfKmJAnIjBItCZ9oT5Xi7Le
bzOQhxktsAzKvNyirFfjA4dcY/S5diXzslirouyuDfKusSKuIivIkn86nmObDBDf166c7gmFeVG2
+FjRWGjPalQZgFNcPUfUUfJkQ6gSw91hPGTMmgMS+r5E0afRjwDlYJjcjbJFqhZrOZ1b8nd8xkG5
yBDMi9S0tjZ9rFXa7t9xY6nlvl8rqgAY0HfWxcAem6krUKTaOyuusaiMigC0x0A4soBie6dC72cJ
+GkNf1YxjzzwXa6pH5hmMO8KA/R8H01GNvsDOKNRygWIMUIUhFrhZ8PCW7j3RWOPowP/+O/BZsKx
aPjoEn2QgISfyi32OkHXnROOsH2DVL2Bm+vpX6//ZWAV5x/VQAweHwkkLd3WxrYT/XmZVl3bdYaT
XN4OKO/67odgLWhItc+ldmMPJvrN7CLb/uwEXVlvK/3r4pdb+DPiyqKohWU3BgRKhAsgjfwm284f
uNVCSyAHGz1MEXX6YFm9q0PJczuON8DFCwsWL5X30+ZqkT+H7Kh8CjqMwi7nh4dLQmtsttbo6Ot+
lFUF1YcqwCFy/Hz+GOT2b6wyw68Aw4aUnUcdUj6lwKrwKJ5140iPwmE9QyFyX47/ogyQQR/PSlmb
1QYaNDtoL+fD1jrPuCh8uSmeszOW+7DWr7n/U6c3JJZsbQat5RphxNf0w5V1HZr0SWgLRyK+yRP6
7As2UilNS8NiGk3OT9UC+hvVibEb5S1u1cdggaiN98G+W7KK0Cp/4y6kAw3675cHSkikVtGrTgi+
lWn9CbEFl00ITcXQkWKl8TUcllXfrfsmrbLHwiUiEY8jDPdkGW1/5oa6UT8rFnc/k/N+mDIbUckz
lMbaez2lKZpVt/NNNQFbpmLcp2sY3vtZT8zu601NVIHzekTOci5SkBxKWf4X/5Bmar9GAIxLHp1A
2vA9aVgmElbizEMM1uVw2lOrfQ2KWXUCht7jmaPtd8eCs4B8fMVVojzlPdpb8u2JkTlUQGeheEtP
8m+tapkdsVHH5Wd0TavTBqd0S7iwjoN6RQrNON6sssveSSEBhJkDWpwV7fMDzs3T0A/NnSU3/UYj
S6uvVMgkrx6sfphhWgHwt8C6+CvDPbDnmAPvqlkNwTlV7HesQ+Qcw87/C4LG0ao7Cm+I2xFI5+TA
hkRRdNr6bQ0ye6byn99zTR6c1J8bUwbHsrg5g3BNmgAKuPBNYpTQMZRKvdz8Y9AmyjjcZjUTquON
Q9A9Zyrwtetr0pVZiMujRpoXLw+5lV6Zh3lvik3iZrPpsIvMzzHK8AULrC4nxrGAYQSX31nORWlS
0j3yQ5q2iBOIIpsndH4BECJuDSrueiReN/2ZoldHasa6IfE16th8Va7RZawo67yoeAlJVoa5PavA
C3XBuX41VXd8fchIOBwd5iJ/TlQZM5ZjhJIIjC/XNNEWlFNRcIP0yj1/3r8zpM466bARIFB6r0vV
lGAbJOyu4BdAHfUMk2SCIAJIkqA680Y3D6tHXNVN9AcoDU2Wekx+OJOch5Lo7w385KNJ8jxMhrVa
RDKZC6EAQ7nrFI8BneshCtv9ZfuA/trxzvFJ3CP44ME8B1iVBY55LnPX9N93qg80PRDq+F4JbTZF
X0Me4WXpOkS2+i6cIawcq/Dg00qdjBxQdiQrzpc7qbdSudGj58yQBw5G+YlfojzoI8X4sGQskpoN
61sXT696Zxz/aDEY6TSQkCTJX4Ylo9Pv69vmBREey7w3RZ/1IZIfYyJaonqcKy+c/gr2UJspdafB
kPyH9DLiSjjQoHk+PBpffw3x/Ll1bKRXqL4xYaki7G03D4mqB79TvSPVlcnlhs00qN0oSAL6iVlE
tEsLksjRmpDzDadPXVhKCdwftJZ79h47Z3WDRT4wRKxC/HoAmStkAOdg7lukqPhq7bPHIzF/afkf
na1peb1zpGx4nVphKN7ud6fqWIzLJRAzxUJKiBOQX1l1MTnwtbhiwIIrtckEYA9R4RwcbL5dtt2w
8iCj4Iah1p0NExObA4oHAVIoddkVmXJRJ53evPaB595YzKFqk4EB2RyW0Z1NUjlkMx8xk7f5eaC2
fPSw0mcCmEsx7Ktt7YkU7C7KVOjzNswe/RONY0XAsWJrAZe44iXZZ66vlNhFwAqwVUh/wKh5XZa3
8+hln/V4tW+ySIU/MOORchY1pPg2cVNvSicj3oWUgEEjtUrCdn9d8G7eogJ3GMkm8nyLZJocT6n9
+0eEmKotR06q+CNQNKLFGxmweLKReBRu6lT6cTxS0d4uS+yTmyNxAmHsJUScqXQ/4fAVu1H60KUy
bvPx4E8bgdKE51WVInNORYbvQ+/LCHoZ+FgtvdS6Y88i56DaLE/XMN8nDlrOacZPVcHhn0ManXBW
K6Dn5JYgTVWmZcnATIxU5l+0ExCDYndJCrjthS01PaGw6dO0UPo/XLl3sacvS8GCN2C9YyzmJWj7
iVhYP/VjqGiOfrL30d7J0T7BJfpC9eTTluKu/Dgn0X3kO3xC90jmX7g0nAvltK9QENglynq0HWDV
i4+9CH+wpjFo3F5bF/Oe8JyHx9FqcYOC5hSa4UleEVSYY0+abC77z/Bcuj9OwO0yrsGiGFLEuNJs
GnCGFTNfnoDtPUQXMtuXHKb/QJA3xEZuo6rRSCEJbUoK7q0P+k5HRyYo16W07DYYKKxqP2pnRKaM
1o6Yxvv3/oQwO+rXhzoM0J6RMarA8ppdb8/+aDkowyjyPcVzSPclXxkHDMNgqf5OCcwz2F2u5vzE
3p/Yf6Fc0e8KE2SNuLNtMlfzCLusmsg7tbyPDh2y1oErwIsVSClDrA+kdFMXxyynVEf6cSdVSHlF
5i0jzToBS6aBliX3sTLi0KXZfhWxEGez5jdJU522dwfv/Hw8luRrjFA672hUdBUZnSFQr3jtCn6S
ZIaa7nvgqKLvO4L1SUFsJEaU/6+yFxXrTtDZ3+9No550LjHHtYruDyYFw66RMNF8Qw0xVAWxr+am
SLsyDE8WvdcInjzbBD0GD6s6xQBPqCCaQZftahkDtN+wACxo10uavEZwjqkyakljjjT4XxrXMEG6
NlM+lb6O8GCd9oS7sYb20d9aizb3kzR0m23J1iHU4tJIFO+Yj+6UB7s0eHelRA4qVzytSiW/GRTE
SjOxsoHecOKk+pAw8TgLHhbXt5Lx8FRgR+wxe6jMaD+LVe7aeeSW+AsDkCUncbaQWTl9jDta1G22
33YxphyYDTUZyktcXukmHE69ZrPYEE0OKAYWCGW7Le3yNGaiO/1oB1rtK0jr2prc45Ercubt9nlL
6FgIetC14G+nws36+HrFoPvovfrX2oHuaQal2PdfmHNyzWC6POv2G0JI7/1lQWZakl+Y93L+roxQ
Wz9uSGW9jk7NHJ2K2IQimNElh9F6DW0TeZxhZFRmeWF1VLmCEw9AisbWUmMqRL5kdauOs0ThNWv+
QLxMSxdksDeFoQESochmEjoPOxoMmOTfzJ5T4045440HPRbaR/XZPpzgy4/Msm92hbzqUS1wE6ul
4EHyH7Rz7RH18/e5WNcCjief84nGd1vDvkVbYbeHDKDXP2x9aYrBt/vURcigBXoaotUIekxv9K3u
xk1Mtokx+s97hG4EX2WYDp9hA8V88L4V3yCOQIZsHp+kBYdr8fT/ZIbBwjMdvosiuGSiFmZb1JKd
43ev7EOGQ8x95CygHDl0tNGL0Po1TMML7AATELUp1iwZDTvjdvznbyiBeHpS12/9Y973j2EUsZFt
k3XR8jHMZBE8JXa3ulwYyFrnDq9xKyf8zVChQBSF+GAzZlJO5ggwNnka/hkV3f1ssbJ/bbjkYsmh
37geBwfQJb/rMlepXXcTkkpWSJ2CaJ8zuaJHNoHB5CGRyvEWuDTqFoxnSq659PQ640BO6tXExRjx
8amCFRg0LRtu/80qY+QO9ogMIK7thr98I0d78baGzecoNFCoC3ti3fscB6QoF9cfRKGSrAlVlhKo
6+YZwaJvE/hbpkmKKIJv6xA/aoOqM5OGWowlFkcB2/0p7elDMjo9DB9SHO1uqeUCBvpLAa3I0KQv
nl0YLrnToHHDYq7WN8PGXZzFaNJ6nHfZRgFdlJhOfCGclFaVM6vvy/pSiP0JdNkiiaagAEFslaGq
idiFaX+n9CN+Dj3CUQrMEUsdycVJcLwEkhDBgdeL9xfBA297iXBU/XLctNJ7tyzf+Sey6zLDuY1d
oeUGtpnu0oE/lTu5vSKFOVttButjryBIAeW8QlaMT6CpiUvwQcGRar3l7gLSYpbZM0SApkof/W3G
tjDsRSprbzcQrn7vaG1E2AKqh14qBqLojzYlctaPyzOkeWgogYSBin4s2WiDWhuQEmujbDDS+4WV
2Ih0LhJYkA/eujkrJ99YQRKCfiwO6+XQJ4W+X8+mTZC7VxGvZK6czrYt035YvlhwFzoD2no8t/JV
NpJV+VqcMjnClbhT6u89DSot5EMHSVMsafFgmyo0iz0D9hE6oSsJ4DDYX9/syJd8/+0FJWm1PaQG
INI9aUCS5waoPseEqAUFzZTLXwufCnZO0E+oAsPaxM214f+CTg/ogL7wGLRoMTXT+ASuBSO7czuR
jWVapwCDllvqH8I8633ywyM1M58eGNuNlsMEv/fnhCy4lFNpLsLd3vuK5h/1jGNNRiLc59O+DZXt
dT00PvIZgBb32r6jVFnBkvvrwFlXrCektC63Lu6opT1watw2nk4dMlS8z2GBtFTh+6RTK2XNilUy
+OtNjwFLDk3ISZFcvwUHw7FNmrPdAlzs2FrA+7/GthXE5pXZkxC+BDl08zVx1cmI//1fen6h0mrH
mpJJmsxGSnlkPdKZUaTof7R2pfkC1WhBZl4KtyYGh1UXhx+NGQpLKzkPxhScNNYnhWq9BnVxCCVo
r7SvYsQLhcBH+A+72Z0UvhxOZrk+Ul6d+3R6txfDanOjkouWh/DgwCcX/Sgz0fAPjuoGUYt/L8KO
xLPnOUJ6hhiV+Owk1x4m1UoZMtMOPT8Or7U+UNvqpI9oPTFMI7FJgPJuw/Y/aQ2C1li9BnU9QW0Y
ykkwVrivewAZhKwyOkTP85pJmIX4/0hVIveLRxd0VNmpmGOXaYThAX+w7F7xlmqwPJU3tM/Fejq3
6YqL7BqpsRGqrjELyuP5ctqSR4vukRIa1OY/1nhIUH6Llx/+ctMZQ4HxA6MVqeAb+58nxwMXWFgO
jL3Kzoz9AsfOYJrEcJiOaR/iI/hAvD6hG0EW6QbPLoNryDKoFs9GTgiwg1rfUDbVlHTsaC82/gnB
W8YtCuT36HnT2O9AV0xxCkpcNC9t0vPvkoOxWxtgODf7hJoUji8wJ6SZFWQI+DA7TEguejAVPpxb
JoPSYy2K/L9rvydRxANZKhPTS8kpsTQFiHYjQT1pBYfl1Oq+P281GQf9evgkr6s+VUM2HGWTfeZx
4/j1xXOxsMHfnQkUvRgcf0VRNr4iKbeMy19Z4WjIeNQEoW9R7c2tH7sueeGoo/3YXOpeVBRzNqZ9
N/BnvxlDN/Yfyyi0IG+HTbkFnWAjGA1rOTj8Oo+9yUahgfR+ehqriPNsUxGKi/iZ3WRgRd/gS55f
0LX3KJlllOGs/xwIT2w5Mwq91gXehPvmci4+GYuAa2ZXZcVK5NjODrRu/DzAC+05ORnWxV6/eF/K
rABXlKzbSwyU5B3Jd+5ZiE5WAcjBRkp27kI4n2MJjJeuMRjku5TS4xNJM9SVJjOXxWzwSCYiaADj
mMnpJYsucv09BMrTJeIB0eelcydKLLSJo0FxYcwwN3PdJniBOg/9cA/NvtUsjXbrJiId4iWAMcQo
3KfrB/E/mT+yQMPnLEvUEVVBCmCCaBfIDQi3Ak6xruXRv/T68fTouXp03WQckrdrjJgizkTmqP9P
3Kg8rJpMZBzxokoHaluDEW5GE/ozXy1Sfnla8Sqh71aCcGaeS75jiuyFzhYetl2/0yb0OJIQLo0j
WmImecesZzK1OYj7rJkKXwxRjUANguV/iZjNrkRD647MVxGWFO+sw2QufLiu9L/ltcy7AnIeP0CA
zCdkGFkkBqyRckLtQwwYoFo9AqOht9yOrrGli6eTYgpPlB4w5Yo/jvcfEohhXvkDOV+1QsKfl7Nk
loSIeG3zYCqRktFSbb9d7+6HWKKBS4+0F47DPjBaTvbTTdDSjilD7o+ut6pByIFJP4Z+DK0QCekH
MGMczWvcwW8oQPqKjhJ/+Ru+t907ZMprixAN1soXMEX07hVS21bfn2VhH8VfAmh3Y2sQHh03jqPF
tZn22gnWdcS9bbttQmTWY4N7ZgJJF3aD/1fPQatEHyrKI24+iIzxjUKOAD+glFjWmq7mtNl0b2BP
Msecitt+zQH7WAVLZuwu5kFaU2N8Sx12KTUEUmy6/98lHv7Pc/lJNdLY8whPcWR9O7sYlR/h0GuE
qhrIeEh/ARKI/UGwx6K7+kUYKCwn8tNpojngFFWw2sXmuOEdk3cA9B2PTbLg4uspUjtWrdXCAtj+
9A1TGWZXxMmT5l7JWIke+yavKDxuqNmi2IjJDD1c+4k4uCv6cmjN5amFdizKd+z+MAkf33fba6UH
mTrkCy1UJswwcechKDYb/eQ/tV0nkeeam/kbbTDtf2E2rf5EM2EG8HOb6swSxQufaQYdpAUbN2Ja
ZrlUpBqQ2i86FkWpPQnz8qO4SYDdCQab9FaYjkhOirvie15zop5z3ILJkQhD4GsfsD4KeA28KuVn
A5mJgqUc7AWg3RcpAKo6OalU8mX111mfBj7HtVspTmZh2zKldI/ygbApv3iqZciYl9SOh8ihkWJj
At1wIKbYAZ6cmybqtu7jxU69UtBCGe52O59/H4pq12RVn7LyZQN81hoWDUz23VPqgDAbQdSkcM0t
0RkMpFwQQHRKgNEsf7vJwmIjvOex7JZ0f1Z0+OAgjRgdBFDKF/Ygj2HWzvZFCw8lgzhnaRWPWuyQ
T6LiHzNaXl/YCVZd+ZnN+dR94cGE9BEkqtAnxOo++QTiHYctF6fFDmq7mHdcRyoItFSGXOaw/dus
6jyBluRYb3UDIcCfp0gsdCs13lqrd6j0nYpKsa/+Q3iH/7DatnwfC4ZX+NrsIyZawjfDhZdRKNoQ
0o/nUC3chC5HgytfH6KY9cdgG8bm6ZHAqwf4OAApURz8TyuNBBT7rhhnw37ui4ZeOeIPNSzzSf9I
z8mWkMd+io6wIQ1yuyDGnWVK3V7LFWsubJfaom57NPSricIl2YoZhIoH02LPTfwG+HQD/DkHDhcS
zBvBZ1DVM9Behz+OkzwPnBIpulos4d8FvW2/kjPSOY/3DXyeCjAt1K9oX9Hx2D1ZP5EFHWPvhYpH
NIyh69wQRJER+jSk9TsmLwbOs2+cP1eUbBSk3vQJkT/K6P6OD2FbFzCW3qNEvCSn7+PU0pns2zdC
D4nNdPoTISAe1j42C+iBLKq9fgsg3GIybC2XcjOI7cQKvnN8BbWt6k+bCe2lwWGZhhhG/TD/Y3f6
Hw2kY0XN0OUxpaXB9Hmqmfxg2sJ0n5YYkCYHpfWuy9MS/MVpoBa+AQERYZGAwOA6Hv+9pAyXYie1
2hRu0hs2U33cqCAa37nJ0huPnfztpMw8Z7lcfUPqXcgp0gcbeZbynMOWf+pky6EQ5raam/AGDPLc
Xrkoqp9+Rm/vxk9jMda8qSAUhmEsIqQMdE90b8z3ffuOduVqqXWEuR/qc9LZzV8TeLs+rd/vf7Gb
eNzNb24BgE9LP7C33ro9blLm5xTc1rm4np9jIkO2gMXKNKkxI7zO31k6Wj1iZYVzNBGpKRwE4RZf
ZRpN1L+iDzrrRKKdUoF7N0r9LBpkqyVNDgxnylFGyWgDNynE7L52P5Aym1H99mgETNEGQlZWnYF6
/DVslRORWHl4eVjjpGY0kDNoxSR8dHwkZ7zyb4D5xc/d/m5cWm7VpwCPN0MBZ6suhs+3Q+5HaXB1
u6a0hbdqA6cx78SKEpM9FAI96VSdUn+XmHKcEGd7jLkO/GT7SHXybRsPhjHEIkFQ1zjbCUmaYkvP
Lt+FESNfr6OahCNEko2aj4N8Q3ISWDe6Zwy9bQcrZWz4S9GkLN4IMnG5XSswwhqndQce6nX01m7Z
4tYJnnqo4EoOLxwavUgcJzUDrwSZZv/1cg1quq8m/lIqS2wzT4LnoZmctStNCLqvO30MnS9eDTA2
3Lw7PDHUfZktBKjx6jSKa8xK7HbfFkR+gTHMsGrTwKdFme0x0fPMirI8boRyDZCEFf4OwDDNlid7
jaB0uJDO5iIom1thUYTbN1FPo8rImiiYQKGWCVd2rN0kdB7sehyVxRL4ZpVHsWRoVOilNQM9Ha8F
CDSVr2yt1LL1ADE+0oCuAPV/9KVuG7/58J1+j2Pi02+l5Uxpxped9QvKcEmhSq6itW5KXS/fv0V9
T+ZCBwR6+AJ+CkXP9YxbOX+B9CWfhfNQGaQGCw0vDdXNpVWsmj7cmrvgNuITFuCZ0GVd6x64ERQ+
E5qqfbWSrv10AaLFjSfxiPkehom8+pb6ik4a+jhwaeSXiebdTzZr6qFw5NSQuSLxw3/WhRituNMU
8UeVGRWMDqhuWzQSvIvPEXughGgc9GSPLpKFt9kOPpb8TJKb07XQGkto9TCv0NIhm4oNH7PUvPKJ
vw1O1Zs3l+KTMNIsCAYCl8Ykdyn7/VP3eYaThEm209uGI2vxgvKAzkzivF3o+JqnTwWriePfGEde
7drtp/luMspmoql1LQ2vZBlK2qvLmisxuxLnFYCQeVsLO3+LAojyc3Mhn2rR+/DI5jruZY8f7ljL
5XZNXIdiXuE9J5nKSroebCWmpMIRR1ITgf5ZMFEmzfEmpu4Su8qR+koxKL9WJBS2+aqHi/BW7loL
jgGgaE9rEukNfZIbXG7w0iXEZ2fE14X1J7yE+HN+Hhu0m2zIZutAVRXs+bKJwwEsi1qDk1divZsn
RzOoCKputNfT3awYJX95TY1955lnLCk2tEcsoOu5TWwUdmKwf3ZCDsa7PXzBk+Ohw+y8STH7KQHF
ibOqUXabecv1GUp6gS6/pW+2y+ZAX4c4YZV7JZhfFsJm69/PGTu6XXW4Jbo5l2I6GdIJUwvk1ky4
nKZjhzEFurxjgo9zTHlYkYm/yn0XSaf6pFLDj3RUIC1M4tBMjL4Gx6cVraXeEI09Epqm4iIX7cLy
qBObKydH/qNzuQmFyU3Kaen/0/aY4yzcm5UHXp3yKe6suwqGljO8jDMDmCH2joGSJFc8kmFG3I1z
WzRmSPfZ6n8So4KNfhinZXlX8FmCpMGR5YZWlkloyM/eYDsc9QFyzhi44tqSXyFsQCuo4Shj0+K7
D1QqLeUOSG96gcm/yYQLRDcRhbEPat4kZTetAS0KAqRoBIVYEZ81XxhFdFIEys+jz34ueoRGryEA
kvuo8f9gQg/MFBiyTa7WbdnpisljOM+6bLShdXVZWWmmcNhnAeLq6hP6ayIi6zjNtGwGO34Y3H5O
FLEiOebWtVYTrMcNHInk4JU8s8QhwtxA3zlmN77gr4icGcZjY1G4+H1Bzh7YoY4O8YtyLtZELQ5C
SJEk2g8sKKmhBLKUCFcaCSi8HEpOUXtOZcU/YU+3tCqaQP38sqoGsN3FRxc3/vhz+z59q+EbnK9h
DxU19soia6NY88ruxApAOh7cauiDCEDB6tWWutlQN5caoP0VszV8bBCNeiz7zoXBQclqx/hBiw/j
SL0224ogVU+xre6O7t//1G0esnAkUJfuLRPLbhXx81JMhwfSI4i+QqpBNyW1awWkTMHvXMBR0LOD
+y3nTkWWZwJtzNw/9qu42ipuRBEjh7oxc2PAr+ZGUy2foFz3lxTtw3jiZsWxKEakyNruqfMrctO8
J5unAxVuqyRvlmX9XrXdzlwqeoaAOx3xaC7ZXq4PesYspYlhAG8gqmfcMf36JVixWNnmV0AwWZIy
6MY85owXejRkRkY0fgZOpKwcLs0yCV99xafgCtsXnenXdSwB6lZ7cQNHMDN0aKiuONJmSSKcFqYa
CPxVbIbncltoKg00MjUlJ5yyW9+wpQIoT8BhRO5Vgbj/r/CYLU1OQ3oxkh1+X4jM5vkxP+RUquhW
oR8CU+/UdARUVQ6OQ5JJaOJRrRf/5DbP4e989DQW+2ET3XIqaXzPh1l711P9nsR5crPUZV4MZ0Qy
oasFr2TsG+mXlBVav8qUEJbHog4zfo4=
`protect end_protected
