`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
crsuNbGKr2+HGjsnrWAO3ApjaENLE5lmTkmDpqy6wXOqFQIJnrktoh4R9l/TVlY/BEwSOhFtvEbq
RKvf5np1ZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfoL36fNI5DjzIQX15YYPTK98uQI+Z0aMjl+hiAVWq0lzClrfpDjXWaPyQGiPvnYkkUnnCNmSyGP
qGrNm7GOsjezCGzMgQVr0792OKktWuV2kt0zVP1RUZuHk/37eznwh8N2o5rw+1YzW4dGzl1QbJom
tmB1UpBcp868gDBGaIo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nZKDyxkYA9uy2Xb3FwpEri9edMFM6SqsP4Aed0tRsVeeX445M1QANBu8GOl8sJ4QNxr6T3VU33/s
FK93SNbe96iXZq7rd0ZTftDGFn/wlb+m7r0WSjfp5pkNrLXaYMROFr5Y+cSF68dabG3s3COIhufS
z6LjxtxffkVZFl10/p5NYIyhVlCgj28/qTLowb5EYe1tZ0WPUAxBFuTyFKtX6X8Ha+x+nETiYK6i
PAhbV564AhzWOG1ohxDJJcn/sq1JfdeuDFdYSbNKycH1TqhYGY4rODz7EB10q4+UCVziUOr4Tv4R
NCotWnw5vu+fF2mIxu+vVyyYTSX+rhEfPs2iXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZ2XWhB75BM0Dt/9VMCHTjvBqUtECoyfIkFt8UyDN1IrerieLUkQavGMJnAyOgfgB2F9GkPnzVQV
7H9tsdZ87Y+A3ybRmsawN7gt2tqx/GGsvZlikuuSepi3sHN1vWxch8VpcI/SFn7CnlCh0jupM6VR
707+yLDj5AJkQVyH1LA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S4eCKuneguafnmn96ntdnponlGVTmyJu6zrxyF34ICbqsowM9Vhvgm6poU8XDQ/BrjS+RNPc37Fg
G4CZX64FNy0IB8M93ARmuOVvrGN2bYMf3jNRnVO/z1hOqr23u4iXXLcNjJcX+q+ntygTqDn+dkJa
tNf5JDJd7KcZbafDC5iOu1RcjafQnwlpqyaxuvNRdQkJM7f5tDyB/fmqWMaeSiYSf6cbwC2Jk6x0
7wUP2rAkEzcYQjkJqSGT74QQ9ZxpJuO1xNUbfsJDlmWbSmEyg55J46Q3XRBw9O4UV1TNB2XnSxvt
0rRnDIzS8sn75CDPR31VCmG8K+PwSCayofA3ZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15536)
`protect data_block
HGwVbJA7sypyD5yh/+WUmYczAUp9Ilw63ul2foAahIAqxWWNlG860q1IJCvcDi+ST5/TvxcuzPir
qt27wGW80Ur84JcU1ohvXeBLj7wUxE4SSH0YZIS2OeLGptmd6Woi8Jn1Fge00NTnYbclpz/pl2Z5
tH6MrZQ5YNH3C7MpE4g9nfQ3KhEDCIlLawmwB5GKEKYdLSGoZYR1X+d72CfqT8B9WGCcFGZDUuRO
vxC7DFNqRL/7XV9d4CN/wmgi8Hmq9xjz/4Rx4CJPFmOpEu3Nor/43vfLwppLHjGNuU15K/zxpf+M
lUcg79DK0C45qoWNi7BUfANh3mQcT++RpnIeqcTJ364MtsB2IF6B4F7WSh7BQO9kjjwSSdIzAC28
5VgjnECfCYskL57jf+W7xhhdNPlcWzmVogOVaczKoxu1U7jeEXUMADDkTXtIIcD2yoHeeCt8Z0fe
CZ753l1i1WW6lF53WEqKqHeGl2GxRQagNk7sLnLpT04fywYJ1FLSMt8+4yxVLoQQ9glps+K9qLm6
T+bgle8N6vtV+vubvM2R68jZgHlIZ63EeOI7D4JKXrML5SMrTGhTD2dfAAnApjS6z0xL8TkyZ4Ui
RhtoyBHpguv343Kk4G0pU1aeKD+hinJbqudgy/srXcfk2JYhkMS2jG99dOj/d4PwBu44wZaJsmBa
4g2jfcNgWkIkAxuwHSfus9SsZLopAhx8C/u1iwc9otxGchzu9grBIDnOlCQtBsh+xOdcsGJF0rFy
OK2NSkLE/2DYkQaQ6jxBv1kxZXk38m8vJ91MJcfNVA1ZQChOAhDVb5S57g7qhQnym3LhrtUxaT1n
kBgguQBC2c0ljhayUT3ArAmVaRKSipa1ZVs7stkI3Sic8J4WNMaC1KVGeLS4cQx/7D+82CfpXBEs
cxpBnzj+j0hUNx4GnwPU0BvhQuUlEQ5pcjh/Lz8MS58u6uG/88jOjTAXEqypCcnSCweCmy3RjYla
wC0kH1AsN1+wT5y/sN7L4LVItfX91zbohq88CB+ySFUyAiyYIDb1b+Uk5y78DRIFgZaiXKarufuU
9NKCvJ7TTINVVsuTEY4MytwrpHc69qbDMFgYD1Be30k/hTRS2Lau2u59TVQVWywoVDVmT3vIpiWK
PgiYWTZyb/KBqXrmtzLpTlJlf5YlAYYQAipaE5Y+MSARC6wygUZe+bpdIxzDXjFSAv581BK2phz1
xycF3aDTGXp0Qcqhh+em2VsK2GxT8iNMhG6+IOF6SY3xp4gGRt2NHES6dns4JcFvWs2CNSJG/1rc
gEyrB+O2hsyPzphDzJ5/7cSKZZdTUUmJko3GleV5s3x5ngDxIS+TkdRMBMQiXosBv/gDJ9+dcM6u
prOd6wH2gWjzoGH25tuG6sMC4m8lwpR5GfgcYGQgPk3UtxG1nTAJDFY6ZaKmrV4IRuJSy8fFIEsk
C9dYUseF8jT+5k/enbwn9NrWq7G7ZNOac/h+XGMdedmKR3yt1DDj9RS6RjX5wgkZ7brOdhHsYyOE
WRCM4YjxppknQNG2oQUhvG6MXGH9hhGPXoQ3Wulc1dzz4RMyZgei5QIfABiebfvetIWJLZwaeg8i
+x/nriZsijqtehbE4xMemGaOlNghdy+5aZC45UpBBbQfOcJ8gzR8SoT19uAUixrXWegOu9l2BGF4
D8rJ+39+K1E0ZHf11APC2dHOdlR0mcfX71g2inoQ1dlx9gbqE2xucL7ZMOqdm910k6iHCHVbYtpn
XR/f6k8wyz0570Vw33RmBH7hjP5ON0x1/FrqIA1yM+bCOyZwlrJix1/2LugUczLNfNS7xLim6G0X
Q0cbd3Dxpbn7I5V0wSSVIAYkxTlnYhoDLC4kjzgRySLMgh0HpkqwxpklFgsjgHX5lqXQ2yJHso9P
CmghAzESeVd4RUqEpoyxY6ZMxjSCgpHMm0alGm/aOrYxOPYCuoZm2idBdaZGeSNsG7TR4/NMR+7J
Jf/zrYaKOxaEqGF/Zd8UKftRZi0rMpvdg+bXnDkQ8v852iRBndh+byJ7dQ+NGfYx9MaFnDPt3Imq
ZT3r0YyXt+XifiNXCSIUla0WTrS8K3vQBRuzU6GZ44owA1hKykYk5yI45KQiL5jQQ3kYAQNw2QdK
FWKHbYZSh6Ub3skCsCYqqb5QI8q1NwMpQR9MhPr68KdO1evLSFb/q8T/tscTCPEMe3m/gmtSYCqk
ExEimYO/yovmnbjYSpMasFPCOJbxTfHgZTfwPvmm5shiw+TMc+l64xt1MK0obwSoLcW0cezQS0Q8
BXTzOAJcP0MwwqJHr3jtXo4Yx6ZOfuhlYikRo9xfJwKcQZvTZF/ByQzRkkqnkNyfmszAjKY+shvT
F2FgDwBvmxXo8T9xirKCkRpK3JZ1jDofgsf5SHW83uBeihHyPJ85xGKDiBPMvRGsxKKoSvWEcb2m
m1/qoHYNkmMEIzYLbHJZN8pUVP3B8vRMC8p+Vjhrr5DRI9UFmeGgUA/a/BMGwZbqgor3oAQvjEqI
6dg88grtwYLumb9nlU2q235lhomCAkrkgo5FAx2TRRhYh7C4orrXqkYa9QzH/+Z0wNgkxZ4oNp3g
vVRDH6ovgghGP60ijDhBwQo6foctHitDWIkPVcATz3g4+MvdHd0+SFGRylb00XsTll1WQ997NmJF
OUPmSg+RcbF0WAlnskVSn8tnWE27H42oxTh7K6n/cNEAEwQgeL7ukBWR2d4+v1e0s/rjp0NLFFpG
sHfg6oeIaibhX9mVgAbp6+1hxJLYecpApfvu/54+gCT9LDECiBJx0ur4HD9zDMzvISNlR5wBD498
2RKHVqdp+XEQ3sgoyz8lsuW5cr6dGqHJpujUN62iI3zsrTGwtGYSYS/FUsditwwTw/lWIRB17RlL
a63ghxEg1BQ299YYwW94c5Iw6v3Wy076jPLpUpf1yv5Hywj2T3CzuvccWQO1d/VTaNBWAcn4NNDh
DIMcvWSJ+R/NqthgdjHYZYWdfFXyVt+z+aEUH2RetOpu0kCJIHs/r8vyugWpOBwoP32/HIToMBsR
C4lcFH6U0nCagn5DF9GdXFIMdfZiKgs0UyGTSto1DfLvxNxUmzL1zYUt1+GqFOvJe6th9TzDx4SU
sQsdVXX2K5M9wBnSoPdsbCP9Y09sHWt+MQgOmg5xqvAC19J6EOdqGaFN3Cb7C63kvD1GWDEBhbz3
ht7ZlMYu9efq6eLyGXWoMYsSvIzB9mPxxbhZ+uhFdYA8o4taq8iZpxShWFUWumlgaBANoSquSnC/
CErE/L5SQ8AGr1/pLIQzlgwHx/EUEeQW60sBNrI/2pot6ZrGfNUrfyoqgLeNz5mZUk9zqh/sxAJ1
bag3ScQm9cpVNoIUK1yl941JtIgh9nGC8R4nLyXu29jIK1gh3EgOiycqzHc9ATi6SDrNMG5xsjXs
Q9I0ANsOo4H04W3kAhoulgOxX2i/KbDic2INq0ftOv9qR//YRsnNRF/O7RHqZcCimkcLBvtkgngI
Zxs+kskE6Cl9ofklrKId1BEaH0JV1Ft5mz95xTAuO25Z/2XFe7qRE2DR/Bc/1xgWWhUc5pvV0cTi
duD+uxhb+0zNR89PjU+Gvo0n4SRIyFhDFIc+GjDGlIN+h51x+9LLWGChFh8WPYjIwq3pz6F3yV0C
Lo8OyR/FF7fB4Lu6MQKnV/tDhdofJhxNdCeCyebkkylDrX4oWyjE/8LiZnlVkctsxkEEZ7AcbBVh
DsGhGvOQLln8PgAPioxBhdS4Ycd3HSC1Sk4eQY/xMpppatGEvfvZpVfQb2nZQlef3MmqbG+E6hMH
LYXFf7bC/bx9asPqCvEu+aPozChibmwx9F9Hw74EuwbnIZOI914sWm+6vtEHSa0iuQjggaRNgx83
0ewk0es1NRf3GVSYuLghmzclJwtEMGjPhrspYJfIuFMRqU4R4jJwsZWQipuouedpIoykLlrD4LlM
Yxyv19dN2XEL2TwxJBxCSta6xLIzzESeywjjNGMgssS9Jn13HVW5xvyiNGG6+Y8sjHW1bEJrmWVS
eFyFjv/UTHgK05ehuLn8E71qgM78uDZCnqFz9xTQ30AQU3iG0eFTF+SbZve+cu6xVNrliu4OhDHB
MhCL0RBjKq4jpUpaXNWya6CxWdN9I5f0/ob3tfpe5cpgTlgx/LRX6ogp+XpLgOXKNuEJRGY6GXKD
Yy0+nOOoltKcEakTowrZOehx3/ZeWp+Nuz8nwIO/mHP46/6M7C0dytr3di64r1Rtc3sSORSwuMyQ
z+qpFKdWIToGRX7KwB/ZI7tGd4Op6p8L35IRO5b85WI7HYjpkaPA5GoVfmC9xt7s+U6Psv07O4m0
3heBCcml+XfNy1upfisPr+2faMSbT8bV7+qR1Yvd6rerlL7a72IJ0plkZ2NlsuhP18v/EfyeTgw9
CA0JvyQjEeLJX0H8O1gA7UdHQJZkI4RVqjHeBjjsIPZ1qtrDY4bYkJoOe5C0D2KsduEnFgO/o282
zHJ4xz2D5e2vb30fanljA5uw1momaAj3xIbMNYTLxyicFtXI6nBO5ns8XGdStowo4HBowzKDx+UB
AtvaMs1bwdp4B6vVuNbdFjkKb7FF0LgkNyUGm/Rwc65rpzU4PSutiPKr4k5iTyRFpFaGnwdIIXtn
/HE3nEOyUaESh/zkZHYkdFwMVAj7x4iD0/Xwp8G0oAMBnbv+1pHWrlXyKrOvbhvwIyrHvXcCvRcl
CTLWFCOxBJHnsr8OVgRed7QouvrWiQRYzG6MiEWFxAZXRNrJod2R8+fBFgTnvNgDckHmUmaXeWZ6
gaxS5W2HGEGzrllCRWaM74cgida//VKrq/CVwUdryH+fp8HVsZ5y7n+K2lTX4IIkv4hS/8Zdl8tw
hAO4qLLzyUBvDjZQmDZomx5vbcHX58QOiMz1IYeHnq0efUzleyxHWzTMPTDScx5pwZuxQwjIwkp1
e5dYSPMoDW1cMl/H/um39ohRyfTe+qUg1IZ+zk3BPgHzcAr0DHNJkzr31bTISJZKJClbeOnj0tsx
H8b4nlwYneKZFe1Xj95uBWQDXpzGcblnRpFqzEJKMPSB/0pq6z+QD1IxFroBZE0tYfMNYVLVm3+9
8GyFr4gAdzVaApc/YX0IgcAHfCWtijuAQNJeupLbDZ2okxQyopfSp0peSICjUtvRXMVdohEg9SFO
hl3aFzk58PPVyuTGIdYX+Py4gIe3Dq0BJ+Wep63OikyjIHL+q/v5wDP1ns+qaU14svi7cXQ/CqXv
yZb2KOFai8XTvvwdpT/gx9kpXxcpEDfMmDnLi7xS7Y55hjPiSvVwiZ2EBLfpWPqWU456inlXiPcE
3DYTtQKctDtGFTBxKl5EDUYkJQNZRwwrMfSxnwygXfb6d+FTXHVxQtX+zVmSsEPmh76d3x8kRbP9
yi0qXWjGGucU+OwI2XeponWAsLMNJlIMOHgVsG1c5suVsKAr9Rz0BCGbr2FttJb8kG4a32lJ3Dej
TKjGJdjkA8To2N6qitmmlBdVsOj7Vj/WV6HsrlaG7+JcihR5rnoVgbWQR35xVd9QoV6rXtYpPBEO
YqH5v8nZcUtndYDyltlebDuEyZaCj7NqPzTZLLVTkbjYohUOOFFCm/HNZ9LMY627CICucmIrTsl9
pDVN2SWkxeJzEi2duK06URc2Yb4E/YIMmn91d7PfqF8K5l3i3yoGSm9wYflRybOt9yvZp4UQ7IHU
vZTie5F9r2+mwk3DrlYdgi9KSbBrVM3zbDNHaqC/16C1uzas3TwFY+ZDBi5ay62KO7h3UHRvU9X9
2F3uicW0OE1YRuL1eAz9huf3N3tH8CNlGTy7aRmH6WjTM0xz1z075gWEKCNwpCUbONtDqnaysq57
sXMOjNiCVCl7brC3eDZpRFXwv1au31ALqe/9DFYCNDDyh3Gy5uFmSVYxgkhiBtlWEaGqhrt4BJ+M
RS/G4URJ45VOcOA0Ud3SPnNrkjXKVA5rqNpdBIMEeHVTEn326l8pFWNJ2078lb6lx20HPp0/qhsE
6Apo5vp/5BugV5w4Bh4+HqZjrpajthm0GW1/GotykOIkYs2ip5qpTBtCT93TpInXqgSKEU0D2Gap
BiF+twUmkTaZfc5AjyLeYNHCf37tyo41orTUnyZD8cVm/D/TekX3lfQX9q8GbP8nY36NFZ+gjAoh
Tkp/5mcukaPxlg/9bj5T+OIRsdQb8FZH19KfYxRziVTRZwlsgQ1vWoJHHchEOSNRrLrdNIKUxlOC
8nU0hA7ffbzacNh9xjSruK/74UQo4UG8U4/j1W/RexKlchTK1iqEYC8mUQRskmrlNVbOYnBubjjM
Hotyd+qyoMUPde5veOnP6x0g4e8TIJlC+zvJpR8volGqA6rs9rtGbpjrZ5bLMO9w11SgGrTowR0w
HVnA4tZ9wYIHKrQyLznfRyrjCGIIOC90fcilQHZJrV6grtG8gjos5zzh+4VpuhgM24WTkpKOxsbv
swHvrTdUYAxkDxfCf4aYWX8WFOulGfluVd6KxATQ6F1X1widqbN5eTVrvPmFV1q/bw+SitC9048n
pP/PrEhej4Dvt5Bz8Zs8NruxxYCdN8QLQnM46lS/0jNy3DRKuUpSteQhEegonye9vwtte/8Rm/eC
KTcqVIwKtEuOv0RRjR7CTmLJDcSLkFYR38mYJZLi2YHAQltpUa9rVG3JMcZfWTP/C7p7slEUO2gC
Wj9XhB0+5l9pI3zfkjPJawLpzgCXdH19PxmgOmX4m9iZANMO8PTcACPACXZ027x/vNHuXXa/CoS0
SDMWWDlMDc/jQIUnCcLz2daL0EHLsKIGkX582yB1D9+DTe/D/u7p8xGp6kmzIRckcHVBcEHqzsNu
Vtycng6aY+Nx//bP6PkDYlhOOndtswL/RIwxQJ3HcE5WR55Jos9hXMZOrBsp/+Z9fbAmfL6D/0f4
CTdyd1BNUK1FZ2HD8nM3KoCsGgSU4ytgzU992aNQOqZGFM+eCmwxLsYjNPNnonKnIX1HFLH+CFvo
8eFpqBAi++A1cfTvmdyB8NCmbt6VSd6nhvDQEwhgJJflHOACxQVtD2gG2YQuPnR+41RNpaa3kZYg
rcKmRYUt/8dtops1BNMEPkO45jbIudXRypMTLBv4p4o3VyswmGkPBScehn/5vFf8QVirG+qUaWXq
BcgXb7wIvlCyNt+gTjwfVe4k5lZ0QyaSmNmdCeKiWRZzWdRZSyexjIRY0TSd39pn4pQqrn1YFoek
UNPM0DxnxC+0M++tOKEQW/wp3TzRMARVvh+AWl+NZoK7VZd+R0RJ8tPxMXvemk70FMW7Y++PE5T0
d7UbYvvsE+MKHBFB7+3h8FbG+v2FD5WXIRvucj+rsEu1g70N5sTr3bUf4hhUHN2iqFy3BrDD3mQG
Uyr9NGeTIrwHLuZWHnceXpCTdR6umimkDqbJsCRRMq2rIUTQWkdVmRSztXBYAxqx1dNH0bOfrnIX
bpq1JgiRd+vWSrRwgaZBr4097ieyyCxxpoH9Qj1Zrb38QfC4FL0cg9WqkC1cfwE4jz/TQGMbiHtx
lubrdkZYRow/IqVYbqOkC3hLodBHeSfVYbMRj5cHrIIrgl0KQ0A//dQ5C+lM/fk0gA5TLkGLDs+i
SMXCeBavDge7CPIkggdZ2EVEIEJsgPUa3iuN+d3mypjTKtvxL1kjzjbaBrtke0CsEwPpwXu9efAA
4OtodYicVfwO+WyaIzhM8IqCGMqPoJK2CgfdHt3F4aFiyBR+gY9lndIMwhlDp445lHESsmQrOZHX
0cYEWweZluGefNpfvt228yzXQQ/ZHFp57OkdhjDH64MKvZjIVJra+GFk/uX6lujCxKhDpw3UayFv
6oodyvWyMFPKYQmY2c3Oe8Z8poEjOhiLPwvgsVkfbQKssKuI6M2Mg+3Tnr/bQ0Kh9WfI6nfNuPjX
/jGfHD0TtxN57TzMnfEPBYRZ3yb7bM9RcZsxvZE68G61II4kC4B3md5QIb28lwEheEQNVc+EZxfR
M64TTIjGHtrMJ4f6xikT8Oz2JP7HoEtXtKWSo5r9P+oeU0OIekplNzg5VWyvHSADMnCRk9x8Yt+I
MxniQol8mrndWWH8uza29or5btrEEekfSCKcpnmSmHY6x8D90yETIhg/E93erZ6ihriWGWpvB4j6
GBrjHyTNCCyBBKsDNIQ8PbHtTFC15EzfJn01ZldNmbClEqxO8Gg/aBjyZ5ng3lsPVEriIljVhYfr
deOlO6FfX98Earf7tVrckhgp/G9IkvyO/aqtnR/KmhkhCQVSmvKhWS1axmV2+pBoijOamAY2W8Ek
+loBpE+6o6Tz/+Xk64MFVa6kPpYF8UREMzrzyAAR9eX3UEL5g+JH8YNyEGR7zE1SX8g+HeXyjK6i
mViuMDRli9lFBPzXYVbORHtTEkkhjU/5cP8qUwZSn9Shz/DTQm77S+gZiyR2AaZAiULbdNP6I7gc
bVDM300hNT7ABm7hqpjSGGy/6lsYsoXxsuifwCN2HwjL+/5zdf3Xn5rUIyoZXrVnL7DujIMKaxrA
dI9agzrxzbwUBfDL3jWtpNRcH1cM9w6cfvfE0MELAd/T9AsSsSq+OF7jIMoAEnu0A14Ny62/gN5i
7u44UrjF1fhNv9/+8nxZee0sWJ8J1DLhVp+tkaTZ0rGxouBU/avtFxKa7ScAKL/5l++ESnUjoKXx
MKtL6VD586fM+Zirc5FbsW1je4e6M/ya9EvKc/+PqgTiPErjk+NsKqAJGeXcypm93ULHfU92E6sw
jhFi4tmR+AOVAq7ZZHpq76N1twgNVYZ+aDWm1iApbJWPKbpWYep+EDPPvXOVkYXaP+RzPxD2mMt4
GAbfxEJCY9AaZMlSSHhjiF49NpSJKZ74ftxrctUZvr4wvxGAV0ebE0IDxJNXQx1ESBNTt/YiBJ9A
UBFzsxRWjCDahLV4CWA0qclC95W63W3/Wihun/INP2AlKGWaxAVFT5AB7+QGvJQ9PbRrI4sp/xFS
pWzlXyxDmU6dlyp2xbw7ZnGBQeHbaMpZJrM/j1MEUSD2jiI+KCi9HY1KQWw4540ETCjDchcIndtE
kN3DxXruLtzAR2saWNxdzVApBrp+zB725LXTLqhmPplDVkUsUuPsLMlF29f/k/N3T8K87YsEMaPC
/62RTCTWTVSYa5/0Tke3AyagUhosHAKSvS/q4H0shDKujbYoao73g2lr3wSaiWw8BdArh1g4V63b
sD+xTLsAHjFVtKqPa8YyAK8JWCYUfEDm4Fr8q+RCAe1kf1mBreX0XCJR8Bl2DFE3JR7V1GBzDhy2
QqbGSTj7Ql1UtGza8FT2LNwUiaWuc7HNsFyWAT04dkPVD7prXfg7qhJjU1ymhUMK8H6OR6WKM2Fq
awY2iDd2NUsEKFCLm79h/cizDFAluTZK34VlQ3VFZWRhN38cM4oRrqYYC6Hk0mGyk+JwUDn84VJZ
39zD91klbSnKCU7CYZ183axyOI9chMHQH0dzjQJnf8Uu3FZ+qAY5sbgBXSTL0mtl9HDttwcLuIck
4EAVx/1hPNdY3o3dkUEGXImrUQTnTVdARD+p4NMb0HomHZ6lsYwmfMbOgZVIVDNCi6rPeltBUle7
J+xy+zylWGQKEmGkLLBRiLDDZehrwJYPQxcp95CLSesyn3TKjsNenAQj99zNq0SCGZSuQZi9AGo4
S+bvKKFH/HdUZL6pTOYySUbzzjrUgJObjez2iS2sagcNl7v3QYlF4XuAEdQ0pwAfxSNGxsY1hGTl
i4o6fiD659xDInaLm6gyplRtCJBOW79XQyfRNjnqIv1rEm8aDjUA3BgBnAIH01xpB+hj5UX9Gnf2
xKTD66lHVpyCyDyO471MEo+umd1RTocSt8bo6hLJHKXKMy1hfNqaS0+UrgA7+9Lt+smOUibl1wCT
884tVRcf8XWg6n5UlJwK1PlGeUDvCNVKYnm4hCIAE40avE0V5zpc3BNbxXcEOYhMCRwwgtxT0Qik
ixyKa6hZba92UDMxn51GOmx32jC4Tq7ikS8RCZNrZvkvtM34fsLT0BadBJeve0hKy7KUATUOCRNi
KYNSF2VsxZ2+SS+raulg4xCYQNebsrHhnWn3iwd+ka4Y5PdzU++s+tfG1pHghoGG4uubc+/Jclyb
D17tw+gRB9mOP/wixo+xtBJV6eUWT5q2AD7U+EtcGLNjq0eK+m1/zabIWuvNMqlFaKLAqt5WWLLY
iy8ph6YKM33/3WI5yaEvxNLK6LYBNmJSG+avpcjXF8NPass2DpqJ8eqJjb/e7Zb4znubhMy/HG8q
Jf77rkYRD3vV+VaRFpXu9T6vRsQDbOpfobd4KKdQKLPiu3CnON3KpmeIrwLdUDkeLoDs2wbSkEwI
TyAU37ovLuwbuwLyzupKJSnztsSB+3b4KVBPYjl0xAKCtVKOt0MhTMMUEVgy/Y9rgL7YdkGYeF09
P3Nkyo3S0dzmkr9t2jePNMtr1o5R2T6w3dSXhHYugjwIDrZFQq+QJK8F8VyZ5B4dxqFoD0NMozkH
0XGwuifMjmv86DAcMcprPOtsoe2R5YgP7+jzvzqT/oX4+C3vggdfykGY12j8K4ykoalYlAtgtMR8
E7yldG3He7FnWSlzKIrL39rAe6QXKFc9exdghVgnP8gIz1Mp0SEm9mgjzPMaVYpHAUAqDVuqUX0k
B3lQKAKFNZsauXsiQdWxJ0MXwBnS45VHtlMgWh5irvmbUdHpBIXD50ZvFoQBP6Tj2XbCHmhjY5KP
QRIlnR7wHd3JxY3LM8OzGkUE0Eb+jtZLM0ZEPYdqzbmkID4wBQgYvEmWR0QJZghAXfNqyf39ftbr
2FguEz5oH3lUo+EJmkK7+S15Mh+82dTo4FbAq4gyWnPWTloPisK8ZD7f2590NdY/IZM6kIDbOK4G
Y6Za3AUdpv94dzBddYueDxwYUvKHRPxaw3o5caaZ/Y3IplFUX8+Ym6hmFc0ltsJUJRMMB/Ogp5gd
aGJMbbyBBWzrEflgloarYdors+omU+ISsAX5mSrZGxMMb0ys6t+ukokaEV/EsBDtzpFNROoK3++I
rWjoXbgvZnUDYY4oz4k/H76a07P5nRp+qRDYAEXL4SF0wMfsUMhO1lg0VrrMTissWYBlhc8j2Qhm
tPig/MVb7Vd5rOfgGmo8nmRIWMRfw15EDePg4fltlVqzn+QK5ftTWJ4ykJJmXy7BfoMS4tKUTEic
+sKK/q6ijVGs/OSAk1cq0PsWmrulaNK9FtsbmXiyMQ521/GJ7q/HcfOFJyIFRHOpHtPIg8Xo7hrj
9pyk8UQmwD7JyzuiBBNGKxNILecn5YpATYPsq/aw9OlMwyBsCwQ4MK3uOkchk8C3sDx9bRvMkZBA
qaIXP5rzipusAEDzQHuedvvwmqE+iz/fYqFGJKR+1Db0jrfo34FrXJAt3JObm4HB51ZLZu5mG8yP
r5lebel8dMRl6CvaS7M1d6o2zAKedh/1gBiHzQdOl9CpMFpRkRRoBfkph+Ujdo0+NKBlA/pn+oXl
sJPU0heK+CG/xwQcC0Ryperj+DIJSAnwpLTR5EY4SXwd5XXIaACose50E1Aj01BDKjubJnjpaxpu
0ArL4ItmgLfXwXK1xbtVamKMw4/d/MPCzjVSsObPAN1cVXXeU4ye1Yy6I3cCqqZ93QupZ07cVE9x
WHAFjr3jAUT8x/8/E+YTrdrHcKh+CP/aEGX3G+2B4MNNkFDOQyXF+2GRS2r8QI+B3xi67Dut77dK
/yStSgm/tUBhyocbtxIlaNy0GMpSo6um2vkIXNWhb1u6gzVldWLBcFOaX5oaIdJbqRkGmSzm60gO
q2N+aj3TTI7b+qh3hFElUdRGpXVhzPOOeN6Gu7vt1lbQEB25c238QUw2pBsYjSz01xvGI64HF5Hv
G7Ap7CGQIvBy5RgBYoNYPMXbmz2BoJlrMDdQ6gMcQEiyuvChlCUZOhdo6hQ+5JblD9RMgvf0R2Qf
P+rIh/6c6h2LlIUzXc+A5vc34ZuS+URqCf5jyG7oCX3J5WcrQmV14qM/b0RYwp8eeyPsj4hZiJEy
sRU8uk126IaEvTE0Z+0I5SRpKIaY8fOvZf7ufH9xSDY2Z5AuhZZA6HNkKimufRNaZbh1e9xRZwY4
BKv6gE4CdwLUmgDYjnvEQ9/NAkKJrXrgvt6nVfTC9mZ5cKtr7I5ZCUCAlSSYGpnniK0ykw2L2EDy
MQgStux3tAC5+ekg7AxGES7fpcrXh0dCBscsj231TKcbO3ObiFKh/ebB0zHq007/nRIjIQVgbdT5
rDplGMQe/80c6sczA8pNdB+CFV3GiHzZaMvBYvW6InYRJ6lXXYZwvkKQq7HA7wGPitYKOHTPWF06
MeDbncxc3qIwzYRF4dVmZ/pzVa0ksN2mF4n/e8C0sTn5snoo29+L+kwspcOUmGcivzfwUjlixDuB
xmQ2IMd/1G5O4XClKCPNcfQHwdjSMjMOKCa6BRNZkXTbZgr3joEBK2kNlOM9l90cOiOQlx7xNjx/
4fFwBvVIrvdQu86SHg+mvuUU376YI4t7Qr9uxlaUsYxeoIoX4JBzc58S7YkDdVtaKKTPKo7tLAmN
xx1BtKpm/L5bhJaPN7p/PBsYoB/PYzouWEZUbauZco+gh26HmuhX9y5btnP8THXyE+GlgLoEDlEN
ChZwx5KpV7PUABKOphbUxRY7VZxpD4OTEe+S71w7pQXNCPKbXHXtvVoJxG2uQw4X2Bz2iXig3kTI
66mkwsrPYt5vVORZRYeTqRG9FWN0PxswBNL8UqR/wt/5wC8HjP4OwigwQ1O3JGzlHiK74iXYinw+
P0K15iLKPkfmr7R4xxrkoBICAGnaWnX7RLa6kN70gWUtrVP8SlDt7xUqdjU36gxd1TIgIdeu+0gD
vnt+n0Adqo9bOagDKw9te8mzPb+dQdUOuG8cqLJYaDCdC97btYGcGp9Aos5TTQ9+mNcNrrzEp+h9
ZavQ3Vzn4PTmfh/EOGtKFu2TiYHd+ApuxmnRPYc4nNbjd1f2K/zLGTsOpY60sfLu79DohXVPFKxm
j8t4Fg7GHFnMNmVLAfHXLbRJ8aSKm2QByOKumP9hsvLUDkLDDJAiM7ODmeeVx1FZDdzY/qqIZnTr
JQflQ7djtmTsT+BNQgznBOAxUxd+V780DnchdgEgctVojVXb4CukaAicqpy7CYdJZcPcaBt+qWe6
LVHLlhdssGGUktH9BNaDxkNRhYma9wCFEuc085CqC/fi13NRonOxFPrJVip5f5q1lHOaRsI0rMHV
vvjUx8hug5KD85X5DhhXoeSpvD+SR8VY1naMQwACG2vx6VJaWrcyRnCYCp59AeiIPPUeVIOWAlFI
La+AlTAUQE7HZHLSMIjhIaFVPRuzAGv0+VaD4WH7inYu9MAzQddtou0xqxzviVKE6TUWDjfWUnZm
HrXTnXSkwfzMtkkm8e/RFGatj3DKjzo38cI0gqX4u0WgqerBF2aGhPKk0I+pnW74OTbLpf4kWuki
ve8wynDpek7Zz9mn+yW3AeGuHpwk4tj07YVbc21XN6rmMHrF08IOUqldzKbzBfyjIHC+D5awMVK5
7vW/GBQPutGTiRSd/TclQdcn2Mkd3b18M48ZLo+TNaXbCurJ3qqUlII2Gb4xdzfdC/cMUeDv8hWg
Gj90AQEGatFhTasXeIy+TDQh09PS7qXyvj9fhUoUSNukHfxSeq6K5ZHvxdSlrr8GzqPMjBieAyML
UTeCxNzYtTXXCYQSeFrm1iIWjhAPxGDpJ62U4Ku7t3XngtZ811wqKo8HSTGMA5RrsLxxvTkgG0sg
IGUU78jXnHmajXWVUW/jTsTAmHki7drIyE0RymL47MQYDonS3PJvugbVCrMcYMqmLz+zWop5/mBL
AyiJ3DQhAIeshOcOTtkAkm2DbmhUoNAiBJSxG6SNrZWrIvG1Wcff1G6SnwgM0uDES3tpYzPdLBqg
a5KBnpt4gG2OEa0Psk1EFkkkhuMcmw2AB+SkH58/wDlYj9/+ostVqYTe9uCNDo6yJhXL3AUu+YXS
j6u0fe64BSJGhkBIYTMvRCl+/iHhP/cvjuNt44W3rSKZVPqgEkgxezkr5euebwCVJK7N5LZ8gQAv
BN22rcMjilE88M/IviPFe+UnL5veLOuxcNoaRRblFh5supSNFvwSKOnIjWbb9Ol9NVES+oAxg5v0
leRjxoeV7v128R+KNB7yVPssxBLJMTGYXjNeSnRYbQS8QaTffEQBhJIwgIU7iRRWK+TukCSxCk91
Hp3Uf9MauBiz5+kOBpQyfWeDOv5oKig3ltix1J3eiwp9GX1zPvzFMvjoBVSvJsK70ihRr1t/i0Na
OX5d1AbWTQ+It37AcoSFFCUeMpHFxIvnP11DRAwH0NgKKE8YQ1D8xX7NcqtG3EjQu7tdrJMZqF4F
IPOYyfyjMHgQUmNVhh5Wc4rs3bfUBonb0pFzLPrMIgvNxafwZiMJeKr3WK3knvL9BgRYE64VONVB
K9TxkFpigEaKEoj9zsGCQ6vMMJFRzezCvlVxAMu8jbO38Xnp/eMwAFBNnclHgzj8cleo6poKXZt+
WCDf64zOYbxb66cnFrjPfUPBPh5XYrZI5VAF/eySazh6wl2MaQ0XqKLksJqR5hmjNmUNoAZpnCkj
udyEXiWJ82N6igD6s2/vPghAyS01CAZ1AD1ooSWXzmVy6YnbDwKIM3QxFpFV0HUBNtw1xbW1mbrT
v19irq/ssD+HrwqORFDrEW8+Capvq6LpW7enNtoRtivGkZYfbsuDeDIBRDLMa9EUAm84QBSIRZNg
YXQ2SiIfx1YwrcQFG1BEf+j052IbVQxzM8cQm3bmq6jH5W/SDQ03k2xGLT6iB2+3/KuscG7O3301
pYcF2L1uEzEtz9S1/sF8gOaWDg0grJSHxMAx75DDJ/sequKkYdUtK5Z36X5MhUdWGS9bpNnnWZCM
vNVlh6i4gBvj4E7gW3NM7DqITt5PBRbonW4N8v2XSOXJGWFtw0u7efgNZdxTmzG5eWl7WxpgSQ1f
mq61IZJko12J372gpGQ3AfY8TVm2pfjjpr01wVfO4DbRGKP5xCijxIXQ8k5FGBYeEiV4ykrfsd7M
Jr17syyoDrhUn0zg7XJcMjhOJWgjk8QoPsnETlaoC4LOjm8tZnU/s3oTyOSqXYgTiseBeGC42doa
2dE+iK+KMduJOM2KbMDNXxEU3I4QeGNynCktv2p1o6tmDJR6I52tGJPgyatPJlqKp6loS2nfU1ke
AHwXWvWMVnjFYnJD6KCA1ouohGuiMw1OM/OoHogAoOX4M9bzQ5lO6rtYsJNdu3IbnluOta1Vl0/0
0HrnK0hOxEfzHyfrb/0eDzOudh/zVd5U4QVnFMmEb6smwnm2quldtPBwpJZzJelaWziaeoSQY6Xr
Mun+xAnU41TlNCwey4tC0V3a5erPha786G4ISpW7ExhA9owgwgofFcMEI5nEC/hUhE81SPDYbqUL
5fj/INnXF2evl07496jfHwTbjo7U1QarT7J0/MyAM2L+sbE0lhGHCEsIlrGWCKXfY+L/mFU1k6t4
Wi430yWupZNjVK1M5T4LbVHld6jvPddYIpBIIvgJld8CIeUDrtntUncwz5AFLKWxt7Vss5TpRnRE
sazZ+Hc2sXSGGkvHxldtIhDYGkkEnAugJkD9E+kccJPlcZ28yrg6V6QyehA9ZrDkvz1G9MrSaU3V
Oo5D/IEG4w+8oI7bSHMzUiVcAZw9jwNj/7D8XLIOZWVZ9LUK97+Ni+j+0wv5dcpmOs4mZRXazTfk
c9MUbj1zl25sV3yFulkT0m7iYmQ4TVU+77RkPVyQeO+mAhZdsSoRp2XYWJqgFCfcLcdonfa/cpXF
wsvXfunjuEhkmnY4fF180v+x6KWZjg0OhBlTIgxaqfnczmeq36eRku1BjkCKYdo8ut7CX7EP6zPo
mnMVwq1eLA1SbmMZQQEa/UZ/6agzhsx9mYkWm0w4ZVbcnsshhQsvJToqOMCvSul6vyivrp7HogFZ
6MJ02P+WT5EOjFdol23NNLVAl7FHF0ezTjpImz5Tch12uXlKQHehVTRXriDvOfihSvGJQrkx2cDd
9CyMzWMM3Ef2/tZmq0817XyTZ8E2MuS/mL1H4GVYl+2BetZU5NE2T+Dc9kgCbvzyPs+WPsCrVvU8
JRUw5ksPbAYuiBGnxrl2tJWsy/w52MDlEjj3SOx2+TNVbLgcY8gQOUZiklvEqSeH5aKLh/o0xwB0
SCJVduK8h3epXIVsjj9dORxk7PEexHSZEG7uYFLWdIc2T0NTX8K3Vmn395vxVHkyk0tH09C0KzyQ
asXsfR0zsZxE0BNSMEhs6Jd7/o99iPBZstaQL30I8/HtDQhSa1LzXkJKLfRPU3bqlipDJIum1bqQ
hgn69wNJDMDAr/u7PtIDyg4eMXBubTD/Pb6ZNWIEgDma7xvJIs+HknpvkxZpkqjnI10IKGVzM/gR
iX0nfJxdff4OwwxMIM+RtaHy3lTxt9HiRC7wyseizEeBYR39uUgkWhV49H0Vx2E2zXPTdF49DENI
aOZLc/IxaJSLM97Vnym2Y2cR1ofy4sPlL89CWpHys9tmqzjhqxvXOKLH+3CQAWuwE5L7q80QQBUS
8Bi9UAOS2FNwaBv3tQDqKuI9m2mhHuHa6e834j12tbA1OSyPxfGVYVUEDIDVDYLVAORBwfeBpmOL
giCiMhcm7+E+2RVezvVg/Q7tyGLRwAg5n3nupnb9iZBJcVPLVmiPOJ0EV8DJ0FeUWJNb+ss35P07
jaZyuYr7a1lXXy1QJaX/xwnA5COu/UVh+G0hvc3V3a+dRXLPjK1xwpFJHC8u/On/Cn8ZimKa+oLu
R4akDw4beeJg7UoCBV6VzTyoPdGTW5fD/n04R2HjWAbh7mlkj44VVRk5pmHHXZ0bAHkT2FbObCok
tps13TaCw6DHmER3PHn+ffw9r4DTiiyQt7+q/UAF0StUfLWWEif/ZE0JDaPdWxcuKoPjxX3DalU6
XI2Yn30gKgAyZq9KZshkXBAQo7+L6aURM7KwcxnBAKfjIF6Id5fOvI9/ViTTXBQtkrN3jO1AKSy6
+aDi+2qaUumz2P05zTv5nRkvcQ8pqt7sO/8MDd2TIQaYyPXuDNVFPt4l6iekrpGc2eqrVBIWshkq
z49Vdu1jNRTK4XZaT2It9pthwZy3BcQ8z8jt+jdBkv0AaVJ9QOgNX8MV7JNN/XoWGlJR2EJplzqf
i1VQX0UWLxEJFpEJ16XHfjRw2YHSpesofrjJLnbsI0m8LLLx2HBNanFd2uPe7mEkgjKIqkyyjqMM
O3O7+p0Mq5Fbj4e93N1b0Wljv5kOSDg6qT4t5ZtiEQrJL0fX5UD6HjhmWSuKNJKEOlVkzuiJswKS
nQTwryhObdIoc7I9tHE2rKLl0z07vCBk9GQWQY9UCNR7RJpKIy61dTXoA0CPlfkiNZv1NsuglHMx
jG/OtMU0spgZvzGXxJgDdiRLL4y1mkISgkxSob0i2KnOFJ9ZBg44PDyvPRT3ufLJICWrNfcQLYxZ
azdOnb5+7x+TQj6QHu39dvpI2IYjRW5Bk0NO5iIy/GpFFN3bVvFAOKQTmyYzs5CoeUnDlHzcTKZ7
KAt4Hhqt380PmJuTmlUwhhS9L5ywZsa3pqTq84zuX1dLVapMtaf4Pz4ajoVkjzWQ52qaB9Lw5VbH
3yXJCy6v2K58ueLqD1c7uTmmYmsn88tPzGp1Nxls1ThxLtENnEptsichvbpAyAGve0Hq3dnXghFP
4gZ+bKbMM+A/bGG1oyoOfgh6+fP86wW0aXetyU/CZgRstbs6qw8k14Mc71BwBLKqLNy04BrO16Pr
ctOPb6YCX0fvJRpbuXsR1/oOSdbu+vFsNdGr6J95Qf5q6tdLq9z0Co1cUYGtbyculvqWJYBSCjmk
FZoAsp0SUe03FWYMF9tzbaI4/R2JlWAjtJEVgSB1FPjbItMBs1lQ1yQGf3et5VXpJH2+sT6mDkyd
nSA9oqEHhIE50+5nipoJIho7c/xfbWuydw9kzBaPNnktO9d85crIx92S+OwWn4kyBTooDihK17Bx
ch5R1hOvTe5Iu6Cn7ebOQt3YanosOSnu3sOe/gbbHw+QCeVkuiKD2oc7QAabTgl4swQkMjvcYadx
GY62kTleLSjMoOxc3eQj6HoDJr/fu9sBKpUUJGnhZ6iG4d97sAPxC7cUhyCXGDF9s9z/KveG08Vk
eSAqY54crjmwsWT3U+Luy6oCiksqziOiIHLxbuwBoIF0jQJGaGNNeQjsTGufGpGsFI8egdt/pzmf
5xDmxj1wwWCnsAaDaNsuAnMtduSo8kFqHpY3C81FAJYZWx5poOhi2+vDlIqzVYoz7t739doLA8bA
2iYmYF0y8ZvXX3E7DHItSbKCf+E4hDCcI2Wy2evCSbG2u290jvoRVPs1tSBzlKQBr7YjqqpLYsGT
G08kBCXN94LDBER9QOcLH9gY+v1VSXkW0XTvAYZDPfi9gUGqyb3Y6qN9hJKwTgrwDxGAMkEBeFC5
xFO+eGg2SiV+jOtse/MoKlCVuaFwwcokFolo4xdAaHFrrLirKHnNJIaf70Apj/1MvR78kKBuU3B5
cdADcX8f+z86aySZPfTiJekImP11Dqx5IchA862Ndl8ogGU40h/cLS0jt4ym0ri0WmgJIbW6UnBw
TTFBmLUSeYoScMuzJZvWO9wW1nXQBu5o8gSuIHM+YYTD6gHnG+X77jDj6CObfLwyLUrGPlVsWije
tt9JlRBzsl7H21adsSJG1wSpg4IEc8adIhN7VlAb36BD72j5TXRpHLi+oxJUHdNXFCsFuV3tgvmB
vdovC6yaoysuy3KTpRJ+XN2Bd/hKUX6mOnFk+ULnaa9hJDGrLyG+vCis10RvkCn7/awLD7esl7g+
OyEUB9h07tiOfyIZOu15dB6CxPDoDbB1pSRt6FcdCWxx3yU7LX/IH93DoxIiwFp2t3AW0iD+uBAe
pVkFV9C92hevwW6Sjh4/6HkZjA3UHUpIeIHdmgkvODhf9OMhhKY5Ju3GOK4NZvW5eIS2pVrlnQiP
GR3mCIj3hvYT0RLw5loeA1mTiTqepDqYpKw8LVXPjxOuxWCmJnBkHPToEuLn++OPhiAWgWc7ykNZ
W7NOxjFAjM3vxZqLTHxlrjA3cBJKxie3K7jgsJZf5dL1brvrsOdit6bHJmD29IctfVcxKRhWy5Yh
oQTpYpxQFsr1HwdgwE9bLL23XZZBoaYGK5HQ8tEuryr1BDB4JEgy5Rq0OeDAAcvPQsIRYRkHG8Ss
GwHXQzgNjw1cQSvvFfBVYCxlPvaqNl+hl8k5rONw6u6BoC8Zj1UVrUkjfXKKBvkS1oyyHZiOKBAh
PMs9q+UTIy3COCn4LShuw9TtjTpOxN8Ec/Vre/cvZcH5Kg5FgzJKRDqKVd3iH8rOJBl+Ba13E7W1
eh6yGsI+hNA402LmlIZhrnvYeop1WJDCckJULmREq0UND/Rlb2PByKFouiaXv96nog8Oelm2iR7R
0zAbIosEW7gm7ku+5qmmyX58zIVdPBKl7Z5Vnqw4xvy0ATG/SEeveizyyAyardHV42q1fqnhD6JP
xaXtqFK+wA+fUbb9DyDzkQhly1PAgP172x1N5QT55TTF59NT6ojIx0K55+XoiynA69doV1SedW9Q
VqPCVQDOUCUFYs2qfKl5eAXn9Bsu+C26yHDZQuVWCUSsodjBBZTh0DiVCqC5Gfmsr7g90vV31Ide
n7IM0A1zyVJ6Iywq4STKk9N9RhABfSJtm2LGoayNfoB+RpYrDeOMWNJnrAUMZ3S2wcC3sXLLp9AD
+0s8SfVK+3GOR6Vobm/tYh/OWqtcpRWNnBiXPSJzeyKTOoGnSsJs6YiXkdzgnj8Bm69MxeTOoNj/
xtsEDd28Av5agx5g6wKEs3wxP+EGyKUeiiA2JiA6cqfWNKFBOUIe/rblN1XPaLJnHed53EcUhTaS
PGVgc7QvI/lMPdElD3/r0pVqHviFLwwyJZvJ2E7TZ4TVYy5Wh3LdRCVBWubzEJXZTfqp+np43lfL
GXPbG4h2qd5ZZDUOO7d+2fTDHb/Bya0UO3QTQtbqzgKBMopiaKVq83kqUZDKkTwIUfiuG4K1Bn07
xYEDLjqA5/qsMhrH19vicUutQic7wC00UyeU7IkTwGv+Okv86eahyOKNazRYl3mYIZG7EnKt3k0a
/373sJkY/oZrlGCvqAYp2c42iBFro3OrQC651de/GAuHUG1eNntMT3X41MFk0QZFjdXze29pS2+i
2ZwE6EYDkdM6oU3/AboEXKaEzxfVT7sD7fWAKJb84t1u90g7HGZMOvE0xU/SuKIvNllO4ZjOlpyF
JOR2jsJTFD+Dt50rlg3byVEG/kMxC1BliQ9k8ihOJfsMHNsp6JqtK+vduI9Ifs9gJ6tqRkE/QBFr
PGofmIMt6k6yPISLG2HnMFHw6AYV7tt+IvuvZNi42eYZraPCG80vzy/H60CPxEACWGwtnRJjKmBD
L0VYmZWo49uZJ6lA6Af9HhDAb1//wUNm26k4x0JTgAwZ+KPELDLi6V/fUtzwJAIO4cg8tHc3mQpo
YsfEDEG62U+G3+575xLgvsBY0DE0XPVfP9hl1HdzMZBKM+9AdtFREp/huxqaautLDcO6oWegP0P8
UfZ9R7knY5XHt58EaolrM6rvSGj0N1Iqvq7R9MwDvUDWQL80zagtUtEYBrytqbfkoXZgUclYTu20
YEaGwtv3l4yNfG8bmfWmAHUtFP45mmmv1FOP69NYvl4=
`protect end_protected
