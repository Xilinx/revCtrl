`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45792)
`protect data_block
hTX64IeLyHzfa3tJyS5Dfs45/kVXz4SgZWvyCoI+GaBt/ajB1uarMzYwraP4bzTsEtY9azSypdEp
uMJyMTXqOnV1lJafqt+04VMWhtgOPNjvYx0tpIk7nW7G4hpM4kLNrnENZhsHqae9vQHdDyy7d5gR
+3OS1PcyGSJl+zkymRX3rUzUpMqV3ps+9lol26l66kI7nb0CSe8anWmsAesfWebQoIF59BTfAr9C
xnyzucg+GMIkOss4CgWrkf5MWBeb+eFYYi6o3GAIwx0ovIPwmNPqxveLzHqfFUrdOUHzbTqlYWIG
q8Kt2X/t45pJacYo4KvYqbDfGc3+sn3ne3JDby17iRxnxX1dHoz/+hO9YZEFHXpSfdIxlLVnVROA
38+hBmzFlGfFmdokAICOkPej6Oxda0UrgVwrc/QkL7E81VKXRlpDHwJUR8cuc629fNoJoN9y2xVz
3e/uxq12ZZAetVXUhw+Gy3iQiOQkAkwnuuTlsyB1qUMEglo5fc4cdRFvvJTMZuDIHp9kv6SxrYBd
ew2FOZxumtC5Y/FwXWiaLmByNRDoWvtwrhukL7FN0a1MYo2hx+PxAL3gI/y3/ndB/yIbteBr2sZH
dbuzXDde4Kcyi8LkEs4ldCGH9FvV/gDKTQkFqUhYKGGlug7BJWxNKyST7b6SZbAh6DRchnhJFfln
CGjrI7pX52bXTqw8rLCWhY0/V1kWCdgIkQxF+v1sIY9Von//YgfIvKMIzXJk7eS76LwEcKv0H+Fy
R29LG5Asm3lns037N/Ux5XxshJczgiebdgWKzxEDOmfHlN/yZnK4f1i6RIYbHEAHLW22SbsH81/0
y51SSnzIpefeWoiWtayg0Evd8S8zh8xTXXRdAYSfUlCSOHFWzvhWkQEPkH5rGQ+iQafAgpUfMtaQ
w7xDB7Pe63b33yLKhQvkV4hukrukp8dFFOaPeT0r4tKcQia9BkJDu7PPDArXlHgCJNG+F2vm27Xd
sBsNJ9ansd8Un1wZ5WqveTlZT18UlG/It48BPiihND+FIUqRyfzTthvelgjsxvOYJAJjOJDRnAf+
18MZ6PgSQEwV3lo04dY2U9pKYnwSQ3FsTHf3rtSwzZtIrx0BAs8+iW0O68i0Mu2plGvDIQ22pn1q
PQPTU7i9SenukvjfuLXOcl+fR3y+H3AkIdjcrHbqijO5HZJBFySlsSze4U1Knxs8wU19O5a4Tdde
He7Aer0QnNoSO3s6lf09MZ6xAbiH+ScvohpXF6gaZSq+dLEEqQjnOC9fR1iQBb6a6nv4G9lXOuac
zSm0UNhv1CdFmUavGT45wZLl/rrZfNTDG9oUpqTDLryUgadJ5Y6X4hJCgKuYFZtG/m5RA/cFGjlq
l35eWyS0lCO/aVA5w9ruScPGyz6ievJbY2a8uLFcJlAp1GUgp8DP3nUUPSwcDyy6bli8oJpHpPFw
nW8KuQIz/9MsUpODO8Jhi+4uZ5WyiTdGrASPpumAcRTs8O1WDd4n15jut54otjIuDFxGE7eNYKVS
qtw2bmBm3awXp9JLtsNbIhpNXwbBx3tEo4kDVzEYM7P2QYrUaevJ4ZlzrAaXbbq6smyngzm6zkiM
yh7UYYJZRsX0+jI56hj9GJMKtUWW2uMCyWowNvD9xqy+BoiuO1rBEdcVrVcboMr5EtFrP/hNOtlX
X98SH9xvQCLh9VYamBw0a698xkw7MkWMSGwYz1Imzozklnokh3neFLxtABgmcQJc/vajNmhSDa5u
gCgIZdLisPrm7LUwBNimv1KsN6GWil0/PTQTQ7QP2ZA0/bGMFqHS3/LLV8XOqiEIS/BNdoHQdaJ7
79AFlsJ6+sPfWz5Kzu4FStqSyxxTPYfUv/2pOn3Ggs3Li8m0Mwg+8jhaMrbhXwkQkuVj0LXMRniW
q6rpgIFrvQOTYGQvxPSOZkl6bv0fdPA7em4ZPRvNpZ1hVFu7zIha4LS0doYaeVD3HA8z4vl9093W
xGaA4p6Ldlh6TFbfqz8Dsv80dYbbUREU/7Wve7INYasR7uRJn/ebpTYiQu3gv/yygv81S7NijEPX
BEZfK/jL7oeivtDkogvE4T+BkoSEaQSy5HDjrrxmzQqhMhngdfKlzSpYE+L1zb7NsUZlCjDDK1YZ
dQEnMZNioURyMFnJ0hLQ5STaOFNroxuyaVFh8L3CFcj2Fl/sM0Ufb4lrMHbBINu06n+3hqT+yofO
OhdRwD2Ws2SDoXOjXebBmlVHX7ly2FId1RAJLpY+SYqR0SHJDkBV4HWFEKL5kFfxnAWGNcmgZhDk
K1/mVoQT18uAyyA1ISZGatxnwIjoJ+QKDLqZZHbqH44nc7/Ta+vfChNY23EinPaiBJGlgDNiIdXp
rnCS90IHyiz1qIBjfegYSlq4TB1aou4zv8CngKBrmFwHRTOEk1bixwm1P+GdbCtHDoHlyn1BVSe+
/YxsulQBKG7qJp6Iq1Q4N0IcASRGUQ4mGFZCTO1256OGFMmzlx0wvaGgH3sufpNxo5TyrB5tdpKQ
Lfd08wKQTVZzX5iko5p7NaAL6u6dEMDUjzgkGmxivWl9TMx9e2HTsx0B/2TCWaqIpsUrIIE/+txP
F051TjMgM2gtDdMdBgFoTlzeX4YZWb3LEAuzoudyokxcc03pVWRIMwrrx6hKw7Dutxop0SYUnK4t
IIvUU1ppnXvzXobPu+aJ5+BoBbL7hMBteEaQiR/qsVJfSx3qsiHAPQXuAlRhd1pXEAFS83qhD0y+
I/NOorWHfhPhBWxW8By90q0f62MaGegGk3ab+4IkQncw+pBzzQaVyeuQPEX8oIsD4EEuWBdYnOQt
unHPjfOO08JEUnP1/8VK2Y7aUfG5nqDussLtGVH8JGpt6YLLNZ6eXTK10gos3NT+wWNMBdnI1/Yz
j+mmhuSE/Yswdftb8tvQAg9vcI/HZXxr+rb5XxCwL24dEDGnSJyaVLmNw7mO5pGPKzBX4N2IUJx4
9LX2DFLAVEI4lFPR/6x8IPMqnmBRlMQ4czJfW++Yn5E0LG83Kh1hMdJsXBV2VuBnpYbCrmLfo4YO
Gpcm4UXyQcV+mUUpNNsLN6WH97WYNz7XF/yKqqkEV6c/5i3ZGPP0I819XtifYEltlf3mqCJecu90
pyT0xmTj7NRROuTHIdhVoz38UPG6w9QfTNNqU0w+D/EBhnJzMQKnmGMvSh9S588FALYGhvAG5nDE
CNfghZBaps216m393OwS4Gruk4AVxQMKVKCsmJFSXEPyS6VpJt5muQFy1cHqsyzKIJHAEm4wKqd6
rBPMgPHwQ0w4jqi3IWW56QVS/ZQ26D8ZxpTKsw4Y2K42CkI1tAiYco6JjVU0JnjE5W6Y4vKdWV2f
2o0H48Ny3uxMnMmvH99xKj7p74VzK7uW+u5abvi6+x18J0HLM+200O6uJMAfcbxmatxY2q57/bdb
++QFehU6p32rTxNsgk//WRHpZNAAdWGwU+gLLxoZt07/otQ3hpn0CBOC15Lmxj+8LLYWYsXaEBru
37HOzT7W/5CLpqcFet9H9GMRKYulaw5QU+O/JeoVKLZvhUzuCIHMyq+FjYcOxHj8lctqkSb1bZrW
/BjsVtWhY1+aW4NCybgpok6L1OUjBFBjcohtYgVVn9bb76Gj9hmZ19iP17n/ltwPU99o71hmIg5a
8AcpbiPD0L7nIARJ307JWP3eGwJ8V1QHUBWyXp489Ud2JQoIJ3/EgF5gXvNWNtwPd/k3+RKOWWkF
vMSKdzeU7eqQC5Bx1P+F66y/oeINzFQFcTZG0+0hyNm7lKOo2h36VOI8E+vGp9m3XblAz3dVRA2r
rfKcKqbiTQ060CFXhwWoaWdzbo0juF6sjaLBkaywz/r3aeqM1zMZ/dG48+jZhtCp/ZAD+eu7iV/o
yhEGXdYGzIZp84GxHnaQ8PMwivOGpvbFbLJs/Gik4anS9jYF7NPYaiN52Pc+GZmxwwT4LnuddsUM
/up5t4iXh90YeJjf9oh4xNeS2ulLFSXKmgnAxe+hdfguIC3hGHkZ1OEDqGj1ox3QpZvK+oI5QozL
e33EyWhnqvBflxLGjbZVvQM6R8kE26kEtWiiK40NDfhEvGFY+OPvksWkDFHPSxMTmgXZoJXdy6/k
3pZ31Vq1EWML7rFGnsoSu13lEhXjW7Se6vfOCMVAxiYmiYqX+O5QgyzKHYU27MrWpKs4D556++Mn
zQ2X9NzstZ6cj/nngqQdbDz6G14vdULYCK0fVcmpfOuswNIIORsOa/KctpCt4WU1gh5vLVgta8dJ
rOZMsLqtxMhY+EfPRsFREJmRA9y7bIOrao5mz5bk+WeterIlElfi7xkeXD8TmoJE6bBG1D+w563B
ApNOllUDQyMd46VsvyxflOKAFVSrVQW43qcCL4DpHcHiZCCQno30lMaiD7wtJyLlpgZH1ulimCZg
7IL81kFNaBfb1fJs0X3/6fA0c39BAE2PjbLTdtnbTynDgLAlqVxmCwASvoArtetelUJaplngRwmM
uNZJ+ix0jKfPk/D6ceBls2XaNzcQy8G/W+Peja0HfeaKOCbxEPJ3O1vlUt9+7oM0xpETPVcEh4Sp
raPf3lwY98GaS3VSyRnObOhsetxlBF/5qi5sH7s3TIyH+Raa8FMzIruLrV65vHfodlExXkzDUhVo
2hW2mjWqBTlF0CsyFknmbxJHGpK7gtyrTxLZc3bDp3xRgXn5/upk1P902nftAxuNxxuBBJWTyNru
0wRPdD+DG4pbSCLHxN9+4HQsa0JKYKUQQpmqEr1Br3HjQVlhU6VvchLWpDjny62iXF+L3hNBJAFu
YJoUlWe3Hf5BhsTTsteoMzTd2Wjk4nMganbXc1hU9AaftlqJB4U5Z48wZQ9SJj2uZwlNhiV1OETS
ArE3Hfrj3ROewP024mmkYhgqSuhq1Umg8vhB+YN74vt6Q16xMwiy+/RpV9i4X31QhzPpU+2PBhDw
cTmFH0ZDTsm9aTlb5qf1jGlhkRLbu+fl7Ba78/8KCvbR5HGviJ1QmWx6RjD5D1N8pUSWzRhDLdeX
ScInQ/wRdwRYuv5N5iHUkiYExhxrfj1J5nOUlQ5TRqOhF4dr7TamLtCnxgAfIzFQjd3Edm1r+d3T
dLXxPEzjfMrfXeTGyEjd8LECj4h+9Gaf1PKqpJzYzp28tG8UWonoxhdfEDuYLhngHE/GKRTVLDWF
0BDue3zuGTGHSRtnr8srppDRsX0j/Ahzkvblq9Kp9WwwDpbhUIHObBl3ADPGc01tw2QZJGAoNSPC
gb6kCn4MOsBuYrl+XWqVuFp+w8X2lfgW6KcOM+bgRI26lspgUGhYXt2gJxn3NmLCMNgEEBwE3GI4
sKiugXVoh1nG7arsfONozcSs6z0RkZnAQ3mGQ2Q2n084heXOxoJopp3dX1xCbNdW/ZZwd1xneTw8
i/nT2+f5Ss81jAfudBZ2wsU0hwX32f8ZG3NHBaRa8+YEZTTdgoTPd/RbU8xA5lO9QLjXnbKi4X22
dcbeuvna/yMpbrg40mMRssJLET5H0Io6084Is2SdK2DV7arxR8qniWiWPYgS8/eIlh3tUAJkepgK
KJQP9B2ym6y1ddHjX+n0DP/yCly1jR6+/kpEgajWkmmfm+t3XQneXfqq1F402A5mNiM0Cj45YB31
PtJ68G+vZvLhGKRNm3YRx1AQZ1PJvhItifBWW2yk81ktSav9ILJyyc9rW9MVgcZbu/Hj2JoO1t19
rzjVHZvF/jLMppXp3WWrtmG4ZhqeCgGAlEOcSYLCFBtM6u85YQvo5CmyJuDHWyfhZmJdFWrbAvGR
RHAttO1Ap4HK1u6+xWvmq6jfk7Gu1Jqk2d+Serrn5X2AGxpri+iWTSX6LRtqYIQ/DhvcW0y996ED
TtfLwwr+te4Dr2ljvFONn5Z9HYq5Zf/ngBOu5ndlM9GDCs08ttuDCJLf954+bBI9Ag+YY/5PO9Di
0MrlSgvrXLpsIcGqTQD1G852PGGkWc9zARWbJfa2noQDs8Z1HhMEGv69HMs6F5ZBJr1/qFPsO5bf
DSuLXMoTnGBZq1xg0DzZgaHqAqMi40RXh/SVLZl8fIFhdHPl9U5BaAD0w8r8khOxszldSers0S+h
IBQ5othdpXicg2/njNxzpSwpLyDGLhhuCsFr5xiSCwaMbmTPDshSNR1dqy5GyFE55zE9KIlOy3MT
z6NvvP5WUOIjSJomSoK6jgIO9JLiJwtYSZRyJN97cKj7sJ7d4J/HGWDfua+9sC/SKkDV8amj1IZI
fSq8fZbGn2jnYmCOwSA8v278TPhbdQUN/A5WhDpU0e1MqRp9SSuOvZqgYOSTeHSlR0NmK+ysHozd
5vnQETFqmQgk6PFTP71KLDu/bbZYnGwEaJ6ig4FCFHQmhaaoutx3gcaXpxSk2LuWIaBrkioXG/SL
dEC9Q1KX/vcPmPmE6cWMzes3fE9ZzVtdhtcsLkLyXNqp6n4AT2E1M6+8YRkpf28xZez2nIVeLzda
1RRTiXFdp8avZzKNqZgzXJk3ZVi3qOepTKcbryVLI7nz2eRzX4rl0ZtrDISgTBxBT7aPV2RToftN
GVaxBwRuBrpukUjN7pRXSmDuloZ0NyL7cZkB6FYE8gO/yXvfM0qEin/qLW4XzYl/a7qtoul8db+k
m9Zt1f1vhLjKMEaYFRRkcOXtDx1cjIhi1GenqSg5wZXRvqLMLnNIlGpIdquJ702j/IwrBtzaNm6k
+bErsKmNov2pXWIMZJgDBcNVi7lHkc1j2kvVqdLt4nFHnN4nmeIE5AA6X/ZZgKNWyW0hF8u6CQ89
oFe5iZ75Bt1Ibwk4r50Rlb115F0iW64oGJ6L0U1adhon5eqtgrk7DOkIORS6U5QFXiIJvgXkrcck
lgIBd5ybKnyZWQofgJ0htpmxmFD3pIK9jmeRm0/mqhZc2mqINdXrkCcZsAB/EP8EqlioX7GveMG5
HuXAxVffgc8zkEnBUotJp8oIgmbNqsdZNtb47qKCW+VUx3Qw7oEMxKwFGlddlrTHvpiq8KaZPvTC
FXNWKq0rMQ1slBJAL6TOdhEAXbo0KIcJMtUJ2LYpn9Nzus1YeSEPJ8Z3Br4pEnsbCucQJR1BqQcH
of+teuN+Z7HhOd/IkRdFQoh10a4+VVJaSRaoFVHKupE40sIBwZ5E7wXNJTa6YYMvz6wgK7AeoOOh
ve4D0nyQDZVqvDB/2WeHQjzIpnjqXNYHa03He0GlDng2JRJjgy+4DKAcyzVVh49y5KupG9kVUX7R
oTSn3GPAVwTZc3ruvrleIBh3kpYJ860Ibo3y3dQKnPi2Bafzq+RZJV+l/+I6Mbm7gJBZrYhyGq89
oEm7WVcqjH9GnLcaQ+8ByqnX4ZwJLKyErr/E1QKaYkxDXOjdAr7+B8bhOEE/6axxpbVZ3rV/RBjZ
T0reyGBTLKpqkKqd9xaISWfmV9eZJP4eHB3fQAPsAVBoo6UvYwjjtkE7Y5sZAt+n3EDwOH+xQPMs
OpQum232zy7dYCvvRpGI4SaP6KbAQuMGGO28QJ7FSx0OxwdGSIfkJTC5L2nFv2Caze6bLV7naY0f
UF02n8LIbt/8xX7oe8pdpsdgNzLqpJlNNq+JwmqIAaze1yewEoW6aXNDeuBLZ7Dy3TP6zs2XWflL
TfJON5VHN0ENE8ZFfCHEuv+hVsO2bmH48m4aHCoRiQFSElnYrkL2igypNRabfb4WQPjfqDTZGtbS
oXozahzLRy+JwSSZ0B/6HcaFceb7gziczhKs64tvhhOskMLg++ebyTm7y76h1/VHFyho9fCBUWeA
8ecggT/W84lNmrMI/TbLs3ETDp+uGgJZSmhHsUDOyErwgQCcKdF2r0TEyi6Cnv4BIjWuIED7PqUZ
A5ehCLZ0eWIsuSu7zbZTOtqsHjBFE4h2FuCyr0DBdytfyDmpBFA4aSlB9yietI2aJF2spowh6vPK
Gvl2+3P7JNorPpmNqeP+YP0ACclzY8sHOxJstGbqrHwdplto+GIMcss55VISjTZzGCWgQt2x4W4t
VMGr5uO9oEmqE51bYGCN9Q76pL37tbNsXvaT/y9EkgAE2t03b/zxVG+NUtiyvmQa7uiPO8UrP+fv
yWVPme23GAv1MaxjPTlGgUGS6b6VWJYgPcUZCabZ7lKQylMY/RuRYgwObgJ9w+vpmpvbTiTYTf95
AZsC6WxsRgGeta0vOMKFhsq7IM+ypXbwmTevGxqKFzMf/ZJFhvwtA7PmhVBMtaZ+uAsZKxrcozZT
gha4TARPHaam2R6nkpneX/WOSvZ6YFxQZQxgstzbun9a0v/WJyJTn/unX/0odFu0Fn39tW4JQZPL
OF4N3/uzAGiWqf3ZVJG3JVbMZtG84wSmDh5neaEHSAEc8a88KZZsdau05Rn7KTFMqDeah89a7ReL
raEPtXyHLew4YNoCPnGAgJHVCC1zrMazn0g6r+GYJNubKr4sokSSAkcnqJHnBikNg82gGfX3eiYM
PO5qfNXCNq7gt4Kt4vVhb0oIiAvv2rqPBh1Hz4Vd//MuUdLNJ+hoDub7vcB+SU36ydO2EzRximwM
OF3sXuQhNRsSmQoe4KSwL9H9MCw/Q5I1c2FpJ6ZvWEFbNPFXkzP9SoBpi9MRoXSxz/m6xvN3/f1s
f/LkDZjCx1ShFoNh1Tn37R8sRwCnc0XrWGM/P+1KcKJ5qVA8ZZn5vJQa1Hgww4+pPZiEpftMBupR
QG8GqX0l5XJW/JDxm9Mpl1zJSyCkLMZG5Hg85TRky+Ti1vS0dci3mZVd/OJvg/zG9Z+fcO+rcAkA
Tjjc2GHc3z0Rz638H4rb8UnAK/lu/OR2QwqsAyl/kynSpeoxJYuBpwYHhIevF2jZiZMWZuHYYYq+
HlQaEYJvKPT2IohMaOaBlbEyJFEKjkmRNd8gaa4sWXRudM3TBvsXaseenio5VK7RTejeQM5SNLx/
f3a2WRKtHwujiihW3hu1sJdjrAUNH21myzPYFlgz6XJKU4ZvQaLq8TaW6eFc8krN2Mut0xOea2qk
KFNqHyPrr3ASsqVCXpwIbZEYqUGxwgQNjaLfutw1CxqRNwiUFEJlOZ0luTWwvnVQoBix8bLjP424
zMAjD7mMCrGjVh13Y7NilUaf0+p/Z0kw2FDlYtLLbnujQazUKYBhciQyYnceNGHm3nJwTjRPJz7q
SnG3TdnokcKv3FYSAO3H4vdRmJOwocC++3DABJlO2lOzPCM+sLQU6AFAwUdRLfH6CQ9k8aE5a4+Q
BtC+bOV8k+XdtOncgrsMD8bUw6emvvWJtwB+KXkfDc63H3wkMR/MEKRAaUYMATvTjZlssifmHKNp
jfSD/3XkKmjFjV+8QqakWA10kUZc+R0rveBcenXGdelL1KB0doUXQFdW3/sZlaMW63r2K/K+El3i
uHf7hpNhdcekRTZYsMjBQjY/sBnqxZZGUU2jXOF7AiNBayNBJIKkCXdfIF7xvUiyPE+PvNb+JYoP
fWKDFMXnEggj+pknRK+APNca0J8UMBWtQYPwj9yTdOd83DGYe+3g15H/zD4hkz3DjKHfKQ1s8aCe
51yk/cE8hiOwUCTloL+iY9aBWeo4efgf60Gy+m42bveSOEG03lqJiwHcpD0sZbkpo2MtuCO9fH1M
ysxHwFYZNJHRbT0/YRWgXMiq8WcGjzbh4UQizJSKnqy4A2r5J2rEHodmjdcdLagzhWweo6zYYx6v
unVCysWL5Fqup3ySuth1HTXpOGQgsxONsbZn6Nm0RYUM43zON36zn9sS55oOtRtQfNiU3jz6tPYn
PWqxt12s+Z1rJYtMj+jNVC/3veSVp5hvWXugiWYjanUTNXsb4Ma/6Own67AS/9kNI7IdDwDJKMSO
GkPCIq11pDXswa3nOJkigFG7GIv/qviEOpgXK1PqNN/SD2CW+bdK/bQw0oDZWI/fLuWhWFSXX3Oa
ff4v+pg7SJp+l/7QqFdHUPaOkOnAcyjB8xWxQ2lAVbhgNGeyaxOSukTX8XnflR8H67Hy3lzF1hyr
FzW8Fd8CCHiyDASZpJDjrJdFwNqEGqF/6Ze7cL5Bd5AlrHO3uJudQ5JiZbCtbwRyzOrMp/zzu8F6
csy/8AlcLxebwAIsZp2i+FhqlEJLIA97GZ229fg/sZTRjH0Dx5J6xZfUIlbBCB9mSZc2Kz5JM+d6
4AcLlU34hvQYrzJ9NMAsOvli7o4bOE0z2Ra3U/Hy+WsuPfmNJc6+fr8Fjg8MCBcNdrBQMn3ddiR3
xIfWSfqM0rpp75gMZ66q/QOD+DZDExD8RHPHTq2ftIpu32cG2k9GbOmWL2H52vPSovaWNGr0lB+N
m+vOS6CTapszJNcwns5g4/NXMgck2iNhSdUuFzLOgmk6stWKizyL5wgOElRB3yTLH3QxADDoPbLk
UOlM9+JX0zx5+9Uo4iQkKPwBcHXw2c39ZD5teW0B3oGTWX/IDexzVf8Hjgb03U4eJ+yiQuvLEojC
FbhyYlgB5UQueZinUyjSv/XDdvQc7P2UKDumEysZs0UZb/zZBr+qo2KN+S9AjOqwVR2VVmB0W1bm
bCFcLC1nEbbRVoRaKYYz9iTkah9mU8AAixjWMQ3fWlYrEOxX7oDiPuFC7n1emVkrs0sseIjl3yzO
igeDbNms7dkCZ0gYikk3NtJmFNWBFW+WM/wnKyPdXj2Xm6I2J6bRww8pi2578qj4MZAM4o0gPr9r
IEjj1IIo0KyM1s8+ETmuuj64FWOpLthyTKuyeBGfTuWbpN8cMCnQpHvlaFly4023FzdKdkfiwg0l
h9mjAqAmgbYh/csPjyCTcYQnRJeUzzIPtogMh/o1/datVAkflRql5cwAhy/yW6bGuT+n2zM/z5R7
ZtgLfDoUklR4a21DEc+FY0gC649a9rVuQBAeZs8iybbAgyR6y807MnvKQeYXfrf+dZ9FvXAPrOMP
zFONr2jHecn5QWsUysrAN1tW63KtGMOTwbjJBORWQYVvg5qjFzFzCkGvYUbmqlbavUetd+nRIAv5
JlcvhCW7Oy3NuN0Gu8cqHblcBCn8u7wwgCH4oBqtNy1YOfkhDGljBq8G3nPqx5vI/yCnAgwzKC3g
a6zTTtUnaRRxkESJlD4LwZfj9GI0RAXz3g+MMfTBjxxjQIToBtKshfvxACUWvEaZzRcIAZ4lz6Az
5vpWXcK7N8N5OpztHMEt4FmDkIfpTbwd1vE8XAfP2W+Wg9MacNXVRQg+L+E9xdBNFgDN7W3R8Da2
sScc+YQrtkcPqjSazFEk85A7zDAYfzxuSknv6NS029TKogVycwlQEibODQCgi+JP0iRTmfFK3F1e
rXJb/RfZ/bx08IzHyxAEMXGrQTIGWa8KU4+7bE5z6238UsvAmrGbmKDOveAWF68WFOd+ohW28gJ1
VF6QFpE11MAYtrpNyDpL+gVXBE63nAZlHov7OXoCfmpbRStYq2T+dZY4MVj6GNSdy+5KwRceJ10q
TJGJ4UnVlfHeb3kwtInx//fdN9DfqbFTq1nZmu6+Q2ASJhHxAkynaKH8vGTEWGV+3APz95utSJhY
WUEu53rEkkXwtRe91O57zfEzysrtMEN/8acVb5PuIdvUsk8ptLoQUzhKxlgtULXeX5wNVe/ZW3JX
cVUjfKGyTBr0B3Galqk39DV/Ujf9q/wjIkdMcJdAYW9VjrBBQiCerXppxI/u8yVD23LJpJUs5bJy
GLiuFnBXDwl+OvqLe6N40IMgnEQGRz1wOPV1gDpmBsccj2UColSTvr2BZ7c5jmOW1rfY3pLIiDZD
Rxa+W7uVEt91GzO1U++WAZS8sbI56bnNWLm8dwTqIbj3hS+eSdCeXT+ax9EGF+3OeKjGsyVGR5LC
Cti6gknZAe831tVtrX0atHaKuBtKGCqCTHAd65ZFy4QJE/HawLA9xrAgbtngh1vDqRO+r5WTQiTP
97CLPtXkNpBqw3bLk03vs+tRioQtw0HnQnLOOjuVsSmsq6+UMpAlmfHNuiH6QBTxgytQ6hjnh4Cn
eNcIlYb/gKmAO2kdbmlY3S0LT6hxLjCOOasFrGtg3rYTs6BnLN6oGtnwrbif8jF7FSEuhHKfOsde
/JhIM9Fkl6JGfLVgZU+EVs0v4DCiZW9nvHctd1sFc+UWzKS+yD+nPVn6eGR8Tpi1inwDSpio00nK
UTgLFYJ/quAZgNBFa5sFLYlYXNIh1nzzGW+H9/Neza1QTHRkZ3tv/QXC/c4otEXNlIsJPddutLIL
gtum/0EROcaYOd1+xMfHNEaDVVa0n38uPROwFPRwvdBZ4lWpFSYjMwDh3+WEF4PP+hKABZmSip2C
vyvufXi+TdUduCfE0YdnXU0QinmZBae+UgYilRNyjR9MRUBMPaolRwe5b/HdUcFXHByf8ZRA2D1W
6/i/Hp8D/36n1H6zf1w+kVywmgPtyz02FC7+rMc6/fz9UjHYYvcyBEfGWBxxzS/e/MqCvGfLfz9h
znuUmkySj3SELlhGOfiAPi+QfsAgrDT5/B6Ij0uTFm664vHnRcudOru7iBFbgsESMqZqGTZZ1ADn
+pEHSB07rKa29kuNBRlK4OFvlKvEPCwJyw+ELSmtSExO1+eRx8F4ei48/xUrG4ryvg21ZqQ0ROGy
K4tLLiWMPHKwGmcwUbOaYm3+x4wwxOvC1rmQzZ0V7OyDaWvyh8l2OEp8dc3Z7oOwEiJD1wZp16hU
JMc/pgWfMS66vu8mL6fdb7UxWFS5HJlaQ7nc+6Bej5Z6FztGbM7zmXgiFOeopjeuex0nIiyISxWL
V62VpzdoO8lxstjHDiDMPmOgZb5Sn/iDNbO6DVeHxts0h391hcMrFOwqvG5Yvr0lUn8XxWj7iLCL
I2dKY6/dh2xOEK4JRXaZn68Ro9h2ZSiABoW06W+u+nKrYJRV0eAUIHiK80CV/rSZ0+F6cdH+Cl19
ifH6LecxNDWmNvNskrXpNW4Kb8+37hrLQ9LyuC2dQ8UzB3K5HeRmOLinieMNqJEsHEebCyb+Lonf
AvgOBIYEQUyxKL/UK4zHC8JMD6GjiOmgX7j5aE9YZ6pT+W+mj6U30ksHPPm9HHPrQEaOMMDavgvj
BRnSOsrJ0p5Qnn6zHf8xNA5Fa6u9AM/pmyydn6Xz/60T40VGELe9MfH++mqSXKULUf0ULZztHy56
+jZN61T3WZ1ZUcWnczUwbv7kGmmdwUiy1mPDSDt9Gg7+BxRxGvcoqhPM2h1xgVUIcNgejvpC2bvS
/pfHmbTurt9FdNUnD1gBKo9ltzKy+r+j7bSPTtTIaE8o/R/++vvlS+fFcQn0d4fuh65BjJocxkWX
/NOHvbp+Z9LQov2Ck760vyp99SfsaK7EI0JCUUGAkD0GQZdiDZF3+4b6Bl1nPVRnPkqgGvHk33Ri
5+8Bfxy/Ye7PRVKlL7Jq+gs9lYr+NsDJPog3Y1LQyF6RMvfBGeu/LCem+5Xm0QCK2rSidBYl+SeL
CH1b40dywyiKc+lxsIaPmu4FLlcmODtC1v0QUoWiGZaFPPS9iGe6UKR5ImaY01KTM7fs8CqyNI4T
Go6XlU9e74yhPlHYpdEcOrH0a5Nn69kUYVhliffX+S013+qo8YzwxAcXnkuXFinUnj6ic3ctLtbb
AMtveR69O6HO6nfefoTjR6wEshBXwVZS9llbIStqg2YAnme7praeoUBWIff7mpYFoIPS6f0QVGKf
vOUOvJLzGzhedrru1yXGj+ldGOdl7TKLeNvoJ2YPzkV886f6B7il1n6zHorxVB1znzZbm5xIk02l
XhWCYy9nDo12NLKa3f/IZPjgaqMdUB5k3LMSWadHXYnOWMGMgkJYFvALLsrIo08+IlCrs3oosZ5U
PM7wBlCI6CeGeLAlCRGo/Ta6kP8/fzTXX2CweCt2N5YOTrLULanIFu1TLb1Rar+R5tQBbIE3oNXP
2kGaSCX5+B1A9g7DXInH0nCsqA4uTlq716U+jRNPrOqeVVkXFKfYZTLqvfrZp4RCyRb3lnBmzV/2
iwwQCJ6l/KwzO8HCKf6I9po4aXWVtrm4+xy5oALVj6iSdsxGgdj5HTThi471GYQTtPBmuYYpdQp2
aeN9N92hmm4Ve2gP5okUUv/6Id6NOoaOliUM/5rxsgbQNplYrClOCrH3KC3+mLBiaE1Ioe9Y5j73
rUUTdpwvKlgroHm07yJ0OOy+I/eldiOhV4Y2ADr/XAqAH6T6GcZJaW8uxHi7m4oMwfgb6i7up1qf
v4Dnruo5BKiKKQOMFHWrYSwggSa85I54siGH08xJR8SDbIZGir9462BOhpTXx9UfNP0yTJafY6h6
CqfEYuOkUNNIgyeRejXMzUOhKrm6TjGAPkRC51InnREwLNzO9p32J67gCWZCQewGmq2+x87jvORp
mjhWOwbjwU4WsMjvGpT16KK0hAboQ2azfg6LEesqeM9qE80o7aJTPeClecObJ4VOoeQLPgvXMxhM
zbuVzZrClZQZLa0+S5fYsFfT5/fVy0jrPBRLNnKuX8GDVmNgJPzvdEbbJUvGflvcLgghhIt0gsRu
CIfcf3xqk5+03uHeDEHlbFK37MbZjFsIFYzhfarKPRxqva4t7WNwGDH6NYCJYwbdoSm/6d3/ZOjI
mn3FOVZ4v0+6JNqVoOKheMKeyk/tjROA6A0g8uDhKty80JlfwocEuMn4VUtSWsSZsQfWlnqaTHxq
cNx/kc5AOIW5JW2b6+X8rBPWGY8Skl9iDMmwo/6RmljhFW8gEvfYDWLFogDjz0nI4vpLLXwOFP51
nWMBl1UG1/6KvbTnJJC0d3CT7cHKD49kVKXJPQF64+5NLyvISsggFvHf8v3NyrVgU/mP/fcvIWYZ
fQBNVn7lYr16aX64eJYr9eJgr9dC7Hnmt0vfWh9FdGQwDffp3mpzhXC5DgYtQEpHXyGxz5bIOyzI
PSISnG3BPkZoTudLNX+IX3/c4vrWUJpE5urROHH+Fev2N6FJQCqwB2wbZrpoAlmAtIpvM5HQTqhP
32WtHaLHNCFQkp7uEJEfbVlurN5RqbkuQCpYKah4LfcMiT4BNN3j5qkNpcda12y3Z8jOpRhiIm2+
eREISBqVGXcvkVGYJksxSHOu907v1FBhqKyBqFhNZVP7IzPRdTvJU1io+/JdEHCEQrPAxQCYKkJN
sJf+QPvsP4ndBCF9q6C5bLh5kFk7k7YHYJh2l+lOlp/A/n48x+8JIpPH6Vw0u7uTJ4/kEUHerFUQ
pwanBU1ejA32MEQNi5yZ8HUqMnljqRIQFsAZ5hd4sZWGRqvVG5f+vuNu5tzWRFsG6Rbpo1RcY6/B
pRp/PqxY0kNulSM10+YSlTQnGQTjAxnBs1eJEE2g9IzkYuCAYOsCAgNymOnd+Ip+z865Rtlhw7MA
pZSjaMPyHWQtMkV6amaOuWGqZTHNBSmCi95JoXIHwxYxkufas9sOlxdiMMUPkbNDH5Edzi9tN//2
E9nJ7/a0PMl+p8/4BKnFeR/XNPvx4MtlYtvlbO6RwXSOK8KYU73KcgqPpuwch7g88HoeLL69E7Vw
XE7vfmRcGPx6cfypU646f+367r6PQ2sWJw2A3LOoi3/l6VJqhDl2I/TvcVUW+k9iIVbH6uisRWaG
ZmDw0W5dKkAsbKhf19mCb+H5e65iBBHeW4sy9C1jiaxQFM+b/f1dwDkFZF/G3pHrBYoE/zDHFpVI
FN+uTQnrNH99zZbyRFHV16CNml3HDkaSx3QSjZOjUNHuW+o9+y3A36bpYhBYlI4/B1Gb+XmQBcGP
Xn4xkpSXiUKiPu3y16YlFEKlna5mYntqQ9MccYITgRHme/eJJfyAlv7c0xXUbNo40zh0Ihemttw/
wRU7dDbCh1SLZRwqyF2ErkuOZG2fbPsQNeSj4YgA2KfOsejuO5bGKrVDXX0VP1Qa4BzZHcTjdkhe
27KOEhjitV9qeCPMZzZKMMOavWqcbFh7Cn822+MKM9brnyQiEnsip7UbMJus5qkCARM9QWx0plQt
MpQN2h8U4H5n50Qat3mLzsEdNTBLqMsq/BiWBV50vPjDrm3URl+vApnAfgchQ8wxzAsSqL+INiAZ
YQOfQFifuUSn4X+TaAWi3jG7ZqxHVZ/IxofQRaJoQAIX6JQ8dhx4TcUY6IJDJwLhLsSOlYNGrmUI
ND1EAe0L6G5UTvF3v2OaBK+KI2puRUJDC7xDDIwGDuxmucpyO5lXj+bESXwDxD+mx7cUHLO/BD4W
+kHkPF7jHJ4dwiv8E6nTIC/uoa2Ihi28YQVQgUcAmr7w1GPijD73PtY7k3qJqPJ1fzTxCOLr9V1r
5nRbkRrY+16wCVZVjnYtW4HJ6nkNZD2s0OzPqEltyi+9StFz+ylrTAiyXsXfCePfEhxvtvkoTH7o
9ue+QyZv2x2SgejYWHAk2SosHZr5u4/YDmgACzNZ4wk53K5EdkNPi9NE1uRMZ/LMTzpIIQ51kxho
ThKY5KKaktI8Cbjyw9wVi1PFnF7gw5y3DM/D3JEJ3qi/XF8pCggZsPYqMbB67+vn8DOndU9vZAY3
10ATaEdkbC0B+PTlWbnLuS6qfllJxrUi+TCXAGch57qECA43ZUanBIhzTauW5kR1xuDEDSA5b9kh
oEfY6xKGt4K2LbZ54Oc8B/PX1F+yqcsXF6M9seMvLpYuWQ6ti17gsE93lQtsKnNygB4bCsrkd8wO
3rxeOGqRHkqdCKNyotwUENKw5FDa2ivep/6JnMS6SE0PsJ8nmZPbNbgGSZCfNj8NrjtysIxBy3ma
CV1KT9LIH2Fz+m925gHxL9R+Kn7w1K6NwfewpACZJZxVaswQEKMRVd3pEi6MODDG8wJ5+y/bRQ43
l/Z5Y8YnziMOfDuyQ1bW4IEMdMnTqLpvg5EYrb+154DuEzdxhTQ5KjFaERx4xvZZT8MXbIf46Jj5
PNs/Bb0ry4mTKkBlBEGFbPieaSGo7iQctvTHQPH5ylne+NIQz6KPGLQZNfuGtUkdZtYJs+/uy52D
FPGX9V1SERaaCVmsltwa05JFU6hmGPMVi8e1Fz9kaxirmyxWHR7efTtFCyr/VcibpDnZezmHDYXR
l+5rPDQX8DyncSPLONZFtj/8TR/wqRb95Y0jvvON30rjKVh9t2KDmRqcEA8I5v4TTdnbAlH9MB2M
aI7sOupVrXsEWyaiPRclPiqwmbdH9ua8ScQznpTE0HX9tgVkTdLRvMXHHdZJrs80sjuZYx10C4QL
u17/ZB/k8Wm7KPHk7XcgOgzgt0cnqay8RwSyR8+NivjUI40TlvivwLe73NMvqAV+gWMXMettM3dZ
403jEuVy5IUhdbMyDQOuOfTIZsuLWMiwPWoAeOECtS4Meh2TjvwdW6rE2SdH1MNf29jyIDmJ1Cqn
FsVGTagJj2EWEjFHzSqM0kiAEVkWatlH9YzfsGAUf7IkVKT4pyEAo+QU90m7R/yz+RxHrIbL5Uap
FJL4lU5stC/6ASbZ97OSXEbY7KLNR+XgSMS59XSrrvXCVegIxYTTp2S59KRRjxpB68JodxcdRMDn
K7uHRNAAPKQv4iYTf4T70lKkYly8pH/0dgStKzOOppXFx32zOH2rtTPdTlanFjaxHVikkc78yDVK
CHGoHrVv+yFzCPYktcFkRvPsgY0jDcPQMbLrE7b97fZv40/gSJfnCMBUp2oSlDPyMKLko8HfYoxT
iBHEMgZhLhk6MCUSNkIQELot+cSJw/9QXeqN6FFYXa003vq4kW91lXSqGc9yxtQZmoZaJSWkd2Op
Zyi5sUSD++aOc2e1b6Hit2jdMv9Y68kkzlfvQwyuwe5YZBnU/ZqUe7/GGbX34YnFaSKil7QjWf7l
w8y8KKTIvwQauOwvvnzIRUXNqXkG4Q5WaEiHgE+eK2M8pgp658uIrAf2Iz/MPwyx8wvOWEDFmvDH
zWXNZFjuCgfSlW1LKxcvtq1RhnqJtJK5gJUtxHY/E7g3q0fuZ+QMaa6odrvhuo/COpmUyY5ZBuS0
93MWBaUE4FlZANTF7bZlK33MuhIX2RxokARn+FyW1xzLyuGhL8URs/Xa+rBDWQGAk7dJCAOpsmWK
U4PAAsxr5aW/rIkX7ThpL/u1hF4F+vfJb8WKQee77avtQjRlOaWjbQZj78JGrLLJpCoyqKF3Ql8x
1/72YNL7lHiB4EUpL6MjmqkumzVFGXVORZbAPlnV8tWP/tV/GnNmOAh/UvpoVaG7tmjIFh9417h0
pD4zqtgx6EAeLQ2PonrcnG6ggz1Dp6RMTsPvcSvlEgR0G0OXmkNuy4riyA3ER/POOjXgjzKZY9LV
kGKNkOKkcESil+j1X6r6mCH7lD152qFE1KjIJnKJFduwklMktYcJ9FcSbS2tipTkspoaASnsXtu3
WmG4SyZYqJ047wGeYRyyxHyrx1Hq43LpG8GCwaQ+xNYB4HtmXsoEgyuEqc6LXEmDWT8BS27TR8pt
yD+msuXjsGa3xETzk2IxNO79F2M0QgbTVhrg6MvuEiGUPBBDRxIMejmesKD9V1372eEjAtQMctwD
coyz5Bj1HK57zQItRni1AvONR4MI5hhI9wr2A12zgCfzjbeaEA2U6ybvByIjw6uH+Cu/knCCEz+e
1zvK0oBXgzt3ASMhWv9pz2yqw2JG3ptbBwFLdk6j7wG7PEFEMy0J5xgFDnO+OHR+PmObEy9jMrDx
mQSDOMdElkXA113429jbXUuiXfw+RAhgrqrhqDwUUUQwZUCwuWxaL+AS/QMm6C2+ZAp4yMUbW+4a
02+9PgKAO3zzXT+rA8nynIh9tWcMVa2iShJ9M+68TCyQyZWK+FeFv7z1dKxW0fC2i0dnNQuqwwJz
H2lMrjzZM+Jr1klD1caBpkGQ0JsykF0ehiLjdTrCXQxo1/0yPfh5wQU8HRTY18B6RgPOswx74EZ0
rSfeC/zK7O4Myq2MYLZN6+v1WqO3AXH0Zs9KYnCKPYiUAiG4U33Z/vm2uVsRA2FjjoOhZMyRVi3m
e5SIxlQ/r6qNx0Pv8PjrdvkuH2k4xMStGTkqs7qzi9D37sDt5/itGdD/0Fwxe6rjPri/YsDG2cu+
N1WCbe8PMeZSLJ6+sYSau25XfyUCQAFP9TFkwbZob+Zm8gDiGs02gATwIuT4z3EHl86ZLgXCHvxe
2uTEoVKLjNGKv78vNWCWoUIzqQEFGVMPJFwFuF27pi9KosgiRFXxLbPT2yjH9XDlOZt0GWWYaYU6
jxw7SO+obF1pcdk8UtYH8YsLcDPXSVUMo0xZBty7fkyxdWXJQIDsuJGI4FTYEh4D38HE2wfGUQpF
nzf59wxmmu/+tKYmsZ02ithe6UC1wI++QmZfzSnu0Ifj7yBMGWinpKD3jO44NJkPwIrL/7tP3D8Q
o19MP6MQF+N3al4NMFb9M8gBFtl+/VgmS0xeWX9qXXZQYlT7mQBFmIxZw8LhAFSbLlTFZF4TWXxJ
LfnDyXHpHzPZitsH6ABsWZxCKpEX1uWKaI+dyo67AtDFEHvzX1ZUUXYqEuhfs/1+5Rpsqwxk4h9R
63HU7pIohPzLVUoPWDNlXv5lxIuS60p2IX1m0EkoreWt3mtcaWCyKLJkmUFktAL3o5O2pyQUqHZt
zbjd9h0VKYCXwSTYUglRzPZxW5Ixogf+ABm+iwIxEIbpsWU6l5RkVExsIXouPTIQTzlhvWAW8Kxc
SUQbeuZahg898Q7ylbqIRPuHRvoy17bho+loJw/6LJ4MF82SLTuh1uRW0v2rDJ1CVMJHtKu6T1HR
DE+hglzQ7WqWkIvkzJagUrtyBrbvy4etKSaArS8PUWQIowa1JbTMKej66lwf1h2I6wQlEm6LFjxD
HeJabswYDgQ8j3snAXLbsz3fLZAFjenJSI1QzvSucZ86XZG2V/u5EmYdNTgGruSqEqKUbi+PdxKL
KTmlwY1sbO/8QLGmwBRfnFLQoU185D0FI7e6FwLdB95r9BS91lrCLhk0+OrdTXd+qOja9whb8hHR
XoU1OzfSKtsXv3/mxrvzrQYC9eIi89Cbqe2W8pCwJ2DGVXgeviPJMmDvE4NNRAAaT0iBdvzxb37Q
hKRSGwI6nD0yL+xi3FwfBHcciolGbpgP2aM5p2sk0VgmC4klmrfzDkbSM+vKxv0u5p+N0xFybaST
mU+pXTRnKTHkwc6z6eLLzg6g1/MeQc3Xucp4ruFI8XDbJaaPXJW6jHWbxQu42v+cbCe1QjnzmsY2
9SebvguR+TBgu07hwJeAjq1F/t7Hd1DCeJHer1r0DmJgvnF4NYPeYfH6+ESMFZjutXIICXJnXF29
4L90NP4UJMJgpcKgDIzQSA5z0vsGrGB21DhqdKBD05e3dc1I62zQC6mdrdafFCn0i+BzXXxrmfsp
w+AhweQdl1Nfftxgkmko+UGQg18GwBaI+sEVeg4/3nw/TLrCa5zK7zPTomfd4aYj1LoYpDDbiD8s
hfkQXn15ThpVjh/x9i3P5QwF71Fu3yjGRGbCNilUSQ6ysXeDUrwv38sIbgGrXte54LVJgvXI6wRg
EIdUvcamDMQQifnD3kWqGTamkFQbyqQm8NIdH71zdJzpsqNYix1K7BdEqt0ie1Ezx/YD/DVML3th
jbv0qwRLHKhj8RtmwbXiIxsVgBM2DzMuYArnB7cZFg9qJfy5+9g8YlnUVbeb5C1eY5PUwE1jtUB0
bbmkmRTdJbU1BiyCY/xkbSXWamAw6QSDqdpyw8nFx5QtJUWT2RKu1dLoEfxe2pQrxDg9QSMyT+WI
eAGvHy321cROw2Ci0pXnZXs7GZyRso37ugKE8GGWSrYH0U5Vlxl4lVTp2yOyc64ifQ1we+CDMPsX
Ktl7zDNk14KEEjJYI8PnogQDceQS/yF4II0n1jDJZs2yQtvtx6GUHDL8FEbE1ef9VHpeVrHclWPI
DpXY1HxIgmFBvI2Id1pLCkrh0/o+zJHa75kKzBR9l5ruVOVSJb5Nen0QbMkx1l6twLPHFYNM2Cu/
HbP8Aa/eCWf4JeUmp1J07NFndUzmf+zjt+Dr/K3LpkrUL4QW1qLWnKQ50Uos8GC8N4BdVwfGprCf
Rzjc9142Iz2PdEFAnPjrZAHdmTIrxHYKAllT4b9VEdkAjhlKRX7OlLdenbJ5u7psXKYbI9acGFZl
y4iRfLNlc38x7XSpAuk8ECfSGIT0s2NvnGPcSSg2RDSshhGsTz1UDTt1WzNx4WTcFdU9byfIA5lF
oQ1BjlZJkajNpHC3g0oC7NY1e/4C07cLwFfQxfIg4JMcvbiXl0U18XNr0dn6sEOAe+8uwuc+Ujs2
zYdYe0exPpejhwUUqDu9Ya5DzMHkkDr4n6t2BzU3YzhRMS0zkyrFbNK5UJi6Etgxb+jjW6Q/Zvnk
+x7cDBRmhui78qgvuS/GNDt0zKPxKzwkSAA3LU/VVCp16VbVQBsK3Lm5LvSjoXp+ev/7bO5QJsip
4vFDvSjWpJJvjieBUUidRXCM+yfOtzK9Yu7arh9H2LYNkRQ6sQYabAMU1tVBpJHo9znzmSyCDWMu
DetQuw0jO+SLkrLQlRL4xndmRW/7wnVmGLyBZ4a0P2vuRSzVtYRJsh9QGe8v70HqE2b9z3zNuCNE
Q6P6x3zqJOqSp/XsLxiEf9IeRJAMDvPubMGMZqnCKio4d//ylvNt+4XMsf+8r82ac22C07dhDUXR
Wlk0GviLqT74sdtjgN1CKvFTQhZSU7iEw8o60JBXjYKeyNEh1ZvznsobHIrwiXR1xbGcEroaUbYQ
Ou2XeWIvBQFyZ3RFBeMpFPaPNYyLC6p57zmUU/LWjg0XWoT9k7L9do5FTrWA0V3EkF/aPQzONVQv
/+FTilYxdJzG95J+ymuNG3UGDmuBZDoNGYD2pVBt2KCsZkebyh5Qe9WIp2OU20TgwUdhTAYCbLFa
sOftGyneO1dliuqDlYnw3NNVC5Xazgv9PE3HzEJpj5JGVM4NYMDrc/JzWxyVrrm8b1Dw2SvI39W1
d88tzONA07q6w8Eoaw/rLdjas+6AMmEQZYYJGnAlJVji6SIZPMO/q0Arxz9/46CIswCOM+odfwXI
cmmb+iAOo1WBVpxslh21HWhOBjd4/gP7VHITeBAkczlofojwcH5MBKYeYRJstNPGLuvPyXqN8Ys7
HWxOMiLqcjTEX0nV37h1ZVLvfPFDWTiTu0KOV3+Ui1adBjDQqqKyv4JwenA6a3SdsIvvBuCydcLn
hDhWNGDK8ROrGfz5Cs9RbfOdiOxhYS+W68hpXsTyjUB8e8v6oLxzfJpEkBT2OoSSnBUyIfaxTcCF
+A+3kdibNIbANYGYON3m91ATj25BNm6q6Zh6qCWOTnll13ZVS+vQxPVKN5eHStthO5jP0J+o20TU
p3bQhEQBqFo13tYwNjYiGwto+BzlaHyQhnXFdvsC/As4LJiZaz0y6CJXstF+oEZ3wglFnfnvD/aa
cr+3SbQ6MT1RQfq2p+NzdqoExwH6AYr9HBh2viUoZzFxfi9ATazmER1Nnw44VAM4EZEzYhAuz0DI
G3VmYdWeeJeq72Kno1hPBPAySrps046ASC6SJ/Pg+VNBj3dmDf0obx2aPu/DYYXKQWBi923NifWu
X1hLPIelJ2cBeD7r7zMQ8eHXA0dwZPV7ZVT/YXeufbF7zOoVjdZTfn0Jc7sZCWCdpcXpNPyrdrVZ
vAhQqVhYijlu79Y8DqDO6dN1biIthn+TRDvZ8SF3Ncs7btX2Cp4EzIr4AC2Ubh0ByQNrjuC4bw0L
xmXnNqhvDnc0LH+djXFY6+TCaHmqeI/mmtQjIMdDcBT3ScuWi5dObWbNREH4In0IOehJ0rQ0Y+S9
AmNSdY90zhkaLyu/Iz4m3GyNjD9YkIjPKR5DiMAmMiwejrJ7dT2985Aa0TWdnpf/Ri//jq/lqxdB
z8wwbHEbyrg51yhMOpYWtWcSaT+gGiIBjul0gsRX7PYlvwMqiTg+mJYKfpa0kMb13h/zMVR/uTk/
xHtuZsRHgWpiWoMtSfn1qgXF+2F7LBpFq0mStlmxtQEPqY8LGmaBWfarHtJK1jNjFdpKNJfogouL
nHPF1QQNjHEADN6RwQC8G8FkFe8PmnmCygxsLgYG5kckuwsehZGz2UbWrcCMt24yO5ODnNdOunrb
02Z2x8ZNDgW6mlZrMlAzpcrqvnUOopeB3DKPpVTuOOGHG1Uh1hVkt8izy/Cf41hjGIytJ7UAPIuN
Hb6UOaCt8ei61Ga97+3+EAMyCfI94JNztIaUg4SO4WnU78eij3xkkWNIT2Infdss4QlwodpfNiR0
OzX7IOMUJ3BDZ9uJQCcnLQ3EoyHjwj1XyM7a58kVQL8HIey98HiLfLebWpk28TqHRGUFDop5L/O9
F7wFnD46E1ocfI2r9tz2sin/DCdNOy3VspAry9r9susOxcDT6Z2nea/fUl1MnLuhhIa2YYEZfH/U
IclxXHgYqu7Cg05gt06I/vKP84s+vJ+mKQYdKn6Ptry4owYfv0NRvhYf1zrpE/3496AnxfNfZkIq
sknYhw+EtLmqeRfbTwUEFLDmtM1UcX9ZYDr52xZ6/5RWqi7jiYK8XA6hmvJCnm4yHwPufFNRp6bD
Z7uHOOk/f4ImsAnVTx5OxXgV3LCkKJcyeO2xyNYFuvCewFcDVpmymcsisjwWP+5K6nGpR4mZdHaz
hw8uqUsDaOOuSK9MmoaD9wSo+wFkXJQoclOwlE4F0nUrnv0l/ZZSGCbdIKafJdB1JGUYmVc57VTb
1mavdJqLWCLCDU4fHCKUqmpYgtbwjJiAqQYdthTsXWg4nPzvLYbUu0+DSnCFX+kHNz1H0RvNPUdE
ISwhzAtkIjwwl9PQf9v2Y/x4m9sP4atseMkgkCAIBbskVOQnS4AKaQ+5pIaNWtefdLJ3mOwgm4D7
Cz6nxEa5FdVyAE3k7haWIGX/gDYVBEex+/Z8sxx2Q0kLUdr6hQcdNHf1LcSmWu8a0upy4OuWNLOX
ykeTUBgPQZifXswbXhp0WQ1f+L5pG9EM3wccowvHIwpCspZ2qkDIfNhvjJF85t8uyNk6WxoNOVHz
feklz7AkGlPF79z2FVwlDfLr2SPf78Hi6zuq4XEbNKCOsuT+cMhwxeALhOQCEnPD/eyyW9EYW7jt
O+Aau3iP+EBIMUcmer0RTJ4rNSDndrB4W4S5/5nmI6YLKZZI69ucMhjHAD7QpocujlD/MsmNDjsV
iU2yI3QiMx3nT/zBbb7aKqDTyaRh4+Y/xvrjcuj5IHH3Zs1OTSDjYxvfBLnD53SXhbCqacUJJ8fB
GamiDI+JbeL1yUHlriovQnRQPlhQ8Ter3+FZWNzwNAbv3YrIjzMt94S40s06qZFJigiYil2KpmrO
XjPrQMioIsgi4cdj9troUJz0UrWVNeRJV3OlBzOcKPbon9kKMY68f5YrI66Y3pyTttvQn4m8n1UO
qFzRBESWzUd7eb0g1AmN7HBPUgZ6gnpQI1GxMRbPw11P94lQVAoo/3IY0thWRSO2Nx05cRb6qt2k
tzqqK3Y9muc0BLbbiwnaQAxf5W/VPh2apBdKM4dp87j5LchBfvSr0+iehlmbfIJhepbhEsahhLdf
p83iDh2JOpKg4lBHKjQWvocT0TtBJXbsEHrq1aIhQBIbtE16YOOm+ZcdvozGMmgOrHYrri8BEuwi
J3ZFmj4lQXGom9DK7GIsAGCPosM0zCJ5ZE8eE4ttgOwLizElKdjD0KEeLAGqv+zrNDwTqmRbnead
ZkoLiZrkr5YdtYWgss3gjAcDrKxEQsu9Zyy4u3aCnrUwGUmjd0ZzmzuelA8xM+AOLUt+oP/hk77W
KQGQrEEq96jplFNun3jQszT4iNe7L0xg68kN3JJpDr5oynLd/2/QjtF6zUIKipvpwYmjhqU+Xn5A
a5rPE/2niBglOqaa3ntomP9DCBE4FXcc8UM3vJDfd26zYoHOTfMDXHkHmsGx6J2A7iFhPWuZ9IUv
RaYDqRLhenI1lX7xgSP4kkzZGnPW+7Z70ZXfUasj8iX50KYFNGEJ3oQP1wjGLWY3Tvy9X7EUHe9n
ISTyU/KRleuy/7eNqHJvv28eWLgl3w1FdYq4lhfEM8snJRFI6aUxCF3sfcIyCKkdwiKf0RVKn9KM
lYzMP6NIyLw6aO99QevTzMscAj4PDd+O8eD8pr59qkFASZSaKpjVNbqrOMOT5hbpW6yUPbTNiQPk
Bt7NG/yFcjSUZmkM/sORh/BkLUrnr8wsjO+2Y7btpcd844ay3uo4OK4xdNbMkErqVMrFI40o0KYV
0EA21DidbCYoC6LXi8r/E4CFFLa+txkJ0RWptc3DNOUEUGIf/Slz6sjcJgci55/XUCyRQCPBNlvG
K8axhDWWUOMVjLHUzvsaKvqAfVFUQbsHSPt9VUgDxUSyturHqc6n3Jdc7txg/Rnn7rxMQUbeUTxo
Ow5JnHTke9ir++adha+ZLc7C3GGj6G21MapNSXgm9Tq0vabN5DSLCm/P91jwGuAREecKtksNBT7j
wVQLoHlODscK4HnW2v2gGNIh6vXkFc6OqRNRDAe6OxeLP0Ib9BBBY8B8kKAirCfv1LtAH9rwSHeF
8jTOR0rcz7JdJg+YltAXlB167b3f81ei0a8759Y8c+nE4SouLqy3T+HsN5riV2TB9yKWn7dUZUb1
b7Q4fBV2C2/i8a55QPSQ0HYxv5OTymHDSsEW5mzIRck7yLi2kf9wszmRto4SE5tj+x95tTjFMALV
8TPf+uClko2wfzkhe/tfDJjFy5aD8xOIeuy6j843GNkvpwxfH3BT1laTn/uq5BfofoZnPSjirPMx
6egAKBuDJyvEXYXZ9JjQ34XoLiED1S40EgRjqvM26+5o/q/GkiJCimUwGnHHe5U6XILY3DNEdvAi
aMw8nLWXZP3IGQpev87DqQcePLdD78COKTMd0hKZFCtRjrcbjYgrN/NHzMLdEsW5LlJ4GHYQc+dE
ncI4YkPvUwSD1fnp8q0JbmOkVu3BNDlZb2kkMTSYPSCClL00QY9RKrWyPSxtvDoJkt02V8Wv8xlS
QvHJz6Bar71vnZiAAiY90yfuoIOzVzTzZq8Xof/uXIup/Mx9688xischeSxrAgfqAByKRYNxmRar
4nMum9Ra2ulQ/YgoU0g3ijQChgRIOCRfr3vRmxvCABIQFsRPbIVJQQPo3WrRave6rkmp0rk0fvcd
QxwSu26FXw+fibfdQytwDP9L0g6sSGUrW0mKqKCS3ybA5ypD7oVxUgdCu2u4N/kOALe9JqB0XJOj
vw8dNqG66A19sdauF7ASPRAMW21ATwFDcVcRomsnS7PVd993ImrIVc5o6WdTZVodPwnerGryehEB
49T38CJHBx7qjghwZKgcVJyNMS9xNaWbbly4WrP7O8T6ebuKcesQrzQPfPWlwIqRQkqHXavxCFYU
IMSyMVxif/tvrP9Rjt0SI+Co2DvUPO/TtXH5TTceVMcqymyJHHaP/S38gAypk7aflZJwTcRjTCFv
tkB3ehg/oVYcCzvW/Fx1xiOIfR7fble6vD9Jx3Iv5yUSZ2TnxzpOpRkVpqvCT1KfjW/PM0T4jRE1
4IovV2m8TMRIeff/t4gzeEDrLXJRmMtOEZI5b0JdSez5cl++iH4Qqnqioi+Bc9BjQlDAlAggK2C8
Ej53jG7nT3yBEjpWyJkrNAwrSSGvtqGahRSp5QHVRkkxD+/kyus8VtXZyBr5DnW0Hpr+kFvkxoen
MvZoqjP7lirEUQeNHJkdZCh33xoEaU4rB+9r/mFTcFTU9RTDfwJ6QzLcLjdUvvi4keMGlc2wIDdj
3Kx0l2n366Kwe5OAS2koKMkvHAnytuG6Wd8+agn5WVEjpVtk+uGo2+1HHpe/TJ3RxaEZoNGdoFCD
3RKB5r0C/LGmO+kUi3CLfHm5ctItE2gV5Y0sX9/xc1w+h3OiVTAawWG/FJqrBJi53nJpHWuFvdjr
0wqPITMzq5bTaevxiXt+of6lAyQVjkdOFU0+BMTRe89xqzjfJgwV4U6e8HfsfgXqKEDWEmZaCsmH
4D2wafDUTVEZVKvGy15VtoJQP5QLwbsF/iykMRMvOspbAZ0trkEVlzjhNFfhexyK1W2++Adp97fN
tz6/9UwaKB3oRc09aqFIXwVKvCVHEqEkcMYfCcsvowc4F8dptCgIWAXZIFm0PAY040OFafkIlAAk
bv261ECl/0+aURCQwPJkNMj0qnuBk/7iKhin0D57Y77Hp9L82pPmQMbJW/JqPsGUhj091zxwW9QP
miYNsaYGrJFt5PqazqHYcgaXoJ23MkvADQdfd1Wu4G1N15zKjOfZCaFwqzfUZypof0NhU/ic4YWn
/oPvK5w6Xz3aZ0gfCebcXIFuxXo+Wo4L0ElNy6mkulvZYr/qtw1uhLq1GD+k9pNkX6DGre+ZC+gi
kkt/eyLcty2O3debq3B8rzLN3rwLCBnpQIwxLcvbDgwhsC9/R8uHpF6QXcqFSiTFi40QYpvgNUQD
B4vrJTEyRYBKnfAV9iXFMn6PqTsOFHztPmIUeHaw6lH2dwYTiObhhozRvOOxJ9zcpg/a51HUi3IV
F93OS0zzIV6xcKfvdsMbVZtqv5XkJBPmmU2QdKftPdXrrZ+UjWpHF4Ma65TsrJmfrKwXvzrKiCzA
Pr/h59DGoD+/4rZ5VJWiuMH9LQHyyR5U15K4VVt2gUbTDDwH4ABVkxtVcpbBhCX5AX2ylanuL7uG
UJJPbPWuFd9fuZSHFRp21Q0bKPSSN+hyV94PXBNnDeUScNszhwqi3GwKopOEo47isYgtxBthsdQN
sk0o5hJRJk6XJlB8hr6DGmtlcEP1iBZDqSd+xT1hszdCEVfQOwSICTSOpXoOWV75Vsqkjc3Q+c8Z
aOIVUIvQyOebHLgC6SB56VHta+vjSh8VyK/Q5Dex/N2ovlt3aPlP7f5Lug89QLxJi/HbN/mhPi3I
4I8V5ZN85yty6mOEPtruo4zwRfqn5A9sKmsN6djtgcT4Sz8GML2yRzwHSk44KDVlnzwDPvvV7mda
4zFb8/hn/cJLzN/0PPnwVML+mD7AREZun38AMdQuQ5QTJnzPI/ei3J17V+lTt3smBCY0LhFb6Cju
PWcuwkZ7zkMkwrjrkyZsFXfzm/ZHCyv0eC+TtPBzLsoBPGiufjtQgiidamaUHgvK0g2G1eCy+W/Y
qrYzpnMf95iKKx3vjMhQ9E8jPTqzR1CPfVNSHFkGd5IGLqzIe5fbPjxiuA3IecjEV0d/tdDKbawS
17BoQl7Afze6iJNI2i2jrESPW7noygR1d3rGgTdR5MmTc17Txky9BCZj8/hMbNdQIhHMqglquqgO
NjZCuKwVBuMQbdgNk8Och1RNyPa8Ns5xOGsRE8mPikOtZCHlAMucnKWC1CYqWCOG8rxf6JRtIqB/
bFk0PkEmtsCdw/6O2R/3M8ybppJmjfptTn4r1Q00w2xOk/aA6UAtpEweArCIMhp0RKmtzBx58693
71mS5wC1KXh+fuyw8Nb9OymNpmSR0l8K+u73FhOZ1tl6tXLCnjKsS+eZE22eUZrPHz/NroiR1nq1
BBcTy1JuznTiMLzA4ckSfzX9D7F+vVXrPxTFqP+ZdE8FmMWIOzxbNPu+oi9cW3OsYwCOXfi6vKqA
whf9wQiWV5amWw5S4vVDrTcLXvkl6V3eewR6TWdN6k30cRaGWEdJH5JRFS+RqTWh9cNsQ/ZsTYFn
nzFdRe2INaeMWDWqNBDjExiKh1l4e/1M2eIX1M+7LgA+cKG2y+4xL58vkO3Z2qoN1kVTLcmuIVwA
w4cvwnB7zyDd68N43TdwbhM09NGAta8H0wncnmCVLcPoTJgPnHKatDxaRmqcQun0RXofobyHlUc5
L5HyZZxegKGdLYDw+iOSFguxoveh4GAGRrs/SLZoe2RHTWMfQEFaGtLPGsdOFgL8gGmbEC9TsAQl
5O6wQxx879gOwwu6dxzZTAO7VQC6KCY0+xprsc77aDqeBK1zWg215FTFmrWurnhqiPwRHQQpgSJR
rkh+H1QHHICldYaShnCNFdzz1LWM87yola3IPQsa8NxU+8U0uEevBKwD0UmznW2sSotAjoBdeOOi
CuxUvLX+9nlYuGL7VfIN1jnuoulWB/9Erzn96XbhbYz7Yvpp3+/Z4uZQIsg1ZfsvRclgO2VepOll
vFqjtUrpS59KjCYkAcxbgLNmrq6fsZY1Zr2ZiUc0SWXTIkMQkbriuxW0KLt7tyEBJPjHX/pzvkFb
Sa5g2L8ZiCTMEKW+Ws1a8mMsXlSufKtJLSfekNXy2f4AGkhXJBVU24gNw9YrnOVuCNI658MNV2hw
HoGo2wAkAbJ8ozFqmg5ocSzeIrKWNixdHhEMJxj8IaZp5aFipdVNeGnHMt4dqudUSAl3v3p7nTaY
ca2snnZdyM/4P/efk+an+v9BtGPZ1Yi15SRLJGx4R91kz8WA2gqG83EomFZkM/Yg4qHHzH+mZK5J
jbZLyGHIdt7ZHLEcbNXFb1eKAblRESBo6wFU2yEq0k4szpiS1CmiiWf2x5c3jid86I87DdowBR29
UHdPYBA53zJWe3/WyUCzfLH8YbFr8I66ARQ7MF96To7TT8aU7TccUzHV4C5it+J/8QrTzIaUyRVx
hncGgSUdUBh1Lz9cqjoch5OjghVrikF4ykh57ycR1GGSF2hWzWqRQVsHNq3uUa88WFQqVOH6W0Df
B6ECFt4ZS6aK6trEPfr5QblRQfUC6PAos3cKlwI5Ppl0c/bYp/DtIJwHhnSRA6CaMS4e4qQJSYK6
Z9EcJU0r8AF1ZLIiMixQ39j4ywdMMK6tTayRTqijj52veMDul/C9FTLU7uxvYucvXCJzaY3bdnB0
EburSSTKKy0NGRPaJ1r9W78jkmb6NMDpdDdqKWjog2lbwiEEVUC4Ec4ibpG1lfA6/uw9f2ER7HPi
Xcga6DtQP4MEf/b06taKoOX86Bzu+ekz/QmlZ8agvTZoPW927LRWaQ78P939z4BQtZANXBoOJgze
FmIkZ9loLClK3tFhpgxzXLI2j3Hzs+BXOSJcxvkf+o+9Rh4e56Kyq2jhUb3zifpNv8SfPBil1V/y
BFpgsEZU1gbtnc6vV4lYv9UBrMupJp27PdGrJfl0dDVpb8awZ7BG90gJRxwFULDrYnkbQrvHBcKQ
1IQrNSThmYHjHQFc0ECJeuMgMl3rKkUhlMEUZxJUYKN+Ud+7A98zjOjlXcabFtHieSTuzk7GRdV5
nmAW/zqsQYoKM5yjpVgJTAvFQafS5xDO0TFJJsNLsCLOns36+nnvcrNBDNDeMZnI5hPgRM6FSx6V
y5+lFK+2xHCdkjbDDVfYios5atWc0zngoxcOeUXUeiHJas54EGlA+4cwCXAerIv74UnsI/zVQvcp
5r5Qi1BRaGtyl7P8NZrlam3NO6+7ts3xmoTHVHtEpBkJ3DMcvvQsKixTC4f5uI+wI3r5X6vBg/aM
RvB9Gh6a7o6uPnQmV0hapCGaPd0rTDKuDAn42DP1Zy2rOkNluh33xlgiQCc+a5geKp9+0ccaucrI
r2InhEEFAKJWBJ3UZlo47k3wVLFEpW1r9egxgzm5exDzGnDznZn4TnHcGgpVmvcpJHzeNCXQfh53
fML2U/bPxeyh7TLy0nNDtpTcHACP6eZ7sIq2rCztAjkDVZIjkAilNWWhXwNcFTIYnj+O12G2ywkA
doTINdSfq+AX8mgriub0zmOOY/HVKCGVmQy7c2AxQbtYhFdtXIYnpPbUxj4x9NItLgTsNzfx8ty2
L55rDYWJGfr1JFw7TuTg6j+Pd+yzdHnkRdEOju2qxgahiUtBXrUVk6B6YmhtuTqrUEpElqxW4wQA
6jJSAIvqJTWJ+oAWR4CQYT8q5rvqRCf2ko3obqSVUE37yjG5xhC26svR1ER64m3j6Ng+1/gEf60y
aUoWWyK0hxStsYLqR/tOPzDb+jY/bFjBiUKnxnLg2duDl6qQQjGfSyAcSopXw0WNIbcp+Se8mw5W
Eyf7SQdFJwucyDF8XpBpquHN3kFdFCvH3qmKwIwzvggUGxqE03kQcW1Jeg+0EW4X5w4NXq9J1yt9
25GlRDuXonO33p2jDURe/oSs9wXBheA+Xmfn4ly/ysz+Z8FBqnObpyAcHA2dXqarnv5IKoHNVskY
IAlRb5jCOpC+9qn7HHbiWLQSFzRg7y0LlopPWMlQEx0xVQcDqw+TNHEh3pM1fWQT5NTm+KTcq8rv
ucyPhDeK/VpCjRwwPqIWgSxi9TDme5PjSVgzqjf+uEcE0LPG7lRevUdahuhH87awd93Qo+L4wfog
jqIw+O1BOTCU7Icoq/D73Ic4SVQIQzUwLfPlJcGFGjmBlf16xxZoSno8i+C5zwe1bs/9aTA3s6wA
aCgmQgqpwrJBE053brmqBlFURhzP/IdxhqDj9phHt9kKdkSTWwJ1qsWFXioP7eea/0iE4+26+L59
MWJFO0O6s11Wl4auJ06I2PVOnLdIt5rGDAfWI1dcFRB41Z2ZReBeGJ+25g6GD7mswS6jZlqb4K5I
06WHO++O/rQJrVwKQpsHkNmeBOF+tSx5KygYCiE0gjmFOWD95S9SzNnSyn4rU59kmHbrk6YHSrVG
yTuX4NFZKYcoPs1XbuGaejiNTuq6YFLvnawObwP5JXB4WE6wB8QRMC/1k4qt/8OSEBnOzocoZGKv
7vF538y2Uf+/6KoG1xIXL6TQFMFLqJJM4+hr7DgMRLRprjKH30bqI1yErNznxg9MkOyPz8AOh+8N
qupnQcOfDrjzWg/WujS69omxYnnT+rBHOtYDPFkk9T2Tbk6kLM89AWQOFAh9tJ/OOoWNW3j5Thzz
v2KI3zIIEpYEsSns+QMgtB4nfuf3pegzVnRzlEAVVfAyX2KLa0hUDtqgIEaAiu74fnbQq6y62bNu
TDr1B9Ss+LROZoy125aAp3NLnE+TBmMmDofiVAy9KiPfXOdzZ/60U/EoNKo51Vcxv8YHutHlru0y
wYIMfi1vWImmYMzqCWMU5u4AZP6Mb/43fAHOw4WpwSEO4R9oixzbKeS84vx4Hh/qmdE4+SfLW15p
s39pJ/3lMaBbnlUrrkOXNgf1dAyiJZ6nmUK83TcNV+RGW6/e5ryAGBtaMvOqsLufwSCzJ7Xtr3Xh
Xf5R3O0+dtcigxZvT8bcB5G5I+x2H32QyGdr4e3xf7XvWeEkF2ER+lwBx1qpL+t5Tc+53Jk039gO
7VVL6IwgXBkzzNK3lzTP65fm96IW55LcFpIEqDFba/ScEfi6b1LJsso0DuvIXamsGdPwj2e80e0P
FFG8qObne63D/FhuELmlwUTV6+/C1gdpwr6EjM57v11ZItJzsN8RvZiWOGouQXBzeQiI4aZBlk2f
LZ6Bh5V5X1XISD4V3Pn1yut4M/32NUIMu3ep07K8BrFsS8p51RyCZhAH6MQ590keKLHL7vbq0z/3
Izw9XgnwLk/xFts5ZWLLKhpcWiO+EZXlc3azvCuf28PBZnfK7IrEnfpO5WGuKTeFaZELTsvT7+aJ
TiHf3u7evDd3GFy87WiCtsOXL108PumSFrEP0AZ1a1wCwgHqgqQmGgx+Spot/scHUDN1Cw9nvXcr
kq1Dpo8z60ik5Eq+v7twYplPvK+DHAVty4zgHICq9pyt36PcbKFyL1k/JTo8nf8ypR3AcsR/qSBm
ZY1utLwWC0r36fx1xMsZNSCgZtNFTalLVnXsBXjsq9B+Ly2iHzrsWLu5rW/uJkjWnfxerwCDvYPp
+Hgh2PG7YSwmStDODN6EwJKCycX5Z/WijEnk48PGamEI10KgKxXCO+GNRXYyvjjlAqtJNhpcN17u
EykZhEdJp6nBZJfNkFdxQQKYrnwiZWj5SghhlA4ot0wmJhCCaBrQPYEI7l/1B/Re84eC8FFZBvcY
PL7jEvFs0nUQcN2KyM9Y8nAKa383VGBSbBkbFypF9u51M+4QfZ10O1t65nIKp+M90FbTC1+0//Mo
opYjL3eT8/RJdslBhtB8ZUM6u0cgpO/QRwXmSWd7f6usX9qBTYHwvK0gcTPnyrB3BAKeyAf/4hPu
tQwWsoJ0U74m0/lMN4OTSQHYLisjkM1PQh0S4SyxVDLYyvKaHlfqfArxKDpQ5j9Hq73/jY2Pf0OZ
S0Cejr3y6aG2BtPizb7+1TukwtUj0j48wpjQmATga0qXsuntAbGEOVk79Vq93jtyaFgYGiicySHu
LUpa/X5qrrpgPhXn8Eay81dDJhi25S2O/vOBqtwNNVsT9oeKkAuwQxPQDKVsNcdCv/usuG54PHnn
ETXCcenHzzTBa3KoycNCC9ARgCkydRfKnA/T0urHu8k3Je8S7bMGtVVHlgetraM3XQsg2Pq4jSu+
raT9A+Ku0KxfbwVBr/YP6gaDR++bPxCtVNyLMAMYopE3yk/z9VTE/Ob3fvdVpb3dMyk5HWalyEMR
9mq0Sgh/TU+OToX66wYmVlet1s1t8Ykdc9tANQ5KTgN8rog8oJUb5k+zTUiGphEcWW0hOy+aT0yP
0dOQJL9gVZ2w4uHA7IBEEmdfp2CvQOnm4VV/RmjizhwCH/aC8y302qi2iQ6wBow/nbbhyq0pBT/I
BR4z9XMd44cTU5/mhRlE18lWzmLnSwv0eHnF1WKBdUdvRw1DwBpQtY1kD2J2UcodawNCr+gG0EQ9
xfX5yBRYqVaXu9PmLK80lz+wReRbfIh5vULr+rJ6gUaPrURUCNitUPaRCbiMZ9jIZ+86OWnGj/fG
0bVwvjNevbK4VbcoR1le8A4Y5aFIic92O9WFf9C5Lxhv46lfxweO8zQ6ZcaC/OY+2m8FZiQaEzQP
6GwCCdq9ghosu6M8P3gN90HzGXHOTIgAALMIuAaL+g9esu1zmQikcbvyUZexfDI3xTW3e4DNAtXz
tl6GYfLQFWO0+O4KGs2k3RSNXfGLcAuIIqkPQex5wD24nnMJY5NTd60nX9UOdPninDdYf/hL9vg+
pN7WWohgBi0ZS4Am5dlonYy6Qrk3EMIWuwOy9D2UxIK0UQW2onP08lrTM/8XLqINxmQ3f3Lz5qZP
m+kJAiPkhD3aRWx5Yfic7BTg59lNfbosd7P9Z6o/ESwPQlQxNE8Fo7XbF8lM13URRS+/aFqfjGOZ
yD8uhvnAG2GRtFUfDN+pY4ZkzHmD9ZbASF2j07o3622/YgDlwplgTCmIJDyuq6LqtkmscTg/9uH1
vOnGaC/s3PD7tb6Li2WzdE05rmXWniGbqyaJ2akp3usLzGd0aTbnRucM1/Eqm/Y8rKt3BHda9xQk
vuQppI5Bj12z6zafMBHlXkirpQA8I1E1zVTE5GI6nX4vLQajVmlrLC2Wtdb6dUXUkMTOLz9ywUj9
BAue8NUGHg+l70vhu2jpbkJvRQwpBgBfauAFRJa/6yQ0FfzetBlbbQHpaFU9dPOlwOwgRiXIKlY0
XTxxIwhvK86/dQCVeb0HWnzaWGkSiBzgO6v74kis59A9lpt3HLBvtS45dkVL1fh5YgaQuDeojGw2
ARH3YYwCwsGTEdiE9cIFprnA7uOAfprOUfULTVIKdgqGLs8R6S3n+9/7H4K3TsNGKgylwv/D6gY+
cqyR5xaGKxpoCcnTBVRoc6W/e1YrBQISvpMPJ4TTh+i/EqMAOZmW9iLJV9bcL0mFT2TUvSuQFQ+O
zVeDSGLsitXToy24zrTq06aP4c1q3VhjhXk7s4MWSm8+CT/YlO9QcSOjG0lN97wMc6ezzP8M0dul
7Ig2P09yGRsqxNOT+XibE6Ud1Q4Xyke5SQ/ZctF8ru2hGSPXRRMfCvMV6SuBcfe2A5tl6b8TF03t
UXPfUiXtdj+rhPT/vMO91r1Xt+S+oaiJGuwGi9KBDIXpGZL1YV0SXsIcdlTAN1pP6TYSxeFvvt6u
SWqUtoE1MDqrqEBqAPclQcGZqCswRypxBax+5saaOPQFh/TILAXaLvTSTlJDF+MsILJp0TU5jPeA
n2ejtGf9szd2uoLpAPaXXcvchI3GROec06C/BhdLCEZRuqB0x0uLdqRp6ZdwP6q0ETVKaKK/bQ5r
hKS2PFPO95mleNkgRek/EJXq3d+TvPweBeSB6GDaSMeZB/1tTrHHJIF+BWay3n6cCM0GH7pNlcBa
PONRkdGZXxmFOEBJd3Yw6udtxig6uNNkn1ZijDvSfFctYn4Rlpa4IxKOIS4DFKJT1jjh3ippT5qt
Xd8GHBczumehTgeyxZsDMCqueTx/PL7s01+bj+E7GY+626ABkvJPmNShnso4lsFQe0A4zjp7eYxW
Ysd30xBh8ZJ36MGjB7anq2MZJaNdY0pqUojc6BSzUBiuDdtqLNTnM81g/w98fzh8ZdapxkSZxNkM
AQHO9ksCxRXSD5YliKxDXO2mZNbGiwCbmeHoPzfFqdJrLENwtfeGU0YgCWoImm4GkpD3dXkxsMiW
qXXObp4KiNmdldXRc7rjLr4y+ATVyYBBT6InnRKWY8DKpffzCNflk06EW/36q6JTH3eETsbmENHa
sT975/MMDZpiz8mFvBI4/Jbr2MPFXjm2JX22ukccGYQwqaWNMW1D5jp5PqeZz06E3DragHaObH8k
u5H+2YmrfG+Jm7by723h+6wdHAFtggC4CYpZs8ZomCpFltEunX/Oj7QVDO7joTLTProEte9GOKVp
9sxwh2E2vF1Ta2fdC8vxaTDW5P4LBfiK46qLlQQpw8nu/FaWC9dCfWTw7UXugZpKhMaH9yOdplH2
by9Vf1DRJlL+iJTYHphWAN59Y+0X7AcVOQ9+wqK6F9zoibWxJrlItAz2Vt434hQ9AfN7QeG19Qzp
giEK1EZlXvm+AnoN5Ej27ddZ5rFhInV3jOZE+psC02g3IAACSpkHmT1+Q1Ul/5635SCvwAH8Mmwn
zKgblSjz3034gDRGJuXHmw1lvP1LjbNxBnqBCheBJIOwCPRUTAEOVMFIDvkTLlkpLgeg09sDP5KR
QndgMYiuOc271vi6UtsKYoGwa4i3Mh1pKjz+z2jxgc1Jj4MxVYd13vuWU6HB4AcmmSXDscEV4yhm
+TZV7PCpWmCGm8M/P4muaBjkFeXdBBWyaqc5B89AOCABNv+qRqyvKENEbluNBe5lvI+TUF8LpzVd
XQZc0dITzkNgHePlvdWT5odyC7+8CFepfrhEMR7XkqEOY8gsVnNLrjsD89HUjamhEtAdwXMK8m04
CTNiC9mff2elNKa7ArNPzR5NzqzfXRk9Px11JjRNEnPFPF8TzZgc+F8g3BpwQ7H6oBXb/VqiReW6
H9+Lp6ztKdMm046/pNacH/FyGf7QZoD2IHBCWGwUCdJcK+h0EZZOYbpAnzTq8941QIsPoP+tZUz9
C/haK6XH5AaRxfS+6fj58++e3wBrAwhNO52YFDX5m1LltN4p4LeX9028IqJ+ZKQZmmw2MgqziW83
2pOCzTZ9EO0yUypu53qA18EXwhY9jqJjXYdXX3O78xVbeb+BB7QstzOyn25ILZXFFJfyN8nFRtba
/+NhuU28lI3Yhd9vNFuW10R+XU5wc6nMh1NP8PNOxq21iACzD0wr8C+TAG3eNKTanbRIiFfx1Ggb
id2DrsuQs1MbuWWajG6XKUUIL0ocTKymiH/sqsU6xxA0rWuC6JkBsmaZVCUGiTG/MmTY727cq3XO
oYPiJIKeUswui92J4tLTTuY7Poe1KxIAu6McY+dCaGQCZXPTjZM5BWzFPgq7+lNz9tlPM7KDE2Tl
qNL2O5YZua0zOteKA7rdBSB0R+9gk1nh8d9xRzMY7u1Z65PUiGNE0TwcDYnzUt84ImbEl9Wk6ZD+
CiYEr386Z5MAr5vYSIYPo0Aiq7k24GipTffxRmTalT/EttY1bIGVBYvAu781gXBhfYD8DndJxD9f
R4gLeshv4PjgFR7XOo9hl4/F7/Td7aVE05YVyJgQPyK8TR/cpI2yBcVbTR3ZagEwZnfDD0jQzz4E
NYn4tvADksdGiHxgDcbvtYXxo/6UX9M28P6rct69ql/IOW1GaFlFkanFGo7nGQSKNsxjHlRnnBrT
XBXW9a8+7eXPEk+kdz2bJXiNg3UCkSnB3TOCCQA5fBmfZ+W5LaoRPbPVYxFDvKe9+iLbliRbFOmF
moLbciv+2psVgzlVmDzX2HdJBTohpC6qEHBPGk2RVlrb9tESpmTQIyAJfMPJ9TEplzoKu8JKs9eM
lkLJkqtRx3uTE5KkQCZBy8Tld/MGEXK5ns5AisjuXaTmkNg4XPNmRY0QLVmBCR1vis4XjKuuD9kt
QhadF9XThihziqHq2nLjEmacB5ngjpL/ncNAyzw2eSQa0h5DN8hJaOq2wqg+6jcUs7yKhK8tQ5up
d8zGscoHKqrn+HhB1AG0X6PJD3R1o+pHoG5ELk4G7ydWNTC5jDH0KFrYIi9gzVsOVh5/7hMP1GXD
7FYhMVrwZRwvMU9ZII7PULRYQRdJqhNUBuUb9nGZ3H6e4wczuslxKwthaPFJ0jzTjNq3elD6fLlt
ZPJln/4qWhhTGMtwMkubu7s3SOM0uF5er167X6KyEplK26DhqzD5OocgAZD/DXck9rJZ+52f6aju
boBRfeQ9DQR4uInBqNgBIGTKuRsxjzWqpkyjDQQEzhkMnhh4hCdRxTpvGlZBokABjpxjoxVP24yX
BXUI6UEEp4+YlWe3G2Iod00Xau6D2zKUy8RagcNIK+PVKOX8igRhDTRL7Zh8uItTQ67J+0kI7CNV
Jy8YN7TbxSLBFQt6uqLMCyMbihMHKGaE7nuIj+vb180k5ReBTX6W5kTePYFQCFD4ajCa0fWIuaaD
a+C1L1Ay8hDmyQhDYECWYqGCMb98QCUIOqe6omGMKqJF/I+KAQDguwq3XaH20b4aCo5EYgVwPw71
tWHTRJ6OTl4WmP6WnrCPHxlgo6WBwAjCNF1rLC65VyyLmV3PS6A1i1ryjAl32Wx6kO2EGMo/XxE8
CjnXUSDgM/F3Mj7A/GUAElLVZ5hH6komiFE8BAVBn3preoMFF3H8Vel5FPMxz9Ldn6zpEcldcbAz
cFv6tBOUg6YP3idsyKxSZp4jzUXVUE2OR46Mwl8PwuxSCtTSkeR1NI/bQ0VTN9RLcMkuBxmj7OPc
U6CM0kOnS+XjlW8fOPULRMmSPoZaQmoKUXC5sUKK0c+efVlLB8uw+u42FDl0n52mPJbOh9TlsYZm
MluFIT2jVxNLFcw3RiwEpH/yR8YWNTSJ6B1s/CwRPd2+1Ee4PcskboF/YmqnRxe2A4ZNAxrxnBa7
cSCGFPi573lHyNr96zTMlskDRAGOShmDtOAehG2qptEKlry5jK8D9fEVxVggpe+Iw4tyVg/FRjd6
Vo4xNlHP0KReVc772rrBB8tZiY56PWH4DaCbJ1ICt0AgHWSfwH3LhAgycUJN3j3CaJqOF81fKObG
B0fzXHQblYbFuV+xaSBWFNTH9dVcXghpU40RjN7DSbPalpx5bG/3QWaaOJYcSS4Z6vtB1pEbMTNJ
IWHrJaqfsaMvqGqKTqOiM//TPZYxo2x8Z5Y0a6sTAGWpJNaMhHX1wa6M20X3KCI3FSPnvqMKhm6q
Ujo28KBXN4LVkb1oXC+ZHwy0xs2qXR9FukOLTJwmamZKez0Z8oMNihmbpY66OnUtJKt2co+7q/wu
+jScNwk4hp33dOpNOu+C8qSPboBC+fF7DGrR69PA0Rvb0WFGp+CBFwjZn3uHCFMwNS9Ym4EDMt9X
XGgxOSrfRni3OoRAUfwMcygFjMAsPqS4d6duhOWE5k4XHt/thDiRB3gdySUogBbieu+r5uVxqKg/
zrr39Mnn9ra2xC4KlhyIC02A5CZNki6UisLBBss6iv7luwFZomyyURcxNRggkJ7k+V//2kHZdXT0
5+zG+bAztYslhyjPlXCIGqs21k+WzigrJO9Nm8X4WmmJKEtnzNUwwJOuMy5dUD+hEKlbVkNuaRZF
Pfz4cR0b42Z2lsyCxYEQ06g265Ia29slJenQOoBHHsuq+Fv0l1d0D9+BOXkSrUHYdhKmvjdHjZHw
SmaDudrKQ7HLpuY7ewTb8XPIWwP49iZCGzlVHWW9g/GVFoOd8lSfZhONhurnPYkewNR1L+Rme4Tw
XsM5ZDDw6Nrhy2PGZKJgXt4gs+tIsBElsokgtVL0667c8Vr4X6Gia3A0ZEQz56Xdzh+OQ167ZRzh
CTpQRLHhwpbze3C6zXM/tL4DFP8+AicIcAAb3QymSdSFLu3KT/SPLNE7WyXEc3VTFxHWPt/fBYi+
bAnIsGMJzjXbaq2UAmhKyj/0K8BE40raT9sVLPZxjLgbgF4D6ijjT/RnjvcEPqt+otors/VRE4Se
iNuTz4yqRTgZr/WIT3lM8nO9X8fAMGxiMVE1vlc5ejbRXbCxEAzl2z4ZsC2PbJRyx66+ENg2Ne9f
j0zxALnqWaDnRCfd8R4MLOT8u6flkcWuYo1Wla8cIN0ra3edTlTI1LJgmOv4pYKG+FCqocDr4LVA
jcF9PAo52ViPYILXFLCWYAaC0AoktO9OBBq+a2rVXzWHuSk3VdA9a9XjNZidmiZIUjX19KBdleZ0
JtJq8VFMArxFmldT/DlqkLvhCwA687WqwEav6FDdz12Tcgxf5tijCxl8Ugixfb7M9l0mxdSm27k3
y1Pjuz5dN9YbO8/VgKZK5y4+YvlLE2bytKCsu2K3TFMW0Qx+yr+wbJyhSGe6UCuGfhmMelsQlBBd
3HTbxZc04KgLTrcKGBisZxmmeCoIBicDu5fbLokpY7+QqHDhA3SAhbltiD/croGPt85VkSJ3Rh3L
EtjnPHofIn4y5nc72D0SjUIkIp8fNmFQH7KV+G99c3omD9WXxYegmsa4CE1uUtRt4rBgWniaBE17
PI5r2AaMD8dc16jBbQk+WM4PH1M/OHTK6aF17+IFGIwAJLfngXuz5xcbpvbgxISwRm97YjrxeNaE
I+ep+DH2vyIOLkWvkzl38JHdYcsX2BtQxQTwuE3EBlCt5vDUmh2MOqOuYpi2fDFjHOsWQ9fHr1QD
DY8nTwk550kz/HSYkrZ9dHnQ1uKcF79R9VLGoaWvNTM26I4Enm+454/42szTASQgBUY34GBbC3IK
6dmiu7Z3JRWpeU0pFAreimiqH8sAzCeCGAl9/DiKjat1V0u8e/H/YYLZz6pMmXtSsjZtx1CkxM4v
fH6h4XZkYZn+FAeDB6LOd/7gVsrcN55JphlakIczbsU0k2tEfy3aF5Z6XF1UB0HXrlXOyBtnpIHE
7NhyxLtl1IPSn1bP8qRcEkUabZ1tt1DQcyPofVCv2hrDXo80x4BWfsc+MH1+NcnZowunGkkhsv2a
X40xURoOKsIXaiTKLiM1PZbSUMlvVvXR8fa2p3OoRkorvt1aW2yRrdcI5czvOqXa9ePr/wClhsct
H0sd+bTRSQQ8kplcv/59qgJMeMNzbmRBCcTtM6VAfahBT1rmvJ9MjJrcHSZUWO4DOspJbqHRn0AF
ZXgIfXA6+XyHfYoa23L0KwOG8AvbU6v3CqmxJxynI6aBPwFyvnishCLQu1gmBjn3J8LUHSvHDFWx
aa8pssb2jIh9fCKSFeYDn1aEwJc9eq2sq3q5/3z1dcSwaecPQW1bFO81abPgef5TsChtQZz50pSU
2b2mI0sB36rzwQcYDHxzK5oOY/5mgz6/0E1wK4AE1ksWBtuhn1kYCEBjkacQuXBYuAP0NozQnuAw
CmP54iOaScu1ObZNb0Qd+khI1R45xjl1lIU2RBG4lorzeKM6NV+qkHBG6lrg5socncJQCDjdis23
FTWLhnQp0sTHeoyq/DvzgSrCsC+FKxJJ2RWV6jQboxWx62h1mY2R2Zva5utelw2RZGxxaSTuABsq
GgIn61ujLYmatgzx3XRa4hZeiDdHM4T381CwJ+TdcD6i51LY5fZ18KV4qMMZjhVp3LYocQ2Wj2c4
NwHbUOi71PhK1C2IapY2lWf58yPTMsyVDOjyJo3tqJJIQJsdsmqwBXLivCQhLEFsZsic3Rhnebau
DA1TxYj9culIKsi8vYmaDhjDYOFOgkEtcr9xAaEN1fCLKJaSsAphsDrZyEmlP6tfglnhjO1EFUi/
rYzK5xqQeIIV1i/4v9CKrAqjIIc2TqBZaXEg+Tw1YqrR4v3qWIQLLYI9TttrWULXy58boiomLOMd
Jgu3ify8EuBlP0woQELp8DKgT/sHCnL+U0CiUiy6VMlA0gqZGO+L02ZpljdGS/YDQjFpZVrqSbJM
Fjd/BBt6LZqd4d0XVpAI5c/ZRzTbGjhD5ZwXcNp6kJeVLvDv6vYKumIq7ZvEl3xT/+pOBt3QRRRI
QaZmA0RRut66TacXTYn9rSxZHCk2iWM3gzJG8wC8g3FWDCn5q7dLOmCDxIw/MTCWZgQ2YN3u1xjj
LuPdXErrWo1icdcy0Pp/WjR9KAMXBUn7ep8glL6bjJxN74WNBDfNXiZCJKwwt3+bwvxWfVDMzVD5
60R1n3hCQgD36O0LxvU6aJA1y9iRg//L6lMASTrM/zJ0thIOXTNYD1NOJLfW0fcjmujNs/qWwD3j
VqzNlByRlIy7F+QQiCm8Cnz4qvgn2+gGSiBiijSmRGXvYUmFkQJ8YWdyZIzTtssbs8ouTmWlu8xg
CpHfCpZq32kfUhAGhWH8GwMnXHhGQsd/ZXBDIcZh3sF0COFtDWbzdCWisaRkGw1Uo7FFfHgAJ1hM
yQpUaawUgSt6fH6vhpmAsK8t0R9OEhBF96k0R9qtOpjDLGXPJhSEdZFHxQo48orTzNN5SFXomsHb
LiTTy27hwp3q/uvHkEVRdCK8qUa8d9HOjIV3P6GnYMjPpk9uw9VH+gLJRFZt8XfT0JkJ0CgpkDQG
qxe9YzS0x+xDgyl2Mr3CbrIEtD7md3yYTUBroOOPj2HOXT1kCEvJtuLPhZYkX8T3PoL1x1dsNjin
jT9sDniaxbfBa/fkpsterqVJfLBWdqCglxEpspIlNTyhzXR11cp1r3kn5y3A8l9g0OFP8OlHiNb5
hkRdDCbCZDCTdGOisclwbEjlCw2U3JWw5H/T9MuTnKAe9Q/vOKh8nDv78J3VA3rbSNC6hSsFCHkl
hjYesLhiqj/2r+HalwEfu5nP1SVncc5J9dyEl74bfbnYv56rk8WCn3diaxeoUjQEXftGyp/vnxym
S9ySBMnxwm8g0tW16EHAfYM924Yy/ElLLBYlGkkRyNbDaWs8X80YpC0E7jaVGZ1gfs+cCdcrVIiV
RNLUQSs2u7ELqpLQ2oZVJ1j4dbU6wXBmI04I46T29k4RBEO5zZ7DnqhyYvR3icF/y7S4eSsLY+qH
Xxf6+/ny9Bf7l64gV8ghyWcjkz5oNv0CyQ4R3AR9MfpJM/Z+CNE7Oqe00tN8IyKgA17nNttM0TOD
GHFP7x3vU/y36qcTtPtABUosFPO7emwiu36p9eoUoU8epUPHKg5Kcdfr3qc2Cdo++nMY/nBSD9He
rVWOug7+lS6GR8wHulpoKdd5WTdFI/Ojgoe/zFPxF6Vtq96lK1P4MsKZDGwsyHCFwlJunGtyWInz
zTXilYsKJj8YcS79217P9EEsgTcVlTGRjB+BKHlrMtB+skngr7VrUl7+U5IIWy8wvgpfyJm5PyLy
z0M1oeEBYT8ZdIuuLeotYjwULx3RF75salzJTiJJ/TTu5NETUBl5Oi2cG5+8QAbcDGqqrjwk8JR5
5GhPgC2+sMQXwR5NnYigbSbBHEGA6IHNf8G/0znX0vIlgp6H87OKpDOyTDIcP2OKIGViajOX6dbT
dTghOEE0f3aa5G1MqgBOqTYLonzGsa+5pM+Q5L8/GLSKVDL7D+fbqff7WR8eNU6O2+J2uMxTlH+M
qYbnRi5v6hZarMzZMyBMgaXTtCaadqvw14NtYPsG/up0W8EYYA8A1uZHik5qcPDv3WS+LTr/PSDS
tyXuiCc7uJVTHdDJkvMw7V41p3ZjNDMFAYHlouJlJQ4dT/98ABQF1fNcusigtqhWMMuGY3sxwFU4
cdH/SdabQOK2waUcH37sioMpayW0gWAVjmkc3+wBq9gHi3sdVRJEG5+daV4QCzTz1FrQk2j2pSJa
lQVyaVDWZm3f/Od3n6wgW1ZiWa1DRLJ7xStVX95Yx/o3IvlmtEdfoGAe6vUCBVcyKVQReRQ89IDH
XsXJq5qJIw44jVmwDRf7slokqA8duX6GQhr1BvXk8+5En3ho9Thz1TrO0yr6cS11s7sgwWow8ISo
mAUwGXJjBgbO3ZhPEJ3pD9I6PJtvvEbiVA9cqEcRYoDYRMRds+DH+cJpQzjnf0HfwAoNK0TVvqOv
/v3jVAmkX/mlTuIS5A/VY3AectttpP4JfuryFnKJp6qIADXUVbm5G6W0R+64GYRCn+fJ/kodY/EQ
C0TxSt5CSDfiv78sgxgf9/Zk/u/tpEYskBEhQWu9K+edc8h5kRbjUaPM1W1qdGQohNdAJqxFqwqY
9wUljr+tW/bOZZgg61EfUweIxTK0B25ZvzPcY75CjYtyi6g9i6iLPQ6a2pgFIymugS5Vo8taq8bV
lqq2VNVIRiGjpd5raK8gXOLXODE1DoRyFn0ciHD7iWiyQs9F2ZWmM0TTttyMnn9SMNJEWGM7FCFr
fYa1xG0nQIu4YHgPzUExnpRScaLLY8z3OsNQPgYKMmN7ysjILzssGMI4SJwkMPN5FfJT419dJeD8
kc37f+iQR7pdajHPeeEyfIP4Ttorq4YBMijZutmtA/iQXjdyhVL08Q5J/OtrUP4rwJBqn7ckiREg
qzx7Irr1OEaZ8G2Ds1s4nuYw0hZ6/B3/U41jWnM649yXwumCogh9NIjXVV2L+sZ7n1qA4mUq2Q9T
v67Z7FJFTBZa6XX5doSI7XTcxtt0GIITTM4WkwOUzN5UDUCnG5W2xOjP6DRCh/uJZ/r591nZmQ+B
MS5PJQPtkhntPjcYHBMujvnPTLEFtGMligD2xMtMmEfLOtnXwFWvu/ex8jwaA9peNyPalk4Fryly
apunGZFibqpxt56I4y3krGDMaQChMaAp+oMBZkXPg/M0dUzaqJumQ2HRCcnJhveXcPcnKcTy4hvS
he98x+44giKrH1jX59a/muUoXMJJjAFY9vCoie+ZpXJ1HopMzZVdTupGwYMYHwhqO5BIqvAmqEn8
dOX6JZxSLspACz00dUOhiwevAQHEVYYAxYS8XbNfUVGtkFZyCSWh5HJVndDosJHv0aCP/VkqI7uc
ShK/u/spQ73919o9/tmmk8Y44jyVNX/eJ2vxNv5EcS/CyMmA4UOoLdVw9axG8N41gSRQDm/h/ULU
sxpuglQPaIEp0Tlqz6Zo/sTEqkxqij/hS15x6NUxnBmSN/JHyn4HFJBzDW7Gf89DCjieV8Cf/uCW
Tz6zDLUhD1pUdiKXlUgD4iaQrExO3fSm5t39Ok3TqA9DntH6d5RMhl6aY1fNSHR387lIzIgKyIh+
cl/IS+ytgMfoO/bYyWmDHHQY2gCUAcG4FssqVwK93kitidLfKu1tDga3dlWISjB+Ae08wKkqj9Ei
6k/k/Q1FZ3i9/cZFV4Li/5ZVlcqNjp7ee7aDjAteDjcRMUS9rzoAkxV9mwVsFL/Gy5C3vUQnlghU
KX+7QlGxmutg95Jp20ipW5fd23pc4veCMRC3s9KSx71TrSAgLh9HKuK1ixlszT6orq+/hwxbqYDA
5vAMj3/nPY//30YgogN39LKgTMIEP4GZGYzgiDuMH54jXOWYHz5kMnnXeMPHWSOC8TgtbDKRxy63
G5RqiI8zp8d2jMEl7ArEgpWV3Zh3wNErqW3DbrPE5zkJFTY8AItqeE8HN7FAousWoDz4fu6t/Uke
x2pqo6nHPQBo9ZyUst2I0ctPxsnkNmJwUffSry+OYk0n4lwaOpJbibsX1cRcDuQQwzcqlG8BaHrG
NFEAf6jecA7YVWO9SaKxyMl+HKu7TP2wfjybq/ZheZnDtC7XQMvzUu/i/ESjLfJXJAEkKWj7U3FM
5n8IK1fC8PjzFxYvWOJvIVJ2jd7/uRtfviRAbk2S0Vq8kdiehwxWcERObax/dov0Wu36TTFi9KfE
y5qrqD51VfnCUbUbexOTatwrwQ5MSWGxwbVkTiX2BKxX/xH8razMaT7MI23WnurW0rEh86se4nTl
5wiRi/y6Kv76UXiEmBsaVvqyX4Lanrs8KC9PCFUNhNROKAjd2mHPKYAgF4LJ2GOajwi89rZhXb+I
WUnQeZHo0Tr/jfJFCZsmTWjTH9TKZkUuxkWtB6HjlvIOkpPsldBUFUe+M2uwgei+8tBk1iY2YGx1
ao9zYcJndlfWc3UZzTry37WeQzBd2ah2eNWM4gfWppJqDngRLOb6hfC4N3cTjeWROLnlMRpIOtVx
+ndDlFFQk5OcCYPEG3E7jNi0D7gdok8sMJ7WlahcPCgbyJvDG0ZQtiatzRrsmIhpN0tN/sapMmxK
pZ0Kwoe7XzMk620SSgX2SduCACDgS9fquO5woP6XDCEgD+iU4qt4zTjEm4rTOAusI15XUN+LKN6q
5seoWXDYsckau+OKgQ2LnmKTSM5GPzpCcE++KSvor1Z4C6K9aVVqbiCKiY7MZzHzN/daMGGlNcsT
N8A1lNa/1tG6DhWwOEpW6FzfFKxhKb05r5C2Mj3Npi6NJan0OEXy1qZcYzULIHkh7jKVY7R4mn27
ccoosHQ9n85o4ewCAIKwQ/lVXjjO4uL5J0DzmBfJ1BdZs3GeJa7llupwUpQtDwjZLPaENpbSKFul
bOzAsMFT7FaxtugGXCoZCFjmaZzobItZckM0QCLEHkyAFRvUVsf/tuHNxZn1jw4QbTh1SFW/ryr7
x9IHShgTsiJ68se4QLvQgMhQD+8tEZUmNuEW93PwE8HamZKfbMbpOPF3dBTJkGRrCnnWyii8ctRs
HCBZG542enKabvKrGBiAe+vpHSdk6Ra3z3sGr6fZ33VDDvb4ZYQ+kreEXJz1bOfS99kwihmtmvY8
Fvv7/IVJ5nXlw/GBToWmrCLhw+Ztjq7okaJtgCtvNjH4ImDY3IK1uAW5u+ULp6iRCUYBSHA2Jugm
0Cj4OYxwrd5m2ZFPaFGaOXH3IV1JVQQc9YC+aGrbeFfRIiLqIE4cZsbI7cOOl96LRS7SCUB1RB2R
Z6nZ41e70OOqcbwJ9oejacqcuU+xRykIWBCjrb1O3kLvA6UsvD2L6ATSAZI4GWv3Y4njsShtspIf
Lc2OwmG1gj6m3AbroucPUoKpthn1qIIMTUk1NhzzeqbAhViA8HhKUFm1zIBudX6RQn8mkSf8byc8
uzHTFmGXoV5iuk7xDO+MYERb1NvCt8OfxdgROOCxwybOZ7rUTxrHBz1LN2m1/bsqq/5uCt7mQ87F
FTvgC9AwVRIFaVhCGovrrehjhPvwv32tPOPjVJ/yDfUTzf5zDR8VxA2Lc4bbrlmdXSSWm3d2uLiQ
kb0xquTWwKp/FyJbge3ELXOr8Ddfeo3tsJM6+40dtAa4BvGU4UHbnAeCZY51/GWt8fOH6DDP0pQ7
DktephSQvs0E/oyQZ8cj34e2zpP3oq0PfQ933ujZNbKWiVGs+mfYJ8cr1tRYB4ig+dkwOn4pLN7+
VJ0buGyoaqs5HqqSScgWPaLYD3q/Ex+LHOVGNEGlRX8L7kjCZfNT+ZUrhooMT8HCwsaJiNIGzKJH
0bye1vzz8boMHbhrpFINDcfEvAZQ3lLylmQlI66+GwfjTau2YMRoQV/jW5qVMa/i2E9BWhZNXpvV
pe+VogOlfGhhhsnGSFVltPSmDNd0JaQVF23mNhhHo7PzoELmTeffOBdbsNvGBA5dz5Y6rPsSZtGb
fuLJgw0GUssNFlO3E1ORzsaEenau5jkP2dfrNninTg6EpSHR7xYxyzSZn4ZpT2EWFLAGVfyfZkHN
74n0gJrwATS5f/VEZxdbdsj2yQzRD2/5nWU7CMxQVinp13Q0qU7UAGLfG8jVC0Gtx9h3BQqsVsTg
3fp2G4RCHjSiR62evcn/QvF88smlhwyXTtaeEG38/+oTj3W0uC+AXgV/rgH/N2yhXVrypJFcgFmz
G5Rnd3gBwqUKT1tLDvZzg9eXSXkjmg+GtFIe7gq/9/LzwPwBJVwQisSzIi4aMiarwKyueT2x+6wE
wRZifobvhb+laTrmJHwMWkqcVH0g6FDfqvu+LMFnJtC18hdRRdlpplYcENYitfmKpsJ+FRJz+5np
raAhe83NbWxchgfgUVWl3tpvcFEeZj3drDV1hrlXz/lp5Z+VO6/ZtlAoyqLpNFUfM3uxok59VaX4
l4rIerHm5ud/9h5YfhTX7RafmoUgrFuqSqBQlLFTjDSijEH6lrgVgMWmAzUJcBx4nAGQ8b2vEs/r
nJIUXgiLSkoZRS7GqenQ76xd5Tcd/BLQVHhaFV3GVYBjKBUVFOC0BPK4mhTF45m5MDNysfzhl3k+
r6wa6PK6RF4RQJjGXH+k6z+e1QPQMTF24SpdjljVpZQyy22R7dGT1TNYeVJsKgjPBuCK7MXKQ3l3
RLa/XEta3umEMKVu5jFyV/GtLWqhCxdNcwZBhLnI6FrKnDeTjokv3p1a0oSqZK8YfL/ylCMjVqoC
lYcqHKz0DGoNUi5wQlBOLq1GMBr3l7GUNNRiDth5DEi3eFaGqy3uH5s7hX1LbMIGCkaxBLWfkj5Z
Kcx2nOnSzyNzzSa7UQysmsZiBl1Xw7QTJ16AAzu7NvBklduGoJgsrwTbkHYJd+h0Dig52GTeLqgC
4pYV680eQ2zAmR1BLnFAirJvJ/wdRES+8bQVfH2JqDvi7UWZHRNDgHihmzE67gLVBQWlLCxDR8qy
SNgdcw9liRS7y2CMRyo5aWU+bEjedmO5U/aAoGwCNly8gV64USacwasaSHcdIRKWZqm6ToKt4jZk
rXzUCEn0Cli9uryVtqTrWmO6XIrfpu5om2trLdN6hT9kHLIMWQXMGYEoTqHDT/G9ECsRdH2yGhgY
C9yDnJ9zA6jciJv/RFQu+QomyymRGvtxvn3gVD8JfZm/FkJke2ZlhA710b5sJJs3yco/CP8Tz3ta
WXknGyegmskC4JB+BAdypW7qwtVV1/Zps/ZThKCZQHogK/62h34lG23IpY8rwtq5XA8u2dMV319u
mYb894gh/+vApVMlYcrVnkzAEY5DfwewHfHODP0X5M3b1LBW8g3OlkxV55spW71VA6g6DCYfU/jt
AyXSh9mMkMVdXpVhg8dzP2aPGtlFLOGuT7zC2j/cBxsFc39bePDoV62POYAyUAy2EbV/dycBPBKW
Mg6wFvNStO0EVjLIA9IPK22wyzsscFmuNjcOwguWTe5RUZbj+BHEGIXdjUfQE5P6NwDqH3UqFZaz
msS5W4OjVPYCslYv44H/OkvchCPwyf+OVVzkOgi7ILeQ3vLDc9MASYPfMQvslxnWVlXYP0WqAfjy
g0Ok4uOqn0OgagF5uIuqqzCM1tzbsbr9W2wfxbgMVgpdzwqG2JLMhyHwnWQmOSEdgixe2KDcCE3Q
rTF+14507KFPadCs92O3hwhnZbZyeF3MDuH872xwfbZU6Vo1KGxOFO+VJfWQUYw4bf4JPKBNK+ib
yNpoC3E48a886Um4W3UnVXJj6AdyNEQLVfwgI9TUla0RzMBfilK7zGob4zMEPg6x7Dl9hZMsYMUf
AI+YVOtZKgZEdheGDMsESR2sKu6RqwNYlYRbQy1t8bZxwCUWZI0CPkaC9dhDbW5ITbnewEmPFqXE
uW88t/9b9cl1joPdtFraVQdQG3unTQcOcFCblCRF9sEZBBpmQzFedBFFXvq7tyFv1XOL8iSf+k0T
gNAf0NCZXCOwG8lXCKdhhM23G13+pam/qcfz/IdoTWGFHg4mN4Qhno0xeyQM2EZy3aPHSjJB7gvg
7oQnnPpA5IYNMY7sBAEP8sQHpl84jXf+M1x+hlCqMLssRIA7TLebRIhAr5y5xRWavh7sf5FfwSzk
8HasBheMZsibMGsrcJlCZxeWnDh6pIn8tdwzsa+THRiMB6u+xRq0b08dUnLA1r8EoGHTezegctgg
cXzKhllqOuAOe6XI6ZYde1cZI0x4PQ1xpjhh/FT6zmRFUGl1ZS3Q7msoXzDxZupugcFpC1toZGBj
wZKVyNrycmg/S537a8Mu9KXUxcCqZqia7fmbHUwj/EOO7BcZ8lwVbCR7IGJbJemB/A2oaSl7cAg0
gAEDASocAFIAFTIjjMVawG7M8vespXa9fTFBrsis26qS71bIIxRZNgREfA7yA/tUiM/KHWMkxu+N
JM1rLx3uf6EZEOGOCVWkNfBiu3Ngr7OahAdSTYsjUbE9E8IUSsTphVdB5Y0IC5R6Z5elPvxch/GT
vBcC+TSJyTHMYVSjNoNOU0JkyWL02RDl97oK/zRtmEclCF8doMSamkSFBhWPBPSWWHWCkyYTM/2d
GD3rbUtbA6onbsKf5lfeFho6FWC2Ipk2npaT8SbuI6rh6NGO4WIj57bB215jjYiIiMMeVIJPeLgg
tM4VwjpEhRmapDRVbldhXFilWBVmdNz1+MZxvINUeup98/IKzjL/OPve9GQBDx1LrhpZwNk17ANU
fiFKA4uIUy1U4yEyT3tuxvjMfhJpB6PeIUK7mQHCsYyB0u8sc59QLey9gEj47ah543ENTI0TZEf+
pjepOuEi7OjxXYzWFvnYFWXGPtmkltzrJ4BYD9u6bAQq4L5zdJFm8sYDnk5qDxuv10c/4JtgQHRd
X5ELdoPJKvogOq82pxdLr+jpwcMLLzXUyV7/yXk3Pr0x8Q4ZP58cfOSaxQZnnA/2S3F5WpOKNlbF
J78krovhQkDDbjlPK3O++5j+jlOtnudYIWd1JkcLqC8DC9Hk5VYwfZW1Jp0BR2zpd5GxIg40uRFr
Bw1vyIS6w+0SGN21yRc9j5J9vlyI+s5+LMI3U5fF9wlusOS+fZbvfv5ms8l1KGTqe0g/z8R0AVnf
png3nJpX3+UOEc41MpJxSg9WFe0HS7u6MmXBkYZcwJD8bwsLgq5hioa3RWqgBMwbNbiELgrY7j78
oB/2YqBS/P67Om8Oo/1h6N7gs/2NduCY8PrBH1fmciKU2xy6772FRsDCbe84/P7VjIUyIVFTI8EY
SFZDWpvzxB+PrX6wnKDCbHUHKbdgkYWE7b7n/q0JLZpUPSxtH9NdKC2vx2dCjNWVqvNRjGfqjjTv
5oZ9s4plpPAJcAE2557tbxh51TPNq9F9sJtZ7/VdLq5WHeW0k8w25yCtD0BZc/a5G3AV8El1vlT6
SMuoBAqgc/kQVaovzFLlYZ1FsICepEDYlh8d91rbT37ZxSN1e0UmrZw0T0Vh1CqmH1EhVgx13XYB
XnuXbjLp5tLKiiWksHkcT/gArT3e3N4lzMMqTGmuaUTEoYPIh+iVWkUPhKEzlH1YJcUA45J5AkFJ
Rw3tbJJMPbwaxfoFbxG+qxVlykAV/Aro8kurZNj+QJRvQv3+1bvHmYHjzMn8ERKwICUb/3XNdQLt
q/iCPH3uTneY2pdpe42nFwj+CdanWCwgStWyTJ3n/Ath/1t7MRjB8TI8GrUPqVXEX7KwK7XxGtSD
TTpNVt4kyNIziGbPR3wE4zoovpApFL76NzRPIQWG5v81lLTdNZz8Z6rMnggh49wgdSUcdAeBL6QB
ZaD1hwDmBkhoxuPFQQj0mDPtya6KW/j8S1KzL8pSv+KvRig82bX2mXyBvgbC+6FpQmLrhHRlJTRA
nHbVsgCTqXdcYfoaOAz9fza2vgZZ/wmlZJvydg6SpFPSzJmK5iCLLDvmg/jwBzWB4ikhsTTYQrPB
y6GjAgYJmlaA5+afaYP6zpQFU6YZsqUWJgmv2owrW3YZBRpmxsm5MrQVM+MO2b2I5fsvd4ncZUDS
7r5SEzviSz/LfXy+YX4n+rCX7K8zvzvPPnRlyr21/iplQAZTAI2ACqOABkaCJtgt09oFbJpOSHrr
yS9GaWmnrm4b6zT/QdJAhgO56qP5uUYJzZYcfJhkhu91HneNDTdnVL3H9F6DXF/JItu/lP/vja71
Ucw471j4Q3XEtcfHqEJ/Woc88AlXRD9jonRoxOkJEYxW4cNwbtDKTRcAc8Mkyi4QKWsvVBL5DQ6A
BKBv75jBwjTYDDbE2KoJtLMRoib7P0kKUUrwmPODXrzo+R2v/pajdEfZCIRdYlizreMtRfqv4Uvu
Ie1QEcLToDMwW4/wWDNAF1GjeJ14fO3pyNhACJO2d3cIyIyB1mc/cMWBLUG1J6Rcq4UIkhYZQ15e
WpJA1gebG8YgR+bmRg00ytK/i1YpSSa4w/lj/YgLjubKvU4Ptv3+os0ux7oDZKelx5wbio0Gv2Sh
0i2ivQAWrdFfaMIpLps66yLrwj5jgQMvwUmgVDqR7K6Rd2eVADvp8ivoisnvDdJkHhRdBr8bgVaf
lDwhbQEXDrMfF1r2KXaDeCwQzwHQTUma3rDZcfeLKIg/SoY7OweRXeZ7P6lY0Sd+vIRxAzacq7RE
JsjJVNQbP0piIs3OqGL+Sob+H7+rZcFGDBh3OB6hv/KoK7ukRp8ddmMptojNZ9fkgk20ITFt5xfr
y+2k34a7HJU4+vySxaIJdcUOcF9QLcz/+WUlevrFWAap1a3LwuIWEXRyuj9+K2giQX4IoQGS0DE5
/U+qHVvGuSsBF3Gm9+ojgWkzxMk/PAdA2PCLbM+BONlsEtVRlgifvTxLitxWvfNNND/3HUoupoVK
iBebazIdfvE5KYg/Xg1rx6Gtgpu98H4LOLvFpkWtviPfbBsxZPIPmzeaNh/zgibE5jV4RQ5aTkbb
VXSbt6HLzOCWMqdO0yc78xtMK1GNJB2ZtiYx7QBtz1EJAF19AQSPkSkPW1voygtRGqMY+6/A+oQV
gsKAKDUwGB6JkiWwkf1hgZU2N1u6EG0hVKlpiBMCgYNb1vWiSShKFV9yWMb5OEFAeClnEsKxz8OJ
JyATiKj4xb+twGIOdotvviSC1X3cqGDW9m0r3Mo6XrH8/jYoeSn6lCdbNRl8bxx8XuTy6I5Uh3s2
2RlpyjIOHo51vsqA2Zaic8XxUfutxMQ7TbhzsfggRS1TtapG/3j2H0ZZOqOMX8uUAE4/H/B+8RcI
6+3RhNC1EslEqy68BAcAq9tPQY2v+gU6Yd8PEGi36rrnnmHqT/leFywFkL6XdYrc9bMqjIJjkou6
W3ix88uvYYpSS41gX5EUqRWB9IeUU8vyg7QeGlDnLL34WKOA4eUIOXx/DNl1VO/e/61cVtPPhsIe
xPv8FK8a2X5D1LHL8Ssv6kMXPSbG8WeEpMm/lYfhATfoQzVVmjlNA1oUA4WOVsIdTDc1UIwLScEZ
lMVFQHNTNd1wMmTOpLV2iJcDstkyjJUKA9dNyY9iVAWi0+UiJ1PVw5at522NVvdHXEZ72pbLJv/i
laLAvUGWwCRMffjW7SCgxCLoP28PwCymIy1tTkOIecVOYgq7wM61T6Y3/NCNihVg1WPrByzK/itx
rPUNdOozXqyyDK6l170Gj845B4G07i35eR3sEbmefAb0NIbX1A16kYpSL4YDfDBwuu0ArR+lEClB
+QHBpHM2ei01t903yTCkpzFUzgqs8RL71AMrGOPQmKERzsL060TDmjsuvH/WKQFQoZI5iC4vFvyO
bBrt+BUjBJyifdOLHYdkYmPgvEGPo0a8T7nbaPxmRFKctxVD+kc2HC6MAy9h7fS81uyKKa+SDAm5
X84WE94REvvqOQ6h7Yp1g4nc7I/8PrvOt1oW8HEhF3Nk5cbHsPAV9JEyrXlHKcQUMegwCEKBmYdE
H9WKt7DpS4N/rCtneuH/Lk61aYzZUC34SPvI0e/OKThgGqwEfpkrJ6E9NUsDskzaVmvFw+sZ67gr
QLYRJ1btjbl2VsF1LlnNLlnUhutR8O+8gPbn3S+FQYCcHF73A+Z+NeAJL4RriQqqB2wXsD0B47h3
fSBV0NQxOzoL6mg5Y3DWjTuYpN2Dbjn4mjrIkd/dz5GFWBX3w1vXDJn9elR/I+0q7Zn08xhjEAth
EYlhfUzY7hVtu1FyPA2OE+JFKLQP371ZBJCbKOGSegHzkOXehns41fLYk3xbei0yHpsrYHKHT3SM
vo4q6oslalXJI0ruR6+tfDQOecZqVnzxfj8k+nq8e1wqPOJGCHzDxOgAS3/HHz1QpSTR92P7z2gR
jnID5YjjTb73WmhGsLE+zi8nKlsQCgVpVK/H50VPXP/A1lkZDMF0bBJbrrHxhVD/srzVRH4Hi1Yq
7z+heSSPgHq3vhTYuH5/Q2PVYymR4q5V7Jw6skQCmIaXRV4BeZJtf5u+Cjsm3py3fk8aV2tCW2Qk
GttrYpWgfHvr4bJTFy3dUSyFeT3lQjCmIDZoYMIgeskx8lgQBzFjZrvVoYNjIgvbec5mPme2BtN2
weWmNDQIoHxZy1ozar/NxN4sG8P2zBn2U/OYOoTVaAAL0JSH/DCKL1ea6+IxePIoMdbqaIwfelr/
kRQ1QimzGtpKAgAqr9JEO2Gk10VwAwI9/SDhBdvubISJwC7sM4cJoLwrQjdsJeiiy4VfC+joYINO
aAVJBrR+IM54mXnYxixvRCk6gBaxgD9dGukL/T4PgLuoEu/I2U+uwG0c2tbSfJT36xrOV92VewY8
iJ4W/G24vKKBID8PmjjcwYF0/oxRLAcEIOk18YHBgBY0ihaUJBMGaFF2U3MRXtOich+HDUG7Mvyd
Jv43Tr/HP5yLsXkf2zFRKE8oAJ8ZXylqRCr6gp4tfX0NbZ0si5kBRgEuIZZYRTzbyyY9g5TIqddm
FQSkN+9uYtz9We1Z2j/37DZqsvgWQegzrjeaziEidb59cSJDeLdUsJ1gD7nHdmU7cZqSNYcFhliR
EkykDWtABZ9LI7y5dq226IAa+CysbWwB/og9bq0IIYUJy8bodkmaoy1ejzeM67Rc5ntC9geYgcIz
kQWE9ECh4FlIRw+XfZtaSShVHU92veutvqQFqfVlUijp02aPW8U4lNTtJny+eSMizV2jnO56iRCU
ufzOIoJTJvgSlH4BHwiwJRYJm4Ozcr/mWL0EbM8dBTpzw5qzBaQUuVIHopaHSpHI9NQs2GWxl6TF
IgbiM6UiJTRRs7LTqpoCyUsjfa3YMBI7FlPbou7u/UhJF/VrGzfKVG7OmMnXhALJ9kJC739fMGAy
Fl6c4q6h9BPrPQHH6wHau9Ix2Gv6IMx2DEEFwKlfbWULTv8H/tbYwkkFZ0WTt8Qo/ZlaZm9b36C9
f6WXKxvB7cKahOU/fotrncY38czp4ASRXxrt//e+KPizowoObDZoc8GiO0XprGb5uDi3ZbUAxQeE
1yt65KHoXU1LGPYSq2wkRenH6zRyN5n825uyuiyLQ/JHqmDe1DWesUYJfsDhjc2BWWqNMGhiBSHM
+33rBiw4h7IoKf+xGumjq9wvKxdqP+qTrVLLxJ1btkXpQ/a9/1v7os8Z1bnuCBhwnLjw82lF1e/E
YLKVNHU9Q8898mBzfb6wIA+seMa0lHmKQ2pCzU/aZv3rgSnPQdss7L3ERIxseinWKlE8F+WhAMPT
C8ubN7+cfsBUBta6OXusn4eXhTwM3DRHjRf2F76iGcDy+QbgInimnj9RQmF1IjCVy651QidV1xqM
lPZSCLWh0wx6+it6p27unKyDInBjAOI9/kNl75o98PQPBocBQQzrXGFzSmXk71EdhTskb8kd1xiT
McJXVJfGk1enDcHUM3AWf5LAvkx3CDOcQ+6dw+zmoDt3FD0UKbsbqNuHj/QqNFCMZB0KTGYuDskN
OBOLKEShdmZgwJ0UBb8Wji+PeXH8qh0H551DTs77H1UntCoLa+H8LOqtnLf7CAUrWHGtGwzgSwgP
pORttqlsA7xoGZIjcE5fWLvCE1Gf0JZXB5+9CnRZI9fi1Vp2VXsH/DJkgu+TpNJrOWlyzP58Fhul
9gIuqoSyGJGo6rbzC9n0wbbCXwgasDCymS2TBOriM28HbyfI+e8jlNN8xPnG9hX4AA4GCWuCOTvv
4Fr2vKNUiw3NFJfw5q0DMkpVpFgA3H/EYGz2Y24r9DCyzOYqlixmwvLjz4nh193eZZuwiHwl2qPH
3sXuANGS403AugimjtlaGJTOnt3+/Lr3OD7A3Q8GsLd/Lg4XHBTjd9W/8vQbmtTZT7jf8K5ZTTbz
NeXyoSmvM+NklEsjk6PVAtJ7uGO6/goRcd4l2HoJJvXA9gQMkw14Y3Ue5GFCcC+U/DnucaT+8ArU
58/muWUKqZ9lhHBJLKNyGGh8oyfshenl83JsKQvEhoxu0ggZauhdOEisTy01kg4lNnUOqBdFXe3e
I8Z8q3B1ArVr39A9c9LY5aPsgdSrj1g9Lqcr5upGwHokTI6Y8WVIXYUn9HP1z56Uz8FHcS3P69kJ
ioMelWO7R0pYKjAXpf07zqz8baj/I/sRyfivsZ/+1OuaVARgm4/qLJ0u0ku/GdXSENYmaEevihvJ
RCzc8yNVSuiyx+RrfeaiDN1rQsJ7JvZhDBXgFVddLr2rSuHIlcox3vkq6QonVTq6a4v5KEl86k9t
74GfeyxxtmiT9aNLKDwVVooq3Zeqod2rdqyqJQsO6MO9alW/jl04gcLVXPOOTuZKUiR60dUfjRha
I+0dNrAUaibgrqaKL06wWagBB7t3Hf5uJj4JXGfKQyUleRvlXz1FthP/SALNeKTo3vo21ErI00Y+
C6NfmZWpVngXg2W9NW0Ynwp3u9kMmlXtkgy+opFJsTFnC4e1fAAHJ1BtieJVE8ZQNLOc4sGlBgcn
O4N0/g/30/QFEIpZxkFriz4erwMrAZXuxPAFV8uACwKA5qM+NH18yzQN7Z8V/Auj09i1u4kvWE0r
hmoni0fr0JWq8uozIwkPeUsHjrRrfWonC9OJr0sM0b2tdle1fa+nTvo90oTsK7L9VzYIivJFzn17
XkM8COKy6BkIM3GSOim17KdcmdYTC5tRbIo7AFt2SQ0Yx7KbJ8ecYQXFJngHMuI17yui+kk7LwOJ
9WQCnutiUmipXuQfdEl0OaQC9poHNXUKXI2yQ0rkzcb85/EnWGNhuQuf4lLZ3Hy9GoQ+JHDjyEFA
etnwEj5s9IJWZYF2SWloraL5em+jjcpPULVlCr7Gd0yEYlZ9OjoT1u/U3w4EbWlpJV3BiFcvBYDL
3AfFiPfHxjKRH6cvaTX4MA459pEuzVG4pZ2lYkXudGI4w7LRS6qwefAuVWJCV21I3Msx2vj1YTUd
1AFZpNx2VzZ0Ad2vVmyTlkhiHJjTxS3cmgs2Cy0/OltQqAi1bLMlWD8KBxVUSKnOqEjSkxTY94Fd
bJcE4SZLEAQHF4HUpY+GcfafgEqpC/Q5ehkw44Mvivd69dEm0Saw1TzLxBEGHg5nLNySLWO3b0Nv
dBYs9ZxAUn6hUvMAjdAKxydmPDqWG0qS+65yjTBNMHLJGd1uqhpUurhKBn1sy2xKfJZRN+VsQQ+R
sz+hONWaOtzR5eAfPvSS12imC+YoylERHveYXjF9HOqEDc6y8Q4OTADQ6we1I8qsrwskdIT3+G7d
ber9hG1Nz+fG5zEfEzEpgT73GzmTK3S5ytjEe2GAO1Ge3G4ugtth9a25PYRnF8H8Xm7/MoVDzZN5
eXEsNkkgJYAT1yy/6ETpUSDCOHkCvyWfbO2qzCxxz1lIeZf02HEf8K9yvy09KubIkWrewrjPOuZd
tXkKm1PnzyQ7f/eygBN7rWMJlxodsA5Lw7iD3xOWVAsG4btcNPr9YtM484BJ2yRZuwtRy6bE8bRJ
GocTV+afqSytEnOSKIQxvMnJ5BeLLylghlwFaVNaQdKj0dZMMYiBKiwwcn2Au80uz/Ofq3GVR2Uq
zFwAIGFNTJhhMAoLQ1ALnsUTfkuVtKnu0fv46fUhkLV9VkIiEBB8FM2lB3AIawQJKhjfMSF0Q5Nl
bKpd4X/jY8+n1Bs5RmtWkLQcGpfTl2kfG0oOInb4JtirUoOsitx2BmvkxLOcffUsxiJ6eux19o9f
WRWPATq7JgU6mfLf8Cx4oRTJBd9uL+GaTB67Ph3iOctQd+7F+RMFvQgPU+TDd9WucQdg19Qww5aC
uKWeaTkY+9+GORmOHFZ1pUPgf/b1m0MsDlv/UHzCQTX3Rv5NBRosbMvlO4oZ3lqc3H5yAHucd4tk
Sn+KYAyoh6rfbJqBnBH2kjaTJvwJ60TdzTyuTvVn394MyhGAT5OGwpUap9XyVfWW1PAIZiknGXI8
renNHgby4pAZjRwTCggGHzZ4WohrjhAigcRo6UKu4IEYQope+Ct9+QfpV7GwKXPXyJIB2qDW3xBd
ncWyEPzr4S/W2J189mMyBkg9vQhLSxTIeGYMpSUvh+1UkI0urOziYxorvHAf4nLE5gj/8M58eyvq
QgQDpwlekEhS4p1Rz+pnoSQ3x5rirjkbvd7KIsTfjbI8NGFr3L9ULEg30kIM6erKjR6fTuDbhuDM
PzbhxZzVo9xFZgtTn6v9bGdPuVC1tBAwO+SXDLN4Y/++C+hp3DlD+EH0SUwo4Dla8mImM8TQPdGf
Itz+RjYVlXpWnpCWOs2rgpav9v10e2NWbrBWX+ENpKsXELEPtmkUYApqepaent9qV2FyRhNjkRNY
sXlx6mwBoVNqBM/sf6MNsDxcPQlJab61bHFbNg/6OEf3GTqMTrgAJWQ+BEKzh+CRVCgkGSCePvIA
6Oec8M9mD1J8Wl6rkDhXr65m+Mo/xywQqn2sU6zr51osWM5jdcuIHcELRau9yQhvot3MfjhdmIDj
5iMY2NXStyd+mntiFg/S1q5AGKncuQxdLLIUllAFd5LgVIKkq8bR3KLTvOh9B7iaAzkAWdHGxkxg
UTb56lhYx62pJE94r03MzmXJukhbQ/uAto+Gqp2bd5D1W3KU/Km4zmr97ZETsWf+Ik/bS5ugi4eM
RPhiiUtAy/VOJ2Y91o8nQodDD23uU18+1lmrH8f2faiN/w2+BDIJUpKOXiL9KtsvhKo46tjtgjn1
cBy57ECrEBgcFKeoRsTBw5NHqX3XXmRZrSCKI5Dg4ANKHjFkXwJty74YgACjLSlWBX7hhIvkBp03
Dao+iVWxIOIPdBQEJhOoFLolR9nWy6b3j8q9ZUihxUXbeSyMz8BUnLrJac7V7FEB0rsRm+TkaOcZ
UwETkLy/hKhz4WrU3WBXn9CMWtKY6llr6nrEo5PuHXDnrKEtzYAwvwNs2MngwqhyG/dA/kX2hr60
CJjP0jkFlHMjMTlfLNfe3gJC0xxepF9sn745PYip8Y0AIXdyVCCIhTaGGn26vfJJw/Z7Feq//2yg
T7PVXpg9QkpteV678Gfh+eDBemVpfEuRZYmXqvjTTiqmsm2hqx6YyXUPiTe1mrR9x5g6PzgKU+SG
hD8fp9QWDaa1Lhc4HkgnOXz1XeG2Bk/cJjT4+syrN5lOI8T7W3fmTRglGWOYyttTOlPMfagCEjyt
qTNSzxLxtv6WpVsK6mXRNt9G0s/FRVZnBmNiCq/373nCbCeCyRvcrEz83jqM4oeBCj7U3CGbLzzj
VSEhwuTZuV3enX8QUTBQppqbpUfnwSN6iYJ0DjTMGlik7MTG2n+NzzMZ7FtZgbcz7SHvl5CYrgXy
WIVLUT61IjdLGYypta6tZbNitj9TOQsP4+XEbDeOuBz5Tsr+fKfIY8VflAfUdYcgp7D1ApjnF9nh
TcjdFmZQigJg8JBVtkELs2JpY85FpBaqqTD7mOLzNlA5QpB79YDD5YMQ12GNqvLhTn0haAutvnAM
8gxAiJHR65xrmhHIZK6lh18wDXwy/HpXmnX7zxLZ2Cr7klUxMTuBhuH86I0kElhy0VRhrDbsWDbB
a04/BjuzMI6PszUr/sDylJMrei2NnHeu0SZgtEOieTm0GOSkyvmynq8wEIUTdd1cvUHVT+M0P84e
kiU0ecawJmViZ47e1IM1ZW8J0ov+I/5Oa+0+L0BtWzvAjxpZayxhnkqb7gZAXgJil1YSd65Q1fMT
ChgpGKJ2TIgqVSQUsjlH0FdF4D8EKQxeMJksGrhicX8JWVfCs9YTidSGi14tM87Q5ix6SsTT7oz7
GSTBjjdAx51kwCnJF8xpjvDNnMMKx1byZ8swnKoGgYtFBgF+ijlKELHszELxQZBda2X7C91nuw+p
qK2iu3h5/aJuZqXhN5Rjev104fmo7UTe93JqJtogjP1VDvl8pL53CPT7NUTaa0xH3aEWMcBr0oO4
8XJupTArLE5fwDMkYvYS8PwzoqtLrGdiABJl3VbIsQO8+3/q6kFOG/al4ih5b4fkviy52pKuhHjL
Z6b4SjMRb6ZiGhHFuAuhMjuXXuVdpXPVKNBrdDrfoXhKXJgBxxLM8S3Emsp8mtxp++wCq+IjoOHc
2U7NdwmAMwamKTWxrfxWOfoa3fKvumUWV/X7FsUOvMVtTBMXquW+YITxxgK/3ShQwgZKKgq+yEnC
5InSa7bqjX30XR1BGHFTwXZXMZtTq2xhrZxwv1/1ThF5faKBB6NYc3e7ZaNbdP2amIF7ndhfKF9d
YUaZ9bgUcjzmg6wWAjPl8NrhRpYcA+raUMezGQreqqb+Bte7s8EccTDZTccsThDEPJFcmEhdsesE
Fitxl0tz6n/UtX1cCSdbRrL4F2vlKwPzT9QGX8YSq+Qz8wasPBQI5nWvR0VRgzdr/MOnEjQANOLR
OFsKRv6EMTpMMmtv514VC4SwDQMgIYv8b/UqtijQD4k2TPTGBn0h3QuRf9cCI300gl8wKMOXWu3P
r+mMTcZsp6J3q8tCPaJOTNzGLDRKcSqpIt8e7ax3+iVQhG2xvZIwTBMZv6SKf7tpWBLCpnHnace7
+oYLmsyG7+p/iPRMUtcES34/Vf8TrY7Oq+UPdSpuj26LUxwyuZuYvBuIeOVCweznaTSVuyx3e3b8
Hjo5W8ggY/JrMatC9E523AwX+gj9lYs8pFf8rcObPZVYCzwzZZS3mDuyFzarxvMid+KmdVUMzY2/
UAIRENcG5xVS1xOYvwsVY2g0nTGIM1CFxMgw63QpYeLAdl3iL9wkp2+MU+uzpF5hj6CNmdx59Xjc
dzxAUQlwWRZw5caGwbowQ9uIgZhzgRiCaFrIPp6qfvyGCX0viFCMnLNudi/txzFUIBjBSsJogO8f
XFMXDPn8S9UfCJR6AAa91FRHVz3+fEeoPskQQd1rl/c3UyMTgxYtNTCz4K6PSe0Us9q+S426ZVjx
mBFA8lW2DnPnIMR7DteO2MSeM80qFpwk4ySiifdc4ykmXOwqaueq7dBld1eJcSz2H164FAHPWaXP
KmYl6UuZAn915HS41P4EQKrCfAs0ZJhh/9nObUGYdF8nq6Ainrl73t3PQ8GQjhfMxAYf8LiKDDId
M0H94tilppSrSa5Y2C8B0iWLidUSEu5rok3gyhfJghYu017D5VpYI0l0IsEseWX35TnkNRtGZFgW
Peb9EU7Txu+cQaP0PZWubAz5zLli5lqt83DzmHSyE6U834vrjTCJceohTCarb1jtI0cGzjcZZU4l
o1WNNzcz0XYUTjQ1rPDFQRYbOjhlML32EPWXIBh4XPAyNXf1VeNCDg8+BDCFNb+VxTYNqtQTIzOd
7A7RFAl9clTB//PxKumYwCJTEXRGe+nyTYwBo45PC/QgSl4bf/Ft6SzswSm7BXb5pzFXys3Yy7r3
81mkkjxWJkEn/mFMXvn8cJ8lcDZzkRcxfKZwDl6vKEVXoutacYVafQV1ORMw1/OvfuFf56N1wnx7
iD3uKKPDz4V9jw7q1BaOWuCB3p/Cmf9dGK4PxjjYe2DGs/XMO0y1ut/ZDXxvvBIFyKAqKA2cPz4p
Rbfg5gYzGJkD/j5rV0Q1/j02WvQtUXQRs/+NHskGHMHdC+EfNnRBvc1Y0ZxqA3sLOoCHt815G+A5
IwjUX7G/B9TVEyQv0jytRYxQCssGQXaFnT7Gz2B3V0V3p/25F0cKCKUgbbas4ZeHKpq1YiHaON2E
WI1LsEfm6VUg1uUSwh8c3M/Ao+2LQQ8XlDecHl26UndAfDXe+TZQ8r2UkYYEv7ka/1hx5bFX1w8R
QGqOJKCSAZOJLyr8qi4o7Sx/rj73FNw8DzwNSjzw5M+57dZ/n+gQpeOaO1XajxAxvFLJmDlKttgx
OIYnxRCl3R0lZc8ErUlQojSwZlhj313kb1anSMAKEL2iBrYhjJy/tlEdaOe3YpNMJImO1O2JN/hp
Wjs+a1NLa0NNHhXMFmTiqPi1xXqEayNBi2YeU2Rzex7tpN5pDbFg7iRsfhu3OM9+yqIkqk0cJOaW
Jnb9b4rghxA9dX0OdvjYQKpWL2dAph2ouUf8f766auhgnu/ACUQHSgYuskmh9O7QahBi0fQirWD6
o8nnkNcO6AEcg8gm1RZ2IzP2gvT9Zyr3eDbWmSXydjpSilR/qWvd3+VrYYzReiVZyfoGq4Tzbina
wfYNllIsCqxhy4Zd+ZO7mISf/Me5
`protect end_protected
