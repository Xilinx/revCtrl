`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43328)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAMJI7Wddo63tya2Pu8fbyFW3PSexWbEycAV7UoDuXZGyxHBgasA/bK6J
fOmk7MCD7mZYjez4D1lapkB0Ko9EQaJSiJ3ICr1XCxhZqHdR0eO6Nt5dfJd8gg3qoAfGNihc2VLJ
3cz5vizDo+C1vdJrghG7pPKn96DNfL5kIfbqwEgzTcN6Iz0aIV3wTsZr8u8KdrpoqavLNzdgW6M0
lqdnDcxizApJroVC+gxce0FVFnwhSJ3ikp7MgW8NepER8LmtI3LEOA4vWcjOQVGRfkWOAuXJYmFO
WgGGO7vC/UnGZ+UXqszUJBjGy3zRsizg25wvSagEFzjioID22alxnqi9X4kt+ZtFFJzL1UDsaFvw
orhorbVJurAEgGDYkh1ynhjqdSctrUZxhlzjfw5YLDkULACLs5RK4k2Nc1an6IJ/LdX1ENHQ3r+J
HHXXyGIcHXyhU2X/6v2Dp3dBQIy9sJUT1m6t/vuIFPEvHON4h1okYD1GSDMJCnqvp4Aly+X3MXS4
Oz/6KEhxfWceyonJZInnR+Fc0UAIsIdgZamib7zteqm4Wxh7/nYSsLl4DEdLlA8T4rwAbpCw8Eo0
tXPqvuMeUNvJW+ZgrNckOqYWS3b3+5zaLnzmfCymCSh3IWiBi9LmLwP1F0AqhXF8dBT8bHK9KKWE
0I2fRyrlhYZTSZsbWr0SDZJaHCOfY6aL30ccVGMtZ/4et8x06p6jMwb+0+zuITdp3BWE5Np7ukGE
oe34cdgJOjdmVkn0s7qJeMAUHJ/U3fn8QQg5Xcki/GHWUboXuKjpl53lz5wGK0FQbP0Fm1vGuw0/
7rDzhK3c4W/AmRkm2KlI1pqAzaLQIxtsXu0oD3aFoNyH1UUSXbPrDWUJeu+posHRU46aGN8uItIk
oc+ep1cxcIawfqsESqkfMRF+6NwF24WCgCHrjQoaoAWvrnBPxiO5HgbAoxo46MKSq+LNTO8yioHI
v0WsgcwPUiJe51f+4qLV2I5VeO9vh+8q4gcy52PT13NMZ2nxo4LYG84PEfN012d/ax/oGdPcaWsg
z4wt+Q/xxYrHmVyJIKVgK9TIoJLk/3xwf8HPGC0NzebOVMtOhGkCoR8n+K913ihdcxJI0wu2ylw/
iDXWhL4mAztnegSPrOgFt4JhNngLCVvCGT1lDryhwb5Zvsee3PPjGhuV6FHi2rUzKpP0N2hAGF2M
zwKPkpJEvzzT9t78105BKuKfUH4bv1HOr1l3B/bQVgdBEnGGop29WoLTSjI2ziZB41U4AJCZ69ki
EaeCTyh0kTfTrwi84A3a/2TPeWEHKRsHrg2tMKplvz8hQjK4FreIOUvIenut9xPyPdxl7qinOPEA
BNuO4EvHWbqmouE5W2tZgXf1DE/ITSZ96GTEzUrli8AIW8ZgJjv/ovS9VwnP/jdt9mV/jiejojg3
btpY2l23FUh6QG3TbqprjuHEvr10Cu9R+w034ee4g/0VUiFoGt0W5AiPeGiwQJoz2qTpm30mDlxv
UrWsNPCbEYkeUYQ9v2Vmpt8cUGKeTs92NBKhFpElOJgpXFnLjdX3AB/MHHaLeVo6Uu39X7rXRDst
AeDApMN+T1MNfhLoskkOzvekbauNSLpcrLcMrdILbB2xNl18wpmWQzzDtEr0mi0kvW2/KFgOzCLQ
Vgvb0MiTcmumY5IRnMpEXwPsY/Pnxv5nO6C4+ayVrcTrm1xiBmzxtwgYjjcOVJ/YGV2YSIg2JkFz
lRBV8grQth+S6etYNxOyU/TpO4WdjibyWU6PQJuLZZ8vJ9SSvtgpDC8GW9N3inc5T+CzQIjqgMXM
nRN5jl0rhAc5DYCRTgTLG+wlJquqaVh4lU+n5Rz+GPoZ0OVh54UEKMsWY73TJQDr8LDuCx1NJMRa
okRY8xEwgZFMpUakHRQzF5xcBAOfBeYgMI6AXcaks01KH4amvzeopFDpKbFDM4BBeNLiPfVXwF0l
B2wnQaOb+VRF32mo850Shs+QsInQnwd+sWQSO9+PHKbX1Y01ar7IAjIEXNifhDG3zjKSylVSILOa
mMG4zgYhpSSBz7kv57Bme8DwfoDEbqBqKRAEwzxycvMzER54tBcVwueb6z2NE1eV+zP1B+wY4w9x
LtbYlErDHZsO6q99bbOGrQVk5jvB6kH5apmvw5F7gf+0cgtXbDRvzY3RE02tXEAEvph1ebLS3gZZ
aUjIHb4WcQHCCWNHmPZ11EUlUu5Veg9A4y0jHyg38XSWgajEZ4bV+IgJNNQzBDFfYfjTzbCvm0w/
yE0PqEkj9exAGKRhDBFnyViDqyuv1xJvzw7qpf1jPPTSHrgGJ8HlszIl53h7t1M9pyGv6HtXw1+V
b536AC+YG3eEPotq8WVLk4CSaIEIjHvRqMC6VzFkTHcDhXu34ao5dMgw7wRENeODpfj3q1peHjG1
lRODygcu5U0du2tLTeyccwQQYjA/WrlJUZonZVhdxDg34BfKw66j6666fHae+INGRqsdHMRxY7jY
EffRuS9F5SGS3OIHiwE/Ei1lcXOZS76WVevT8I2ZJWW8lJO1qMrVf+YqCvJT43eF0yWj5a6sLYF/
akzbIp7NV7Ffzil9EjW9aBtqn/mLBSGR7MZKtpU69pBoYJxAKX1tIEqsLPgxjixV3JaT/uCj8j83
Bn4Gg4FsTaKO3MTEIqWfKPDgvEuc9/OHWdnr3tUSW3cr+xb3Ur5ZAnLm5Wsx/wAaQHSnNhcgf3iZ
qHucmvtUiZsKgjfvhtwLTSqvlq4TIKq4GyptwUroKwd3itoyi4Lj9qcWHzOC8PvI/rQBBVBQgMCi
5ULUzIFWuoKXFxe6pgsja6XU25Qa8bd4t/uUDjh5QGhO1RJPZ8SbgAheDSoL4OoKm/wEakynannZ
hC1WbkA2ZJQx1asRjD/SLuBJ+4Pjyd5TpKHAUxutpIIE/LSP7nXH2CkVeZXhXSaiOwEJkGpa/8Fs
kcXj9JS6muxuGwgxsbIqwWeXBmq3dZuTBc+BJOT5ANo6/0NsuYpwO9B/ffIQ06e/Xj0jYlaEQfAW
omNcYMlSziNDuQnShCtlvMs1nev6YyFbW12eFNKdsgkEojW8qEOxzjze3O/Rwjj3XloidXJtaa3z
UYUyTMuAGUwFGkzjy7V+Qd4giNDzPsBbZSRiS+DucqndIyqYE3AyR/Z7vCV0D82flIZW4qxg6fVo
GrxIenjS8DpcEZrLMV8P9pZ5EIG6eOKvDfd1W1D+tRSsTTHRFftcWJv1i8owmingoO+eqLKsG9RO
mK0hzMXUpxQZ/6uUSnqsXnb8fOA6OQQlKnWvpiip8l+D8moeKxbNWJXgwltoNpH/TQsEZmKyM+49
vW3UrnS9bzzB1CIkjhxRfPN+3PVS1VYxZaxYUBcTfTc3nLGSgegBxBqNhcXfJBTLBh21+P4FlsIr
ODhsrJJzgDH09Mp6qtyqUw4FN0jZGBSFEZ/IZRD05Y1r0FFUu1f2fLD9R6qhxDHdwkHgzQzVckb+
2iSld1+F7PQFRC3EqseCsVwrNOPYk6bc17pjXR7PHeW60t19gM5dDoChNCMY8VxV97v/i9T9PdvJ
Zgu0go0pBk6L3wpY6J8AyO3uc1a7DGd486gwdT+44ml4btCy/Ix2zqpjW9uUpBQP7o8/G1a5tx6r
4MmkARfDWgOZPUFUR+w18N+dW0c51lCNZvaCnWeqUM2kIZey7R5wyOkbCA0bLkoA3oOLkX67cCDk
MEHavIPGfXtL6F2fWYzdxj6as7pcvtLgdddRyzs/v8Efgn5iyYAjhOGxnrLRn7ZkwruTAXBbljLY
2ntfNSFm+wEybfp9/5/c7JS//7THMpNeHTQzz67sl17iwSAZ2dWswpBP4pW4NZrIsYmyiXi4eoF1
zB3spuIqj8Vlk4LpCQzydCqMAE+23TLkWPHePkK+U/f4IRg9dcWg83Ja8W9qSwO+YoI+9pG7uMFq
BnwqBb9rYAHlgcbTKvLN7xwJ8AXehtu7Gw47YzLm4//PON80Mjrcw6s2kkKysSXRLhbPh758PHj7
HMA7/PeUzjrdShzouneQ+ZrMzMy2IolubGqauXOSCkxKNANBeKqI0t740hWQnDMu9KpQMD4PHjp/
a++8Pe0nZKGLUDMCM656vfXMW6c/raaAr+ijVjxh7pU2BzchQWNC7HKdn+slASY6WqnYZVjnf2TL
uGuIQ3H7tF7BB7coAXMRisNy2Wme8dkA+/qO8WIviB0/N7oFdzsCvLtCLFy/amJRCVdbbKmJYslM
EqIfQ3AAxYSfZdqk9/N9xCrsi1JsrX7fYviARgntDDBqhhMp4esGSa1KH+iJkBG9xAWu/OE9PE5h
Ipo8jS2GGpBKva18yoCAOQ7wKCz1Qj0auOOYQgaDRAOz6a2HKLgr6tHSqaNHQfRPt+MjTvWiSkRk
gBaP9vWIwa57fFM4zxqesNqI9+STHZyi4AuA0D11/76Gv6bkOMFfH8KW95Hg+hChoR4177Zll6Iu
gocnhqXeNn3/g5VPJrSrB1W3/6z+NxkA32p184uBIuiU4pWBCUqOrL1UkaWOetYGcrEmyBU87851
TWo7blS1bLPYB5dQg9Fj7TQe2MbIOVHL/E8y6+YSLIfL3I9px5DNCVj3VwUxv3UOXdSlbnDZCH7W
qJudPiT+A1zv6/0GVHHA3xkGutQEG2fqoFHciBMV9lmFHhtTims1tMYOSfeK+t63GvxyfIo7yq6j
XVa4+rfhE5RGxILLPFstt1i31p0cMSgTu5NyhKHUuZFDXAuuJi2o4JYmUiHKk10sA+hYLQVgwT4C
FXMpbSr2vfLsol0ZpIm+a+HDbu5ly+aOzki3d/PagWMXI5FhtHCLXRJgwQyMvmTp/DldEBkI4ByW
hjRt7k8sAa+mk7sGjxlSw7inwNN+35W1PsNG/NgFIvjefDtrigizAubopPtmH5+wGJ9rR4IOOufP
zvqRz0e6bdgZrlGc9uGlgQR5t2RjBISQ1Pvmu/Z3nFYZmyNZHYWaPjA0OSc82wnbReKWJ2VaOtUc
midOAF8uw0k4i7+mjtFsCQf5Gj3arm0O5Zfk9r4N1tr3q+P0hn7xNIHxX2w0Kt4An9BM/C6y13Kl
mTlHyHyF4LDF2KRBDADovSE8J9jPAxVi1nkV4k246xyJNFULAsjc4yb6Zb7jalqVqfBXhRIRJGiU
+Bs7smC6FidlNvDgWlEEKzMUGdu5aaN5EzPIpyh40reLxaMOhHZVRrrgNINSwoNM6ZoDHbG/Wp0m
7Vk+K7YGkzZifrHhp06zgVmR8D0mOUxVNTfLVRJFfS7n2mI0qp5fCHkxoKyEKU6aXIQSoDpf9gC7
HKROdS7LBiirpKk8k8cS5KTP3kjBHMmsPWborcsPKiz0iflkaLYMhJX/9vBkxQ9caeHc+zkThY7q
Kmmlce3ceSAU5UKV9I2XWEvr1SgJmNttsuT/Zmr+wmGBDaKeNFCAIqRJ9oRjchF+HomSWRA2vQuT
E8Gp2KrkJnL263vC/c/i8OiltThde51d0MUdvugmOOaKN45LEopKgEOCfwIn8BDpwlgXqheMF1PL
go/B0PWyLeOgPACdh62CrI3uVv9Utc2WocL52PQj7eHhokVoBYv0Ku2q7zBn9lspjpBhdQ63yuVE
I5RfxVV3tgBrikkSqFHevNGck3CFcpVBGZ021IKucvpgmFflX6JC9yB/atLdiz5MfK6DHpMT6JKX
AZ83jC63JbQhyDhGye6t4gpzpSKesPQy8IU6dTLQwnGPFPHlM3613xaRT8E7UdvXhJc8FFZKubS/
Yv/2R9OE+webdCXwsDvp7FZKPZwHI1cf2g/t90hQaiJ2Bb6rn7T6VaU9zGXe/4OI0ser3h3Sdv3k
YtOPWfRqRrqx6iSFYmwHB9BR2G/KrYwjAIeHHa8v7yFsGc2OW6tA7zZtEGB7ePFBeI8T8/Pj3ag1
0BDnXplbqtJ8C1qDntxb4A7LkYDt2lFQ3c1C/fcIGAdIZFzdNbJz2yQXYp3zXY+dUBhdK3JISSGC
4tOrSERlNP5ZOPQHDZrbMS2VmYQUHhJvmKTeU6HPdg2FYEyLLWsD8VVZjvY7HBxiPp44BvjvtrSX
UmRrmFIBQXfKczUyaGTjM/Dyq58eMmhTLLAqoBHToVC+JCJiMpXMHgUmUhi2U7wlr6Fb5y0CgNIj
solh4SoDg95ymP/9e1/LuHSRezo35ydu6iAmkb+qw9Jp7YXak5/CzPbIrrTCPLCmNQwc+GM7VEV8
Sq+/iMdNTcxzsxhwvrrIlycpuERdRMf7AOWWm1rlJPRmqeoOGrtm9u07nEmNkTTNjogjB+P4YmEy
3p8J7yiDC+3wB6cbovDVsxwplrFw6Vbqlcr6rG6Kd7OZf0MobRICo34npHPz63Ry0ph/SLmSUb0p
ZSGmHRu7ayGCL68BnNFTYRBcuL3WBWVz49vjgF0jEHOLqM+PHUbvy8ntweUdHhXUv7SuZ9NjUQFd
yb8p1Pg5/0PxUMfFREDSfCN0Kq3wYOL3I6z4kjmW7nTKiyGoR+ci+zWgArXDEVmVwaoKNi5uOKl+
NeD22zxaX7KfZNPYBa4PXcJi8N2ahnJqthomg1ae4xmP2XnfjcyaSEo5aC7V5GtHQ1FBPz/EXfft
XPuER//RdJfzH8Ouwg3GuJCFOGkwI1qT49OrczEW6ybWx/SyyB3idd2/XAmWxn36su9FnaNu6Djb
AGFIta/FAEeRYPC7iz0YgEa6e6RvPLjDXXSeSjoeW5YkYqo2k7p3uh7qu0/+h+QQ3/7Qqz/6+JHo
4Cb2CEdIEYxwdNkxnNkFhrMMEp8dR7ic9vCJpriZxfbEHFbpoUXHQAceGGauaHNTGMSjJgFmyljE
X86y/ER6UGwly7tZ0ptxWRZ1bs/Fn1OEdMeMR5OGee9tHe+4/HEn831Nwd48u4GOR4wusJgq3DRx
WFupzz4uTZSIVfbNcvHg060Yu22Bi6SRMksFFIy/QhVphyG7ZFoEG786E2JWARWpbxtmLDTqjtUu
YTFsSWLw2PYC/E4WS8wdxK6Km41PWqca/Z34E2I4b4E3bR8zqRXGw+6CWzbpkcAQysETzyYJpgBI
VPVTaKsAlAham7Eut31sUVRfNbCG0YUEXBF62E1UojwoGo9xnwA2ywR0DdwqDilqSTfPydAw4dRa
Sn57mFyMPRly5Z9wahxoEm/IYh1kQCC/OBt60i0dgcOv34Oq/8njNY3d1kUCihKCzLiq9raksynu
XnzHL7hZpicgz6gTf3ktaAjMvC0NcPmShop9XIPoocXn1XK6kfXrjdAjTsBkELWVp2npiCCR92Z6
KkSXqfb/5+jSWXih6MofpOvjcohbCzIdfczDpQ5bduZYIe5pou89LX4N+caC1lo4pFkidM/DFh4U
9c1Erd7g+x6Z6i9PKqeyZ87P55YO7YnSngNrP+dEXmPyAoTBBPBgPm8fxMlC9BHgoSzValCxOmVj
XTcwWMu/lAgBvDRzwsOkyQwIBStWgyVj3wVgZhYZhw5brZyu6jbdzWMYOfoVLFTLqMpH9OKKmrMS
kwDhDRZneZiH1hr1rIPj24YSA9nTt6IHDDc6rYUWmnYDDrI3jMovfcSBAqnCunonzTRiyLO0rA2i
H/r68pflPQi4LzFmEupKCLM7vdNbqwy5pvKvdUx6aNY4n+1u50vSNFXEwgoRsPc9mGzNIyUx3ts0
Had55RSHjLLD0UowzcWL7wmNoiV8QreyC4lWQ7pUJtwmQlGhngOEY3dv26CpRv1JEK03HtqXZ1PG
Q/tRHDFsqp0ZLH9EwVtKRvLgyA5XbFcoVnPNsKfo8a3RLL2o1DW+o5IeA7Ly8JEzMA0LRKyY/HDO
fCjKrnBY7zF3uwLAeZtPDk7XhHydgjPaatT/enrWsq64wvLOzLKd27fyLVRuu0/ZkwT5UuLJkZjf
MQuLUlKYNnO8Qz6Ij/QN18jiw0whu7RWk3886d5wnwmPv0KDh2Oa1nA9sM1vsYO3D5AtF5JXyilK
K7TdBHTqhumWdY+XMTjpEkYITg2K8yAQYU9vYZK5hhL68oT2/WeO6u6dVM4ksKiJJHy59ApvgE8V
ZAqS1hMFncaJBoTH75ewf8M2UvlnTbpV8dIw/oUi425xVmAbenfSDWg3kKZJhtpqDGFj0PwaIDzq
uj0q9IT2+uaf5oVQMPnSwO4i58cp+qigXeR32Ne0plKBiX6uQUqalUyYWXBrDr8kYT1XF5RG+ABs
1keFoND/DRpXZUoxmzfBGO+RFvvMDsz2XAHa6GmG8wnANcuEIUyrtS5nW8fp3LfWW26O5eI5/9DW
1LKRrhhroGZPs5VW4hv6bo+/kNmJQtPxtUKJgoPmxwt33i8HozpK1qXshNIES6V8JshbS6RMJ3w6
bjdu7GBJZWNePEJZGo5P1AlAxmKwVCQRxz1MGqOvlcfWrB115eQgrHugMF9TtuhN+ur5TpV5S2A3
yznxwRoVh+nTJM4LlCW810yXLozJE8UJNgb8vO5qXHCXumBK5NRAfsmebjMIfabmm4PeiYPN22Bv
08HqaExGt10kDJqa3Scl94GXg3hzrqrKGT2xQy9lxAE4zYbGtBtGf9YauSuF/oe3ij2e6V90RMbt
ZVS/b9Avf2pWGmVtlKFJtfFecNrHTk5qZSBMCZIVlA1IeqP1cLJw2OXFEvh+3+tP09mDd4/a15pI
e+XmT04ZqSZ8KgrbI8NArHkqxpkuw0LrbHNvIEbAiwC/rtaL4HuZLoBBir1+2Q39dVlGhW5UNov8
nTQuk+mgLQ/cALB8hIvKoPK1LVK6WLa8uC2MsaNa+vmFC47jj05miRxiqpNwvSjx0hyKXiPRLPat
X/BCTyjCuCfc9bPMGOpZUTwBqHCECXTzgi2GnQf8WbEaAjo3Wsw/xGZXBUWbq1yYARvJ+JP8r3HQ
ccuD1PygsF0u1wX/YnN9AhVGVyTv+iyt6GRaoFFcDyxEaHM1RlgEM4acVfNRL+hbm3zd0bsWnspF
3pfjW/yXA3yo3wKYZB+8lWQr/ceXPfGUwu7GwfZ3PtE4DDoNKqE72LJ9cvU/Axs8ErUX0wzAqaz/
vwlN2ZyrU3MoeYOAeAOnVOMSNruGFeP7wOPAYIFhgVSKZWqBLP7O9INexv1gf+xyC+48lbNgaWa6
EmekL4zSBY6g/5qkSDAHvP7g48ysyOByG7VTFkMy+Eg6PIZpOoA3JTK2WRCSQEYPk75Uv2I038p3
durbZyf2hCngXRI2waLhOm76lKlULUkp5nKNykcngqPJdiHl+LJyxoDv6J3CQ3R87ZdF7UlZfVEu
EbANkjzoSR86wnCdjwY9ArOusOyTXWy06U8s6bJZlI7kXFPeqpAigukhaA9dr+cAFQIAIx+URIQt
VXMr8OtbunxrYm2E1NBc24qjGjhWVBYnkixOPCHpL1MEICitWer1fzv7IVxrFWuI+Phx7XNERxC1
mmx8ACWlQBOUnt+lAACHD6zZqKrnASxJ5NslG78Izc5UQqcQLr80rPKI48dvYWYjLzdZFWzsiX/y
XVZrZg5o0P3wfkqoYaM0McyIXE5qcDcgpGjH9lZnSMwxFfmPc2b6lg6Qir98kIwBw9sEOC6/ywty
bFpNgoDJwUKsp6L8ECYFklnsJsZ8q8i390ZeUzFTQ8//TjmGG/sx7aBGNcNed/FjRkAf1fsGBZmW
RCLZys2S7khfJYD6wS2rl897PbdOQxbrigt7Ypq+4REGZjv3cqd0Bp1xxUZfqqKgfYmSmz6oIL/c
75Daqj+bd6abxWLIP5ClmHq2UnFPYEOTY/k0TlvpHvo4hg0YJlu68nxZVbfcN1EZgm/38hRF5dws
kP/6NP51KQ1R/rQZm3c6BZcdWXVvMcB1RAPSmuXBkuMWGxvgbggpBgn83dp83YAn4jqiOeJuYw+G
Qzymh7EcvuevRHFf7N4+bIqPbYLSgHeTfQOdT927ERQZ955AD6g3raSywk9ITwz2xoFEJgjZoooy
h0F31VMHXWYyk85vIJy87wvcpmqaqK+QlOAbG7jV3V/HG/VKlldYaw3hV/Bf3jt4ANqN8yfFIa80
ljwTy58Y1h8Fv2T5vz5L7LuXkINH/Xl+GjPgHWZGEwC55nbWoJjdKxBbVKFsRCF6gnS5oIN5ivfA
eVz/95lFLPrzd5jqwuGl0a9s9zsUQfzBwRXiwM4CpIWRCMJPC6TY7mRrt+HMAdptuTCKi31IYKmb
d+umTFXXul5KrFUOQZBE2ufRWfsjGMd7nTZo4xPEr9e9ccGu7IlSXwUS5WXOpJsw+Z7vBOZzTbDQ
33fpNfOhi549FWXVzevRanueC0ZYrvxWWn1PzZ6PPJVIqiFx6VLXwc1TAXk12OTPX2Dq0E0XK4KG
XcgexnIpyTPeid03pQGHQjY60a9MCD8r/gBfKOjPJeSvGIRB7vHdXU1XVupTvIU5tbfWBp4I+POg
KBFZBrkTEvuLInlNX3XViWw//tUhcjkDOVIX/bO8+wrRJ79FOIoTlj/x5hvTFhDkIwsqj/5TeivV
H1YwSkXl2o+WwYSwd1mAcW7xY+dne113JCdb2LyJIQO3sa6jhyA2+eZx1t2A1ZOM0Tp3NOjAgp8i
mqeC4IcNaby6jbOWM5eYVUCBYO4IXSCvyWp6YzORmzHzb60QmDn14ulNUcAQuOkWPc2y6Qu3vbo5
97XH+HG6YD8xJSzrSSG+VH14cailCGsPiJOmiq/E9qSPVz0dp0Tyv+hM11sLOMRi/peRF39UCAUl
1oM+CzuvIWftdOSlZ/RKg3JAYH8sOvtCI2fV/cncxWzwi1JB+2F3G9S7c/LC88akEcUBs0FyE357
NjFe0AJOI/vv2wek9dxN/l8AqekdAPzwASEo2VjZoMsm9Q6ytzZbdC16SXFJ1qP81Ae5pyf6LX9n
3Xks/UWYz+RNS4V6zFRnGcl77kmboU1k+bJ2o4fDU2iYa2Ym2FajpgiofDW7Rh6NBx1fVXIlCbGO
/UVyD8tZCBQ2NbpQ31gjPWXhpnz4MSy3GcaxJpXuVZswtc+02JIxxM4ZmUUaySH5HSeUR8ODkVkw
519rEcfDlLH34wfAyBJBd0hxMPZwZoUUELCwY/6EkJsHVoRHWFu2Cu9GhJqI6uhbxwVdjjUjSSf6
meyZkiUIR4GAHgktruUptFUqIDZHKz5ZWqp3kNutCo2T6BdbJMqqoIbe+Hmn6qNXXqgGbp2of/IF
3spGO1GlVA7RwWbT+IOLhXtIbMZKT/0KSYf9xhGYLYO+ox4Alg1tqP52mLHlqOZZSWg02a3Ge2aJ
iQwTdJWvIGA4NBUKH6zkKLgfHREz+pEDvLaMuFcn7iufKciUfnJLzkjT6VHnpVJgNFrewasobRgF
drWrVyb6w+BPCHGD418UmWSCYVFySyxblEMjHQT+pavrNGfEUs1JKOOvRSny9cOfR2P9HD61WYbu
ELfNko12lWfpk8cqQ34nm5Rodw/De6bRENGtPc4aOkHBJf3Zppj+gkM5A0ZFbo18069liD8YO6Gv
KPdHXzffF+XUBXxSnk6nhySsA4gpDmFiIHHd4cMBezQmKkdCtWtt77DDKk4H4DHctXSGVGb3+fc3
Z5So9YvSr21Kw7bjkNss2gGhGs/I6zT8u7JqxJJr/jyHPmmRlFZIIJdZlUOOzgy6RqV/BxJFrooS
lUb74gWgmLzRzZZhXCrWbMFgMlOXFVrOU4feW3RxS6wJXUJljMzVhPgnEWhaHZqtUCdKBdDmAqaH
p1ml0xwdM2ReFgn/a7N4lBZZPYUYa8w+putluxigJsCunU7DpJFgcQnn35KLWGaw5VPudirqaOL+
2d1r98cAGsvzkH9i8tDslSZMCHJgjsBtGSQ6NJ3W1e+nz9kw5PHBosWcqwjW7S3Rswa2VJCo+Ewi
p2Dvgj4374+wgJcbo9mGmiyI+frJ//SKO8ZNBUtxK3O5/ZVT5m2uLvL23d+fi9JMjbfLsm+Oc+Zx
VH7o1U+nlTKMRA/RKCJaDsDMgBKXnppWpb+VSpMds0sOpYn7emvFtmT2ub30G2TjLfJ4cR1FaBLU
hULG5m7jm0ISM+hN0j3cIe1zOWxvYLqOtIGFrC1EpWr2tdfPKcb7hLHHlwkaGWHUPwPeawTnOez8
k8ZDrGo4WnNMFrqprr2W2/lqFYQWUEZWBXG+3j2jzhFZZgdZIGP2I2+H2kPrhNzQ5E6afS4sbLIf
BwhSNnhP3GIIRPTMMl/5zYaRZwdYStBQSJDZo2OYqE3viWc1ahk0K+ykBSgqwxwbor+2dfSnOBR8
xiZv7p9sg6QjbTFUqWQOS8D7CC1aq/MTN1gJHIG2mHrduBV2YKPDR+CxwWYiLw2ai8NUsgRLn48l
MwApI4ChIeO6alm2XkRYRE9lVzgQ7LsRJ+aqqugPamyghToLMXT/shpGL7htAARtbvtYDqXAyLDh
U+P7ZciQr5aH2eT2DlFHHntapIlUEAOTzqPz2OM+HD/XS1L2fkrYC9lW4I3olZrP0DkVsQN3SpkM
cPAmbNFHjRU+hmIqBZi0CbTpHITBlVKAodkFzBZAxpXojABYRAn/Y9KdQNNRmkjdO0qMUo0tloyO
zsaKE7+DuGQKkdCPLvBqidbXLls5aSBcFWuBju8mIgP1gzm1mkag9LXARhuNF1XUa7aNwQdx5dBH
yJqsKaqoWGHgT6pArTKEr7gZyFtyPkIV7nVvvEUS7bm02xKPAC72RBAamtiJGBqMYtC1LNdLx3ML
7oyzQSCFIRW43EGUYZNvUBQLPr3sKYCf6x5AjiA70SJ6Yc0OjX8LQkxffL+BTU5yQoX34Itf8aHP
YZLAfY7ncdxhIU+2cxKrBwQd4dExVvFBKv8I5QhVkrCJteYEZUa2lGRx6HOK9GvoPlq7dw4ba8W7
o0QcLn8NRIfcV8m+T2wdI3cyRA3fGbknIUo2wiSOMxnk+Vo3Dz4nYbflKSVY9SrHPirrj7TNPH0H
wFjZfw5HhiCFe93PktFLtxvObPxI3A5Y2k4eRYD7riTrXq08zRpTImlG7LzNmf1KBVlANd1zhXbS
rJ+90goQh6hs7AC6G7vNaM5BOZlesYoloUVtIVVPDjESTFsG7BFK8TTh1HjQSZ0pXpAs0GUvbFai
kP9GknKdddG9aRcZSVOfyd+ikblDoa8PeNxBwlOBufhj8XAcp1uOOQEeKVuVNzVtHk5xz5Ka+GCv
vBAwqA7Qt3oYjjHuQkwLZgQudWtSxKTew6T72y45k/DdKH6WsOByridk4VyO8ZgdB1oYh7ENSfG3
FyUoXRRzR9EGlF8JqshmhaTJbbAW5zWE5t0TxaVoOWYLfmtMJwMGglFDQlka8JNQHvIHqvfFq0is
3Jb7AxonMuH25bhTHCi7SeyUk8LhgY0ETL2m+dLG5YKbQ0I9Hym+6dkMesNMDzRTTzYUDCh3LqtZ
kmzusNJ2NkZIhryOss/Afru2u6XzHw7zVjj+GBKOCE/xGzYe9fqnvIAj8fLok1kqJu12f24HbggY
dAbGnDWPFFL1GlL9Roq9M97TKOsNwz9T4RjsnW6quIYSSVmbr+niTmmv0tslVVnkWyAA6eJPIv3Y
A+i2j+PBx1hKGKKVzQFGu96m40BT5kQOBZJi8LRe07aJ0G0v37t/P7OG/dnqjgW5EsFnewr9Ream
uzgCI6CEra5oJddk+ctHtyQ3R7j2syT8jNU6fnjXydXNOVMJlE5S91i5KHb0TaGO9Hgpdzh4XSgM
NwNnqcaY0t7wWaNWW2em3JVKAu0HyUOUmg7mTb8rdDLJ91szmHJdw07eFAX73QRdLAnSu1+nqxsx
MFr4HWnOrer68Z6Rt3vLM1xTetsKbGX2PGG6vk2lNbtYGteRu/zBKkirZFeFQlOd+D8yUuYfwIWE
q5hgxJnDvZyR7k683XSg4bxUg0dXo9TA0KgyKqnKowyywkVp3RJvatfA0S7xK3pDrVaZ1K/ZUFhw
taDATE1k068J1RJNCagAl0QKCiG3a+Xahy0feFP5/GbePEqeRzT1+H5Ulb/DoeeTZE+7JLV9ToLZ
oEXy5lULcvyik7NXwCxEyb8672wbYPzM4EuTKlRfUONL6/eUsUVDcw3dHkaMph+8EZ27LlxYTyq+
2qzra5wC+4m4dLzt004nWvHqZlwLSjQ5f95prMNb8LRHObFJpOg1EBbQlNyt5h3LkiFrHucv6lo9
2ypFRt/PTPOdtRgLD32jLtWCvEasUzVFYTzZqiuZHH9B/ZAMigsTdOtsfQuc21BuE8SnzghwvjXE
yir3gRMVO9mh1grD65aS13gwCxZG0sSB0Qn4Oj/ogrrjw1sUVD5oM9v5lR9GbKbpyRa3y6fakuM5
f9257EXB5Sv2Gga7XVmHrZfivH4sS/NWORmAYfy/m1Vwf+cRjBeCiOhDBoBJvL+pC7l6eslOpLGq
zKag8fX97XHxNJJbdx5BsXPVEn0yqHxOnGJ4DX5h+TL7l8Em9Z51QUxwJ5RG5uHGP/DOLVorxJAj
jIAzHGokSbZHI2/8Cp3O3R/ezHYaSiW9Lbt2+DTA04UeGckJyoOTGIAtFpMocj84Xut///Kkk68R
9+iCIEbUsKyyBb2Axu+QC0kokqhTMqTf4DM6zg2hE80NMjx+ogg+04lftvSvKFfPlI5bPeyjQyxH
sUjEO2SUJVqyxos7pMWbsvNlCgjHz28DIWcUyHMEBMSyp55mY2Q297pv2GU44kDL6gP0YBzkdcYx
ipeX5hgqqEJbb1GTQJrvODOQNQHH1RLkTGxSFheMUTGMyDWOgjb3sqtjLHNB7ws76+dHl0Ww3c9x
yZJUtOheAbIseeVaR2nbtFFS8/SnaK2XEI9eHNdrgA7ywWfyETEkVTb0GEHHPBW2OySkAHhq52CK
d8hTs7XoxYyWHpZxqt8eCug4n/RAuA0P6yTuzwQYytmtnzXECZMAtCj+JuKOgDUYfSaevOxId5Wy
sAXMLavGieeGtuw/izz+aLiDvz5glAApuOwuNv/VnMQAnXbJre2V+0vCtZ959UimUYj69uV6MCP/
RRjqpd1wYmW4kkerndSa5OfjyHsp6ay+XldoXleTV5wKOSCWBesi4p82PIzZjUmXWa5hQuyQCz0t
WNFKr5eLobwofCJT7hdThwOynSohEAH1jfVJ9CgUZGMQgH5l8PfmEbDOuW3VMPYWBw9/LahgLK99
s1pULo6nZ+qqs1TOzVyX89+t29NFnzbzmp9qYSgR21H1cQTqkEqpEBaUV6Mu624wyh6B/EzNm0c/
Ts/FwiB7Yf9X8lNIqUoYXYLJZacYyYLuT2m5lYOzVM27zQ/GAg9CCQJxqY/XUjoTTAzrZZBfxtFp
F0IDC3HsZsGD9U/n7Sh+AZJdQZLLJm6XQVyqoXer6v6i0Ozwt2wMIIzUmEtHqFVFjxUCZTT1A2JW
yR/5BnKo+PbkkBmR+Jn23zYMIhUKOYDSU/TJ5M5HhGuJUlTp+91M2C5qIHC/47mseosHQguT0lnh
L4qH2jnXPMBkemQcBlR6ILp0r74R5gzrFScF2D3I31KoJVwplW1mUmNNKZzO+3h68jew28qqmQzu
Hng50unsmqYwyKqt8V6MCA4p6BkN/mAkbLHrW8TN50+E2A9fnnSqonleR4v01+YK/mzrhrSo3NCq
U1PleHsmTbcy2sYD4ADtz/vmYfyP0szYDhJWm2XcY44woRtrmzdTi7gMqzTVgmUukL0BgYm+rZfw
2YXbwom3cofz1y4EGUOVve0SOXrsQ1aRR/OAdb9pUVM4H1HGXI2f1WMP58P1sDgvQz6suJtS0fK9
et7BwHFicg7k5jI3CBdm+XKDMJXAmYhacB4sZZcvh3kmU46QIbsFUJQnS3M4I/NKWN9+tNHNyFTU
7vkrTJ7e3yOmL/BlhzbU6pd1VLSoJlJen1lhSukuRar2Dg5nXgLKtK6mO1M8hg5bf07To9YYk1J8
nnLAeYZigbOTDPVqGrWrGs3u8n6kTq/l7jM8kwrqyPFrYl+/GtfsJwAG6OnXo88uDsPb4wsByyH+
Xk20zTWn44MZB5aqcD0IzNimDvQoESrxmrTYgDhcVWO1uxETdSKHACGN+RxLj9kECU2tYCuSPzpO
9EWGmIc+/0uYCRbw75zCwoejyXBKfx92N0UpighVyXJ+SRUZ5zipXynja2GWvS9XctI9skPgVAgw
lrGGfTcJeleMCXWVDvHSXdRW4nOsEuggSeqOsXjqTwpmg4JiNB7VrhcJMc4I69KQ/lqOsMgRmTLm
rYZK9MYwVbTx2/UinBioaUaJec2MtXzQBBCfjSy/QQFmXO36CCZjZrE8S5CgwwryeKI5asqocg63
bGjzO2R0cOz0UcmI6wtpYAYuW1syTwPv8E1N4p741+L08ZhAaugOpI9UmVx1iYDnNjOrOZ3S0bUS
f0az49PB2a/iDsIScRqdV+sUSErBBgYFfdnQEwIUVhv7DpBc+NBOHkKyq7fXpDOgAF/Ipa/7x9Oh
8Qbt5gTJfBEkAo8elNYrYWF7PNVsIZbVjKovk7muG9jwLBnlDYHOMVnTpMK5Ahc5mGRp7yQ4eN0K
JgsoS9C0yEVoYsrTR0wqdUgknXkxt4z+X/pXY8BNuD/6Y8HAJExEa5SMBHX/OS0BzgnAg8uQZiG7
NuARocWNEK21JjlwZc7ugwCBJz+tM9zlQ38Ysr3BYMS6PiEYPQaObNTVziMxt1AcLgo9S9dvZ9xf
v2tnE/xosQKGdbjW3xGu4ukIiqBVjMxWhbtP0tUOjPlfZ+BrhHXt7r1feCkFJyhTUsjVPxJSquba
Mbk6GG4LmHvDI6rUG0X48/4BrsH5BlO5Bmo8i9jNOpu00j/exOJXKcHaMV+XCrTriErZ53jPRod9
+fBFGt0NW2fo8mtKSund2YhLbUIBNlAz2mddAkp3qkzblsbb2gEmohH4GbAM5dx4GAwSrekF296H
jn4woGdYBh/wgtpeSffrEHvlExXY184xWMrcg/yiM1fsiIcJ+I40Br3mAiWdasx9bo1xIdTdlghG
1XWPQ0Kg88gnTCNp5lyMotLhLzeTbIBxQmwUYvwdUHSRN68O8RescnqwOwcPrYBvyNtNRiCZPDWj
G4acMQ7dAxwC7Lte3Y1cDvyIYyfyEHMLIT6l6QrNyD9ETtXWXw0IJ2TpWx/oxZH8CstC4jGwGvM9
/fNYhW5io2JMXQoLKBkhC3saO76DQeYPz4k5eOv3EY+QFqmSq3zVKCbb9r7oChELmv7RyXgLfrXh
gNXSQ6sPlp7yjAbohYJG4lSXpqaIqAcvHmZUAz9sx628pVCpfHgU3ivKvihdUM2Ymhd0ZulH4Fx2
xAW0NZjLOC1B3JSVf2qj7RQOWTeuAGIGP83QbQbsKCUjsE4qVy86blsIV5uf9kLqkMdNYGk5U56o
pZH3D/RJYD6W2XY3DarGrKTFvwG87d1uHsmGABew7E721JFww79pRhcGibnkStQvFyMHNkeQVIL1
bwScGy/j4PCGUqeejKwmyCTHLRaDCqwZikhNiGVCk3RWcKFuhmktyVwN98HspG91BByzV5TLSpCU
LhXeDUGc1/4LZw/wlzkZng9+9nBWB84bkQuVBNGkYCQU3UJglgQh5ojzWLhunvnBqytS9wT6vrf0
GWRqrsjqcZRdExUTP8dhyK71kGtGsPbXqlSDkxl0AyZx6YQ9aO1rpgj++4CV9WmGb65R4/IPIbmV
OLDf65fNbfdL1Xmcj7dJMpcogwWiIfJ2QPsJquuDMvQwAUCC0rGQO+XC8n4qp47gwgyvuUtx2p0a
iBVlyd8YHkqFffN21Af7jy5F/AljM+Ar2ODVRvOusPuaXtwRtigHh4REtebt+1+wyojXIAmmNgTK
j4Av+GwddOd8AT91DP91DMQjOzn/5dnW/mtV/nGu6+5V0MqX+y2nRLxMwPhgVdkvVGhESzV4SOGb
WcKD+e++UqAWN5rDoc1NQeNwh3bXkEJ2XdnI6Gmgfy2H5tcJ8qyprn7K38f405Arx3D5v1BQhg73
AiXNGJbx0hvHu9v7Hzxp+EowGf3qnFTnq5dbyDugOpusa2qnxfl7gZivkRkvtgSldvZetUHruiH8
j7rdpOdXmLfsQPZvGBiyDfcUgx2dayLyS0A8sHFUKXAUSkgIpnKSQzU/I+OZLGHo7Ok6+JBdAO3H
NuL+MmLP22NKaSYlBbTBl5ikaXk/GxOaTxJx8jXQg8PSQM29MKtd0+97/bBez6SZm0hJO0BRbG7g
haL2NEzM5S0QktOBXgQEZ0+6Eq5qsYPb/RUsXHcBQj1VzLNMdOi2eLvJbAgPRLsVY4Y1QRYrt1oz
8GiW78F6V09U0bNeoCMEMwarkDEcRUWRFtKRYE2AaEOLBYQsc/BKpgmadKlzl9gwWZWHDLoFsE2C
aN6MGNFPyke6P0CkoNnCNCUoG3BiyHtOyRSoJACdxXcS2jfIiDUWK4iS6S8PY94yqCP9qHX8Fz9k
yjeaoTq+vNBWq9ceanwI45FnYAwfCbaPpQEg1kVRQL9iPI2uMICLNgfTDQLrxgkgFXP5p3XUut+j
SARGgEl2EJbuyaNFMukfYjhNM9L96Wau+Q5bVGd+XVQ8Sd/606V69YlugP8EOJckDm6FvNZowhsL
tBeiZgHlr/Sns40NfLm6dBGURnMlstoD0VX7EhlORIxqJYXxysLUdAoR9jhYPprXSQtyiqUMppi+
C9wqbdbfGjbq4rw9fMWtlkOHn1ZWOBzrt19OOqZ36eQx1mSfEQ0taDk1F8USVlXIlhdxr6yEwcTd
PPMyiqIlwmoOFDSGymJyXSq04CAQcvCvsLJ/0n3w52iYKdttK8gNO4S/TywJdjoyq7EZFbFPbrt9
Mho+AzVLNufHpNrNniWF2lpBtnc5MaSq4KzX5nY0APVX1a2hRfmx+hmzOEIshfBNvulVb6m0xoR0
XM7eiCRfi/BlpFNIRIOB1rJwf6R+NJIcWLzMjE3U8grod8Stq7pFHBGBILvO5hbe16PQFOICEUb4
YTOfKGGkD4bl5IOGAFaMHojkXnETA861tinbvBCVC0b5XZWLdD8zNlH029aOddkPpn8WYf8+Fj2l
u5wDruyKTUnud+djsIec19H8bXDPfubd9f0H4ZBoBIbJkz+gdJAWQTb6U3J8Swqd+q5MmN2dEUkB
IzJNSyzUKuh7c9brnNgICskRwlRuX4mLC1VUjMBcnGYndfnixN1io12OYMiKczG2ibeTE9HMsYVT
t/abcsYQbYC0FRxWaDgFyNc4En8t8fGA3Ni62xlch7gcvnmEIp5V8Ivm9qvLF+POFtl6ZIu5Z2Cg
cBGFUM0jYhEQJEghhhzufNjWx4Eg5ziNknsyHUaORtK1qVLEgvbKQQ7TcSzE9dS3FKORdbHavyWz
Qvvk18pAyhTTsRY3r8nhieJ0Qs2HvKwDptSmhVUUqr18qifDlibopAHk2A37boT7FpXl/Hn3jEgN
ggIYf37JvGV02aToZ8ML5Ao3KXf+noaXo0MXiKoaigS9QysK6mAE15BglsxjKdDmzwk39flUGnYg
WSZ5FVNKIcR8LOZuxXMoAqX6fmeEGGoXnPyPVbud57WNj/FfTKdJuJ81uy41JShDtDO6soimfI4X
tV6u58EE+ZmaugdHZI5GVBWcqnwN7fRcx2PsPUOl6DnUUZhsFXmUpUmtMMwOacCUup06Fymn8VER
l19TTNXBTHYvgSjjJg+tEdrmR6DfIExKT1xKoaWZTq+EDD55pkOVaWBR3VQzu/ArfZAJnSZTeOEy
Ktm42B4Nw2KmAiMXUstOw1Hlt++D7JMQpwq7FTQo5bhwfBnHpgomAIfGO3SqTQnCkW8nbwE41cFQ
jb82G44X1SYfAJOiK69kWmb65LfxVCaqAKGcO0EJaLyibkf71ENORSjlH/VMFvGs2fRFsT5JN2z6
5GioZmzKAY4RJkrud3fvVjVRLETUFyxoD51QuXl0bf53e+gXPnogu+aNraJ6Zaj4AO7bKHbVafSi
WjVQEbnK8exuTYy1mBAdeLNQSL8163Tjqt2I0VAOuykgD6C8w+rqZZagB0/078Av9UQ+l6nMqmwo
2z2k+wFmqm0uy7GIpPcAtno5uKJUVZlKRvQJI1kEbl8kVK26wUXhLGDSZBEAU98c0VUb5Zm0T3wW
FzCXtQtm4+U9MMXtT5nzULassjTonjdCoCE/7VqhCZXGC71DyTmzrQYAXQtKzLFc6eGLwqS9YXL1
8fkxqE08MdlPoIyyYh+8F7ld2K9bteaErLis6cqNd5ia1UjlsNroUt4dXG7qMSUUZb0a0XeKZQuC
9GEue05bwWXDOT1em9U1qPgycUSrDs0alq6XAhuFxL5kO0irocKb19vTsIodT2z56jHC9cjLm8jy
wRsw51EmeUcfob8YbVA6KuWoz0xNOmb7rNxcjeXWMqQLoBD/VqUgwU72/BGyc4BanOLwx3Hl/gRv
ZAVZGpCZWlMWuKRV8th1mn8jZ/AMlyHXtuiqQynEGzpRvUH+GMWyicb2WY9MYI7dmsTz03Z9b42f
KEqRKpo30IFUbVacVYbIj4Jn+Fbo7SuErMU0lrUGnpGYNA6Gd1b0JsVfgVEIdXlqZQFoeuEResYf
wxNU1pTpUZUlwyY3iCFKZgzAfjlsSZ0zLzz+W10FK0vY7qulhqcXBGR2wmTU6eNusCyFokFjTvXf
GmlnJEPVYj2fdJtGMvmM6D2tGDeHd6Z+kUSsj0pzbzZZTA1y2ZFFEcJoYv7C1A37VgvPAb6jSIDl
gFZDa6D4n4MQ0nU3HfN59Fb0yfCjp3NkLE0sxS8xNnD/tz/Qczd0VluJ7vjYzsSIWQpPvHUSHg+B
dTBqNP41XUcfzp3xkrIGh4rAUap/+s6T98D2Lj4KIivJ32l3+z4d04VChbWx0GmiXlkOJLEUlEMH
ZhS3kxrt4FmEM+xNldMswV+utxmnLZPtxFJrdj3Xt85bXndMYECRR7AUxRidt3QTp6/MJ4Be+La8
KvMhwrUe5TcTQcE/uI9lYfBI1R8racRRKRsQOGHnFVhsAJeUDlfU+JSFs37aHmYB6DCYB8liNTyE
V77TEYPu2j2PNFpn7UkSiJV2HjJj3g3HvflfZHE/rZ2LrPzlLK2YHesoxUR6c5csiU6uczuqf/uK
gPCjNIrDXNKwnMf/tERHLUtdqgXgUbro8ceCkoTN+ZhbVwMvRc2yzAjT/IrZ6MKQWdBnjRBRpw4H
xhX8OlWf0dQjM07Xy3247MA/ZLqPVCmAwzPy5/bOoUevs140auw9Pe13+Z/BPkDIuuRVnxGWa/5V
to0AHo/B6Nal0W0ZzuM/79ubQPw882oqhcT7kQhdG+ORRc3cy1QWns2QS6JWkk5vlKDMyV/Y3Mdj
dLvaCk6beYtFrb8n/qDnRY7cjFfaZJS7GFXStlILjfeDDYd4SqNCYFkl+OT0cRA/mVmnx/BsAqN8
UxlmBpHY5PiAs43mN4k9yB+JFS3ugnyCvlC6P0wR+IR1BVs+IqIZ1yMSRmtU0uahI2KBGmF8iymW
gxuMXjj3M0KAF7w863i02411v3vLeyvVqTAJSEQyJQv13oqBdV0UrVcJh2NKOvvo9GVZLRYDoTSL
lkOktl3ZSnpiBPIGW6z9SMg7zIxGBjnuzmMtc2L3fk12kxH5dnqVRdGz5utueAsFAYjtjASvB85G
HdQnKOj1tTkcg1awp2AHcWViV+rvlc4J2vZeJNuRsovKsDzvraesPvJu8W4IGd5FhBXhjkXIyC+0
TcOTVFlfr4v7oAzl+9BQA8oOnznD0sNouVXXx9zEe1gMinrdYVtGmGrzip+bKNOk8Exen6eAKGYO
6P/0s0yy+47vWVJp2XHgfP3Cpi6C8DnuEdZbKXTftbKhNFOXWSIwSxmy3DM4DoVVY3nYiEPIhmYJ
fxCtG4CGPhbBnTPx7BDPby4a4C3r99DZKGKr+4v3NHJ+JCnfj1Qsq1eGXSjNNugz7m0SG5zax4OO
s+lLz0k9T06o7dkhaZCOuuoXu4TZCxepGBp4tuF0LLHRq5Bm6tp5hcpHc7FKJqM/k78/T6Jaq81D
M91d6x5VI+8X9xRs6XKC+hVQLghtnJy94e5ehCO6hySDGtaFM7+pdm/E8eVRG1BVvHtII2n84d4E
PYKeT3oKHKV1oZCGmdNkAtkghOBE/FA8P8w8kM7f9xtsqpritwLFv6gZjenvAWMDlMZ0nPNnIHiW
h6jgXcM181436HAzqAaLecJTgjxxu2dk7YGDiMhRq/9fG9FrjoccS5TkVLgYUfJuNDXXlMCZqXP+
ja6ueRVu0jyjgLFGnLByKSB+nGZsQIEfSeKFfOxE68fCw+2EfKx0ADgS77zUTiyWEbsYTh12ghDf
pfiWpKsRMttgaii30fIWvsOtZZ0ScItW5Esc8Y/GNjsVaORZ3Ip0ZqkF0wEXvLlDQntQgskHaSMy
iqeKHHY4YeHJMhDFzvDTQ0HOEhNAm+s7Irmh+7tot9rqaIimf+GKWf5nCvEZFGiZBVmiaIjjo7/j
gcaOlN4FU2kYmIJXDcu0/NBxJwcJMlr+9wdQaHzDulVICuXBqmP/NUpmRlQeFYtXwji4vooGk4KQ
SDODcSlq2CgnescaFdK+18s2e0j48Ke55svHSTymP5Oo9iAyILgxvgDZPBo49iDh6xek32VeXUT2
wc5s+8TrDWBWScvp7iUiMdMxUt/o74ulM1xv4AsfAlo1vQzRvtXU746496vIszsOufixHEPkXOJE
/8sHp8fSvGkg2v/755lZAnIPrZNTxp2r2ASnZbMhfqPWH0wtpt7228I2v0ZU8GYXjwjWq689PPFh
cwZw2dke9ch9PPn5e0sqFkkZF4SXzEW6QGJSEr1XdiEUz69wl0ozTYlqpuf5lSTNGJ5FGvqmh4OZ
tmL3U/HwmjlkfDvHRIEQK7lxmPWyZwWTDE/NytFRScsPf/NJ2/CH0Jargbv2kbZSyvx0TX55cCZ1
bwLLNd6AYJ+j/vAYHhaeFsbqs/+jrkuyL5MFG8OGZ645s1/xuhIfJ3+3lrg9RUfJgJnPhaxzIDdN
yRLCEYggrEhDaBNl/Bw2zzJCYnmW85jFpxhh3N+/kDr2QasYmAe7afeS0Y1S/gr2SRkQpixLDEED
FvZywTNU8dz/43HkIaU3kXGmG9OufPXQfwOcqM5WU5iPEsNm8zdaSKBox9/yeXI2BCZhrBO4V6ji
ECerNje4OZFXElzBWygSooBRhTNQhTEHw3TcgDqKl+tQUmbR1Xzu+9jEleUNTM4W9cS7L7mvMQZa
7kh4eAcbv1U7X0/Cqn+tGN+ANRq8K0EI486uMUnrtI9bGtKHzddPXTNQWKE6yoYGM6xnebvKFVN+
HKojWQNNtOe4IZn1ry/MeH1tyG+RHqHTTZMpRmly3ahYLtdFUGu+sq0+bj3+idLngX12onGAtJMB
BcUgY1GPzLB8Mm8qeosd2z05eyCwx9qiQK1dSU899foSyjDg9kUPBNQ2tpzQW6YWGHcs080eWuPW
6KJweZ0J9qfovwdqPSXgXKObcDA33ysiWU44dLdePg94bEHcV7g/3eCrGauHuJ2O69iEx7t4puEB
PB1FyZnyeX43AFYJjuQZoyMHklrOrtusqGlI0TRqmrAlGkn3Tzxgd66hZkkK+DTQINq6uER9rkUE
BSXozVY2s5PDVO22UMq+Mfk0fG5Wax6EuQB6l+Hfszwry3buw1PTAmCaRVWdviT//a4L3uVBQtHs
utt09V5q+r7ZSp1jgJOwE4drEf5SYgzX6KC564jZyOToXOWT6oy+Ixbuu+5fXkKg0lj8riBdfIsT
NiAOYFgaWSAwciDnvNkZl4zzMyR4h44RhiO4kqNp8VFoj1uVrmIL1bSF0N9IJjt0Bas/eMSqCBBh
aUqU34X7misVDcGAlGma5yoWt6Gf+sOeRziMWC1phUEI2vLMPmbhOWpLLDZ5iUuMM7CA5SkLjcmb
yY6lkzgN1Cjpu/UJNkBlo4t0U5lohkEiNS8+NZ7G00oK8/xETd7UlR3x1J8XsCxJ8zTeab5YHi6Y
e+rkCFm9ZcR4usEQL7GGmZR+MEN8JPQSd4apIXiUEBniJk1Yc0qkMwaDVwBdSe4gt+ZNRDA5FEYS
cjbClTPjLbvl9tRKqa9TRZ6nPwrk2mxvy8JqvcwQWRL197AJtH16GHsg4ZdQQiuhi3zU7+GGn16D
cjxQFcLNRNiZq8yl3HOc73FQ+zlmx5xkuk+aBvBx9etbFqXyvADM1Eq+zmayCLgMY+5czK/mCeC1
g7UQA9bQUMDIfMElr4Zzmzh0o83XhxYgL0zYRJmJjVd0F+0GVo4BAmPxOZBRn0cFeSpKpQAZ5+0e
YKBpdMgK8D59oxcA4Kj6Shxzllm54CBZ5C3ELAtFVDSSromWPIqrEjeObBqqJXIbq/RyJ5lzu2uD
hDXGYYwlNEqw4ClENXRfeD0tOsKe5QpEPdPBQR7jneexJCfGvHnusyLLKJJLaEILbOkg/KvHh2bK
+K5SIDZU5THOPu/rArcyv+OLKIQH8DwGGuKE8TjZN0rxe2puTBWUsADqvtCbE9uNITzIc2wSb2LD
mKpuZ/04yF2aiwRKz0i+mIYnHK1E2mDnP1hqMdhe1nbi+SMfdrIX5DrA7gQR9ki38j6EKB3LtnPn
dM2TnCHLVIFz85gYieLE/nmZJ3fJqLouJ4d7g1uXWyoOUeolMwm18PkzeN4NVudjdO6yHJmQ4lo9
pG9gbB6hehuceAf7ZfJtHD4s7QEcs5tikHWuuwWoxRxAIRA8g9Bf9M784xcw/8EnymDXOgogNtGN
Tv8HgOzinypiJXEUZpqAqT8sARpmYxE6+Do7HR6WQ09gwc303FQSRVm+P17BQm5iKKvnXV2CMsQR
FCV+EPqU1ED4c2mCxQYXWuZNkUgeCDUkRosLSgO4YDFyDc6vg9iDsUUUrLjGLeTTd1iRof85wGI/
k+h6jIBYpnNlWRTmfvfIk0asFocf3xAEYMio+xWc19r6bFnjW7f+87o9tgIU3xW4+pUsFx7nWdMk
g2fxHnqVP6O1BZaHxNm53FRdpj/vx5dxusdRXDvWcyIlcvJJOf2BxyAR1peRrubJPF9xdTUC00f4
n1MySsZd9P9YyU0CAK07s71e8y6d8i3EYwGX7jBlViAzOoHS7eFqsEmvCLQh0mDORXNQ07ws5pjs
gBArhSHAk9+Ngf+oiV8OrHccK8tabQtT2LM/yFoRmLHlQJO5FeoSXFXQV8i+BBAzVpvp/p5S4MQu
E7w3jLaR4qpLzWNVpy2VhJAmKU6LPd/AWe6hF7H+9VJX2Gfe1zGzqYb3qRRgYGwsffnx9dWvefFf
+QvsaBSRqDxdC/4K1dvYM8Pxc2UskqewlsPRHCNiyr8NH3wmLJFYwTum56RrSWm75Sz7l9QaCnnB
pCQEdr3oHRwfwDkLWSdYZ3EtZ7tCxbWpRUR33Cp+qG8lOf5diH5dOCrsYZkTLRKQzg9dF9nhbcEx
IVUmdDtHRU2dI0rGozelaf6++BNBrhsTluOPLrCYWsu3eu8vx/7ujorSgP2U68Hog4WHZZaGuZ5p
j4E2uor7ywMVDTDXRABFC2a06QohF4cn3CX1tZa4vDPEDYcUJvjFGJV+8NJgdJqGhuWNn8xKpdX0
wPEYENo6nDxlmP9a1InGk9hk/7lNfde8AZYwoTI4cVraswkH5IciQa0nwFPD3SphLbrMlYvyIMtN
huxGLWEqvCbvrDdy3l/58iZUweyND22OV5nukcdkJSefN6bSS6vcUsX/fTHhZvDk1qRx73H7sVAD
AcdKv8g6Y9QvGtgRAc1M8I4yYtS0lCKnPtCWLjGnheuDk+c8x6+JseHFWUkiwJEPV4XAjjkmmv+F
WGx9geICOFlTuFL2knSJ841jY7BVmI2N4mu/TazC9Cn7nWUoFJF5JiBW5txmicGRKIiDu90ycGy0
TJAWmHW7/Zr6wdSEXaNBFSmBbms9kLQZRevYueJirl6ay4McwJRYlQLOAPLZyt5mSwug4yetyhGd
AJZWTnaaee8VlEsTHJaSTIaE3Wa52kMY0Ij8/eW+phDcC2LjPOipGkcQppVxIhQ9IItSGdAL0Xdq
PBkqh/C9HueeCDzvQz5B+Dzisxf7Rv0ThHzhdlmn56jU9FSup7z7V5RNql6W+gXoSM2L5VJwXsP8
5ICJ309xngfMnpBWi1R9uMVFvpykx+qzzjHfZs4dwywroezLc17pErXCqXz9g85C5Ld7xzMoxBDw
DZiWCsrPo3VJ/+/cBBY0acPS1eaLno1wX1liJfLWAeBB1pDKyRvLh3mOuUNpHWynRfu7x5hgZVRY
Wgc5qgPKaN8WGjvhIyT32erxldwb7fvhDPqc6RGHtl8CmXFppY+dXyQFEy6uKVWHJ81fCRgG1UPr
CSDcU18P6SmSY2CK/MbiDrUyrw55iSGzBCbyDjFYhHEII2DQDkh/LLdPTZNqrSVWaqLQsYis572I
1v1JG4AlykfIcWZoHNm97MeHjl8pSuhYdO60wV1wtMZlPCOWLVlcgCKzq+2A2ypUuAJEep7uFSdm
DSPcPK/FwX40EXeOIL4InyGFe/Xm2WWU3cIbnt3jTWe5Qoexk2LZN3whR3d81LwCL9SP0Na13lId
lSHJA8qMeYP/IEGSODm1rI/al3imKBZ+v42KllS/9PnHnDUI7hBWg8B041pW1OJUqeQ53JMdAPXW
gaZb6q8WiLAA8p0wDEAjH6DrDuUCSuPbdCmgu0r5VKIrFCokeJdvFmSSCeeM9GVZeksGSQ0JEpZT
ggZrkEfEw4dM3i/TU7xwTjg+S/xQMg6O6VinG1AeEiBfCQRa7SF8DG768p1cwlIKjNEh7S/tz8Or
d4rQzpgC6QlQCvuW7U8yePMUa6a2kq1xMsGmVtAXNJDywg9+uGImKAzu2CbMgNsHfJImuWJrCbEJ
ZcKhygfpOVdszfbT9wDKptm1ZAa0doHp3TJa9tnH+RybJTOul3SsLsqiqM5McGlW4+puSvxOyDDD
P7OAQA8Kp6gEBiq5VH9NuOM16ncO2Ia1liSj88kU+Sf66STAjRK3Uf29NK4SzlwEz0AYZkSPYuhH
DP60kMgnYAkVx5srrYMkllS3wHnvZGCzk7Sgt57FOPOM+sUA4e4VDvEw3f3Z7Ohujmv3G+9yqfgE
+eZyePHqJFQcJqoGcrvreF+mXv2Xnilm1SMFgWCLEJAy1Djf21dqyhmm/e9aVpegpW9TNr3Bmgia
3DCNORFTVwEVyqmWJCilU+A+hhiP53cNRG8s2lh7FHrb6eq/VhlKwDi1KWhlXbMW8FWjgLH32u1l
2sDxG44eBXhHDGxRiC578JaTqr57WNounUGAunuQpDOEBJhjE8lVILHnzGUB1XLlPyfd9xWY7ULo
O0Vz6Zbaw7itQgQOtfqx5UzSZeELFa7yfDcqPtNWyljsgJy28kvctvF01aWqVkW/YiNUi54NKUv/
RRv6C6wXLDq0n15uL2cGuT9GO9a60TXP11u4ctGiv8pGBF8aABDcnC8HpsU28GSoX5y5cz7zJ+xm
M1mnZmhWo58RTVhyJnFWd/LjzsvyqUIw0aKKEH1DBw40Kcx2HbRqDld7swnnBpgWC23P3FTzHkX4
tfBLCxA+tW4F5lVUKf3V8oJgwf8OXKA0zxEbQhJy1FXshB7HQbJBB/yIJiVoSxmnT1i0VyZewfj2
Hod6jXSvzExxtjliGI03y1W8z9g8zVLte7iys7DTciiVFP2lUzB/G6r8zjhAcubabnA5KuCfAzUg
GnF47uRVmj/PI0bJI0QWAyjKlh8EBvR2c3UxU3Q9kANUkeJhzAmjK0BD40ryInDWOjsKR9fd6yFb
VNb1rJbUxGNaYpz0bn7Ta6HROB+uIPZO0fgfgieWRRs8xCoGajvYR82DJRl+6X3JEnNd50T+/biG
yUoDkgFKMKeL9V4gcau/5kzNOBb7nFUsLm08TSCAQbutnzvI9IH94eWE8xMKcvVq9YRfxI/YLee3
RhKKVezcwRozcdvxLw5X/Dc2qXcG8A8LOwBrlug2AiLOSMGAfjIKbXIv/BPJ1mAsId50VINzahKa
OC/GMaI2IPmEgDSUw3vNkZlnwXEvyNMToLjzGlGCKKjb5f/D5bYfZ/+UEAEIohS77aCTgBUslmrx
HKWo5IYVDOJQAb3D3dL9NSstfmcXTj2yHVRxKMV9STuzZOztrZ7ZwlxBvLDSt6uZO/uLXm5ekcqC
Hi4OF6D+XMOFo389k+WpoYQbPfCnZv+vkHy7XiBghLgObiZFTc4oABHXiPfqls9vZ8045+0bfDP6
7FIsVmRQ/bK5Q25mlM4TU6IcDMmgH1IRCgogsJ6WTEskfea1ErlrrbvVvpSQzyPT9Jm0WvwCQeMw
k8qCLWSYbT0Q7ffGd+2nyA0WXh7TXxVVWLzksw6m34vWwzynxyyUuc+g7cutA5Vg6N4GD+/s+Wq0
ijYQR9/N2w10z15b2s+zmPDte6ar2sl6RavMY4QlBT3AdW75SowXFwYj+fAh6RsQSRsPH67bK4Wa
odU5r6jjD9yU04lFnad/HMAwhd9rBSavqXnRB5Cr+aw1YUQXke+JQ0qE5fvwjDcdYqgqGTabXrWD
1ZTyS9DL9KA5AWt74YeH8uWcw6Ys/rO4iLRhleA1wnn7JuI2C9iGG7gftqm0H+oNw18za8fIUGG9
vVOr1FgaBmV6uMwfE7hfPTfwdPmRKrh5XpPp/krQIsofRTPsVnz3q9n7zYqpU63Mfo1fWB1Z3Tz6
LkKbFeo1aKIVQP188+w00AkDgLnjSRdXxY5LsGcZV1hboDzwWBIdG5g239TZ/tssxtaVDKZS/5CH
d/NM6P5QxF68MWK5bQ67vTPU0o36hNkbNXZeMjmBm6LoZu5/PcqPGUlbng2vuIbN8b/V70BmfgGk
wEQIEG9tW8CsPK+cXC2OBKlPm7yWEQg4Lxz1CxghfYgCNqLMB2ymf5CNgWS57VwOfTxyYTNU1kde
cwWV6ATPvo8+XuJL3Y8PoyD8N1fWMD0ChsZKx2a+CkvEaYdaSa+JEEOkXUyPHcgtPyAvGLUVzxdQ
Hoz4/j6eMXQ2L5XXBMXydyGclqPT0x0solIUm/J7HCW4RJ8kCr0n30dS88LBSJKOp6x9sJcRrLPF
ex/ZeEPYjG9KyVO0+wNXHLleJNFZGvqVqI2EugB4r/MARXmC4qMlmrmuN7LxYIZ8FrIkxrnjQimO
QfNRN0Cplq4YWwPqdQOmSFHyGAjAHfzDKiogSdAPRQBK0vfMJ2L3VtxjOWZCY8Qf1KbXCrMaOtLc
PNmmkDts7O1sSGbaNW0hE9ekcfhiGdBQuK/Ch2OBHcocbRiXR3DRPzBreOJVjtoDqOLiE1g4wzCi
JOcCJ233YOnreuEcIc2muFh/v5ga597wEvfENca7OSUI6LRb8qd9frzRBcGWHg4K5bieO9sCNKEb
ztnEGbnDcE9Ke839mxG9Im32Qipha15TtIvsaaThIMwGYlwmewg4K2YNeSXFRJr45YaNFbVU4ZTK
xuB1lHFt5Rc9BT+pkEkcTO4hMyqIAXlC0jzmuCHOguoIpr9rofGNSRcOqeEOrcD+UdQyJFyTJ2oJ
IkryX57uycnXSVU506ibL83oe8EUS5aoH4IUJ0vxgDCzSsn7/i8QyIzNAeQFi8XVy7X/OE4WhwaR
BQJKtzDlwKfXT1mc8CaFBoiwDPovmfoIqs5VMeNLVwQvO9q66DwXsds49Kej0sRgBl4nl6KWaWOB
r3RxmvECO/IBijqPiCg7sUYChtFWdJJJCc6Bp00xZN1Vng9IYch0STSbk1nmsZnJbW3szXeTYUF+
Cmgc1zB/RcpbImpAv3VfJtGKIL03nGJ7talZkd2zkLny22HvXme/VfsH+D22MSXKWALoUf6gdQWo
K5rfQYs9xaKbQ1pu4FGFrsmmr7o+BAfEr7EClv7CHiwIrBZ13DKvu8tQXMhS3EQFENOFvJzAwpmO
iFVkXXsRQQL8Dl0BD02WQR5ZMRNDtaJZYNXd0Pj0pHWIazGAaJqHKmDuXt0M1jgyKinus9oxbzZE
em3xf9XA3MUTrPqhM2SG+tU8AqHQyE3rp0sjurvXZXot/Tc383sB4t4gf7XcI6oxUqSjB5bl4MeB
p1c48tYeRBMcu7wV/nbeRkqXJjaz4LtZQuzKwNjuAN/yAyw7ll64A1mAEZNgwMr9GF0euUOqsYMt
ikHsTzsW41CyRmyyo/Kns1elIizmHOKcZ2iuQYuEdnnSjhEZlUcWb/j/ucjwfXOzV4kVjUiHAsQS
rnwAV7UU+5g+yi0Zh2jVl4Yecm/8lvKVpPdTDNhAZYvKajsQpiSORrEGwPhnPJnAQb2CuKjrU5on
zU8/FaP+thjkwP7JNM5toNnh9zoHucgSgqUhvWqlb3bAZSmDi/WUCumo9x/88yQ6slmwazZXUIsx
9SDJiXq8V+d9HlJlo+HKJmb0JnhymsQpQOlk8u5SmR7ufonBvbFho1ilzGMd3Uvv4fd1lM94NWpO
OXPfDKZzcZWxv4U7nV8OtQXme8+g6IXbtFvAjufv7GuN8D32KWg+1nJjZy5fsgXyBijUHbgyDa1h
KqmbA0j9zaXRu5inzaG2v52tUYF7U/Sgdm2p+yMnlLdq6wVi6JKaiCj+TQ81c3m40IFJEbdVRYr3
BM4MmoShTmmc+CkD9wS+CklaehnN1F+qLoiI8j9ggRFoJJFqbUKI6g9zrs9fJVuXswgEZInlZCnY
V6sckzE5fMSwve4x1J3ehsqEnuFEdjdepnkL8VaDKx3uxwVIU+SFffCe5bsTpgIXhCBhJmiClumA
SH2a3+Q9nnID4m432sYubolKjhm6GNIoJyCxolwWlLf4NbLHXV1EL2UHmaN7xmjJfOybk1ICUbVX
EvwLU/cU0z3iannpjJ74iDxNQzBLNozb2nLmL2TPfVQR1hbDXcgSIMrsYfS1xTLPbNtlyvIGNoCX
lqMl+3LNWy4KL9eMxfkWWuCMYU4MwIh0rhKGkLdT4pBTqEh7QzGx5A9vw1Ie81pSwAvDQwdpVjuY
4hvldFyUCrjuMz6w7GAyPVhDIRGkfeUJTnU5I2It95PA4rH3JFDPSp0EMbITv+Mc6YtkXbpomN2W
GNlPhBroKb8FStJGRKysB2Ze82awQ+VxOjI8PtFp66PdILha8oTs8F0BdH+Tg+QF0UZBHmEjNM8O
jKoISQhT5ag1OSdc0OHyavH47SA3CEvnZ9N27dCc6sLZiwOdTSdk/Gsug2Z4fxZkHoY6aQhfz/Gd
8wWvBbrtd9Rg9McDiyL+m2eLwhSb4vUXJiUuXLJH5q2/GY1gGvjMn5eoI6RStLxj+F6az+Ej/qDt
YyTd2rz+EmcWDG16vcwXIzmulrMWts3QEFIZGZRrF0o/uUHTszGmx47eoT11AFUQpdC7vqDDDK0+
FeVL8pQ+Ei0Kl0axsIip3EgbYl54vAD9k3Wgh0J4cEnyAzy7UncTVj3bN6Gyo3GH/ocftme7nIvj
Ly28EAiMz5N4R6pRl05GUeS+f2tqJWa8ZC5aGvnMH+MBTz3sdjBcrvFv+He4+lpKoepggDVfndpT
VJ+KdG42wUo7p4uARfd9COaEzKo7WJMqCTsNDgJCheVjTeaiQfiQrPaonuR/7aBCdw8NtR+tzw2e
gPzo1wPA/yAZij0fbA37cugH1MvCQyFGpsEGvdjPxtvjl2+j2Qii73rluIFBc6EZUfBV2ZWpGzxA
3f3YZu3yERHMtPO6O7SxB6ywyb8Kx3HU4K213PC/H+tvlZaVY6qEuOiXuYx/DvdbGBI/PoAscynf
9WL+52Q9xc1kNakyPjgVNnJL+e0iLVDrRJ0lUWOarmEJjKSe1kfiOj2hXbkbx2C7FrLBOkbcY9vN
M9KuioyrAtL71GpcyDv6cauhlyIgXc4e0qI1nC1BW3wJ8rigyQK2uK/BYQSyw9mwSKG5sOzfGJGF
l0Z6qkvyEloPP2YXqUkKZSB5jV4YO01YT36y6Xl75aqXW5eAofnzqlrZB5MGwb9lSkgx5fVvf0/Z
9ODTav54zw1XrccIZgNnPOJY2WQ9/TXN9pvKUFfp4AiDzBg7yMuYW4KMgi4nZLguwczW/FF/RivI
FsoOBu/GIcA8SaqcSAvORaC6xcDH9Lg/rePS8Vk/Em7LpjtPVbAi00whlziF2WGVTMbaUNOUPBln
i7lAC6Rhgoa2dwJVP+wqgRpPoL2XBiVvzcD/Z2AXn8Wxi89/7OqOfPv1lFLWnfFQYxhanzhvXuK5
itbMFZrQYmkc4/vDayZj36SyyFYB3fURm1JqZmxqOko9ddyUv3tsRWa92HTN06+xy7ZlLTnro5y8
6oJNF0wfYnNY6w+5A5EOTVrIA0zPg+3kPVWrL6sQMeyd/scFA37Wp5xbQTUtHHgOOQ6qkXoezDVD
/y4J1ykqI9by1IBOV8VTuhO86mwgoVJkQfhXvkpte73rrIcCbIZo19adD8CI/h/lhWMl4KMsd/AM
8Z/7+BKRwJt4+iZP2ntYv2DfIbZIuCbiVpXC+6Kh4TgNZZ+Emo9R8cneV7nHIx1K2lmgxkf6dX3C
UBKOvm5lqMApz678JnHGEZ0IEd8CqaOL6u4eauJ3Jpm6Cp11TbWTAnjLn/WZQ2PCouJsS4zowYxn
ozB9uHbkcKZ6B3HXufEX9x7Ia9pQi3cKKllg3XqrE55FTTywlIB2ojMR4hcVb+goDhyOiR6sLlsh
LpfxQB0PHfYbEj5N/uNZNdpwLbo94nNLXWxg96Ru9vkmooZhxJWGCVukWtPE8+/5pQ5MGck2rFSc
WMxhBDPdVd4jqycE2szvlaJalwZimecHMRFSx2pmf6OqbCYtz+z+voL4uZ3rTHeRK615NkCbrWRS
8piO8plWQLAsA9XBErfvWHpCevIx8aGwNRDQiOYsdz1evRXZKprWESOD/CTLWzOmCFClG2+izqh3
IgDFP/QKTq0uDVK2ZlfAyf3GBuIHDVlz/TU6270cl10TN9EDwh6oBnMf4tfKGkCyJEY52y0HAj61
4tlHQyyh82EkCf4Kl3Ja7I4U5Lq2UPlvYVTSqkNM9j40f73Q8UGAJUh2/JoUdcGPfWvKFuujp0jl
fSTGJwEkpZezKAD9ABkKuJz6JML4Kl2iDkA2islM+o5JG3pqTTcOrZVGnQr0qndMODZaA3aFOM7l
c691brLsE+b8J1sk4Zxf5pxDsehwR57F4rBkH+Tqisqh2cKbbBPcGPNo8GC9DcBfwIHOvGEX2ZYS
dfZ84RophDNLo95S35aYyfLT7XsL+4sAM4yzd5h1C+NnVKmXImJFtypVzOsF4I9EsVKIIFHhW5Sm
p+c/B7Xm7FI7SoySrtJKI0eIXlWq/nuUOKkRUhXtIcgY43L8LNq8jsVdvg4x1Rt4TlDZRh/ufLQz
rF/Ahw7DNlV9xYXW6l/1bLUoMSrH3mN0b00nNAC8M9qSwtE34f3XafXuKBgrtIOq1O8te/Mpt6dA
daq0SvDeA69t3yIhybknTKeqXW6S8A9GkESEwxD4CQWUbFgPR+IliRmVJXDh6WvUo+jvtXbh1p85
Zdj51AOpf2zJNSy1cTXCoi7a/0cl9DeA1lqLH5kd7o8g1BQmmM4MlMADniku7AIBkjlKKuJUv5sn
QWt49hvJg5eZmRPXA9t7wO8os3OPWlj9hFDY558io0+RfmKiKiulpzBDULga+vKg91yLa6r4t6gh
3Fgjd9eaWUUyPBHwtv1q0xExyJA7J4dzYh8emHT9Eh83tZa2j1HA/5UEyBvaD9AJSxtpC3vICg8l
hZpFcfzP1L6qKn5PEmEIz4PzCjuX5BFAEAOWS4t9/AvLT4jgR/c/5SlfYHnlk7CnQhc/wn7IqdFX
eevyXQe6iFeh2nkQu6QJury2pKX85Ddhh/kQjL8V6wZMgG7aS9ZQX3lFC5524n1OPKCjNnLpP/Qv
GkTYKUrwRCRVYDljR7sh3sfJZft0kVKAArRZHvOApad9A2vd78yVZyHKosVzO8fnpUbncp8EmVsb
aDiIojCUJMcCQcUuDhz4mZyeCOr1rl6BWF3TgQV/iguGDgD4oRn3Ryd93kYPADPCwhCEPIL5BleH
xQ3QZpJH8SY44/CCJ84PM6g9pe5tiw8Uv7g2K+9y+1+N05dksKBe+5zvtmuSWVXvYrVdaqxQ2Mjc
Jm+RcYAaAX3NlCBaP55Ex4gHwyPoq8t3RPe0hVECO5EkspotBF8oWPAI4Gx/lJJ8RVfoYFwo67u6
6iUrxLXhLcW198TX2wpY93/9rQyOEdxAtL10ub/mfR7Fd+ukmCVviN1f/1Z6u6BfGDToQsmpWOie
d0dMYTG2ITwYtZeOUD7VB+Gw/SckvkQQzI8HjCJU8oVM4UBsH1eIqIiSSy4dsDyHolb5aXP1rO7t
krQSz8/hB/jxFuz70N7T9J3c7TFlrDHikHzc7ujswd7db5pa7QmpZ/neBIuQ9A7YUQ96xeuv7gMw
jI45CUrs285AqyFXN+PHTDQ+GipmKS5aRdzC9aZY0qNSBmScmt3EheEtpRguUL1UlOh9jOJ/ZQJW
lo3Ehi1LbT57mvwVxc4nhGVD3usQnYVvArlglM2kKFBn9vug0LbuS964ulFl/qjBZFHZrH445LfS
P2J+pUy362mh8Kb+s6LP+ZHThpUgqLoZeCzDbdCJxdogU4hCBK3ehJfMZsDMzJoZEp3DmksB1fgU
U89itb0tECxlV5afUakj2q+nWFrxHZCfoOB583GbbPtMsb3i/USpMyrMZWGsDBm4e8jFRPwi49Uh
WOlNCuY8VPUZ90tmrQ44nAU30kAm1G3Oo8qlE4UUM1KCEgXcFn1MRtP0pZoEBBxLNmRmRb7Q/v5c
xpYP6mi4il2IKYYJbhX7u0FqLsDZTqjuZTFTukMzi79IM3JIL/PEJ4nvFPtKPxWCMmWuZwKvAYct
6b4MhqqVHDL9LcTxYdchpOp7G9hPFJtzkF20N8phUaWmXQWsMBoAhgG7DDowqGhvc9t5nbKylWMw
XMr2TgUxUAD3jwdtxwyDiRIqPaABkHT5GcwfqrMqaZD4jyGGglKwCJXZISP9ifp/Hpuozzm9ypIB
qdBesxCro+0tKGmPJlTpAobOGtRgLkwATO65ioGUKC3+mXyNL3LyvoyhsYtVEVQdQmsuqye6q8a3
tQUrXFCGsyro0iJHhiD0yW4Mm0RWbmkcN0xjzDBlSwW++lL+0jgvnXw6IQ3CpBCO2z01hn7o1dQf
nXMeVDmwpyzlu53CHTOYBubHOKWw3Ms3OY7EXG8Jud342ONH6tjU5AHwUGptyWHvYccCJUoe+Pal
+7U2eOwsi3GrF/R5dhkzG8+Vtgj5mEdn3oDYeXnxakMBVKVH4Cau6Jv2WoVsGw8GQ7YnOzrkNoeH
xqI6V4r6BiUGk3WKKSJZzRQ/HYRKOoCuLIBapcLnDG4c06pkH6Oqfne+fmzjkTMgIFYXqDW/WJN9
14oCKIF5ybdkc5aC9b4I7is7PVdl/LatepWo24QXKRwVEDpCm4F+MUpdLyQbKt3guHLqyxxtoT5d
ZtmZbwaDJWsilxh2e4b3LKaFN+440O2BZ/j9nKB2kF3tpoLkoTjRlC9SXxyOGd0sn5ka4qjh+twZ
fjXpTgQHwAp8vH2Zauc0ZfA9BK2wnHyWYMxZ5uV7BAWRL1FYOCR+jcwSqc14es8Qjypfvf0xTlPF
qHfN+MIZ9HvGN1LccGVVIo66rncIeaayaVQmBJD5/+vFMtfY6P+i2xJ+QNJSN9vxuBPQPpadK8/U
3pdU6B30HoxHIlf1XAylGuRasRWVooi/m7kCMwTxP2IDFQyK6uhtRdUaQVarMR4N5VIr3aG6KVW+
Y/wARc/0723OLB8VnZb3EENB/7CNJnC0VquROGvWVQeeLTff2PxtoYBSWum8s3QXR5B3vGWBz8l/
P7zViNFuU1m205WtXJfBOitqDkQ9fkJN4v2pqTmHkLbTw64SWpuzTqGeUjyKYclQO9c0ebYH466A
Dq3Eo2ATqkyTXubpYpXILVxxHlwklKjiiF7W69K5sDtG2BPLtyQPDOjJh1rBQ5HdZmt4GK7Lp7LX
QJUjyBhyRrWxF8BTVvCpUdkljgz+ZNMQj3IVf0YirSPLlr2rtejtGPNZ6lxiBnbOR1aSk4H6iRC5
ajjCyoj/3iUjJpgwPDdtMkDdSiusAU/1r3aJEJn+CsO+a5RrCbHl7m1cLC+/pKiS7DWvJP3D/M/e
GwXRKCnsY6pTeAHi8sOsgQkR2Ho58oCPv+q7vhQIMOtzX3dXr5Ey6N0farR/xyNp+cPuGj84qiQc
eZXTd+sLFjMsFp0w1DIvvI18fiPCdJhiwmuDitgkmt3nBJreR+7gpgP6umMBrYPHk+gwEw/KzXhk
bti6tt66C2/oOuh5cG4t0zwREcmMCXETahw+wdvX3ZFlg5Zs3olIPw7SPCnMNGYS6LNPLkJam1PG
5DW8HroKw43N/QXvwcnxcqbB1eqVVQsoD/qvEn26twglvDhgx4UTU1hvElsjlWMFBecaxAr/bLvp
pTD8EJxa2XuWm/pBwlV1/WDMzhbeJ7k69jLpAyO8/P8vlGi7FQlOBEAKmhVLSkF7f58o2piv7kqd
WvCyxjTI86tAQBf3Y234KUTGmw4HuLPLfrjWQfjJo7tVKR53fzxXI0yzZmUItmF1wEMKTfTuq17Z
DGdQatMpEqFQpCfybySSgjNG4txAjWLDlwONdlRKxE32WlYNAVDklwsv8HUwWYV8/3YgcpbGmGq1
wm0tW+aE/V2yWmIoS/4YfnDymYNtZEDGIYg/BwrGllPXM4lOXt8fc8kk+kDys3m+NalD4vmeS6bl
NyQULQdUOgEq+s8QKlORbiAg+WSBM0kFGcwX9EsxokyuTaMwqTwALYES2VUMKsN+zI782xD0DUS8
yZ8GzGkg6lOKeQDbSF0w3Ee2W3R6y0r90jCsQ1kE8rD3nJCeai5/DwrRyEauZJ0uPuYeOr6ZHlhj
GfiJWrYlNUMGPJ6NL9+SERJi8pkEeXHSo32RZjXJQnjfFm1Dc6F9fnb84LlfLetaMQxysPOaWz5i
n1AgAQhW3M2EVpsU6epNMJAQ6Q2/XZDoFeewOzV+o7YLPrTQgIT7DvDhvVsW2T4nk6coZxGiAzlH
fh/eILiVa+AduhakqVF8albrJzodRN0PUPQUpyUTe509MgqTJ1Yxe+BxejI9x9OBdCVniVQqtYbw
Cn/5zT9Wxe6HUaYql/X8F3NgQS3MKyxDtkekwfq4Szy6MMivvEGR1J0YwKUZV4S+qhfcqkn5bw0K
y0R17VwauTX83H0vt9gBeq0MKeeKV8lTGQXPNmTgHXnEeibOigWEQGFdP9FtJYU+yFVbnUuFOTjB
3gqScXgYBURyG2vOazrF7a8LSTWIYnCJX/V1dJb45BQqfw+CQTa0Wp6+5tBx81q2HwPUcjXxWwg2
T/V5WiqtGCgdVxF/Yb3F56xqKq/g9NvGu70nlpSTBPuDxet3SR3zLvrbKgJkQoQqRuWlggXKn4Vo
1wZ9ruIxNXMW/lheHxALHoZMEXL2whjjL6zW3cRYgO2OuSCRW8IL/d3FG0nviBm8fB2STBErnOp1
Fdo4nAj068RTAQZ4ASzPzSKhE8j41f5xFjOc5i9ptvHA2/dgjrlfGwzi1rMhELB+OcxhG2e7+lIL
QPI0I27BF1mKP/oxjzbvJ6FP6C2yvkO9anu+Vg70sFZTCW0Sv7sP4SLCJK+g+rn1DBMmg1y1SJtB
lSbhNHHUNIRH1DhOm2XfoyR13prgOMU33QDdkIeFRXyYPIznvs7Q+DnA5GglbXiRRvZohUljjpzM
OIIR35u00gfTuy7LK+cs6tPEFhp/eGG+lSl+th+pXuqrF/NVOj4hTokdXYcy/oZTjAPPcshuhw3h
RF019XHbz5IbVETqjNQo/MjsXgHyTDx11S1UHMkAmKC3j5JA8D1dntZfaPdQXnZ7ya/dKewFXpe0
39BV4AxMIyTdBntQEHfNHNyZ4ov9kREoEuqMVB4EXZ19RYWFtDMxhiMCPYxDFYtbAn5f0woUJ63j
4hVhe1guDuS6JJw5Mlk78cemfgIaaUAo9Dvzcaxxfglr579MlVOBhSqh/waKH/3oHCjrC/j/DToj
s/IqfNtasOv5fOQa8sAQWYFdUy8qgVUBRyJiKnW0h9XJzGUdX8Wud3xETOtRl+qw5SeZxhOvi02x
SeIkXx1/EISq81PfpWbB8yELdD0la36QNJK4i7HLr9x6wPYInhUdKqGCz/rI+o1cfpy0MMPEjpmY
SJmektqxFPcbqhc8S8dytyU2S5iWlVtiJ/C2pMcnrqq3PY4weG12qEeggDQufsmPUJ/curVUq5du
Fc3M5eI/jvfgVXW18EfMNOu23Siepk5UC3iH5Ql7m4Tnn4sxNjxpvzGx96G7tdZjyUlceQuphdyl
s01BhMVjC95brwWADdVMVav97/Izk+rGHI/LLiYO3bRaHKAJAzjk/mtnQLHFgbY7dLkdOhRCLh72
FwaFSdM3kA9juKgODxaq9YKnQ4CHravDS7PWlZ9l+5GPmJPmyfQYqMyKOBQ+r5KQhoAaVDulTSoP
RUPO/hvg/gxvjrucagvjSZoeBtKA9PQFTYieOviOQgwhhgJNGFKNU2OoXwwnyYExCfTIWbL3nIYD
spdA3tlx56/iz3Hmno4a4AbxgCB17T0/kflSsMdr65cBoV4Z/gMlty0eVEba1hviOB59/Edne0Ct
FFsSz/5vU5qcMo6RKZbjtvNFYCH+fgj9JqCfxwaObO5ExcBA90WFMQVyn+WVw06PHQoTd7huJ3tN
htOVprIBhQCe79dV4/v7Ga0lHd46hpMxI9zCgwt4Yk4RKQM+Q06VfebIwqtanR2oMP7nb+SKykik
xwtkFKQWgK78YoJ3DX6GQ8lW5cIWY/F1tU6pFOpF+YRV3sMhYcijFTkr1Wt4jtumIKosBucyHT5V
70ZsErpRIOnK5yFONmR5fVwHrfat4oBmT9C4qBGK+MMrRfss1FI2I5RtGE/cX5s7zJNGbgLDX4Q0
e9oNJPI/jOwDEGjLrAdfUkrBAPCfkKKBl8g9xaI/fuJemZG+Gxj5eS6rbFMQFJkiOwAARNS/VHdT
Km+jp3UYWbhC57l2umv9cELob+no/Pt4Rt2gIEIQdFeGpK+5tmzRKuyXpSIPYehfsXG3bw2KY2oN
Xe2xIvBJu2yt9sV9M0MS7mcGdtgC59tYeR6vZCLAaGrHpPpXeKhmE7qtZwsh49x4mnZmcmn/dzf7
L9BhHwuyRPCt08376v8ShaCe2JLGLVLht+mclkNyiIMYEoN6nXXETwffcAudQCIjEwf+Yzp3f0PE
wONSv0Uu/oZ3kSlKTEfEr8PsqTRkhms3UQ/vbzpUnmPIgAwYF+HNfH1wJkP8LXsbHVhT4FAAp7+/
abSsKD3Wv5hP4e3HR8XIOxpFr42LdKTRAzVMG61uXb8Q2ULJcze37/1cxT0vPddqjHZy1L4jrcEF
fX3VMDfXSg/htM46y6fvJiPnK2+ggfFkgjsj1DMQsc2+NvAGzhXwXoNHUkv3Am7WDs7zhOLuIWTL
00HQeLIn5Dy2ZMsnwlGVVcBM1GlxDFx5vg5XHjiqKSF2NO9NCopebDO/3E6ywTjdQEZayF97KuvO
iyt9hKSB2BkoCsLBQWdSyok2On1lGof4kRUByZAFR4diIFwtyAF5SqHNE14TjvHArmV4clD4fo4S
1ZZbRhJDLwQ0VYK5vjV4uCcyFQyzHQUOCoMOb3PTj8FOLkWdPd4W9hc+bKqjh2Zlnwm75NTa3SbL
zH0p9c9b48Af0/Lsi1eRpmLHvs6lv7NwX2iYrqbibJ2RzSKnWRZAESqwiva2dVPiYBp3J75T83GV
NeN6igx0+Nsx+yF0W2/QO9gdBQEvAg+YgtRlK/YBk2RaJMFJQoMWFNFkJxXH+KxeHNj31ospCgjL
35xBv6soy/WxEn89CyJyAfQ8RdJqvdcS9Vv87yod1Abys3lpbEsCj8Q+znm4v+zdqvFhRr0ZwPxH
2sVXKIayxGTZw3iJq0QkQFo9hZ5xtsXM9daFZmCHTY/4joy9GTzaJINtGMf4842IYOa30bejTyiS
EYtteuJpWyUgALky9vKN5GOhacEBNxkdQ2nELd1bCyRflO5M7487gWeoSc8nMwi1Dt3DqRxwo6oQ
RvE++F1s+dr+vpyYoht/MqKXwveMOymyDJz/Cw4tV18uSlptwDHGM3muJD+cpFg6u6ri4TWDyK6a
bcnvFuNF1Pz0UmuschmJEwDrsumH/t+wTPcLMPZHSNqF67qW4zjFH0chVLgeQA0O/XQLdNDBxavZ
NblU5HMAPb01WAQ4iJKQLai8nVFcqrp/RehQp34/6LA4p6D4rfQ5s5oQlYr27NOg/5M1OqTF33EA
g0yGKo1r16QL8tHVXWsXj2FHN5X7fMik1z+MTwmqTv7FBSeBiA4gMa2XyPSyJTfkO0i9h0Phn2LP
CmwBesq9RHGrHwLEN54DYOJvq4dQDIickuc4/iAbaVMfcUFNO8c0pOQJRTJMuN/Wh7RTn3pO/hNi
zL2I+x6FB7RPKGJ6Urre2eqPsqWScS4EWs/D/r3di9m+C3D/ntFKrWhPlGODUEUO7DS+CnXGidoF
ZicUpC8R34Yn+/z60IsjxGm5wbbBdilW0DDCwJ351zQsExZyRO8vs25Cn1kuEaQq4yqpYrje577l
A9Ux4S7IkVA4WqL3YeB3gRIx1ffYJ9sm4qoqDxiXth7CWNdHmFsQKt5u4nNRokKj0gORYnWu1qiW
TDmCtza0bFANMecBkMWy54/1ZADyeIRxQ4WiGblgFlHq84JSxaGrTb2pay/GfglZ4JhICrpmEoab
HJHYxPu8qhnQNcoqbdEsBMcz2vA8fSK156hZ1MTYc9ArvDM/xqLAXbC7cpchb/sZjGmjbYN1qzOo
+QBKazEFsiMpxUvxCINqXyIqCX6CPl76DcUHme54mNeQb13ODJXR1iS+thjWFxfoEHtmjtaLHN+U
O0AsCcIRlVN/eLdvMlKt/0qCE87eW4eRUERTtbjCHhg1VH/0VwNogz5Wa5ktMcukilruwmw8GCxe
4su9/U1/ftsvNwFc29uWJDHGd/GGRpB+JGbkFGrkaWzZEEDemzoQw9dPDqgJnuNxg2cWJWjcxyhv
QuLo9ywwEO3w/vQkbjTso8SrQtOryIrOs7OcrDejxQKVZFPhoGvDeRuoon1GmKQlDpmQ5hu44uCl
C311Yyzeji1WQXXu/Wo92IMf1K5Bk3dCwteyPO9MlZHheYi+AT/0qK1DgD/FSj0RTKgdKpQDdanA
pXPn/nM8pjcfD2MaBjpLAXnAR9/FDeqn7ORf4MqT2MCU9QxHwm3pg8/euAWalI5yvweHEGxMvTvL
ngWkSWzTo4UwNm0y0bLfswYXyjnUZY4i5nEcTvyPLq4S2/ujAo59SHGsowHX9xTvQZmIbV5BWFM7
CjTndgOHB1OqFH3haz/ayYtjPrnJ1ey8SN0uJffAwhJrdq3AoP9PnWsLZIZy+OHckyicFuugkW5q
j1EgdtWrFK65hc7nPAFH1JfqR1M0ghXA/e4ty1XzZSifioGSQltP+lmgo9jzZPSRWizC8XiL9/No
kF0KBATGqAtsJ2QMk9GtXw9nQFxxdnH2SDKcUUdBxBs6YnMzbjPSGRYWgN3ZCR36bPSaCbkijAgD
bIETtLT2d0y2kUI+bZ0InJqS19S9D5wwV+Juf2wXas6/af+QPYzHbSSw2q6NMqjVfNflSS1Q4YoH
QCXhrxUV/oadXymGYT6qigqaMvPW1kjy4asdUke8SzhnXp0R3dQ/gUc7qRHME4lbDsatMcroLObw
lxwbqHymTkg/kwpzlHcqzc6Av5tCTtxyFi6rsZNX+8m2yD4a83MWVXXfMWZzdWork9164hVmLw48
pgsicMDPGkypO4mvyKckTikzx01RElLK68+yFfkN2F+WVbltENCWgOB7Buu1ZNHrY59o5e5GA4MR
pZmI5cS7kALJEylvzs+x9LokbBoc9zEB/MuYQiFBwzWcJKWqgDTIeWITFP6X5wwCx6pzZxqAIBGE
mP1TEBX4PccgqBiY4QaeJmV/fkQLT3AGrBbdtpP15c2Ju3vsIPbYerNPEYkEds3U9/B3co6shKPe
dPSZ/+4tRaTpcCQtjsJUhJ5kwwxTCpc2PvYxirB3IzmqfvvNpYz1VtK7T0Vieb26AV/JFUcHWvSU
xVlf7g3WQxTLbIpvVO2d/wuUmR78gL5LgotO3U3PNpiUPjLKKSzCV2ha98P0Potd10iLS2hcGMLe
mfGR3hAomu95q7Vl7mXH5daPY2yeCF+iQ6KFo/gkXKm+901XqqCVdZxJQE4tita9IlVQ2fUUZ7sw
TWpZDDxiSHkfeH/r864ZoI559kgmwrCo06hkBjUoxxVSB0DUhZ7rQVfup8GLhI8doUAn8ylt1FDZ
TUTHDS31b32zBCbGF+YNTcYmYUzcijN6apcGMQwADhuyetrinZP6czaF4GD+CYRaSZzKQWIr6Kyx
fxNlrAkZCDlb+TPm3WCoMTFKd2LZOAC9w7zeX1VWO6fYa+ldcVZImwjRdBd7imFC8n/gjGPdDK3e
dLggLCC5JbG2ptrPaJS2+Ch+EdP2FvOEnhILF33WVJurE4L+P8B2JPFlN3huUYOoLteMjwFMoHsE
IWz7n8EUm9Phxwa9Gi8lPTSZxwRJOOgU8v1i2oExW30UtL2z7Zh5065yaHvmCcA7GuaDKL9etSnl
Qc25eqcmEjJxiNHRAKS8nH83nTAYEH6lm7fDDRkC1Gurc/bET/Ko6w/tf+w234Facc5xufRX/HWi
XYNWQLnzGWhShPrflFCzTrA1yIqQAJg1Av1kOzVmCU0jVsdPuc9G4Etp2BvBvtP5WCBvWAC5PjD/
i1Ta27kwNR4GPuJsiSKntW1uoNqkWJkcoWMtQEwyXTxeI3k6ZClpfP7ikQMddVWWtoyEh8ePV5rn
RBH2rvvFh4GRE5T1I/D9HT9cg4wlaVSKzVbIuA08xw/74eFZ+NSsuxzpw3axbc3LnL6LZNpIEC32
4SoOmQbc/pC64TKbGgSfDYFahXjJdn37dQEeAeSegNvhxvaXzx2AQTQaJ40GbPkayROsC56sBCjL
7M4zgLXnC4VXPmf8WWqcXWVEbm7vCHmyKbw0fe/9Mn8IwCTFNnn9iCxCnnMp7XHFU00adPcvpMM3
mJVr2BgOzeaPyfCExicY38eRUfmxdlHTGuo8K6QecOCKFi69lwB6EUI/U6RhnvU+3ZONmwVtTsNh
Sb7BGu96owy9ZK2jxq71TUIcpNrEfkW4sfHjyHaZDGeVdmeUnDFYa7g+rmzvrQE+OZSlQDfYokRu
3KZWIzRi9ap/4kbsKG/R3b+/8qFQ4d/91r2AOkwFxGzuER912axWus4VwOzcKmAPilR6294Me4rF
CZO5M6BP/0RzvK7ljeB73mbZfDkNqplbznSpY+J19S/tSevph8HhhGx6ERvFoh2Vspt0tGO/gwqK
Z66vNvskL04UNNsiW0uvWAFuVnsX23RqbNt+IsYNRssw6sd0RHvE8JIMOhSfSAd5VOgGUWJdm2+j
daWvkGdPknJPKJP8mKG5Kd4NNBUqvMMmCY/4f2giP60yj7oxcryJMHTR7AxEE+Sn3a4leA0K/v2+
l2mqboRW303A+KeieHeejNy3qSM5mwxNZQvZ04iQ6hBE2eaKDyMy8Y6ceTWaEM7JxNkh7yNYkegV
fFqoySDHRURRoSA3HMgFrSHhCgeIBWk+T8gehoT2Pwrqzzr4nydZnUA83nbPYTTfUpz+du4YygpK
gClnvJ2ZxvfZ1OcYUnZ1PBpTxAtK1fAKBNpz1vBjql3T7STf9m8zzIyoUFlnzrQgo0pP6IrHfYct
xw27A06T+ms0GW3uW8kSZ04mVdYRmRFjRh+FejnN06njO0hWwQKHyYrreq4/0Bbg2bm1rJ+UmEJ9
OsmGWyPSeyL4LMwfJvPvxz2XSYf0NhA4bDEPL/WzOEef3qPjOeo/UHDYb/SknGOnshzZziM9SZeu
89/VpmwOV8U8OpVA0x4Ma+ciw6LH0T4low/M+frAgJK5RZ3dJ73OXQDQwWiXjOqhY3JcBrJ6exhM
0888u1b+YOb8JHa4l2Z+lQoQjsBEIBFXJhkFK0MNZf36ejsArD9ZZDCDiQpxDOLMLR+jNr5nuMCl
/cj7O2pDQ9yLJM+hL/YLqIr2DBQXx9qb5u5IMZj9e+kH+KBvdO0Y7xx7l0z7UL98G6Ndc6jmJyWU
utwsm5ABOx3aF6qmMzuFtGHk8Cijn0Zl+5Edg2+dbNty+WgZq3twjr16CfkL2/3aZRRGJ6ffRD44
SmarriDDWGqCW0NfzOtVJE/ej10GT43kYLW0gAp+0cW2SgyX/yxVZUFDttd6CYIRj7UainQKHF4j
mk9Lqt0X4YGYzF3xAgIGw+a7LFdGQT4YYYmWVNmKN6Bim/K7C8PnXhiFU9fgm+FhUWgqHJYRBcpO
GTUs3FubdFoIArtlKXCh3LgLtg9t/E05196vh/z6+tN64IKwMtgnQAaz5ZKsFEi97GdWLaKWjOMQ
L6tlZrWShiTFJ8y1dU/1T4zMt18eiUzK7a+t7/1ba4PICk6cwQuA0bGY4CNmAX2mUTMlZyScacNt
ZnuXpDMChpolyVeD8t0hPZ1bfqW+qjBhHz8UjHOxxsiEw8ZdK8oglwPlCohXehvnZus3jlg1qhjF
VtPYk/xNmFGXjrK8EjtzhnOLu6B/0/y8DKbN0dOgxY8O0CgRyGzgLXv3Z5K91iaSLhi0vD0L4pkF
/KaD6CWFqAPYsRy58ji93Yz2fM+xRYhe8Pnv2siIr9FL5wifc8bjkPZu10gOjTkkUooGsu+ZLI6t
dMP+3uYCT8ssMRf/DBK8J+OK/RakwC1r16b4JfKu13m0O6T6EAlGR6ofBua/GVZ9RWHhgbjbpZjs
f0UmQ3dmDfXCBQ6GnSpar30VKdNvgxoeThiFxfl0PQQwhLBum2vE6Sp5fPOPTmPBZMcQEB8IvtwL
nmltJi/xBH1QThONlLVe2nAP3bAv6fKlLm5h1DU+Sp6S/2Qo7VK5DLD/kRlfz1FH1UlU0De/sZth
q8ZTzr9XHm9ArH3/j82o0O8anOHq7gnWP/Y1hO9C2JobhToRVhCdtXPkKwqcLoBfDA1yBAM7Dkj2
KUM0NubajdRkm2oRF5jrO/8pD3elXmesDArMj9h1Gt7jq9szG+vlaiGKn7LQ8/d3XgbZxgXkqi69
tRDJESJojb2etth1/q7BOuQuaQR8geoAor2DeGYejEOR+ukISd0BMlBfP0StVNEb3HpiIaIVvJ2T
+7fMStpSfyGohrthtknC4QQlSlxOnquh63kz5VILcJFKkbrSmP+TgzY5UjYr+Moc7zCqmE8jdu4l
RM4JHuXfE0tjE/UAd9SpQcAC4LGO/MZ5w67fGKeUuDLw60df8fULMThwE6ZVwrUiHZcRqyp6Vm6i
HkCZJ0F+Zxuy/th+sgh/Hld1J/ESQgfSX2qStRqt7GZP92WfXbfgZiH7GjofpvWOj7WpBHwaMJmI
HECn/VMdHyn3SBZi4YUYbTo3sQvH5uAdVHyBgEeBqN/TLiZseSWACcZcTNL3iibggJlGEduHSnd+
xnJ+xeKRcLVezpnIZSCVmxq8uqhCNAlnCNcu5tIIXj03nKk2ddnYnFsEakoF+bwuXsEezVtoCaoQ
VtyRsBYpyRkLpZh2CkrHVFe2cpDJlgowKpxXr55YCKW4pbjhRTqordRLbrbvEHBR3GOeVEhz/YOo
30pfYR6Tq5j/TCA1elQ0L4/J/lO2sf3/wX6+d91nDgVxYui2NToKvn2L1EzVv1UUWvx5XrhDcCfo
KP0F1tIueAiKbqHaifAoxJBCe1MZ4oNNtC1FTnN4bRmO6gR6QdDYTuq8BRGzZwvrzho9RZE0hGZP
nKZENvWe+duxwvHVBD+79+fml2tITs9k/zPwLWN6ZC4V4p4M5QZB/rYB/4LdLp9Y6XEDdzPrXZkq
BTB5NH5X43JcWobOSzdtFH+VG5kSXwu+lQHsc99lSnpA0T6DRfdo8wWlXy/PpGadPTn1SoOUkbIW
j4vqzRoDLGvgSoIdxOtr0uCUON0Rectg7e9R0zZ3PyduUjtN2bTqeqEzd5qESOz44j+UvcSpkP1j
oghARB4oaqd6ALqu8oasGL74/43lF8L2iFP+c0VCP2s347n0s4keUzWleJuYfv9FKzkDxSoYxdf7
jD+q9Anz88EsRhGfZ0VucFX/o/mgxdyX5RIEFRSxrgZ4cflqkoGLd5siXYwovi0bTMXrDKx29b+7
gHT0ZanIBL7CwRffJTaqTAjHrWssid+MWjYe1+T92LF1N56DQOJbQMKkwAEP1614Nc8Q9gOrwdV3
gMKyeZWKXCXLzmLQ90TEUS2u6vYherBgqUSmuN9ZIsL0IZtUAadAjc4rmeGo9G/2lDMtQch9PZey
Ihr32d6ueIFQxQgEjhlJWqveFYGi7FGnQkwwwjmfc4i+DkUOl2Ugb3LHvafDZ1lPvwk/2OFnDKEI
nc5qfclzEZzefEbGKV/KA1V+wMHMr7xCbcHcBABm/ZYEVK3UiV+buar/Xa+Dz32lV7TS2sEHGlux
I3cXJgfQHmR3V1nMtdXR6891+PcEAWW9WY4ynK+Ma0wI2HJ7OcO10rPZE7+oz5jJfIE2ZYASzzEE
HOrXFbEDp/Hw7/x7Jrr9p6X5ryFT7757K4ZhAgp0oaNk4ddFB54l+lGT2D1rSbNxpND5rtskRjV5
JFR+9JRNh8iuEYS0aeilqrREyDk6DhruphFvEhTO1xt9IdG+6BUKZRpgnFH5hTOD91qvthNtcFPZ
06W+hlVw+RjlUfqn8fcOJb8s4d1LCWuxwNUyQ+7mqE9EZ16E8SL/EGiUozz/nnOT+YQ+6wbmnMZl
zFWwhWSvppYtpaquY81oq5CvIcnC9MKYQ1p2Laoy+cDjxOi/TC31UWEdqRNVFRrt1tet3Rmj9hf1
/YE/5b/p8dByFME/cBBw7/X4S+0uYrbpLj4kQxl2IJT4XUgpMj4ppFrC4JSbbQu8NQmx5mgIky3D
6dkTx4sThYw4EBkZp6tNWN4sNjQxmdYsK7oNtGX6hzTU3y+N/h7wVJt1XrGauNpvmA54PnO5IA+s
KNMoNyQJk+Az2t7qoV3iDDmNBTgKkya8wAJmWszfvU2ceWMEVzlpTqDNdLjQSbrlT+6VDJgPlbAZ
YFn8YvLJxUOuE7jwGMAlMSBHWNEImhLslrpqu/gDdeEAOPsfdaqDFjMBzwjDFjAYLoyMYcGegKIa
LGxIDIRTHDCYIAXh9WN5iBWylUNsmPLdAzZydKlDlNxO6rxpmjg8zzlOjbGdPtk+I472HCJwVri/
PElRoGY1X8c1Q6IMX94Nm98sJBCq1WW3TN3grHNShSLVNfEP8AkZ8rvuzFfZl6EcUz7dQP0RB4qw
U67GWDXWJZJmS/CM46e445Mov3CJXy5D+/4EK+J9H4vChOWbY2TZFfBzBu6Cbenfce5Tq6eudFNk
qsPePE9mGmBn2ujCf+81ImCzjllwsE0WoMz9waDIgrjwiVj5T4UhoPbYo4OV5n9jS+9QQ+6R7wlz
q0K7Xg9tIK78vd9IrU4+qT/DyX7QmSQsupMywTY+Mu2QZ2gV0wxVBQ9Da4u8tOREXglRuzChkSuF
J0EoL37aw/ABVQFxCMtQq9QT+fBbAuUpeOq40gcK4rSFE1kwEmrSZ2zdd/Ca4jZS3VBlMIbfGYUS
6pGRagmhI/bd4AwN7w6h3FS3NC+WHTZiQ2crK0dqEmmV/xDBOrrJuuiHkHCNTGhTwEfjTTwrQebj
c+Or7yb6S9N3R3QVxKot0QYtvq4o++Q1YCsB2mr0X7pbqAEYEnjoqEBJZGlu4cxl3vD60zKat/l/
Dpai0/+2/OI1hDjCL53TtL7HSvtDHfUlYnjNwRikUb8v8p/hVNM8Rhw/rSUTRFZvc3msH72XnoXM
3JtKODXzIIHCgSKEZP4ILSo9/ffbbgNG93h2bfx2OhyuBN003HgF9MiV36pUOZiBA3prPLZ0/rYH
EOid6OriOwpybR4lLUQVgfF6NaldAwvmElj7p/wLEaDfvaASv0mrq74d1/ze7QKO+qC/cFdPPkje
BF7p5jOq9nJfLKHfyHmL7ecbUJCh6O+tdt+MDYSB27vCJ+lXd92wY9ACI0fSvg+o0120Skm1vsVJ
h/E4gu7poHpy/o7MHE65kfvl3jDtiuxMsKa/nX/Tjk0H8bszkBuhOcwjIp/9ETvc2SR7RerQk1En
7hLZJhShb591tl1JTghwt1geBCFZMGRW5vLXz6pqLXfLJOmmAL7rJgNrb/Mne6CPhft+AE0459+s
8h/sznJ71CaKBZZL0sue/Mqoh7AzMLHY90vlxuxAap6KdZebwwCFXeS1N0ETGZT7npQKvHZfAH2r
wYyK638A+UNYCYgHeCkQ4XnQVu85GIHqv5H5YQ+Ajl8+IKHQEYuKaFRLf1Dp9pl1Wy0RznvOSO8W
WdHRyDkL+OVJ+GHdkoDGlxro4LH5rYqMjDx+V0UsluCXXJGrz446Ldna9WE2wNyGzQ8Q0XLP/Ake
lQ7XunSJwf39uxD7bSx5gkhqTJKmFsnVTLoR5CXumjC3mQsE/Wofjkvq1kYdwBhbnUgMaTeW/Bsk
tXN7cBh9C45P2wnUhktxLFHYqT8l5IZe70VfEP4/Gsvj4aHb4QENpNq3+i9CQ9g7FhqjE1kYczgT
9oeJOTQPeZ+/0Y+2PWIS5CR6sYZQEifEQ7iiVVAElP8eqPL69mRkNkzrPrIWUlV7ROGDQFehBHkF
TZZST2JT+bi5VK1ZiYQCp7FYcPSiuUB/VgKFm4hj7nz5c94J+Ruq4x6CqSAwPZQVoPqLUjjyHOhd
u757BhYiikmRdOUJB234NS3jcqH3TkOTprZ8eCnQfeoRCIS4aoePTBkyAgh2LflDSuwSTQiyOsNL
2mxIlBAVxVkTprjmV0hs17vCdXREFRZDSyDAEJBKvggZtw4XsnJ8wHQ6NGKia5mM7/wOMqqGXgu0
lzuD3hS19/gOS+m3N6k5iHETquTi1Ve2REcBA2vkhNOmfFL4Qv2gRDUT/N4V+O/he5Kemq+Ck3Xo
jRJQpyFiISNeDdjMqbrrL1wKwgsmyFqQWxpYDe9RNgQNBMMI0NDykWgzvhxKbJqnDI0Xn9v+UZV5
X7DBOURki0xyRkNccDXOk5tLj/xoHLkKr2faUnMAg4Y31jtqZkilr2iJWf6GItWSl9CXGoc86yfV
Gxdt3D1EEC7yOD7r8HT7btv0+pagf4a+cqGEJdLEN3iArr1/ZJ3Dqt21h+2/am1sj8fNN0DRAf8J
Bxr9oggCZ70IMY1e5bimRCgcaKKP1v5jRavkeDQINCtVcXCA8+tYT1Gi4qSQ7oEDN+wgIx2xBM8+
UWZ9XUxA8hPK0pbRMuE15HcG/V6SddxzgEBbEjO69KczcJ87jUlraopUS6e8kLbq4Z0IGAizAOA7
D9Lt2/3GdUdrBwPNxtUGzMqoXCKhjdHD2jNHfLBPwfX9T+1lLdeO/nLfkWZbmvHYdKPZsr+V4fYi
8jcgDuyiB9Mrr5+ukAmkFmsadQho0dvG9H4T7XuMR7+Ooxn/+45JM22U/akua/Hn/dLDMh/hGt2f
g4rA8t7BwB24C/RsOchr5gmWofu0ZXrsqrruxlmItqLYaw13D9Gn2ntmcdjpPamknKgSyPtVFcK1
XVB4U0tKG4pxzJpST2XoqXTep4eJ5tP1rx2bme7yGuJ+aOvWbjONuEyVJxDq98fR8X+0lzr3IMd8
+/PvjxAILlS+wlDW8SF8hCHZ412DIIHp4CXTfyUEFfVayJ4ka4+TxECkR2hYT9m1Koudb5ctDVhf
9KmSerwHQYcsTK1aE832pVm7J814y0nG6QCbxXxCjIlet0omZ06Oes2HbQBSh9EWghmX3uSl7U3T
HuVj+NkcnmVCTb4hnBbvbB1jeW9a4Fp6CkennglxyhAZI14XAJqd3dv6/1aqfQv5g4X/FkhgTzYc
j4nn/1xKU0ziqYOS1s3yp5khXe3bgZDbbw3ZTxHbKNGsHo5rFXqRjcE4JF0JyE/56pv34uQI7XXt
eGt5tvoTTiLFpkXej/YpgwqCVN/m2zgppP8BeuRiWcI/zPWFbVP46T3/kT4+7X/l6NwxIVHsvwBd
w6qb1rinP3L+kq2/U6nmfytIYry8eKBL3KXM2ulUItjqnCzQkhDmqNTsiMYWlJRITDZ80NmOHLYS
eMCYyLO4odZQswnR7RqDVqLdq5awgANZFU9UNnwxB6BfWrGpslSEYbkSbzWv4s/8CDSinU9NOdiD
B0GBqFnDjwuPhNL4SEN0RL6hKWxsfdA6Mbav4udKXBz2GppTtk1BfwADKOyUQtt+taxX5Hrumjmb
5vCXhEHA6Elhd0RL5TN9UBqym/McizTs3BQX/o6qhcbV6SrCBGG4EQqsfYJfmFnnYvZ9iZJaIp+D
18fO6aXIjwyUDkDHmpbAKk7QrDq7Qx2abmyV3L+QR+k4LM3DObA/VPWeIQ3pkkxhQd+JwXubWBI4
DkA4Kpi749tTI3CXBY+ShQil64NKEdiOtb2jYwgCX+irMSMYmPsk/56del+LbfwEdweA6BGvhzOl
WkpbCLgQ+Q6ZBc2fzbhI7qHwxsVVayYudpqCygzdoe080moTVElv7Pytg/oRPexqZIs8huBu/hOr
+MEaaLLtNLXrN+CbKAeyXAguZ9kioNFJ7bxx4UxlkmjA58cxT48I3i0N8hC4qcrdI+QrQQj/yuUd
mwmZzbzRnCOfvYi52KjVBLlCKNIDKRDq67Awh+qY29mIV+M9cF+Rf8wsJYZ4tQUhXfGLXtT7M8YD
5RePViuG4Ub1ugcSGs0Ra6GEBtWY64C7FB62zFsHU1rpbqIwEv4Uh9mzSVovfiTpUr+5uejqG3sc
gigRfx9gxHa/U2/sJIHOu1UaOgT+cbKfZhGjjoo9BZPW7fxIklWoJcKSZJuuH6zBxMAUFE0/v8ZQ
eSZpbZIP5A7nI2D5M6k3Rg3XNfzUisMzoFuIaQ8wjYA/ZBRpJqzoqxLrdkuTDJ1Umgn/arwbcoSJ
xlhNAHtWlYs3R3R6SBOYhCz1OzX6kCSNlnWkP3YgFnjayuiXWn5EKcdLbpWtdrzsB38aUQ8yTsnJ
BeuvvMiB7HMHqq95OjJu8oVa+vvTgOOVbU3qweK4TjmQfMn0hbsx157BUwRWmaKsjXaOys9hHIIR
TKWtOTWUWRbzzs7wywtG93WLlatmVrpZ643Q5l400+p8741ORyL8TpjPDI0AfowzBDamfOGVtoR1
e2XLyfmOLOMT085MqfM61iE5bcK4gUJqy7jgl/d2+/l3Cepqi/icdwJ62NQ1dxY4FGC2A7+dySeD
N7o5PN0CU30R/RV52Vt+PYMuTDwBb6M8G6Nr7imeSia3L26aPiBAhlHLKX0y44V8oNKCOdJ3JKOZ
6rWPlnZ5bSrhg/EfljcjVHWbT3/3LvZ16o0GIh/8EK0xT6ctbDeT0WMUGltLfa+Z39gYm1wMQqsf
zoRF17nJlUFV8v7R/Io8LIyPHTEbN9Xkmp5Bs4oznA5WdegOE1NnuXTl5VVl2K20+CPHhm8VTW+a
zGSWbbewhVS4vEwuEjzJvpy6IFgv/OCl8QwSskWnrLXh+7rsHcdr74eOqk+SQ8qiKCXgMWeiWIUL
sgc5fTimU2OklVFWdvCOONGp3adperRH3n1s9Ibt4yL29oudYrIcAsCIM3tuNXtmHRjqedDpG3Er
KqsRdyUj4CVJrpyutxa6ASzJ+bbthvUKxpLujIJg13wrq02+KdYIah1b/kwkc2Xb37ua3kbFkTvd
59GN3Yi6YMbFhgsIVnrsGx6Yvu/jX8MiCn/8LQNp1afEGafp0nQzrwfBkAGggCVcBtYQfSvUJkP9
o+arIUcVyYXbBfUuLfzuRyeHUC+jMcfHhaMRl2lfNhNz2ieScK0tyzlGryVXT+cMI5ZJeGu4uuV0
ZvZcTnqc8Q3bqYtui5DsnJoenmgfHRCn1E092IKejuHaLcuFRRrp84g7MRG0unNpsh1D5g3I9s4z
D/L9wvknyQv7yOvPFlO0LOIeDSuYGufNG+hZDPy5LAWHxGe2zjWcFdNwt3nKumugIBhkxTE2g209
i/Hbf5XmufPsXaRigMkbRThesb06FNpLpxo4w+hf29tzICEAI4PmyGOXo/ClvNI4QIOYJ4J5b55D
yniN8hbLjQxz8iri26mR09Wn+rlFxi77adOuEcHpXVqn94hKtxX/VKtKU0ThIEKHpHmKDbisGgQY
VMvVL4TBheYmsh0uvdArd37mx87zfiLeYYKr++OWVLWAbIjBzfn9X2nz+wj4gP2AM0HebtBatYag
P6mmwrRaj4HRhJVZnzpkx+iP9slHi7G3gxlM4l9Bx77O7Uqcs8g0BCtazxUZ2MCkLbDqEZTvPJ+T
WHZHuefZW6ofjuprcMVm39iruQJqbAuUVNFtCfZjSTmv/hLfYvqJvPEtZjDOAOrmTLy0Pm6BO233
AZPtt3SvFG0PfElUaZbfHuiJ3RtUshqwmBeJByBhVFQrIf7DzsXE76K4z0qn5eXj33dLlDkicldW
0PSImJYmZ/c9jOv7EzMqpk8uc2Ocw7ew/fN7VlKheSv/NPvpIwCCP7tP1K1nVxTsnahRkcgyz7W3
GKKfaK3DbNbhrLTsuryC9ox8UQbcrecUdz815E1lhuZ5gX3BJoEPM6vcTICH5CtMvQ7dKr8TE33a
mVgzIie3zkjBdso+THKrGaA8f/nsRjZTBEyVXJ5VDCqgt6gDwV1bZRUCCIRdSmuw9gpebbtyu/81
sP/bJnpi+tQwbYn5B7ZL+km597gcYx8vc6YHoQj7EVSIy0xDzK73WO3udOvfFsHXtzXYmXf0iwEa
0jBc8NAI9Lc6ueRHp5r4ZJh2q4MOzch8Tqzo4j0TNqYkf2PREjdir10KE3Lau+3YIluWMYk94OOz
p3vC/77Hrxf+ehB5z5BPqjiGtYFfzxC6iJhvJlsdi7EGfUwGRschmyW+9cEo1x+pKB1OaZDGTbLQ
bCWrT+TbiF4PVpqWz6PrOMGT1K6kDlf6sJPR6Sl2HBK+qk8wZiRgS3OKgr6L9IERxi+Rnj2xeYeg
XsRsLo4hRL3ZIL855lDiAA9baRDFEj05QAASs0vIzY8/V2GYGNc0zEI8yE4PTnHYTVZkyIISZ0p2
qJmOnRjfriC3XeHTMnMR1Qh7fzOzFRFuOut6+QXhIPRVVenscuXrSRnzlcCnsGyij4RE/lVB80kb
i6q/aZvQg1C5tkdZIklBVk84P194GM0cupXcll/3VZToeTZ4O/KppyHSXYfhLNzLaaxNgdrs64cV
eyMLrPHL8/dLCxhcF9NQHvYdR6DWu2YwzpcWK/F0jV7Fx5DjT2VTLIqYnX5ZBcNSB+lEwNZmuljN
5eAcs+vfG5L3aRjGTD2RW4AjCUxFQ414G7HU5D0XibK5WDUNngUoYkLc2LukdgoJeiuu7X8akMKU
F9Gth/La19G1xnNryAyc5k0y/bFeDdZnGasA5YYPgEiXQEQTyAiME7/7G+T4LxOXDTVbAUEvqeSq
jStWtIjEhFZ+sFj+C6QI5VrOlwFGFStvhx1EIujiYmCEyr6NsZzlPTETiVqG3+Cem/SW2xn+gF5r
Av8YPm0M1n1MS7fZ3KFEE+ou1ijl7L9uCP2dLXQdlXbu73xvOUQOaalJHhReObpSQ3y8imyB+Nwn
QoZQ3YmobUf9Yziv3thSEsJwokJWhYVbr42leAbw4EA5O3XZmWG9p+nP9B9gtL1AGZ53T4ItKUo7
eDvJ89ehA+/rw5t/mV1p2t6clJMwkSHPUxXhGdW3jKY3yLUeu+RZVcVSJRSH+NCT3uGI0gh9dsAR
296WaPErUMv4iOFHJWuYsR+lqjb1S7f9I2ZrHprP8GHf3KV/2V+NmcHIaYsotfJ2mrti1I1NA7lU
wz+uSjtHXPo245i4YrFopFP0SM+AV/TYPHb9prm/YLBcmbZ7jPSI41/nfNxLopLviTQOADMSPG26
ZWvzbK8k9gjesTOqBooWpc+dRvvQ+3xFUwTAYgzcw7KkVC/HOOAuwL3EWV19XzJ1/qxNvTPYpQ3x
dg93Z/VxIq/bQn9LKycgnODKYF2abUKgzlE7lh75wglFgIAXrbjswBcSGVtN9qNbB6P+Z5aT3wCt
Af1hOtP29RaGBXgoBPlUy2Fybub2y4GbPlSwIblzWWiaPy+O3ciTpp/BsNDaw3HopUpohdk29kAQ
Ix8rtq4TnFZgLCHIT470qmFC2x6k5Y0YzUs2ctEFSHD4j4BMuV3Bx1mjzEKBByoRQdw/IY0tO31A
eVGSyvGmROl1OuZhGLZ5IGKj4myGT3wZ48NtYN57nnYZnHSSS0S9iLRqrp2HXFSip1Wx3NbxF/4/
zRBuEgLtEQPIa00fB26iSEsnFxye32Cph3/janpBPrx7Bg6/pmUo8NNNQxyWP0O67qgP0WC3Ytlb
IRsT77o9aXtzUFr9mNlrHFyc7x5RBvw3+tZ099r484Wywleh75B0+SzF4Te6k7KpXnIXRGNXMxoE
BRSTie1//qR5rnywjT/PDDu2yF1mOUS7E2xrRqggddqbEcxFlzbLwB4RpMCUotWVy5joNnx8YI0w
kMyq+Kfl88h0fuvLdXk0KLSxZw2CqEiFtoL2TInU30+ON6k4CSQYP7jQxLSfjC5esYeS3FfwlBZM
zoWV9580V2yzVYq4939yJRMj0QRRxbSKiv9VS8pBfrCWFkZy9AiTIm1BDLBxj8xgaiy0i65fuGDb
w50jRCICkfMJnOUWtQ/MzYuDgVT2legLEl00njaItfBiiPn3Qq1ba19KVNWEg3iRUO3tJ33MolLt
kDRMiUXKOeUk3e4IalEnPBUX3yhN1zhfvzq7A0555aJyHrO2potlwriIcwiqm/U4dvUeFks2Fr9q
jSjQ6k8r+yue7I72at3l0m2Hwo5G3HUNy4Ean1fU0JxiCoQiBofQ2biT31Iz0LlBvnLvFoJjxHJu
P1Lk7mZGDF4ez7404prwKHCWgBNFcpD7cxU6qdfpmCgT7LFFtNVOsY3JOkEAJ9+brIOfxtGeyi9W
D7yeTmhD8WZRvtFU/oMPOW17Sdd2H506mV/imctFCPF73ISpbL741zwYyplqfz38PHK50EeGaE90
ZMGCxfTf95hZOrbZt47gKA6JlmlL4rMD9dFW9bTLs8BXbYVDpN3GQe+2bu2Sw6Jv541GBD5VIUzf
yQoH2A4wroPdWbHk6NTvgBUR4dLpMFTFP3u/I9XGmBygLlBf40jOPuJxdUnS6D9MNSs6BXrmILyM
as9lu0UKYiTnapFA67KjobT6ajKJJrEcXFDaFhAFpfLSS2ZYumW4GeY1X1G7eHry2bJKI8+hEDwZ
sgObVni/ClhWbxT303FFyJdiiDu6AmZxfabffohDmwiM5pu5AGFXBRlmV83Em+/rM+fOSuduTkW5
2my6/h6qaA0b7dc6mhIApWh3fvoR+vjH23mpCkrF2Yao8w8GTGfnzJrx6BiGLvX2BMxn8miSDZyQ
ejJTcupgNhx+KRz9KwbWY0QTgI3GE0Kjy8IK/zl3LZFZndvL+fAnr1bYHxxj1lkDp1y5vmQ+x7ti
lapHT9tQnro1ljjEdfCLclV0s8T4mAZyHYwVpQHMJEsJls41QbTlNN6W+w+bYhrdsjW+Rk16KMzX
O6Xbc5yorF03Gpb55//v5AcWLdI8LuaYbJOL7q0fSNYHmgONfSN7UlaEaHW9mtnGMWNwMlCzlzm1
toRwiCt2Fb6M+UIynaZ+TfBCQGpbKmM26LaXPLMP3P6qR8/wPL4ntcFOFXorEj5EbZ3Xi6Pq/Y+h
LWHCUMikwPo7efqQZRJCZOPkfzqP+EAflx07nrbU4eiopd5j0T3mFhsujzJoqxJGrjhKgV8Pbcoj
7g4KBwjwhjW+bdjYxtICxwvb7TFxtlf62aOaWXhAOc8+I3mnJJfqdUNqnrKUCqmJsnMqDrCTH1pk
+CHlq8eOE5xK3JCSS+s2Va3bwzeJ/TALUBIoPltYJn3BVwqNrqvfksEb664RbSt3FneIi9p/b/W9
F4ujbnTBgf6sjllTVnriAKY1K1J4PSotNxOxYSMY6P27wu1A8hVJiuozVNoLRTMQU9Sxdo1M/bfS
vFhndaVCq/f8qo3FGShG7uzKKZEnL81VErNE/vRZG6DNPLxaW/E9oK5gIYtvIsIqHTL6p3jc8Rmj
Vja5CFiXwmvB18Fm9gId4jlpAoQhblH9LltCPqJnQnF1fWe5HJTCTA7dCQMnEcSUiY881XaNOwsq
vhsjg/zdqgnRedG7r1s+d1RAm/vmy8TO6IO40K7g8eE31Jq6m90MX6njVkdgYFSpiyS8zTaut7iv
eSYF2H50rHZg38S5m8TZ1ukqhsAwF/Rvsur8ZAw+nkbwd6x++wbr80GJxEyMkxSuJUcA4cjwZnuY
SKivV8y9KeCQ8o6X/aP0ptqWOZonglzWzkgrzW3CqOHV/1ifMcwtWT4hqTzfvJiTeWdpStokgwxe
3DL0RD7DJqERU4uJjY/It74vHOV0PEqViHoLQv/iJ8qjmQm1zEUSpo4StIdDCY1Pqz81CIy9rMgu
k2VEAuYBAJAQF7nLibqhvhiIoJuFUkr/xCW/oznPl0zDDHXIhT4fREiZgG2TsAVBMqeDYUbZo0ad
J1Ks08vwo/XfA6yThNSa0zX1izhqvaOk52lXl0S2J1rbnlDDbQC+V88Cko/tRudOlZiZw1uBX719
wSFP/OE7LLeqGTe6FlVZucOarQA7+eWxbrbj+dReAaDqApjMrD3nh4NmtKuBSh0E4wpvXNXR34kR
JqKrmvSIwz3WtVyXD0lgkdSa1Ykmyud3mIFKXtSaNPcm/JYM0cBYu5z3r6zBk0SBYfOT7HMlRWmF
oaz3+hfP+SzjojLNCa+JK1dcfnDY9MRpQfs7Aph6FFgwP7ZhplffU5JhqMXCDR865PO9U1xBb2gK
pQoVjkCw+A0FzqDvg5KYyULDor/guzRNtZ9OhTmxd0bGxwQkmvzjgs6IW0ZOi2rKxwoCuhXFxLab
bD8rv4VFpbqq40YZ7CyM54ELreGCIUeYgowfEsO9ee0H6vLBlZNsWIrXz+v9VNQ7fqd+qGAQUmsp
X0iIdWIKzoySzhTD/NvesVM1RCYDfL1DVA6rAfv39NK6uaUgoINEP0kiQ7szClMZo7nObhFEV60w
O+Qzcs3lcJvj0/JveRBiLitcrz3eiZvjW3eCmEhCTFaFICGYLEUNfTXXX7Uzr6HY93SLS3uiJJKf
DDT8zLwAiRcRrsCWSSUzk91J60uFVW31L7beoLY/GGomTSZJr0yyFIPPEsE7rbmcJRKojo5j7jkd
VZJEAsJf3qOjaynEHIhS3b3akIuoC72wUYs0feqz22WrzCgIO0i+FaI/cYsIUA9SCthX/JNCoVok
+ESt48ignUsNy4fLJucvX6Nzn0ubhani8stBwHOUzoyMe7IirAnF9uvS7rUe3uPHhE7PpRfZkJcm
mBB4ZYIP4G4gkXo6KOpyVviaD22ZpqxyodKDYBryO8OQnLm3EX8kDuC37LmQl0laFE5ta6P5Yl4U
/3WSMEkMcPNxQUnuU1cP8/TutvA57MT/ZQajYIzBqnXpK4RmzQGEgmqnlztoBVZ8RWG3iZblvGTx
rQNT640q5l56rf/prNXHsbyS7+KRREx/h0l1PxfaluhCxaR1C+HYZ+cFkj3mrPm2rCZXUtnX5AdF
qavV1is8PIFAICFPd5LrN3nXPA063Sq74SC/TpqIAH02cX1m353qIyW5eICynXfDrQlUWO91Ke8Y
/m5MfU+SyoI=
`protect end_protected
