`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14416)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf2yj
VPQAmUsAt58mMHMw+w/DT9P3PV2AmIveltBKo5IWsW3CZWsoC0MmLtNx+2L9oMKaH0rrU7MZ4yWE
fdSyGktHrwaAfUSYKDL2iGbtefan95fZsH1ajOfR3rlizQ/AvCS6HNnByGi7gYowmGOJE9U5Ams9
p5juJefe7B+9soAe0ROQLDh/v6ueRjuhh80V400rXc0aqVhF4QVcf6PRvv3rYiHhOJW3wHf41Phu
NUcYC5Yyt7C5N75cInfMsegQaEWKw/hl7bY/DHVnVAAVeYh/hIlohaoNQzDR4YW/Jk8CfLEuunsZ
rSVTf9N223MlGFHGgL2lGV/c/0lco0va1Hui95Nsg3M5BN5D8QNpwgPHMYt/Cv6gysG5XhJRRIUi
HS5z8kInGFyNgr6F7JZUIFeeVVgux0VbXm7nn0elVAKSrEPaL28c0C/RddUp6Rj1CWeCZ9o69F/n
jJQDagAfoy5IVpVLZz4nzSzUufU3U4yCxc/oaHTE2zD0IlLMWj5BFosF3D39GH459SBGAMpgvSIN
FoD57tL48kSu/G3EvFvQPpmkovSyVM+L2nP58i6e1FztTcHCPRvwrDz5Iei6rRnkCAdalScgd2FK
3l2UMyxDnl1T1tXqUcV7I1VdgAm3V2oFcj5owXlyTF40DJvFQSzgljIT5tKMUVCMv6chVcZnMRae
YFI3k+2j0o+h7elQqGl+9Kgx+pYKGm1nHdut7EOfLa9dkwInjKvXJurwgkfkbOoKQeV2xw0Hk4tk
VXjVpXMhq7TZOODK8R9xyNPbGEBo9HtDWACvni+HC3YzagYZ5Roxd3zj58i5q0EejWoAvig1IVsj
xFQORVxQjGdXr3r3dOkuBRvzAXQgTC17v6hB1glCh/TmaPuy4iVwsyUn05C+9MEn2nzTkwYPb/R9
623wz37efWNLj7r7lIEjWDpfP9KrTw4LjCtrkUyLQZdu2UY54Esp7b3YWBRGPs/DOV2tmtcwn7Z9
S78mNA0CicpzEjHU7zwx1uOy8wNA3uCPoeShBIV4dEnGnOE0pBXZF9Q1XhUC+Ef4ujoht3kv//Ow
FVHJejtIRhkjrsxyH1UdGpMEqy2onu13IvV84QCPJkZCBzG0wZPrgf+U73dDvnOmbYp6A0WsEBwV
yX5HfSxuBpDNezloR/IiGCnBp+b2hY6jaMNy8QV9RTFHD+bqcjFd0NE52XL/iy5mzpxu+RzkSJCI
Q9d3uzDmUgRi/FbqvWA5At0JBF0f62nlRvqu8nLp6yv4JoxTJeYhXcFtIv4Lo4hjSibkADsmeiV7
AjfgMX9QdQ6tkuw0+fLbG9Ur+ck+SGQTfzozeiK2z8bLXPhYoR9tNd3RnkWweldsbbaFibFVlrZJ
WIqNQ7fatNdQ5JAJ3H95KRLcQPaA+6P8X0IGdN92yaGtERM8Q2Mfd3xpyKFdpzN/x5ZysVH3O2iP
mKaQ9lL2R6yl2X7w8DN5Wxtgpv8UU0vL7zqWYccWideAKJS3uyLjkYUhGs1pYyt52Tkx4e2CUzOU
vQus2bU8AdTS5d2vQjYqd1ZIoK4AwVNdWhZoNL9TFuAw0X0dbR7/HMoPx4XSliPHMrDXeTPuDmxG
R/rFhMff+n/haqDbjINO9hbtv5LCFhlJ4XhMtpgCH081pWdTb1MbFloJqnpV9YK5L0cWQqtu5wV0
TW2cycaJRKT3YOF5dxi3RJeV42NfWCMtA8QuvdhLJQRaj4oiOgM0xROciGMvpoernd6GTBCKc2el
bkmeCHk0Ne9iM/9P2YWBaNCWNJ19T7MCYuwVwrwMoOKYdxGbWMu+SIv7AMZRfwsri3bpDozukxtK
sF7s7C89IQ5xHw46Fq9rTC+fKfconJdFs+s263Peu8gHpC42U+ym9+HwE7OJAfhTBdc38963b4X6
/BDnkNixTbhRoS29Ks1AEsewAtzLd1zCreizBODbJJ9xf2MEmk/IRNGi9v3Ku/gbbpn1lx6aOQPj
X+wl9QRWeFtExBUqV7ZqTFzjXU29TW8t0K76N9NyVDF2jVTAkuHuDfwC8ayMVzkmLBkB8wh5r8E6
EZgeOxjrCos0sr8G/Zvpkt0xj4VjhsTczmT+nwo0j401QgGHLunwql7tBoHu9A4WG3S362qi73SG
ltB43BrF7VpDRxkTxhVBa6qqGqosfjRu26xaB0iw87WJsz8tJumkI3b9XTH/k9VOsfXvKYcj3Rn3
SmnzrQERvQiqcht6T9EFm3CrcWOmwp9ZddEHBqRc5KoyESCEZ3YLJgrYWL4a7Q5qJrc8PHXWDsos
i88Y6BB1uNYcfZeqrFg8ztdSMpxvf7FAwiYvAhKB6CP4kXX9QnSFPd9eDS1GQ2LwSS2FZzYhKNIJ
bzq7bPBaDQ7VSAclgIRHW9LC2aM9Oa6XourHQspPZjj/2y1QG/Vw4DCnUzRhaEFOkCzIcJ4eYuJ0
2CMEE2lXJds4qge6NrLnzxjgGBxqHqjMNEFDqlkmfHJosbhjmsWKVTZ8A8ZtjTafFiXF9FdwyBzO
eH/cL23spZIJx1Kt9FSUa+XGeVmy6fbkMWDFG0WbJAdOE86OLfDo/pNeZ0MO0HEA5XyCIjsDJKIk
uzLuP5ALET3Fi+nWDVGagNOvz15+6uRnBJ2MAItDc2eloYp0H31wwhpMWSZgnKX03Yeyo+0ARR3Y
16Dl3VBgHoWx0+7ac/X6r+S6Vsrn2HppS0LUROLoV0eny8JGGdMrxhH1lDlYdhFCIH6z4FkXwmGb
4d8ylc4oUWCTHLnC6W+X66SrhgQ4yXFIifk9WJKRNh7UtCKQVtuqo9WsAS8dS+VH/Y/MPn0CYMow
NAIUjqvGXw6RxChCCtG0rtia6+9g+vFVF1+VYSyq6YJBmgZbVVs8v+wi/oN1v6QYCSyDc2fBvfkV
z9wRUXEGpYGMQ9QYWuk1Ij9IIBT8213nauu534fgTpmszdpQm2H7c4tEdlzyoEICstF9AdUjFIP2
33IGZxtZ0X9vWRz6E4wu9tU4ANOURhSiH1ubCexH33yhRv3aUjtKUFzztyRBcjoo4BtUdU1N+ws0
yGuMpzSNf4r9klSUTvqc7VlfrzD+IAVZX9qA+R8y8/9Mg3/WhEDXw0CBMJpqhEwr8isun4aBSWnl
vblb9+qQXoVnQsnXkcsexgB60+Hn6XW2GFw1y/7SU8JED/4yIt/NEFL/tOC3XyIPwTdzyFnFUfGI
SIDXgTqvfzN0OFNPFCuffjzN6QfJtRQV/hSOK70DL1cevyGU6YEcByaUllUOLzsOqe95OTsnLtZk
bQCca+rKE5xDUK72ocQkcwSZ+gmNSRWxjZ170T0+NCc3npnhKOFTWd2rWfDbo1wwmUevl3K/+9Co
3yi5WWZ5XkqSAz2A7UwmS2vVFBtcVhvsvJododuBEGj8sQ8OW20yIgaXD9TdvwHgjDxifghlhotG
gtSJ672xfv20Zi4LtjobIbT4kiqcWAZQXEqsnkVjqNUQNjRXUmqBNeIz3vphsYMEzJ61HuJDbpgL
yz0qAJoqxjjL2r0SeyFpelXMU3KCnUcgzpUbdlWjJhvQ/DRkycEtmwmosXd7bbFb1UFyjoUWkQRU
L6X9kHOsm5I+3MYhi0xzrZcngF8FPEbFVaofggUynsAEfOlB5p8F9gIaDlSSzvJq56H7vJJqIofV
U3wlfcG175ajs9/mNkfWWqDKro1AyrMRhLOa6FHQDe9gNoHQUFObjthGpKSeLdM7pslIW0OLAqzC
CJChpbIJIbf2v0M+77TbNySSDSqjjJGqpRY0P5uvPjYi0PM6RIx6Li66NBY3Fcs0HDRAVDI587Cs
2CCtP5y3NwD76Jf2LrH2aaCPpexKzVtnSIpJ1KN/RA/KTz/gmiIa6YS3L0PtGO6APn/FKr5s8yEo
3VzBQ9pYXGVaTa6zJHX9Cdh1FhWUaQwzvlF4cNsPRNcFHSWyK3T2MDRDr1HaoQ/VQbQdN+B2U3fl
mu3BAIwEWjt1l3g/YalJPhZ1V6cLqWnGIwI4rXycHaxASaH/p6VaE1atgE27s6LCut43ZCdbtKlL
CXi8C104Ce12APoeiwPdQorCOBVBjHf86OWgLAl9dBPgDPR1C3ZTgqrjpKkRI5nQaUQhCz/q3a+U
Hcv5N7V2e2/pb33RgT49EIu+rE+2WnWwulTSZa51dy5xrT3o6Mya1puCLrYNQPrsmL91gEoWfQRB
LOEz/ZlHUl8d4PbbjsHB8rVOkzvddyYhgAFDQUmvmLsELRK4oB5/iFR3X3TBxpivYaEXWIXUhHUR
7wvuetBBXyeB7iXh4bRJgSUW6dGEXC+lYwN44gqgVP6j+bNvYjpdVGsjM5877lAMmtt1v3wlcAw1
f88nyh7uHFWsjoTDeLsAmyetBBlgLWadVY+4silF+pavC2Stiw60CR7kYH4U5xovl9+NDpJsaGhN
upJK6krwVVdV9byvcVLERcokzzxAVDCTRckmMv5DYpDjjg5ns70dWMn4v3y6Tm642jmgIFgeHwRX
YqTHdrIK7V/1Vlo88IybabLcO2ILt/cgrJShOr5yhaC374+xMQmznlKZtID1eGjvCNgVdkJUOyAg
CAxx0yE3ed6BQrWwiPY9iCAFOA6vGlmAm6GFZnGlXZjoc4/5TqsiUexgzi9SByQ+9Eg74/em+0Rv
vWQm2uUUbzOBapEFJI91wlnGT1oI3A/cn8sWsnOUqqSECG/zNvJVlLHCXEX+Fe9AtnYhkuhhLDVq
Cybuh1KtNzPdqvY4Y6MS1x7Tit6faKTufSJwUQg2dlnRwiSmQk1Zsaj/4IfSrLjyV8tkJ4vEcghq
VwRl9AQBGNBpYkLhI8gTWZTqefbScDqRHHYWEe4y6vZ6NIELAdhRk6GWiHGK+djz9QHHkwcX9kYj
Y6qzX52xdHaU2CwL3+HHEVVrN6zssLyqWmvmgLGBpS1SJ05NmD/PTxyISUpFdEGl6obU6wJzgdaq
wLk3E4g3ToOdiL0PGu4szUvg3v0TKPrfvG1+jcNJQCz/iUvWuaMnLcyj1vgK40chHqwnFM7aIIWE
oN1VCRoYKr3oGt2a7+Z4cDqF9Rn53Nwqbh9k7MEf/QEmYbr7vZYt13cqm9cJQpZiuB7ttZEWX65P
f/MgypN+x3ocwGouNc46CLNY67S939f6NZYyaAcnMt5c6EPHWGEpE2qvB/GGwFFqOSObbI5mQl4F
va9BhPKe/XvtKV8dDMo8MDLWMsYnLRh3fI2os1coiS+/LaWx5Jrj0+STtLvUfWwOhhn/W6JUmu/l
ZVdKJMWSN2u8j9kEbLiAzs+CXG+8j7kld+kpENrt66fz4cXDiLwsfmE1Z32QbeN6QB9JYOUNAQex
IKW0oFIDEqS/nuHiq7PZlZ9VOh8dr4EBXsn1S5vSUk8aHivIsFb2dt9R8HGOVhUllwxREphOtPQ8
o2qnKKHyk1vFb6P+LzZTpaMStT6nK0lSNJ//VkRmqc166Z6qUee+V1NIH9rTJ/+59LrC7ercPIr6
xJm/XPxcX/ReH/7cVvALK8MYL3ahjg3uWxdHQKmOwGc3FqecheB8uBVVL4GxfBGWIs7R3dsB67Q1
nuEzmQ6UMov01sDCqDpwFTLmwkCWy2F44IsPcdrPmD0/Xz+LSGEhvNbw8setJDmR5r+BfuvRfvjE
9dGQc1Ujbhn7pmRD5u8Y7MTvAG1fSYd9NDkWsPNmpkf4Ud1R2z1adfgFliwSZQXu5mvYxwqw0imZ
z4GRQqRxzCh5qBzMoCtNgcSmy9zmMM9BnChvH3bVMtCDnOH2kpwJuft3FScp4vf2ob1v1Qba7lam
kyHMQHjwPJkURycQW/+wiWz63L1ADOiW799XzpCUGjxAJxNaxZHt69fU0CVWCAT2EmiIo7cI6B/u
q02kp5LkHVX6msW9yS5mr8pU7JOtKbZFKCjxojKprLIpau0sbZN1AihbJ/QX0CJloPe79oECQFpH
c82bzH8a/xkRieyy5JyaCflfW33rz+99T5AwRkTo2KUSuoFFAtDKRqYvALXqxznruyLZQDNw8INH
xoSn6t+vltHL/F0Wm2UcaQWMxgrxLeRASKaNowA+kFVyPPzo6RlxaIOn5tr+C0Ad6mP5bwU9fioJ
Xp+BQJ69dibpkoe69kpPxDvHT4K2pk8BmdxBvL75sxQdUU5TLSuqsg0FRaeryGWdFgV69Ean6sYR
z11TIKtxj8sSSzXmWLxfwouF7XdRHlXg8b/4+1XH/dxQbzy12IpPdV4kgl7W+Y/lKlxFM+jJtEpP
DphmnNmZhEqhQiPWLnQes/r4gEv9UEJJ6aOAd77OAbj54OcdBQyZy3VCtR0jvb5qxJN06WTDvsTG
E6KmlLVnqZ7OOnlCnA99fLpQSr40hx8kDbdnZciOhNk3+mDfWdhadNj6Q7guwS6aU3O7e1L9d56v
yxpzqnwgf5eB1ccivRW1aS5EHVc++qfWFWQC4DpCWXNubirY+FBuoVaSQhWu5EXb4Tk5VjhAqL6W
KgM6GUVduvhi4qmsYKFx4ZKZ35KWxfDIBcvIBOcBehz+3FhBPPqR9t+1kpFOWesohR4vWle2QQmy
bV487sTtd7ltz2mXS8orv7M/rLqdpy9jTYALLiCC8JSjahGTdrh5+IJyMOT8L+Sl18BcmPGZJ9G/
PTVRGjUx4HfvcZiQTGWqZqHNLo938nGHChCNEjsB71LKq6nEsyj1nO5JiyeHgXZy8XVBKxl50tZD
QuxVlVMPY+YPQNIKUe4qqUqaFupSG82++6yNNw/bsXW+wiXVxGu35/O8vhQ5PZD/Yzhu/1kqzgH/
N5b1mz3cthmZqQKCUmLBIXKiCGFVEGXQxy7t3wKV7JXAQ+flwGhWGcAeVsrPMuFqC/b+y+wsFKdh
S9D45sZR/HpZOCTwLjYz2V9nn8X2JsNISo8oF9oTow0uWtqJ64whhFa/qpu9K/Ke8AWoecZCksRK
VMk2V0kCbBmaIAIMXQ5jkhxPthJUnHbN04ouHdA+Hr4mUftFCa5WgdiVNXlPwlX2I8/VFISQRxPw
CF1P25Ioc3VMArZCp1GUpDeuEfCBb3fIW5za7GxQd0miR4dXzHL8k67hhlurxgbj7HtY2yvnuX9f
JKRv2/Ue/4mGDVX/o93cN0p4FR24l/VNzIWZeoe7s2rdZI4UB16Wc0TaVkqOZ/w1psItuup0y2ck
iP3DoOOXxvrbq8zGnigg+WbX21juliZMXrru2GqY2MS7BLILZcYs/699JBvmDgaKsmrjs7EWAOWg
KDunr+rt/1huyY4f+lKEJW1miPuUFZUELfj8cRfd16oaKBG9GlqY0+utLaRNzWCudFRTJgOYIRAK
YwwtzIn3XgmqOWkZrdSHkrCUgX3Z0odD8l+FlG64CxRSsooayL6btmJTFQ+PQtqDjnDu6hCSNP5k
kwULmLI64pwxyiShYhxp3u80b4bEVlrU611vU7+lEbNp95Er3eguTylE36wtyhLSBcEBYQqRk9Lr
He5PxHIlukFLJS2BpuuqneZt/THKLm/Ss31BfOEoXs2uNH/haqWfQ0T31F98dYlhNfGXM4/KmF6+
xMo+QNgn8ylUHu60NE5CKi5j7wlgyBPC4hdcA5WkVge+TbtgwNq/A/lc2y0zPVFEkDdiNAWqjvPs
ZgNKnvYp4K1pw2BDGlt6IC+lgWayGBjAK6HaS4elHcLPHba/s1Tu6FvupW0A7wt+CJw4rPbbjwm0
1dYeceWAXbWE8wI+lRcyVUYLfogPO1p48XOHS96REczq5tDG/kP3viwh9rHBcXkQLwrEVBCTtWLl
ttNd2sW+EpQ3PFnIaH2XYJVrxECP3DDsrmX0fuSDqq482p+oae09S5DXyhyNZdGyFoeRZ4xooxXo
1Cfmb+g5G61IXgXGJ9J1CLCdzGxYEahD/Uu05ybrJNtEaD/+dzdiA+z4Mzdjdqhtj09rhusiZfzR
VTw0ur2q2Z5962C3ZBUMhBAyUC6FYVLTXFh1kTt8UCOndWAuTT4fPBLTPE2c9t08j1/I5CEmzteV
1TsF43yAPub2zdmxEDGh8U5i8ZgNiK1h1AYqTijBm0YkU04pSWxe08VmgaBMfm7R6oh7e47hRk9L
PpCX3kyWKmSD7iWKRS/r2fJZpWWRgtBwiQRAZ5FEU2w/BJtkbqVK4WoAwk6xJc6EQB3H+9MonlZ6
4pisUbgvLLCH7Nlik2tKt8qiMu+4op4ZBCoU8204sfRef8cX1XquHv4XN96Gx4db2GwzecJmWlCT
FMLv3UH2EZ7qHvCBZSljLqFms+ScY+19Uw8Nz34aKjY2C6tm/tWAeWtFY2kSv4C3EOFWQfO6pf6O
PJ6KS6jiPYTo5Tda7ZvTWoXMljEv8p/skbJP8LX3ROmzuUTrXnvbjPCpoQLCtLs4fAcE6+yFKt/B
2CFfEL3ESj9za7eNw2yGAn28sLiFXLCqHq+MhkZ5MvODrZtsiyGyvDYfUEbe8X9pl9ge3u26cPgG
ITi2esor5Z8cSspWDwL1L147cZDPQ6kO7GQEXiVU8vB8PjVz/gh+l3DLOQDXUyf9NRi3LICw6Qyx
arHes9ncqMI5G70p1bL0FP1BqAEb4AhDn3r84pTD4ik2A5hKyX89CnbWSjycn5y5mnjAFYHUdleb
Fks5wzaRpPCstZytRtc1C05vii0/UxhCQ8Szch/Jh0t6qwJJjrUA2IJBAySa31B5vPk9cJ0trATx
6/c8AJmGZ/xTxIm+a0CQ9s87Sjq/7hMmmCrcYAdunYkG5rHKT8C5n/Hv7pxJkPQni2CBTBtvGhjG
fDxrdWuWW8wByU4rIXGD8/cQ7s+Np3S4e1J7/24iagIrdDjjqu+ryYWdq8n6d4CkYSlRyfuqgp5W
PWUg2KI7yVAMryIZ5Zx9apDgCzQsSWRR3XN9OqKvef71/D/bFg8BEOBbbEGoI1bGeK6056pE/qEd
G+mTSEkJQMvcB4Sy49L/S342hMfepJNUG5y0MoEL3QcZE+QYPGCmeS+/uePIg53/3y6OHJpB7ET5
McdWVKJRTBfI/rptQ0ZK925fwS4NmHBt5zX0DcsCmFZ0iUerqjsyow7BL+RjqU0eAEbruCgFGV6H
56u+hLQ5ob34koWADOeapQqO6y1wJYOIP22MtTJq7w3iWyWC3Z2RG/IXi3ZCTBiHQH/Bs6IzVuVS
LK7IYSSWMEntDnfcRPQxsDm/jyk9c/j7IT3+x4oUCRDoE9PqZLGKnmxNg73VgPoMRodV02VsS5c0
iOxtgjPVl05M75jkLae/NVxKS3wvEwU7LEWc6kPeyxXmNXZa7BkXJJ7XrpgaNjPlicuF8lprF/R7
tjX28d4kPX1QnKTp2y95GZWHC2QFuEgXs0EZQGgQCrYSVka5bvujJcIPSw07uIzSpfNQT6a42tE3
ms7DrpVclfGKQtxcYKdbJsh98DxLWAegaQNdhlIRED754/0WU9XIZ2XxZ2CWPFtZa5ykjVzGueGx
cj+6pUjn+lA+JVV877NkKp7aALZBazomqIatmnkwQTx+oPY45+29oIQhQ4QUNtHiFUmQjDIrMx37
obXP8VbijnagjB32y8t1BfFmqzQZvojQSiS2JH6Ug5aBMaxBQUSOfuLAxeodzzAXS7eOBDtVnLEE
0rzIvflycl3y/ac7JTRNu8VjGtE7OqWUyIL3Nw/JxRd4MqfFICVpREANTY6VeS7688bE6LWQWL51
G5xvcfM/XopbGkILrBqqicz7OvtCySkA2G4BLp0+7DOgMpoOVSt1Vl7qbjNql6Tyrr5BQV5fnXA2
evt3gUzwqMQjYLVMeV+XjRD6izqazDWXau+2HgyT+Ae4bYdKTZeXKRCzFG9CuWmG6MDcJn0KoHgI
h7Hu33kKeVspmlqfuET6bVCF1EDOTE8mtTN2FFGIkkPX110JjbGZBcJcS0FLwk6kkbRKKIYHUa9O
F6il0QnFyw7TYt99C9dGYuyjXuMp83VjDhazWBpTjUrVGXtDQBJpWrPkTDr6nItkhDR4uJgErgDA
YoxTIGXh0AyBQ9C5W5NgORTWXHjIjCziWoy8XknXIF/zUiHAG2ZFkYPFXEuoFGBdX8w0a5M1VAwe
tW5ejy5CQH2xDZz4ezESEwsiOmMy2gVAGmwiRNAYwtXHIJmYIygbij1qbhWZiYjQ3uLW7YgNUJDe
DsgwOKPQ7SPPLHglOVBRyFJ+obyskNaPBp8RNwdfEO6VEIoIh9IsD3PJCjH2ZyYfFoZjjSsDMyrW
E6atdLheGUmipuzTLR+oBj88XnM1Jm/8dItlJhqIV0qwZ8dqcMeC9lAHxbhr43Bz40rF773+75zW
4xisHrIc2+FB8XX0B+6Texq4n8f3fgXZDy4UbqF/1hnIEf4c+F+/z6h+Uqi9K0fegRA58csrHBtI
C0sO9fPCiB9Kwg7ZEGVwRwUlkFaqwO4bXZYIl8nVGb1bLnqNMD1YKZ/i5DQkyswaF7BrOMqjIkko
QrD+goGlACe3KdKyUcxG7YP5XZzt16C45lwcqVc2JyrH9D+k2Uf6slBONyySTqm7lBCyhK7+qAX1
jIGIOhU4PQW2Btss8bLRd4S4HNYqtq1b1qh3EnyP/YAiYiEQ8Uy5EwiF+ESV6BaZ0wyFe4hTv5+m
L9WJKMIPyg80jLwPU8AJXIPqDbeurUjgLMDZnlSZbHIkzNAMP55h0yx9v70ckLHJsyTkXkkMt1fm
ZHl2GyL1T4cmH+StShi8e1geqE2cmQrnNqgMy4WcY+C5jpYvJ1BVkuMO2Z8BYWp3aQFJIkf4cY39
yWl3aPll04coafV2os8IUiqYoiFUL29bbtGEdqiQ9N8DKc4C44Zso5uMozqMDeMFYXGhqFaw07Nh
7WhehNSUSWrSiMt99th9k/OjWfvoyxyTDljahJawDmBEfDM5R6ivEda9VU6SlfMLv0c32lF7MIu2
MGgqSnSUz6Fx+Cq2qxi1lQP1H/hhr9tRJMpT1xku1irU+ARSyI07VdOJP9kx5CKYWWRRcmZOeIwQ
SOrwy5kHADcgHGb3huuoQPOXH1iswTtItoE6H9xIUpPseXWoKrebkm0In3Tg0t98JeVEXn8Zivq5
bAkLaz59WuK7YcjvKreTKv5Fb76w1UJXV911P600PAkv7JKfSgu+JEV66uYRXqtfO5g6M4LgA+jN
+CARP++Gik0qfxfDvSGplb8YGZhwzSvSDzijsp9qunjSHboC6mOTblJ60RGLu0CijmXzrS7F0P/c
qNsirkCFt4UghT53P2Ff/QfzZeOMn1+ZfIo4VpyvigR33lJPDuhD6esBaJrBTNeSpBOKTRIVxX6+
olq++q0U5/0O9dXYczFmxZSSrTjF34nzR3mTxDSnEm9mzitWEPp8gepr/nmVGwsszk6dahNTLGgA
oteKtTweSUvs6Im/xSaly/DMb5iY0HUhyhcY+IImgVh2V+0WT95KtjVNf8gIWFx6PawlUVbIGbMe
8TrfmO5PTDvXAs5mvfq1t0earf05FXqeOCGa57j3sINtAbf7UfHXH6F9XE50L0FYVqn5jNMhBQes
bEcM/ccW8MhpCGZx3VKwvxoKb8SXMzgWhnBJLJAZxhzmZeCZYcF7o3skorUe7OW3R7LyVY2Ru5N+
PnSpo7AmCY3+BC1obuPzv9iRysusZxzt6PXUmp2uHN8DSQFKrjuQzT61v5mQDJ1q6GYRUxha9w9O
QGcQYnF7zN/UEmoLXk+2CAKScJ0Z164wOyn4c9JwqnVJY5GyI+WchQR2Mp+lLEfnK70DE85Ty9tq
H+6B7neEcgjqxqpt7pAQZivPDdcQkgXBBIZBTZogqdDBStnnkXH0pcJnWjtW6X4RRV6+yC6qTMl7
/obJ/J6VOQIpZxJgqW3iWkzL592Z2YBjxdCSuYvS2kMEkKpBPpK2M/7quw6sa4U6qHdDEL9rPSUO
xG0BjuZrgcdAvPWr+9NedtCQRBGBbtafzlL04pA9IjXV6ZnF0KvQw5Woor8t1YirzMVkx4laUPw7
+3HjuiUK6OlDKahh2q+LEmQ5gKoXiitfZB+sP7NnvQH2SDXLeqQ1F84rjseTGMGfmSPF8lLXXfD0
2CpIR+mTe+bIDDwAKdqoro4xFYzAmZNzC6G5r6O9lCe69GEVq8HxkxH5O5i4jAYquLNYeTBkdGgN
2T8bj/v7aQPDaM/8qHz4XMDF7y0czQAe/kfAfgFucdE+kZ16vFXIu/it8W9nD7Gi1lVaJbRp1OlI
6czjUSJLTph7CjCFDdfoXjFIU1mCbIi4q85ur8g5lux4HScYBM+eD3EODCJm//DuefTZuvulDvwW
6A3CrUMhpVm/A8n4eZN8TIqwYLCcSLHYA9Y1okYUBGCLBL+a16bVVv0L/qrm+xZjFOJE7Bpd1ml4
fpoe3pORmYAZSimBNuBxMVZfpSMHpI3KWJTahqgqo9cabAY1YQKljoCBQ9oevpM1rWASKCmyi32x
n2e8/zFuTwMb6+uWOWShvtf4vwvIy00zEtGATDrQO5x80kDBvYjFEZPnIpOiUdJfaqhWZVoazcr0
mXEyYoeuAzseJHRmqlYgJ6xn4jfqu55PTF5/BlD2RxDYmy5x2HE1rOg0QsAxs1sOTjoBgJY9KpAq
IxZ7OArdY4PcmXDD5QA1vw2vooSnHjyQtXnuYt3Fz50KX9JRB07e3Fxe0WWfELL8oE3QYy04BxPM
23BFoKBUn1J9tHr0FcsHUedtSGuI1r58Ec5lt5kbFPad3YL4IjlFRuBHsBdhNrWDclI+vN9DEp/f
hftYOi5hOFqj13EBCM4IzpslsCcckApcJiuVrpAw+fB6MQgcW9QwwjK+6mY6GQZVNLfAT5oCh4M3
hDgHPQpUrYSmzutLO8Yg38ivLIUx8ukPWnODqDvGRFAsK+VlaBQ2vffPIpdCLteO97bH0dAFxM/M
E6er7fTT+feddxCOCKset5u8qH5/tnwYX0KfpVoY6D7McWY5lBMsuhlB1Vw7LGwJLKuiJJQcAO74
IFz0JyHqfjw98grAVbsH+aD2+mDkTbi9GjSTyePpcbU+XD65zYoxMtAWH2mwBj+tv3UXsxVBJ52j
6RUpriBUi8n5VIH2vxEsfYILet3AwP0v8zeXx6JkhXQ2vlF8nbvupkp3/BGHsFyUSNebrfFNDPWp
uuNm7V1o+6Z85DhoaBRdfcTB2p+zpslhgThbO55E326hAQtIcusWxB4U+DRR1CKSKxulDt2bVIkA
yZdx3xxZqULklc09uLmjAeE3w9XsOe1UZdALnYMiRPaW9lsZ2t7eXNTGtcefwaBf5mVMhzUw9gmH
FgbVMHYYoKP6Vil8XoXm5W6H1uGQYPpb9Ewd5rXbch6gZU/+GKB18JBabOx5gwbq2WAkqhqSJhiy
mtXWaflXy2z/igJM/PxN1LDQDCM0jOzepRrVkNhasVXprWuvk+UGV47zVRslzOGYp3KQtPKYUxFj
72U7FVsYzwii6Z7jTu9u5wpQn+itNWoH4u4fIERplNVU2roH0JaO4Ehk+nX5I07rPCfRqsdYX6nx
9PMI8HXPmId/Rm1bCKD9xNoi/yIyHiHtc6ol1+mIo1z3kv2Eq2KgzIAvIsrvRLBrwNwkDG3yul/+
J2B80CELPDCA3dILYIikiKayE0whFtHZY2IOLLqpETxPjQNWG4MVE6UuCIZyyDLYgINfj6iMkI3K
4F+/yAh7syOf6rv3UTQpY5/NEZfKaKIYj/Hqxzz758IgCgMrvZrKrBa1i/V7iL7TbC+NhXaFWcBH
ML5ZpNipMBaEvvyceCtPv7CZd98ojdGmHOFevJ0zUBN7iRnzPXNADRP/gkf+reLpAH4I7EEyYc15
B5Zg2fn5s+aeq9HkSvqRATxC4ACRxknLdp7KhKTKbQfH6dZQ0ruV42hszWNSPsNshCh4eSQOU4Rh
pSTFscEJRVwelI92iRfoGrYA0x9O2AyQV/1v2dX2ZF7hMXS8gBnNod6Kg/DlcdQqqJ/RrWN+LAIW
XIhcOs9wmXYyvG5ogVRDID9FbnR3n41aejlnCkKTlunwsT30hLyxBgNNPITomJwIjD3tImMUzgXC
s5705eo78C2xyICrsY/OGW7sPELeyi4wPqd1uw/ByNMqJNywyUWvX6uRr/O9/9oPD5lOLa2eAR57
GEwFum0Qnp3pd/nfdqON0MXLCk5gV00G0i2tCs+L4R2XSLdPuYNxMyr7CMVVbSTHKO36pUsY+oqK
YSGKeJSeX2eT1EQqToWM+C3UmB12yHQhGBgqw8EB2TzvriXc2To0Z4OT7KvjPzrfw/ntYxz+dTzX
Y9PcA6ogG7RaITxE0KW7I51hUG4h8nmPx7zEcmcdNY9+53RelaeU1Ku6fQ9Py8NcSOyD0MA4P1eW
lVkxiemDQ0iQrZvsZv4DEfKYMMA8mBcxitstKpqveubxThMc5Lfv9q2aD/6XpZGpdIYPvtbnTXYi
FVyje7efoiP3YnWIY2zBt2LAKrCpFoLoSDFgI/4KWS9ZmqzSxXax1lgb1YECcrhQsyqOGgruCvM4
hHz78S74SQGzP78zf4OtzO+UCXuLSgsmeJdIWxyjykoj9TwLfWsEhz4Pqpspzx9J7CTgdP09G3YX
sJuf3AN69giU9aBceP3Dm5nFlqsauR7+a1TgaAOB1g/1AhclqwG8kX3KskbU/Ffm3qWmYEHU0+sW
xElbw6MNCIRTuXwpSPPwbsSox8tYHHTokhV8vPSD/5/WP8a1SfMo1koaIXFYgwNPJGgw61szwfU3
Ksh/M7cZh3rZzdrQS+EdpW6XNrRdGK4+XOkUaOyeEOOJEk2AXjUn/8s54vjQCFM40lmPK3BZtQgd
ltYfKdcl9WeqjSas693PnKacY0qiOjXgUbt5hu09s6i43Yq2d3xlZvvXloVxZl9QdJruPgI+iWyg
C9scsuvXyD9iiA88NlHa+UGEi6+rVL5AOAotzvlo12xAiGrL2GcCMaCl4MRLwfWDAwGxOXnp39m3
l7Jkm+dtXmpRanqTPkLeiHX+wvv/O8kx59pQx3/qUuZlbjuy2flRRVFPo8dTuLGtny74Nh/CtLtH
Ojl1zvIbcn3eT20GQHPlM1MX1WAsVoaxIcevw0Gx/OebLbqyuReo2TIan3sS6+aiG1+Mv88/H44/
vE0NnPQVTHwg6hjRpkHGc5Sz6/eOmCkJCizmc77w/gRD7SPyJUcNAU9lieSTzTdBIRdUWmNooPQX
C00g5OW2yJb9DuaMuv9CrqQKaFaqY3r3TqNvHUe5zy8NE5mjH85YeGnca32w7RWzfahu8BVPmnqa
yz1VHJ5D0bEImfyM0/zZ4q7YC9xcuJ9d+r9R0JdBY85AnX+CYy7XdUZVPsemVgKsIaIsmgDCo0Zh
sdbC5L7XzJiUEG6dHtmT94aZPtuy0fdiLokOo4raWxR5VNOs2QUnIHX49Qx+A/++3215H5flORuO
dM0dekZSxAX5KLx7jgaaWymfm5GxOEZxCfEKroRBKxVv2s1Tqe+mIpBRAbiONhfeyHohv438HWh5
JiZDLJuVfH2mDXF6dTvwy+oJvEifjOWlQBmFAfgpRqqJhlQSrk+s4cZXGPPdGUansjcvUoaVQ1vG
IzHzTNZ2YbaR+oPkZhDCO+u3EEvM54q+vwQggau6DnOluCMUfojB8WxvX2BhqHTFdP1HN9k32u2h
bGci6Fb6zpo+k/t1RbEfPVzxt75FRFbovQUMuIV5mB3V7LvRkT5hYK/cLY6XQGhQcX6fMh/A6izb
miBjCgrJ5sOVlYC148bKdalTe/2ZbtOqwA6+rEIG6uZ10/SJVLt+qzxzY7onVGusqeorfKq58Ncu
6Lpv/yghImup9lNG38mLbiPWhr4Wugw8QEI5lCHvmA+XouhnmnHd7pFXWYmEPbeuow55p0kQegLl
yLcdiafCXwsayzOalS2WnDSkTntmEAgoeRiHCs6DMoRRh6ZnmONarH5E09oAa8zn55veRoCkkdtm
3xWEmC3ESB5YJBZAdPsHnY+870PHm7Zmzt0tUr8+x63gfNQABPyrIkjCuRzLJsez8JXTxSXo06ju
D1XbN+4yzt0M62wTEVcqpNmvihmnlOQD6m69Vf6sq5qI9Hf5M2QhS785qNezfhwHmP3+6I041EMP
QeM2QDWqR5V9PtGyfhoBe/OQtOeWAPBcRRHKoQ13iWgvIEp+q2TplnoePi6vT1vA+V8cnVx9BTzS
iEO5n/2bgMNBA5ylq/PZ4Wqb5rSYrC0D7KOeubSyRlaXepHFecYLK3Ca9rSJwcEJKS5pW6qY+HBS
h/FnSafwnkLUw6x9o9Vp8tjZgY9dz0AvVJxLiM8pIXZucLatbbLUh+ZwdQfPTMSAKoWc4hF1i9un
55KkuA3zUiYXpwYKlWQyVtgcRqOJNI1xfjQlXxesFyuLF4CFWDlFGl1mlLMlsCRqOQPw92SWKNZw
C/x8/VPWw4fZzV3COiW4uL4CRQHWhw+F5urW1teVzX1lVH5voGFOVpcn+Eh+bglOPaIAdbg6/BuS
TKBVld2BG8NfSkKYdJ9HGFgk/W33L4RiK+4ogfN5wTGtYYNtGYKXUdWYXDnXJTh86Y7OFZ1bXOYb
a6crdc5mHydYxr4GLBHb+kauh21J4FvXqSgL8p9z1RqQ9CrdtQB/5w9RKXRyIMB9zCRe/nqpIe6d
KHgP/o3WPxJ0vc8/kYcFqvleqKse2U2mDQyKhA0BNl2PYDGpFwEp8rhLX+/8CIkbebrM+BEyv5gg
P66D8LhVz79YY6/b6yYSH3z/aWMPhiw0HXOLWqsTy4oYK7L2SsdoreC/VyuSpTMt20rd53BC9OUx
1MQ2poFoxgzkjArmzj+paukAtmrMCIm7AFH9RSWOqGz0nQPlsVyCxdRaxfgWaBJ3XZLLrfBUIwCc
bKJSmFwhCFBGql9JcwjlnUCXo+kxLTpXky5zyKf7coTtyyuDy1Lka+qjR7LARdP2aKbK/ALI9D5C
JUIHGTShrW27NoHlt7JaN1uKOsFY6zRnzcbkMvZydqTxRM4XFgPe/6rwSFe/vEe1pUZBX8VB/thI
WZmd1wcWzFD9qZs8B/ldwtH7fNk74tgwsuMFTQfKieQjB4k90iNd4sKQ4av2BAgdFCHMF9u+kY45
jcyVZd+vzmyUSQUJI7CHmux+MLDgrogdiJkuQHeOv+kQ/tVvQ67t9o1epiaqQhTLtsGFu4u43Pmh
1dVOqQ4bEJdNZj9GpSHLB0ZwGRLiLI7dz/V7wiVRpy8wy2HDHOQIH8hdIc8ok7UGsXZLpxzIogJh
lhU65tesZUCXwuE0YNNZmCHzQvp8OewWG2g1CMMmf29MlFl7cVVdwDGgQjwRkQubdq59GeJHyywH
XUgKirmgbzWFiph7h/I8Taxizboj6L+EYb1SX16AxYV8ATmguQGqg/qKDlDXiOIt7QTm0l2OPuof
bKVRDBEmhe+rBMp+QNIkrkL4xI8JRIb6is+zLSoQXcatxxsX22JopDZv45ADzUtZ0SbAhCkN7MFR
6I9J0KagPoFs11CBfKHy9YPbHQivijZDpUCGxdDkykdicTLwWU0WhCFbyKJVKXM8MOfEexJDU6UD
73HgYJkhzMzpmcejJvy3IwODKwpYDFWxcgq5+p8qYJpmZNzamWf8LbWGBBu6lQTRZ/c8NZ4iLzR1
VVVFC8sXFpAxDcV/PbeTbUWRbGx+PYD9w8RUl7AmEkaKecHH5KXO8Ge6lSWIuME7YHhIKyX3ZqQx
yKAJCACJSsnou3f+TIHOqDL7C/scYUgH5dTH12ozLFIS2YVTQ4Hr/ITcty0KIJYV1d6HGM4uzN8T
shHEAWGjYph8Dlw4SAqiSyez2NIbBablmrI96vRteJzDGMiRi0hMuWku80NLJbAlCJeTznOGpcfu
jZwqG+VgPkZnUvh6oXbFBgUVDJD4gQXU4ohjWZQHNoGMzJTsYxgR+T+mdi88SEgX18kwe0Qx+b61
roW29v1Uj+3va4lSW+WJnk6EAiWJSInRUf0Ag1p5vH2UJI+53iNahym0Z4MQK9H7YqRmv/3PnVDz
Kw5ZuT9735D69RbucRLcxolhCu5GfhxVAyGooX5Q/uTUJuywPbOdS0viyJipgahjECEBQhzt/bea
+h+31WK+aufYE7xCahn0Tnt5+8D+0ck7Sek5s6arjDsHKKsEL87qax2lPYAoPgev6OetVONQt7mW
leWZGUU2RGyYNgW1iWQI4X4CBYwhiMXw4NqXXmfbiaA3IpjtcUsaK+X4xa4ptst2LR1vEaUiEedH
2B4D+MuLQUF4wS/X3ODU9metKjoT2cJ8wFE3siJI3G1/TaXOPawiLJwYujVZesNwxHRKKAx3N1Is
YK5QhqKEoq7Y8chi1e/6YsloDPE5TdvSFCc/0r4eT9yqfh6RO+fUe4jSrMbcnqZsWbO7bZP9l6ad
TUHmMaqefbtsxB2PLOvzX2qBYV/Q3MYvmzRHnhMZI0h3tBL65heA5aGRfghTS3nKhBj0+5K/emNy
M8uttGkwMs+A0R6lb5ixHqX6qc+jjr9bXZFCNFpwWjyAea5CM7XZMGzmlTV6DYwSDjCS/gq1n7W7
OCRh9uAcTZBOBNS/CUP8ka4Ga1eNOKedcinu3Vsi7x3pOVnUsb/Swky6DQZ6jCPTrlXzt80QTwzV
oQIJqrEJnctnAgovdmkJuPzHsrL1OHaN4vCoxvqXLHxKn2oTJCWetIfQbBJSUx8CACu3nJU1y0Dn
nzvmEJtRPOX3JxeSaqjWobY+Xj/sL5FzauCnmDl49Q1mtmtDALNVBQjJU7pIyWiywtZ8TpjDJjuM
LdelBqlcbd25XB/LWQQPGRW8ShblyBUpRtLhQ1T1u9E8StBrSxbaTDRDC71SX0Ai3j4gWsmKVHxG
nvYk+zdXPaf52TYzEImZovh7l3rP/A5oNdYNGCOeEkRrc4MiMflfwTqO+uUXeUE49qaZtxl3LczB
P70ivD1KfMrV3LgO13H1hsGm/AokPZxab8VfVGUFqeZiNKTHTsjpoqKrS8KqASCtL9EqWAyPIFbu
lD5Vu3gx43OSpccnArwEsfiDTSVU5TKGM3cqsN5QbEku3pBBSyI6KJbU6IVN2Z3x6OQhqN4LVk15
muDbhnWPSRSgqTDBOFnL5vEyRshX2BBUrH11XqxdbxC9Onp0wWigQ7ML6FCz5cDhdrHORg==
`protect end_protected
