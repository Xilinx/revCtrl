`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 77520)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAN458syUOoHsc7qgUGggC2RocRi7g+E2Cry/RuBcXz3y8POElHmRahky
R1cG6x1SUXAwYUcb44yux20sh71HOz4ygsstMiEPjuLGQRHm6KtuUZ7dRgT3Ru1ORrkJLjoIwWHx
v6DuXhdHtUqEqmrFp0i89F9xHrKLYAh9QpY4vA6EuH46qGnRkg0Xqbn7yXH7ukHYKGrNW/HYzlBo
KodBV8FaAsRPCF5nBNf6+BTE2za4s/8sY6FGK1LBQiKE0BEZAFIuVRl7y8cdCEV6mJ6js0BPI2SJ
fefSXGl8ZJgvz8jVCEKPl5y0Bq3uMf9+7Eeu82DlOFPMs4IxToYfAxkn0wP3jlCcHolLhtZMd30c
s3MPyQp41VymAlCujJQs82n4kXdi3Hobp+ANEdH/HLk2sgpXfMAE05y5mtNaBeQGxabEO39HiTb/
m0FEv+V9sbx64FYOjRg70U3e37L81Ii5ysv0VbjcNLu8bp+GIAS0suwQe7jgNvuix2A3o09eVbKV
Lc7TcmDDH/uf0r+H7AMJ9lcAdPg8MfjbRbzgCMoqB5gElwCR2a5XlKrfevYXLKO6cte9r90dlpZm
Z3EYy7M4oAARtZpzTMPX2qZ5EZVM1Qd1Jv7bcxiVv9oOu5JMGDCK9LqSTmGwzfRHdITmSb5Mj6Bd
Ov/N481nyfEAIXoPpX63hk75qV38ZHAqAynDtZBXgbRxqnMsNRfPj9ZiSzJwnjqu+5Qjp5x7xFj1
O4rs4PNPILrkUKL5NziZNp0IpNH/+lrdzDCUxOCTWtDnKGmFBwCI7x2OKbq1MXKer3s1WzQp38rK
GNjGviOS/VdvZfKIHOHW5QtjiWuvwdoPNA6rrRNW8WtLnLxe0FdcyU7R2WNzguKt2jfF58VQPvjM
/GBfGkdCpjJhvR39W7+Murjh1yJwUK7hoszGQgn60vHzKv1+MDVTrryDA2umLY5os3NuJBeCvRSE
ZvA9hPj2+O/QFLdMNZ9HAAPeFBq1bBT/1u1ScQMWSbLIGfHlfvq2WTtOKkUgPtoMxUO98Vva5IYf
RtOmPfWQadBR0ZEeHo6p2LietM1eYL4UtYudRaVlnsdk/JUucl8Xr0N3QQ7XhP1BVO+G1k/XI3Z8
uWgMH99nKJo6VEkSpuOGpNg+qS26QYc25HSed7jzrdWZCAu6aqX+RhPSQtYksz9q3zBx8R9foDWB
EapoTaDLAbZgKd5T7pVZHG7fTDftls8NPGG4ubwGITdCRgZYnhmPl+aQjnCV83OAaXrhh2O95lU0
u2quoCOks6ns1izz2M6o9OPgBUMoxt2ryg1Wf+/vLP5kyIJlf0VeVg8GtWO7cw2QjyuMurtkNUoK
3RDzL70yshIdpxgboy6GK+iI3DqEqhj2Bt3Cx8YGTUcAjBo3f3fVYzHXW4BtA3JQpmrOAVL9aw1G
W6HcpHhVXtecbhmDI+Ymc6Tsz41ehktp7fkJPUKV5iLpMwpDh8kJFDjuPgTsNnvmWaayxWVkVWE8
FyFpD+tagPf9LsxWxpEmRY+cpRqWkcj7zO/CKkQkbyv5KyAfYB37DOA4IZfozJ44H1akrxYBrX1Q
qUwCEcigf9t7h2Cgrw851KnoZN+q6+reHXV8K0l+S7gMgNHAHeg5jHymS8BIHe7NPAAMXNkOmAvg
9X5quhyxl5DbTgIR0Hhbi7b8AOpCoMD3GtTgFHl+K0LKwSnXS4TYb6dwbUZckyiRyHx2Qj0Cug1Y
7RDbo5iaeXgM07F4fFuCt+vBf1dQtANwB7W0IEqqNLH5q0nSEtRepaC0AfHMyQ7zeIYG9/qJQgR7
Y+61igbZiTC469G6KeBKwfBsXloxCoA2lpgfdZz18ERD5Wg/1Z7F4a7jv+g/WPG6z0YazkPimkF7
+eAlbQt9wSRp0P8v1CPVRkCqNt2ob5j8Pevj6PEclho3c+Fzmd9TgDqG7aNnJpwJG/TwR36jODzC
OH65O75DojYdKnrmIPwjUx2dCAk6sfFWTbQbEE7un/rOaQ+yoS/+z6kKwBQ7qBqMAjoye2fPCPlo
/gIHX5DoPW52KbFjQhxTi3JJKpAEyL8YURrELLAa8JC3kJiCVuyt+iZ4kttUBhf7lMktNOmwJvS5
Z+ZB6a2Rk1MMtE3DALm0Zjx9x+Vcy3jSyUwV8YPQlrjv5sFmaUix8vSOnaSK+M54N0T0e2WFkngI
5bhOlrMJeRYqNNDO2WMXnn1r7MjMcQOCcYmg6McJffVbMn+/jf1+kI96I/8u8RrSEeqUUsSu5HVW
amqjdXxCodtsTEdIAfeied0uJvlKraxR3hyV86pyhZ55o2ToTwW+oG7T364Lhq6bbOzyf9+kO9ob
PRQPhySnnpNm2AL6TctuaCrDv38sT9r3XZaWxVueOLsq/hPxDZt8/6cArN7dGCqqs/OeUHRSS2Q2
0kps63seEn2SipkoEQHKop7pSsXte6R1RgtmG5CZosgHjV6hHYlEFlDEIPVCL+7TOvCcEIkpTR6H
S+yRWoyy7eG34rTxE7dbVLviKUSDmwEotQUJ3IgG6Y/zhfVpnTjvgchWiVeMdM+oIk1LdZA/SCjI
vAqRLUR0TGiKBSrLTU3U+Re9tZfQp6JTmopdl+NqifxHbRklsn/sOHww58yvJhGEbeVfXJ00GCJP
qinjEecHpbdHpZGNjavcYtVReDYWNIy1Fm+2RRAKxxPsmLw6QtfCeKc0URA3AaxbfYgd76S9Wxv9
UlRbKYS5KHOtqrKaaWgJ7P08fAG1yw5v2vyZk3+MkSCNN3hce2X246u3oEAP+CvsZY8m6ivv/SDP
uISA9gvnneg+pEIIZgKdEscsVDsK3ju9oky+npDy4j3zZAigI3t1vU/YDlbayy86pPmlxI9e3SqQ
lXbVJ9y5I6uE7OPrJrZTsVXtwGQT7oEGt6ZnK3MFk9YhnRM48Wyj4DrC5ias6Qwsl92jgm9g7qC7
knV/eMfEeMpZ/PIYlxZJda/7Cb3eEx1iaBThq3TxSq3mOih2FagSoxXMIxJbodPVZuSXrvQhJgmJ
Dd3/PYoqcJkDKVguzoNBMKUUYdS6DS+Ht5iD2MFMVgyjKju+8ehzovRAfUDhmzmCvGmY0YctXtnI
DLBuzfr8SApwFrrlxr2pDnKYucquxvyLb8LKjIKR6iRt/3cttNJg8yCK0NUhC8JFjT8fyNDX+nZK
QBUP4f8defr5Fh+WokgBvF0yUVxYRacLSGYDvNmgr3FNFPNcte/CZ69aMcT0VO4HXV1uuJQ0BXwQ
2apk9LN6d2hZTeq0/PPgFcfU2nSwGzI8lccJ0KxYCwsprxgjY9R7UkJJah0AF7Bu21YefJGSGOPH
jSlarIdcE0gM3DeCSllwRMAKY3G3BAxw8S3Mjlr/HAsS86i09dn4Jii2hdEKCPr0bchFDWvTrmjY
j4dyCHTHU5qkk56EKxuYHX24KFd5l0RA/U3+33BOMZVIUgBq/u7UAE9gLxOjgNLC3ADLAys/KMSr
EtIivDfzW+iyEaOl8E2EVHH06w2Bn5/iE1e/vEVPr1H4b7zSkYK51RzvbJi3lWB78653TXPXsL14
2NN3dUwDvF++X5XR+KTdOhPBFdWuxlNKilSxk2bu5eIJ2JV20byQKeToqCKpXLLT8firVt/MqnSV
yTNs5Qhx3zal+N8xuqedVzy4dX2Gex+bQbOzm2kVmPRVsY6/Ds/qZyuZQ3kqdFVtaqmU5vgdOqsi
DGE6FL7IHiVCzMdibNe/MmYcRUXQfNBLiOeOiq4J/ee6L9t5EFIxxJcitDwju1V3NZQEb5dRNhID
76wKDx0D9MbrTQY/sL8nC0vCWSJB5EBXimhY7/CKBe0/qjfh6knTASiR3hPEuHgJbRphCDJDKhNo
h/6gNYAmjl1dcSUU2YrZgsmB49IaSBSW6Wj2/7m0SQ1hqGvgP6avrnDptzv84hI+s1/roWA4a3kT
tzjPCNoWqehlANWuB2VWXcdxKzsV5shNANOA3DAlsa/RQUjqy4+JzkSoXhlIEJKkS1WoxgDWGaDy
oVk5H28STPJ7UelkKleNHvQS5LXQOX8X5YL7Fq+RzqWXEP/OhNQfIQNGTfJe5T+Mt4bcDOJM3cB/
6N5dc/R/eBxySBUnMf5KNaIVjUtqh4xNpHW5xvLnDlAk679JyJ8t3P4lDvNM7iGczTUyfLhyDIzE
0w2XB37I3/VRQ7E+1X3qUE4A+XAa7ftTCTjDlXx8+3/myYOEZ8oCK1ReNF0TY89hU0NSSa279O3N
hYnP1FKnRejWUQ+7p/MU8Oyxr7DjrYcDYCqDcQCN7GeD8Y2BFeRbyvPBk1LeI87mjLouAMHG9uEA
oZeGoJeBq0EU/liFuG32TNv5aNP0s41nbGzpPYDCWcmkB+/6I5y10otUX7B5eZeCzkPfucT/DGBF
SHtk9dE/CFGHTDqHcvJKGQc/iaRp2sn31Dsc7j+R20iPhypxHdy4OIsQn1udExDo5PZbvT0QmsPa
fPXPECfHyRsS5HQG2gI08e2PmBByoJR1n51y+1qpT9K4kcrvmXi6V19NTaxLdggIA8N6ln7YItEC
0AGa/wLhY8RcazwNgShgbQ94zr6kVSCRJUgh9vsycPYlO6Sisr4EyAS1/144cR5+fwktsmGnEqby
qOxcvYmvHMS/+jSRq2wmbT/4zgSKg1vK9AWgYuWW8BQK0FRmC5liE0sqi/NGSdJOXZrrT/+I/7EZ
H+8YnoaSXX7MVnmD6XaIupMazPBm15vgEFo7vmMhRIsyOrp3Izgvd74Pbh3iBxuKPlg202qatCra
Iywq2ulOiM65SAPKXlMbMeByNKSHcvB6Hapnk/dKxmQpJhLINqWIaVkf15B81Hg+7eam78FI/etD
fUKbOGCJrePNfXZsRcV7i0wINlKU2NlscEWriwKMDS9CXxxNV+3Ugo9WUYB/qoGDszf9b4iwqa6+
CaaFnYxlJEGVSvHcV4uhk5cUKbB3e3tY0B5lIbaI8uJFLAnZRIMMrfdZIICrTLUK/g3R+G9G3RZ+
T7moRwz95rYlYbDD56OIjV2NnhtypGJHZWea5Ln2+UQdq/AfmqfEYz94q1jLuOrm9H5tBHUWTik0
nV7Tp7gxx/aggPznYZMQqgrtOD4dijC14V9FL+5exOCSMk5zIGoJW2wlFBTi0NvM6udOHWKu///Z
/zolxPjWtj3sjl/UV44lz7DCf2d8AG2rms2mWb5g2V42avdFwhbogMRB1y+fuK54CwwoFdm1BJ2L
e4gOtN4QNKbw8l2BCBRTnY1SLPZVq+EProwiLsNhrg/OqqcTDm3RzakMU/ydLRn1VybX0vLKAAUu
cNgNfXOtVkAa/XNdw6ak+EiWWQ4CYLa6sCIfc7Pck65Pw74UnjOoiVExIxDkLlGn+/pVadbdafvO
gY+n+nlIuMQ1fqv7ZOLVGj2jZdj2gfAp9yrt0oimmMdpIjulEMTiVgC7wJj6bxO+YO1x5SLfZa8L
TYZqXYPQDi/Ww8ZAkmkfgLAnb7HTcAAH3wTOSjVbCRBDsfHW5pcHkrCj2NoIj2YK3oFxEjATFdRO
xxoyjokt5R4EVr43QU5GPp3eG9KVGfz5tk6O8RjWIYZ8ZEzDV1Pw83R3/f7ij/9MzhJUnv+p+r1E
9ZhfRncLAoUd/VtlhZm20DtPfjfMYSxCMLzDhcrxUUfga0ySOSrGbl0NLFLxMHvvWvSOrscwM/ue
Pwxyspgd59hPrMjbhyCtMRI5H4qBbYTvOAPEXsuo6JXgxZP6YpLN6AVYwY4pjF+VejO7LriVO4OA
029sUCrzN/2WG3IkBYtChHr8hLga7j03X/1z4TrRXEqSHzO2jNEkQDcS7T67h1TeVnTaTdagdCjM
EFGIRwSib5A/dD77NZi5TSOZRhmvEtYkNVXzZI42tqPAFLKr4N4wnohF677hC2JD3Tz6gmQ8fi+X
LHr2S0pnQdYwaFy2owWKikRLe42HDAaScJ4vJCyH2ivoevsLJGRS6Uy0yNfL4vxMg4hrP6NhWkDr
2uWxSwYcUjYviX7XAkzqv6xeOhPu2oEZNJbiIo/h0TUaBcUFurzjiUpDuiZu4DfwiFjltwBSLdml
At7669VzqQkzvUBhKMAW5HuvYS37Nz0UIDc9t/uNuRtHy775/0ENaR20hB0dn+79UtytP1DKWhYG
zHuiIGnfN10eI7cft18QGjL8zmUmmhomi+QF7prrJSCxIzYI425k/31JaqWZ/cDX9w0VPe2R7vuh
/JT3oxGHd28MmOhJg4QQ/urh6iRxx+mm30jEMm9v1+A5qlKXNMIfRa5gjxIgU7ZSbPwMLcbedD0a
5IAbQrtJLx4URRgVv5J0i9cG5fccTGdJyIxjqxd+lkk1MZxLTRC7TGpnf/lC4S8Lzhyyt2O+COWA
4s+8Wg33bgcMKxQ0C0ritDHQhTEjgARi218WJo1q0vfzZK9OPyXCwAZu2Bc3MPFoxPx/nYwYYHuU
PDCaXMihg1kXqMjhRjpJB43uqz1mvr4Y8HWTS5rblYVD4tnEcBLL/LkbQhiEaYdQs5r/isJUw8RH
bubuK9Tyip3hi4DbqLAFJ7Wm1GfQzDaplWx86QzQG/Fin/amXYs1a5h7rPpbm3RK6QqavGIGZ3a1
YKYZmJhx1Cw+yGeESyPc3n9AOUOxuWKdd0S4OZqdNGPgKPmmxk/E7yhj6iIqn7rES/kqAoCz5Iz/
VKpIiVl+5nZqQx3uHVuK3rIaUofLTGe8cpiORDqgvg/PYB+jV+ZHS6GANZ86JBFRru5rkJr8JyHG
u/S1Fjr+jNsfSWyFlvVeZIX6n0akVMLpLiCbTVHzOQXFjGus2DYDLld7wIIOk9J1BmdZ1shAO7nd
+QmIEEND7MEWghLWi0e+P+nlx58o5hi9StF4sEB/29J9KhJmDaZN8VNhjJNRjeRNIiKVY1f+hUoT
yG7rxsgGsd5nF7qm1c/jkRgrZUbeT6/wGftD0LDeJZ0GWxXy9X7xdpCzMt0SDFOatd3m8AuACnov
IofLQmuaHhRaJrCtlKj51Gyi4udFGaJsV03isWEQF371bZSHmJRswPMsiiN+OfbYsRQw4QNG9RK4
+4pU7n3PsN17PpmtK5GLIZjUvEAWmwcVBdxx6oGeGoDsXeNtSbHi/eebImeMljDrpB+NHBgT9Fr7
DDssQGbv8M3pvOH9f29JWVKXXhA90guqZKz7h/9v9ItiehubcKe5YAoESpxq7C0H95IHo/Vj4SiA
MBuDLqFKEhd2DiqhAzjj+nVXlyXa64JNelDoUGStlgvI/vv8WogA5bt2VYc6rFf5iB5wLRGI2Pyn
4hqcO34VJbS/YT3BI0P5REEc6KidtWvX7tx1g1DGSuDSeiWkpsJtXUFXSft0Os5M3uBl3BM46Bjd
IfkwI2pP1Caa3s3qyvjpFr93a3Dj2z5LIgUzmnuOwCsAiBxCR3ehYZA1BoVGOXC3+3j3Ef8I092P
2FzS2p0lzvn6F3iaWE6sTJMqbO0ESLePaLhNyg5M0qFxKnpJ1Cz7CE9JVUv5eHXwyFBXV3d41cfL
AgPHSsNG6DTlb7Y+FdxvgkcQb1VEDR05AjCCMtoAC6Kqv71p/vRF3s3VkJXljJ0zCUHFMSBPPdlm
Fkf6sHZtcZMvHfqgf41BYbXfYUvhXsbWvrERvAWb1xOJcD/AO3iRkgmb+iL4Gq6siraWnr+JY/Lh
OcZHr5rU9Dc5+SmAw34iOqB1PZeWBsbdph39+Xa47AZoFDbQfuJiPNC1rAGHcc92aFlklnVFNLg4
FFW73m+VgzqdYY5Er2FlqvMU7Vqc0+Z9u1R7Agtvkosyt4bJHgKk39KVC9y0Jn/1efFef7zDsgot
hKpjvfXKfkgPkDcatP4d1bq8+Uz9msK9CF+Uxlt8JYuKUaj5+kfbtq6Qg71C4fJNBX0kHKXaFPs0
ungZTNW3t3VyWVteqCbtQkOhWemmS+gowIDv8nEWpFCwYmGkbmZdlvS8T3z7YTKF77wy9fLCig6v
Zfz64eH+RNGXsFblvLfAuD3YNRytQBPuq/CMlBxDeOZMBz4mEOWfy1LBlxCjiyOR0UqYd0miN+4L
ZHxGjU4/Fep5SjiOWWHRTk3a1oCY7bONXrNcKSv3EnGn86gtd3uTfy8Wa7yZcW9cDvSp4LC8sleN
SDThgQe6S/FYfewWDBdse7JiGPszjHJKmEHJ6nFELW4yFYt4B2q1i06vK3iSbwF10oVYWrUarZmv
AK5QhlB7EgJxuUFGaev2VNL67VGgeb4Vdez88nAZraBIseMT24v20t1r1awsbp+ikIJyw8kEcLPE
GglgFZzUsflqRo3rSj+xKfMdpl+A+BtoZqXa/3gReeEYCsy8c9hyx3VOjW6+zq7GXP5QKMHPMKkw
M6X1kioADyU8oNF37aKR58l+Pi47+jZyGXTxPdZyjMf5HQhVW2OvzOA/k1YpNys5Q5IRJgE85hK8
b6wraghJ8Wb1V4KcnzX//NJ/jxVa+OyZrZqoS6TV0jim5QXIqojI4FkUcrL4fCd203rvTXMEFCK7
Le4kaWnVc6HoJZxL0HcJiviEFY38/ybrv4lkJdWQqYNeJOVzVx7oiV7FGvn+MLAvKjD9cJIKNpaK
uMU9TPTRsM6eCFSrSxFc7GqyMEMazZGpwPiDmJip46g0vH7St9Og223ky0lPJgyYL/zMA1mQ1SCp
O1+J9Dkolpc/+FMJ9Kn10WlErbq+28+YVPDDZYrRwXgXHKSXfTu9rnfx8gdNnon6v1B9A1xvflX+
lRLvffJrs7XcrxBL8XHt/oy8CAlQcLvBa8RvR7VJR5+duGzNJGdSIFptX0OgPuRvZkCsQ5g4dAxh
rYzw1CvPWrLzek4sMX6YSTQkbtJ6EXrOOnDzs4vgVMQKkY+xCHTgAc4/HebiDtBDYU4d0g+MnJ3e
sHiho++eGzZ+ELbpXXR0juXD9Tus77LlWWDvCfR9dAlnF6gSpTG6JNIvhomHgCxz3ZsyAAnCwJgK
FhcVDc8AhSiXaBD/xr8wxeJ7hgN2BmqOu9VljPGHA43YaFC9DvjiAjTH5rD+/8fKBXbwNcve1JPx
bDqWcEQsk1V8YgvMdp4+AFZ5RA4wmoQjyUYvdYAWzEz2bso4xXYfADeZ9/z2MTxu6HVkh7qaZvqA
N5oQFrf2Euca3cbc04kupGKFoNmaRSkt6GFdl3G3NZG6tUJB57dPkiGZ6mffTw9zTftlWQGU/rSc
VTOTTe+sSNUlq/Rb0VLZbRCTUhJgEjZ+fXCw2vZlKXlWbZfAe/jK+YqXVz8fb5vFYXO19O54VrWi
gIPRWk1vd7shdZPF7flVynAbOHoxNhsq0ke5lOE6SryJiHbINs6EjpS/K98YdUu1z7xudvOB5xuW
mjqorvl09CJAGvzhAU9gv7oMm07xqbC459Npjxv1enTrEeMcY7LBICKKLlufxKrp5umIfk7HE6Eq
D48RJUJi4CInno3bvySdvVh+gS+aUBEGbsijtzOi532gQcFTG3OwyHfEBn5k9DzGD0AmwZPB7/K9
STKFa0WWwz6vPaoRH05/8DNwqRLA3znzgcJZOnwVlX7ioioluxwPK9qWRtuBR/1HTkV/1sHXo4LF
EZrwObg1Mmfw58XjdkBPYr1esKva3f7MJa5B6eeqnnsVgxXXTqUp5ct+PPF0/Szk1lZu0Y+QZvPD
5FjrEHw/Z+1w1kxsQU5Vk/aStXWMUj/lE1vOb0xIRG7HC+XhsV47rKpcTSlt96FpQNo3tuezwIoX
WBQWpglg/DpkfFK/TncXnwEThjbvIcEEyQmSFJ/w3euGUEiKZpic+6ugEa23Y/y4Zt78S1WcSEtQ
DjTQxBL5PZiSJp49yoDjQRXHlqGTL9/f02VifDAWAR4wg42Sobv+Th0Y+aF79RpNn2TA7c20rn5y
Nj+vTkuiZcCpPjv3bV1zWJ9eTdy+5Pgd7VbmRSTxASupkH9YYAB2+RE3LW32upR1xElZ/BbknFUm
iUf0N3/ORNk0FjXPXDoFnouEJXGNHSe1gGV0KFNkYhuDYzQMxrHhhPHYyLsXHTlj7ra+M3NVtktr
pfvbIbJ39iezDmlQhO8y7KibxHuDS+JxPGr5bodAHUJl/qA68U/9HXUepBkklNgoO1dkNXjJYdv2
phjY8agUzMy61AzGyN8zqJzIhCfbktnHYa0YWhrq/o+w2XRep6jd1wkJmPnjLt+E2R/c/OsLCAaS
+cddwn0ujHhnEII3o/K8YPWuwKm4Xsx/RtvqYdctd1b3QOB86s16hkLJEZm1MIxXCe/CyALCq8eh
Ma+ulyg3uvJ5pGDArf/nKbIDmcS76WSr2Iotzhr11CCLAX8njfvak4KI2tEZxp2U7ygO95I0/ZbC
MBjjubAE+ln+8HN4UgpUy1xTM8k79/XrLdzQ43sLc/sX7NJgaN071KdXQH7h267fsDGX8LIRybHO
VKGeS1Zw/Rxz92r66PJ9KM10LZzt1TmN8iFogegup4kzgGZpWSOBiQRZ0uZpJZCukj8Nnk4z/hNC
n2NkLkIYTMNP/oRIj0Ov1GQcGQIWROb3g7fcVhBIz0SMOIbXCHga034hT9vnunTbVdokY2ujk0tD
8UVVA3cchTSPCMbqHauNCyoyH08HfC7ZBIUmU+iRIl+Deq53nHYaqr/shk2I6YekymyB0Ny4MVHW
OC+Le4OG4myr0hLrnghTzQ1ytFISNxB7iutVcaHa8fDU+m7rVXGBahGOO0C8EYCw06f2jWQHxxml
Vr14rcU55VbMaZgucSsVPQqdhxiWrt6X1zMkSx5IpXXhqu5Mq7NdAf1XBLr+Dr6zqSsOveSuMpJv
DTl8pq3k9rfCIfrIKcr3+4lrxXeygt6uvdX6W2QiURgjo7W6WKq+FPya5wFDgcigVAOB2R7lYDqy
cWmdheVCzuPhsVGp4J7BhmSQsRElh/inuhsrXCRA1bp+q9709nYM6t8CWkOnkgOaSeRCHRtS8fK3
JUyJcCuNh3UNmUhYdblKYLnolN0O1XyYFIrI/lW4u84e2ZfsdtmXa3rgBsG5bnf32hij97PVIpQv
PClRQJHY358cyHa6F5pIkANqd3p//r9ugawaS419i7adasO2rJjImKNpX8BvKjRe1vd/vsi7aQxM
4c3Am20EcCgJNe63r2U6lL+1zTUKR/a9133o9N+XW27sa8+FElumOXRSOgBCld2Y6EZjIEmlCC0j
iTVdFXnepm+7W/UKyjjtRJWAC9njyC3CeUBKSScuNASKCmKJ3/GG8vKPAw6auoEMvrLK3tHodKvA
Ds9sxDiBXZ84OxLR0Kc/0xR6QMmV7Gd9jJCc67ck5OXLVO448cEwXsG471CdMCwN5GQW1g6Pec3W
9fN+/0AMvNwwpFCr/+j+cIWlvy0sXaIyOTkro0q+OnkHY9qXElNnyPF78FMFkZrF/8vvY9VL43B7
ELVPOgnWRmK+Z9KnYXhJ7NteUZ6PRKiklTZufZdpyl8CSk/aIVGQ/FuI+sLO3zIl2JHc7sv/dyfd
WjPDa2OUfIO2qzWAjGdlmzjYPSmEVkyRh4Ca36XNN8v7OGuvwjIPr9xyAk/DMJVcS4ELARM5Lrdo
sNIPdLzJI+46fPtOuSq4nUeNtEPdyJphEoLjFybi94wmfxx48dNr2jvWDrybJftjB1/ir3747xtD
dleK0xZPH7ZJzmevGoBMW1umoPvcBQ4ITiNTBdYvUdXJgmszihdHmx2gD6HBwJ2KqyzRSfhmuUyK
GWlLrtsfsfv4sxMIBO0+Ii8Fx1h0F36mDJFpFv6hj/Q8P7MMeib71XeWHISkC28iCcCbuJleo+yJ
XiBXX4h1/9jxeT3iMIwk75EKOonlG+MYSEYhP2GXv2PVF1bxNxoGMPD7LErgJJ2+BM4ERVIz5zmH
oR2TnUdP/zjVlq6zDtst8cfDZPOdSs0Ja7tJptsnvoO4rZzFWnqkqrJQMtwoXblfHyrPYYejJci5
3hnrNndOVIl92uQX1By9QaGSPpkdknxVimKhPj8obLSO8vZqGeReV2TEWObt8V9/ltN52RsMhdtI
tTEalt1vMCbIPnIJF6M2w52p14HV8NYxMolW/ZLkTHWcpP5TVSRbwJ/UKu/4irsrOxZeHdT2TfLL
N/1gN2p3yKu5EWrydFgbyzcHXbL9HDB1QGyUg9Ypwta3Ea8H8wi655wtCNyb5XfceY5JZyeAyksr
eG1h8/mhEu4cCXKT+kIXde0KScRsAAKclNRl4Q3AZfbF+HlZfU/K83I74pMIijREJIyD0h7/g/hY
M+n1d6QR36X64vYIEmIRQhXulb+LR1XCyrx/r2cM3lMaFHbeb0bwuxeoK/Gs+F9Kf6siwFKkdM1u
seki5vqZrpqACxvkIOKiRfU6SEp9A1xBji1CqykgpsQdSxaTcCUEU74K0FEPwUp7v/ulZ/mO8KCT
aacTR+AQazyzWgmIAQwQN1onzvRa1Uos+eU7r3o+wwXN3qdGQPdaKOqADEk66otB/dygK1xae5KR
8XMpQwQnVSlOXnyMyIJqGjFwBKCmP0JN3+uIUNPaSd9QF5I4Vw+O9eL30KdzJ36cgG4p6XA4Xo5G
ksYtiu4f93tDs7YUUugLw/o9HqduFGwWMQc+oFW2ladJ6X2VeA1DVYsCd2tFtdIARdDR8qLSyU3K
m7o3DuZG+6avYc3JpTLveqlIn7YpN73n4i3vf8ljNN+IkjmikbcA/mc21kKvCnW6gwwXOwIRdI1c
eyf96UgHxkHe2IzAGSRiAWB5UzKNodTK49BNJKPz2Lmjn8upyJpBBfdZdhbbVZhmEEUjqg/gXH/T
CU5aNh/ngZWWWfn1cvbq23mn4EWUXCdW94offjAmv3YwvZjoPYN3iq8NqOl5yYVMdttFfdGVoSfb
o9LrXOdNKvb4ZqlKiDKbm3JlcP2muog3tgoxTg+0UUQQY0GooXoC9StSddOGhUSSC8dc0LMFpCP/
vjJvE/JwcAGlKShT+7gOar/5uYiyejedMg9IltpOKiVY0/eQeowCa+HECyhOnB+K2y3bUxokgfeB
lhY6Df/YarVzLazijnsJButlMP9dCfMLta9gEgQwXYuWfe8Vce7b94aF4/YMyfEeDauOrSNGVODm
rZ64UtM8vcDMYoHYzVp4IOrs8WcQAcUzbC/eguTpEdPbDXuzvLx4ntEa61HLw6BEypQV+YBpEE0X
FTf7+D8v4+VzKk4ntrisJBKRTROMUQx5Uyl9XMK4klTgTtm/ln2TdThAvBblLKdcWvyZwdoAM+nW
Ses/VKJh9JopC1LLzaX7zHMq4B7DzlPKrjcP9R/HAPkxIoxLkdNTqPhX3pRKv8haERc1CSnbPgZg
RKZe17LqkEoyHHA7g/7Yjb/8j5AM2bgMsP6WXZYgGgYMebhEUqVLox5pTSM8zsPexmq2usHmo9Vn
ZZhxzoA3oC4rN1KiwWqWzvi9fwi0eEkFSob28FS9DwHobp6RMvg4g0wTjJXYRd2LqqFKqn9UErlk
qIM0uFD2qs342CogEYdTx8ppP0G0K8PIOzGWq8jUrcnsMzODr/plaj+Ha+ivpMy60rLaphm70zjS
dAJzdUMUZ0wnRr0GPysN/0lgU3MKfUQwjebr6pacSqXypf6xfWCzTyPAeFK377MGHR82JEpb3cPV
YYpWipoFvfLPXrh9WhSiaxAjuwzi0MAtOprUefYfP+IaxxaKABWpXhWelSOe5QVFqJ04BOTjJqAm
iRON7TJTUvb6+NhXFm5UWdVJSFwuKp5S1BWb6UnKAahBhUD3GPu+XRI30iMTEd3bLq/PcXDHwuES
z/3L25GwPVc3MKPwEm4IO+UFofoEuAlgfbRESOCcznaF3XMRaXnjWfwB3A9n0Epnlo66pKHVeckT
Ylg7wQQPqq8OeNKpaz0BL2mFvrYNNYV62WRNopZ5MF0qgYn4E2faNb4wbIg6EaNLVvRRxDYjwfjT
0W5XGQpuuO+5AyZIkiwI3Q0c07wLiHJaxhtqe+bJZ/ItSvhBRWlksPIUz4KHy88oWb5ixc7pLjkj
Ov9mZq4qwH9xtUDmSO98X4L2zuXOJipo1HccO7KPXj0GRMO/NYW9ZeOjeTONzo5NTf72VUuNax+M
BVNXUwo9PclRbMNjh9XsUbCHVnbURGlBEQZyf151N0JQTtZDMrfutRTHajzB74gvF9D3uw7bFTjv
2ugn3ggaIuWmmF1MdnDUu1MkqMABaNRmOMzDB+I5YAftYdNL2XxZ8SyLGi7I56NHfOpjsx6J4xWg
eEKL1SqSIxNktgelSD0+7zOpIUjwQtj3UsTGQr3LETucblNq3LMKewvQIxOikkkFo4XjFhxKflvY
p+IJuJN1gACAa80d5DsmdGvuf5KOlOJYAYxvUHuKAu/2t7PJy41Nq3DrL9vPe94jwbA4SLAK6B//
PN3hOLGr8Qmy2VAX1LqMh3gqIyOxOHurbeefKTleUvmWUv5bJLF0e5YPDtP5zkhlvxJXgzEC/tcB
YAwjziK3nk5yWLc/DHeIIUefa+sWqQPqKIx8UtpqCQnkaupjtUzt6gocaDhUFzIQayzP+AnW4utg
HaYzz3EzzQjFOya27uHG8a6uD68aEW7UXe/x7P83Jj88ruqk2ENnVyo9PaANGW6SWGc2bswuH5Lf
622p9j/YF6hazzMMLEllteuhTRJZbhi6UCtMU62Q6h0MRVwD+Tf9MTrPH/TtzLWlRjGRpvuqzBly
ZyZMnr7cEonMmEbsfIGWO1CQjtxwNFb+vC2e6PTFCso84nxXrDPcOKtaZNQ1mwoa4KsgwzX26P5F
qCJn+7Z5JO4VVShyrhKAe+ij07dwtavWIyQ3XxFjFG/NTFK/Gnys9CbJk3plCqXu+pFG5gQvKoIE
DiRt4S2Ob981afsE/PZDPlb+f1fEpjJPBsO2VgQCQOuizveQYpWgS3FzvPyMCVifqWomHkUAKCFb
WQsa9Jp+n1roBD2GmDUBR3IJQSAYXegAwxUP5ItnEMHGh5NkqUVPJBQXfbLxYRoWA7ShrEECyyRX
wxkeaE3jTBW65i6V1tvqMaOjSo63LQVsQYR8kIsb4Cge2W1gj0JzNDiNwv1rjlJiWEbJFTU0s4lq
A1PZUzBz+X7qNIkUCgMooKhN0VXWzv6gKM8dKzLpIoIQ4CQLU5/c7B7enlwoxVlIxo/67YZwMgic
N5M2KS729UKtsJiDr9QtFiPwosGHxyvavqsIZG/0shws1jb0/PX1BJKttI8cHyDmzugApmg1vnUa
SXuGf/JQ/+QsfqfY3BxMweXXBuzmvQyCItCNI2/kb4eL5KbqxPWy1NR3lJbPudbi0GPxX9O1vlDq
EJ9+ELjoocHlBunk6NvIBmHKaX/rTMce1hltcCp3bdhomfBEpkjNUY6Mi0t0L2acavNb9OHV4pv3
6XmM0Bxgbs4zerDH5EYAxaMXQKadvvTLy7N72OcMWcVeIA97CbZShnPMRYRRIO8NpAKKlso+S9US
A+puuRWVgUAmgyDLbrW2aofNRS+GR3/a76H2rTeqXqa8X3jkeMpbS0Yrx/bubEnZECXdMofjk5oH
SDur9eaL65lhMboujy7g3pj2mOW8SUNUFgYHW35PqZlPnwicRMYvjEt0UrB4xW2GgxaofL7WVFyN
G7huUEtcuoV90XQSbYldQf4S8oKF+JftkFTmOk0n6baiSTHBfaZK6iYQpU3XzUd0LM8IKBNHbt2v
BlLdJR2m5pG3B4m/4UNNDPNRSxw9979I16WVR5J3+DB1gqt92y3V0PPnuCjDxXS3LfmDd/GVOLFV
VAP7s7VfOTJJruhEv3d/ItvwPZaJhvQdGcQGxS+Ly0pUQ24HEUm4LmKXmGhm4E6X2NqFT09roWHV
7XmATPbWlow2EI7QxCu23g6Khv/uaVetfq5Zr/lOBg2yHdarH/7sIPBigNLBYRj3W1RkenWKU0y1
dIRO2XmTkyTmvcBq/v3fxZBxdOpBS4Gc3NYRRWPIhzTy3XRwo338UDvtodqS0poRpn+/qhs/iTGs
oSS2Lr3YqRwbAXr+/Y/xCA9Qcm1Zul67z3YEgW7ImwAiuM3VJJL01adD6/N6QN2b4bXdT9TUoAqQ
8EUQZwe7WTyvMDCeCnxDH0OF9Rqk5qZ//WwOIzDhCFLPNtkYU9GSEatFhefk8eWoGaZdYENOY7pr
loPYd766cs7m/W9ThsJFqnZJl3h6sM7jrPKs+GPJZ81vhpkdIHfayXOWxBXb+pX61atGiVZZhESq
CfdMHRvAaSFgQnd6JjZDssAnjltPVHM3dnTrAZ7ijqOS8j5HIUN6ihYzmAgr6/V/WlOlRRayFYv7
PWa5RM+lMPQsI4p+4GTftgpEl0FFCG8/Yd66suWt4xMc6bDFaycmV4BRqyY6C1Ls+vBRqtSS7kMF
neMmXtyiDLY7FkFUJ4OxX+gO1zPTXbAZtlrqMYcbgwuY2VgD/eNujixt0S+maftig7hRdNHAWlmo
+vpwEA927Pf/Ptk0uzPYyn7pLGnaNVwJmLcr9xRLMe2MP8AyRPvJU5NLBjFK+LFrNP7c0FVseKLT
Jj0Nu/4T9my/CJiTM3QBPlwuHwY7AS378/FDZ/+Dxekh1oVsJFgjvoomSBUqMrde98S10lx4V19O
E52h3g4MHY25OhWUqYjwDQPzJpT3090GoxUp46L6wze0ibrq1IJZ4GWGM+mEnyQdsp/qE2vvXgBG
4Jw/SPACJkRf042Mmh4Fc51ZVSYuZetCsL8ZUoSDSF3HOgyDDlgijRVTauO1VXqNeznxsieIuqfi
bJ5y911eGDiGRcuDSxFXUGZlOX1ScwybcCWnAVBXRqPznMVyzyab7RnuBG+hlbchQ82gH7cKIndR
TghtlJjLWKZie4P4vloSyoNlQt3O5MZubN898SRtgBKLvvzfdhTtu14EnJEDEZkK7aR4Z1gVPdj3
3ZbZXqdUPpJUV+P0OAf2YSmm6aLH1xDcH4W7miq/6edoRMWsRLrGGZue94e0wSN9WAKf4lCgDAn5
ofNWkEEepuYocFvo29Ba9PW0VxDqOAxlkymhk6lVqopTkz+vK6kM2Q9fTUsquyWvc/GayNthgirs
MXU7ghf8mxbUazSVNiZWBgRTCe0lmHMKNzKxVXiFmTpZCvpBIeYo9gE4gYJbMaAOFQmgG5VrreVo
IDMpB26e4sgxBumPAzQsEdmivesDm2dDcmXnmAH8BUPUOXS9W0nKz1q9umU9TC5v0ICFPc9GNDIu
p4e6jIFTlkX/32KOc4SbhfRQhPCKRDXq2qlLfV/hL6ey2UliKfYY7DkOidvdYIiyTsyt4iASn+LP
vwgMTHfQLZsUucY17qz08QuSh6bU4LLO0luRm8efhIm4wqR2Kt/ycbFjgP8ToLXYfvux4kD8E1MK
4fhX4fnG1y2JPVDIAFVoHTKK6wCpTpN6JGWBaiSj2KwU+0EsQKt2DSKBIOciZ+AQzuIfLVBMCU1n
GgMZO/NV/MeGRNIa9lVhe11l+ih6XNKDBNBtQmI2DIe7svjB/vIjOo0Tg12aeu7vUkBqPNs0++Y5
RHs5TPTxDRA2P+BOSFG+836o1/t6uBpljFAU6I7OlhpWAHIAiqODTo8nJCOdV8mnYfd30/MGhnwT
ew9E+/vmwb2lkNQ+Gf6VOxNJTq1ZcKvS5CCo4oOG6olVhF0HSRsTZGGBZGNjkCfTGuAMwRi6ps7o
t7SWxyFq01OQNlWkzmfhCpnck4wmB8H59F0qaXtMbh6YW0P70/RDv/0iFQpX4dyNrRcL2qe77+cj
MZO4aCh8odGqxC5boZmDJHs/RrRYvs6kN/kL5390uW4lm7inHt2gSEmfRXzHpp8HORZMYfYInWQk
nUbfdpPc/mg1Il8d/E5TjK7W22kNPGb2xL/dPWv/uJhrbfcr4wBCXxWNRnOtE0LXOjRRfPFDHESt
1qg619B81baFD9ush1RlYljP9awnbmNz58eymD1qqA5tn2z+H0wyYntXe/fk35GwDAhs2LS79ZSJ
9gGMXolQcKDoxVQjR+xlXUgPXes0s19h838ZvXQrP73n3NrX5N+hgpNQGnyiXWys+L/P9MV/QEoy
8lV/+hzXJQfun0VniFjjcFvw9F3sVrIgfllFSY0b4jfs8zxhXp/vjUM0JIoedY7pT7/oaPZ0Ya5W
xsKK1xYDQTzkuzwW4GONuJMK/UtsQOh6s0+/ZeHZUo86tLjSW6xJiYTlJw55Vxtw8FE3iv1eHXyF
SSaq0733dhEivjK8EZ2Qv8bvDBiyFpi2qCQExtYaqbBQUU9yU6yKBWT+9Dqp8uzISE4n+UM82J4Z
xaSoC+q3lCs+5jRVhtpTKFQl87n6bK4PWSzNZ2O+A+UY07Qi1W2FGUXUqAsgtJXko2CcLJRUCZDZ
BjbeOYcTF1hC9cJXHeahyV0L/27IS1dswa7Y82J/D2Euij0UOTMPBB78/qxEfpUvOCDTKdSaFULW
EVZRTHyHrcCFkugquh+LMRtHJVsDNr8kYEmKdo3qKKPg/EtYJveXUxW7in8i78JZHr0xG6AddWE7
QDJkDmGDHSsN85G7Y02bqnuhtKN4MSVdZXEUi9mYS2iJqrA01laHpUGj6LyLsS+jCnC8CoFK1dQA
dGNhulOecXC2GCSh1lnP4nkCZk4RVYf4jROI/YJJ09cGSNh76TZsffK3tRycYkwZ4A8Db0Twd2DV
rFTtV73cXIMyYqMg0uePW8SxPt/pq5ToO0KMxgZUMD28K8kZNnQLjbr5/PrCrBBTrcQZTl9Sf15W
gpe6cahDfDBQLvj92HwSFuui9fsyW/F8khxC5OfCweA0o83f+1rjbnHhdLFLssDXUYzztTg5wk4s
RwWiQWhfPp1BwL2+LOYbre4vo6tcD7uzv8LrcXUaerGLUo0ymA500bXa5dqt0DS0WY496QpHZEbI
2EQwTgwQd+FzcBoPGDCyn/70ae6r5x0Je4tpYAYgP7o4fh4egM3KnRNjVGEZHS5KhzgpP/Hcw6Y5
/A4EQT/wj7IEzcgN+ZdnDN/AliXyMzIWAgUcg0V09IsgJcAMjQY7IedNSswIrJChhPDdH9UrhW4I
QAmWPg3H+QoC6somNXPOHPTgQRwk2yPOzavI/8mKQKcbl7xJEY30jZ2l+Eb1sS+y+kNT4tBaUBGr
7ihlYGsSOkZgMgE/a69ce15pD3xuYct9oA1yZC3q6o584YmJllRnxiz/q1Y+dpKn8lfn6wgQtVuE
TmEwU+L51Z5F7suYo+/71aVL7mR+kDyrYZF8JHoxyulb7okg+GhFVpcU4n5CnaF5VIlTBzplqArE
gA9+LoFzwZI3v+/f4wZ9CZyekL07Wfe5rveZCbYl7eyzSiDX7ATG8e8IFmvbUMZxEu6TVDgRcpXH
dGYLzg/KuDtOCTey6ldvxBAn51qMzYB9vM/cjmBsrgJ2ReEf6XHlo0kl7K+M8oegLegnCsBqWSOl
WAIuTiaWWTJSrf0LgvFHTpSUhJ7+SQYfx2nHFroEy/mL01MMZKUbVNevDYL7YXPjWeAyymba0BzV
h8rb8OmEMslMbjc2nrGpcgjklzl8puD9goj0Ox9ob8qSDXVBJb9hcfyoZnUV1buYAzu4MwT9S5ry
hqAW6S8G11HwaRAT9X6Aalj8X6yJTnauLDAzFLElFgeRyOC5FCrwss5UkBWR2MRTyBlQklAgO6jX
QzbigURXx4jlEq0exoU09ZBkIG0+u/S+EmE4ygF0Hu7AW34QwLfoIz2+tlEtua5doL7cVAuW/hH+
YUteE7laLvUpadPjEarQxls4bNHCbLQeRVjbG7OwwamKw0qJKAQ7mw+38JRllN+9K7kCtX5B66o3
SJIQ+0cWt56205kZABq1m9Vnv7boM045yZaOQrbxORqDV6BtC8pTZDsSz9+L0BcrCMgUNkJ4NS6B
uak74qXgKaB3In6irzWTcRXOJ91AfQiH633S4FuiMK849iEDVGZ+QOLK1gPLWpIP3io7LUSGA87o
tvRyHWek6S8ZGWIsLFBTr2mX9Ub7u6nGarkBaWat68uHocoZMwhgEsEceLC1KBZyU63YXCabY+O0
21J2balwOTIp1CtdjRtobrT1Q/dHUd8/P8/Z26XdM24brwy4au32wgH3eEzFojGMgW10cMM4Otrd
dua+6iQZtDo3pdUmElxG8/hb8jlHYk/1VSkkVOMvfpn6M8mhk9kPKtjwSzf0ID8OOjflzP2l2pfT
hElkclVkmDakwOybWukiLiw+snw6knFNimunW4vas2is0MKOVmDQJzqmQc5G8ZtbWv3uUkkzxtyE
aqm7jKctdIvy0LaE7Q78PVXXmjjfNZ9oDVasFRbH4+xjpSA9NvQCiFPMPZVfL77sneyWnAVkyhKg
UYtHjHq/ZS98/vG9IsxtyRpIW2vT8ZLICp9V9AX8P+Q+yJbU/PC2pXzxJ/7OjE3IcTmQHnpNW9VD
rIjKVxeuXojv2ajjeftocf1hyfnCy4enbTkAq5fdiJWbDTRbHkz6sGSNxnZ5okopHvnDwXr4muUp
X+f4mR7Ac6KP6W4qHFpKPK7FweUY4msbLfkVtjlReJRmtm1sI6CGZ+EtwbLOboHLrM24GjsluIkC
gCqgNR2JfdjO6nX3seRd+eqc5wEDfN3aJpruclIcNLT8TJ1cVVtBsoi1eLQU548a/Rgq5tj+rbf3
3NrkvRMqu/LilzDCA+RpDhfYDEQxvh9mrK9nXitRN0nYY0oBdRmjSMtW4/BPPKc8zzil59LYvxL7
95UUjTq/joSM9cIDvGRbcsUc6sbtFO2qipzF2un6HQKlMPSDqxibSxg7V1jaU2ox/0MXGLPHmmw3
T4JxiGyeHdKJagGWB9FAg6mqy0LRHYOZoOOWhLYpbwdjVgC2dmROf+h33mN4e8erNGMXNGzu6Qje
5r04XXn5Nw2QtLX++QnfexL7EDmazwvJmL2e5cS6cDN2XGs27yyegcFhGYVeuy6UMN06r+jz+hNR
mHOARv2PKZSAAgrnnhW6+J7eq0LgnHf5R7RWolOpJ/PFckTh818trAF9l0ydlKEVfPaQrelYpPHH
ALwSNt13tTmadaCOaGvuA8sRkJVHeWQo42JGUOGLBSNck3/0rm/SE+N9yQTb3FnvDD4iaAwJ5vbv
Up3jUj9zcHSfnefMv3PE/WqVlAiLW0r+YQWu17Wko9BH/qlh2DQiq4SXDoCYCQP0BX+wKxMHvzrX
ETK45i1F7sPFhJvFE25u5AIxzyw+0CewJr6EAvhFnU5zz8ypGu5jvCXxUlJ967uoV9j4op39G60V
TFrb8xYQ0fCzoUBLw/UivomvhQJp5Ji7kwLZ4AO1vBn5sJWHevKVyts2nRab6mLrc3PTPb9RW8nP
l3OBBUHpD+hKdlFznWoi8mfOfBJ+rUrsAjixEeZxKR89K9fKcK1sNBc2Dm197zWb7Jl5nOWKjh0H
eR6ze+NtENN8+R+U2xOcwiGm26OpIy7gZz2qbEbLnzqjeqnLZz9Vo5WLJJb2o0jnZYSm3eO5gtsN
N1UewlrUOUOsMcApk0LhnK+ZlK0cctp6//2KFkYL2WXYDwiK3D7fkHwpaP8bAh8fZfHzEqAAJa3c
SoFEBLi7jhzhJc+KesiXRmsJ2V3KVdzJqzi7UknbuD6lTVwnU6ONmr01KChXTbNTsbOal86i1bMD
1rdjOlDTjZcOOIpvgPpgj5850fY3ihDVoG56S09wUAIDxZHb6RiuxKwGiLMc0ORSczdyKoxhppjv
8C9YAAWZ0ABzZxaBY3Sjpk/0sfNRbojI2OHXM8Thhq36h50Pc5tlLsABhYpf8ZQbdkO9IP/xqszy
fQ6aefg9EjaULjGloIlVP9egDtVbFg0HkxoEILtKAmKnx5SnunxQczvvPFxrvXLBEhOe5xNk0JeE
L2zU4+J/4gRweOq7irOL7Ib0DodndJjQR7mjAYQBLBVUKfuxfqxxj0qy3ztyaAKucGv//9F8lld8
y1KFjvAcjkHKzwl+BoPDtedIxXziKnu7XB2ynXNyV1UcKGRfyTyh/BYqzazE6Qm1gAqcAiW0ALYG
Ug8jTPu9okXkrzs0YMD3xBdykPulLvvgBK4JPQQgJhwTVQAavOMPS7qHz/Zw88RM9ad1LCBXhXTn
TS7C5q9VIlyldGDWpalg2z2GXAuOgYXDWkrNgLsyJ7mqGN8sgLjtRcehHjcscsPrvEjiWo10NF2U
soUMjqBHj22+L8rDUP4yOxqU+EwXtUfaMcpiDB7IYT51a/TSMz96XS6PXrZqV7NNnu1WFwcmvWcx
OyjhSpTTc4ikXBm3QvZHpU1jAd3rrY04Q140d5N5drJGqM49omFq0G00FtlYvlvqlq0qWomrNUFc
vK0TZjJuHNXrVQ0ql1hzK5b5+2KF6xwFHDE4XED6VjyE8x3ibKODO1wT03qD8aPppzFhPfHhUUzA
0kG2Grt5kav14uQqlIZtHSpFHgXizgxwwtyToae9MnUcnDIIQ5AeDtnfErb2jVxVaHZK1doTLzXF
gPfzsnVeD8QEb248mtpOC6LBKmAXCZbjs8h+yStiBj8VFqg5ri92CDBoFMDFUdSRJFICp8w7KXcp
p0HVn4yq60qh1YDp00mDzpwlgADABMSiLxaHYnDRmtd7fu2455Ga3lTXlhbToul00HnVTZ/pjb05
0w5LGtIdBb6oWv6GqZSOik2WKBMxj4c3RA28VbGVftQssjEXQoVrNkUKFT+LC/4UlgiCWRC0y4ES
hpD18k9QBWaoNBUHYwd7FfmrqkKP7hUWtMoi0L5nZx/VnfXYF/HASXoAjuFiin71o1ny8jVKmfUv
KT6RxzhaUEzk1pTH9cfI3s3OxBOLMKu/bHvxdBQXHZvgGiQ1xzdL0LfO6MHz0xc4M9JrFEsYM39D
yOLn4DhJd/IOjmndE2lihDgZT2XxW7+DY0y+wqsBng6n0xonpYetDZQqdo6GA9t2mL0WerlMHxo9
scm09+YVJGXK5JcT+/jbAUAwz3bTz6792rKIohRQUWddgmiC6Q2fwypgD2OZS1AxPPsXT+o20oeg
rRD26pWmRibiUd2z9jBUj16YxaQwhFWWm188FihMuNz/tApy1Wy6WpELll/MdXYgJFQjcq02urQ3
diTzIvlTpLnOwNvH9t2XBAOZGQa7KWCf2cfkQ5wo7q04kNtqQfVeV9Vxns9KH3scsoeQESjoyF4L
s1ZQ2Sb6QO+92IQlJ5spg81F/J1yPgye3bQRZUPki5gblLxNUt1VXt0zcruqWQwCEfiT6OUr9BP+
N+hjffzOJtdHfg7yadTI9FFAZzLM+JO8TYUOVo4EWJH8mLpmxiL63aNudH4vCpiCpicbPE+U2/2b
/vp5kUEseOEP5/L7Zi4attkYR6tKolqCxk14kA+xPfolyRdQ7x4P6+irrSVhBf0cw3IGtQ/PrKhr
lVth3Rtn8bg37L6x/Mx4qwL5KJnZLub2OxT/uW06Oub5l80NN6GfXuVqbMVG4qWbof0ih7/Q1VTc
5hwQCmutPOA83QvwlgSsYaWjJBbP+uWz3hcPWA6k0ohmhrm7impfFZyMSdXGC1FN1pp/vNXj3hbA
JL+VO7poXy9nAeSt+v6g9imCHkz2E4XhweM+e5acO63naCSJSS2lSbJsrKQMxrQcSIXrvvi8DBEe
3b5KQoB+soa6t/ln5Pic8cwub9C3ewENYNbSKvDK5Soyh9mycuPBXNp7oHaSh51C6fwy32CYrFUZ
8KGQWMcHibTBJNcJyb/ykC7/cIji7DynXpOiByrRGet2EZaIECMpqQktjaQgPuNHdorlGeAO7OQf
uNskl5VygEag1cCvKgBn8GqJO1760yDyrkEao5P8qDGNWxXG7D2TXn9q2Wle6iAEcHM3M0kavuzL
hFgnwBKC3Xgi7rJ0Cni1oOLjmj6L4tS3sWdtSX9x/xcFbgOSU6X4GQSXuLa6xJZLNwRaB8p5vriU
Ky1D5qkbG+33aLvYUt9KfyNR+E+kKCRMsKmJBkigLQlfIBcWI8QMSF5/XZZzG/jMnGD5BP/yg8z6
gJtssdV+m1LfqjRMspHPNNeHs/Dhjy8enNRrRBDYN9Nuevh06PCha++urRWZiiUEKfDAeaylm+dV
RhZ1/IJbo6DXJgJBEbaqp02edXI2yPiwpt3aCCg+iTXWM01Vwh1gpumYgKwoRAnfT/BYofvUBk6Z
80/EdOfhtG4Co5pnrc3L8Q4yhzC5LBWGvQ5/J6TnClVNDCkdNvi+Z+iRCa4nxAC1FSrjfmIUwyed
cIfR+I3nHDYAFAZyb+4x4USsJXTQbcbxm1kq92YwXliQTke+Hh1CNocf5braQVZWDCWfrRv+laJm
PFBBLW8Q8N269lGq/YjH1dhvnP328E0KHXXvMAFMXCh74KVgTAyc7ldzd+gjTyZ54Zreb0w0B/wA
Zsccr/Xpo21DGRAMv7VhVy7pGvsVK0NO0A0ft2FHymrix4aRswAsyQGCT0JxkpEb9mwGFyFMqUv4
3MZzLsR/NsnUnJzS3CJh1A8G7f4sIV01B81K+zVrd16tPilCMCjfIWgGXMiGDDQLt7rm2i0/nT7W
pZuKsVAW5MArdQLqwp3hsttPdTvoZgz2C8RCgHon/PsNT7GS6bYI8PcMgJ6lrbBP/okSBdolVtMr
vXUlmDdOMNYEc/DYSZ94mpzf8x3UNv9fPdFv3my6Ir2uOvmgBOkoDKQGQV7apDO/UfR2KEotlfma
7V0Utgn/2Tp4vFxnsSl1An1VcBcQsFWWBTVnX12dyUfhxEyE0pyGV75XQ/vQeWohO5nrJQOiRRm/
PeCN5dnSJeK3PJitmnejRcA5nSFSWkPil4B0ntLeDHESJIhjyAEOGrebgjrx4uKSBYb8tzHNw7OT
tEmT6qLijxXvbcP7prUv/lhQRuCtukpGebXExLTBPbAYLWh7NdR2DBC9i5quGkznlkj9IMRVTx++
XDlJnl0g5LwHGNec+yWcgKcP5Mx97UG8Rkrfhb3FsFFVJQdg0jLgDre0//XwPoTIBGcoZ6Gto123
iySKEoao24MK6e70oH8nx/S2h6oziADDk3TW/ckayZIEERWR2KInE3GnLQcJXrM1ZUSZUd2Yiw6W
BLRByKyVVlKeweBQWfJbLfpEffA2OiZHN/l25tXi7fOZDQiBl0w5u/5PnKMARMk7vJCiHBSLOifH
wNemd6reWXD8R0scHxfezthybMovZb2g09OIdsyU5cby8QegRtPaY4vL/jjNw3iqF9sWkZZ4pft4
4kpVGj9hluR9KoJUBXmDBXSdOzcr74wJ+ww4qsrcjVmuz71NVeiBZ7GT9DrHgiem8d7mNYNsjJaq
qbsJljRiUBT69/wSKkD8u8zWF4EqeE1IhVVrpyDKti/6l/dL19cUGaRulTIG5eP+gI4/qEQdxl8p
qmcE75c5ciZ/35qP/e05+jGNhIpAPokvaWf/uS/OfTW7KiWXSUTWdP20D4q/w9dvar7UIxRkTetB
8Hsn1HOpMXLIBfAhFtK20uGzEHePc5sFr5W295SjWcXdEbxMjf4H8044mw1gN5CWxWxFf/ORzsmD
i3eIRP11AMS8ynHB4sDjo0iVIPYu3Pu+f6CPlIOyThbk9OJDD67TTWDAE1hmeStiVWtOKKTOnotK
QifSUMTLZjVOpVU2ZrDR0eeGQlOfy8PtgM1wU664Yyyk3AQl2A6dy/CLWtoFtJSZAtigLqEAHfWW
RClci9heowW/AKyjqhwEnrpf5i7qNEzu4x/JTZKxD9wMaYQDbFa+e3DxRAo8YdRZqc2eWzDra9by
65ddBkhDCd2d+doMg4ZhrYwt6AO7dEbyhZk9XIzB0eCXuSvvGJ6aL9Z/ly1kKkE11iCJ3HRyAe+o
lBrfDc7Bn+fLq05DLy80GH4Q29zudthRpTIvuyc+qhWPFmUGm/wuAtBHsI2IUduuaWs4mSeif2Uv
BBfygvdQmUVmD9aPahVCZgwPF1lzbA2dPZYrXE6/HIqKGJqTnuiBktEokQ7N+CCre53LQ9caCKkV
Eu0zU77CfUZMgZNdxZBIKBrPxTDR6QuingFjIDeRD3JVGEx9Gm0VJnx++bn0lG46JNVJRdT0cpmN
NUNowpl5zTTxwfdJyMto8kSEZNxfSO286ObEpTNDPoK6r9vWjLRftgPs9S+/sV2K6q+lNxnc9T8U
GytrzQa/Q/eaPrkOy06Y1NagNUmTzj4vg2Dg+Gl1+7j5BhqccgJ4AT4LZL9IurLFb4LlEpLyMPkv
a658KB3GNWVJ+DChuKMOfCXC77tHBfjDAxBSPVGn+k/KqXGymNAF0QezWljPV3Umr585/zKiDNYa
Q7hvpIgB4M4oRvktzj526kOnARNxsMJFC8Pe4afO7pMIeoeY2+QmrmozrbEHxt/J4zk3FpMWNpnZ
tqqDhNWjp+4DnQqotlVhL/8F3GVaQMB9xX6fDmyrH9IG8GHlrUea+yJpbokeXgUlrbWjxtunY5Rc
D4RgHBSvFYR0/ZMU4XzJjILivtnJbnnpBmj+Yq4XDDztcwL1DTtHjgTYQmiGnREcQ9uAIzz78K3P
ltbAs36t8A5MoTospONnOZOHMEEC+sz0QeQZpjDXUHi4KWAAi8FpXvbHJHX8apVaf4V4X08JBLX1
L7t6c/98347rhHT1KCvI5eY4YDbQTg972lsZXC5zr5ln8nO++ow0uqFG6OtacbghYt/NNvlIjMgk
iarjkAIhP++mAx+vTpW6dLQfB/bFTP+EMMLK4Vaec8btU3I2HXACHtKpZ99QZTG/3gfQDQIEok0Q
kdfGSz787KfWlUF2e50405IoBNJuMjGeSIEicmbZS5+BzSM+53KQpLisGWlSKLvl+ICeWZyTjIkS
NKljj0MTMF1akNx0hq5aTOUbtys4NZsWfhsAlb8rr82KNP3gUBQWV/a2qWIqGnjoZ7it5F0QZ1g9
0T4aU3WeYhzALG48kOdGZTIB6fxYahtsiMgAqV4dxfDHxwWXzDGhoFtLuJJy79u8L90c2uXmDtrf
ENZW3zZhr/1mhhztbquTeYu7YMUzY5yGcW4ah/aLnBdP3ZKqSdl1D8YfsyOVVbXJtFaTY+WwBbhI
f+X30QeDZV0Dm4bbiHpEjL9gOP0jcK3POR74RcXt+y4mR6CwgmlidyaJb1icnCvf3L5/Me7HxSUj
ra3VU3pIvN0GEm5xsYuuGNV06zT3sVHngRB34G6feyhjkd6G7YrZZiHs1ZsdwVTKG6LDAQBmROIL
nkuQDWbNbYAcxpLT3mMnu3/NC3tW7ePNBnEsWf9QBKOWZm1qUu8lI0DaRu7otzW+Hx1xcHT4Xjbk
pyGiov9fzMc4y+Rmkl+KiGZXw32s4Pvxf2OMyCLdbrHS5KYWffueyxCjBAn4liJe7xNb0u4FLW55
hdxxdJnTipJ2qAHNRV8MOyrlymDFuaxTkajcNrXE2xYHxcW3IglLSllDjGkgBaSUQ/i6lVn3kkIH
8IrSWy1T5QVoJdb2LgGFGLY4L5H15GDL00rZM16LWzKoAfQE2xCXgQYwmLclysGh6eqM3ryOv1oZ
hLoWmEYdPAcOm4huATSY/ikz1ro1lwakdSiSQ2jveDDqOyTnE6UgXOBW5mf64Pt8ut7D4gn6YPqH
UobCFzPCnAOhSLLZq70iVWwtJ/uIxFBRPV7mP6lCz/Omt5Ck8FJOspbjLoWbDsyWIlGlqf0WzLqY
jl6hGgtJHXdt4RY/E1nEGvGQ2ejIC12cnesa8TZSNYHgFcf2S8GnQwddb7XzZfYf9re+lCfLjPY2
f1WnzranQLctVK872AVEp7ODjGHn+JY5VFKzbB6on6gU+pW6Fi72jXULnYz0KMVr+8ZGW+Fp6gUf
Cv91Me+d5L4DlynhYJvsOH54XpqOtY0wot/ryyi5FkAoRM2zz0MwU8wVjl/yr7joefLev/fBvk/n
ktwS6ikTLlFRHTFfrcBUBM44apUMomPOcL2q3STyJXLr2UGaNoh/KTnhY+R9QB1u0MHE6roKD83P
v6o/HwrDGQiH1NEHRMhDi74/p+bTHtlYfk0SR61j5PLC6FYdv04j0KChJ4x9Vw6Y+ceBjFhwVUDS
YukwWWyd+NEQx8pgE1XkU43g0QF5rPNPwtqaEcIdaV6j9A9niAVb2Ul4+P5si+x+QLovdRMIvD9u
HRb+KdE6rhqVGSp3UaAjzQTG86EmB9JzYoxkO6qSrHVDEQLORTOkN/GCwYnc+wbXyHLlUg54/IGO
AvSVYsbqpmmmpI3F78Ml+dMMMWOzIKkVZCl6xrVQybfKrzA6eONCWuNYKFmlk+YQEqWxyM6oGKyu
xqejacRafiBJD5Ir54EdyYy9vaHy42RxZAtm/GRvH0Yofrie/kHUBDW07KS41y7LhZF3CkFGUb5y
M4h8qUgtgAJ7DtHwDYqpG+KI+vZ/G+/K6jCyGiTXeOvfv1ybgJ0fb3yNEBJbqoWDsQ7o2tjWB8ni
+lUVeqsYfz2I9+TcC+UEVqVEZA+lR21K/g1/bjHuaw/n6bulrVJctAjS7Zx5SIj/l9leB2ccdwYP
ZMkWL+W+eehpsRMhjKefbpRjT2fYYM7VVDI9j0KURf8vWoosWPyALexRRiYk2VwvbFEttKx09IuE
0ODXtxdygPFkdaNvkEDbglDAsdPmPaDxOmOlo4KmWIbUACQvUwYl4kSHAVNw+gXx/hhLK9U20uwQ
QSu+zX8asYahlFjaFwR9/2QgjWNXV1m2+N1uacHdnmVSv+4q6KqNpIOl7gI7urfUQW1Rheqw4Lgj
fAMsD1potqF6jhnBEH7DZFrMUfRhaIxKml9RvIo2zYXrO4JD3VbCbwaWPxSkXyF7kj4v/eAqak2s
sERHRyOIPQwSW+hFxomjSCQECNtm7TslK0ZPQ5XRq23t/YZHIXbq1mlQB/cM4flbF72VDKznIWRo
wf7PjHYLScK/ul5Z13m7J/ei9ss8Uxo3NCI87nl8grQQIYDpv+cFuCVGxtihDlFJjA6frXMfjWy/
kVTJXajZvnBt/hzE5It6Yj8dmxvbAW15gzf7fzmmMnipAtmnkWAomhbbOi3RBkDX0magWeS8QSb0
dbNjl2SMK6+bB/ZX4NNR5IOqEPumgz27dDTJkqU8P2ZftqB+3murDUpiPolhpup6Han0BuDXyUQq
hWhj2Eep8YUiYFlxiTdsS6eJ0GaV03mlECMcFHEWWzKWX0G4D6A/I/x7Ywe9UrhXet+SSho+xMxT
5XGwtFHHnQVVvUJWe1Sli71+k38gDXgZxteC2D1NLtmMcMBImKc8QgRD8RlcYgjP66oOmizkthft
6vCHHe1SI7QbrZuIXUSbmYv5PRmfnZiJgzbzSDAwOFy80W4Y7WOQFxcNDLa49WYhLQUfZ5drdjlw
hqsDkPlRYvPxgwsHoi7iJ902TNfOzDvfTua0HwJkgA8UKTWafHCnP3BduQJtKetsTMf4y1ELbON+
6/3sXTJRqYwi3xuJ/44O1rZ49vLeUiVx8h9qGXxYL8E0YJTWgjpmeZsYzRTVCa1EIR79TpP+X4ZY
MQ38/DcwNpy+EA10aQ2/z48aIN717AvM88MyJ2KdvaIJZyZVyNhqnMohkBdgMR2aktFwhIckxLU4
BbELX35ui/5qJJ805cCoovsf1LOVQFJ9sGVDC8uQ16geIWfNU0AtdRwMkhaUsgPqSaAzD3jU2YEF
QGdQ2CJdrZA4omsqwXitd3xTnp1VnTJNHP/fhfC9TbaRkgM3JUQFN8qelm5Pra46CpNzyYRaO7Ac
NGdQ7zyXv3ba0CNWUOVyRI+rwuPMXilqaBVwE9wIlz+hqKK3Bn4MAfKt15uHcV9gWD32FxEwWdTp
HvlC36x0VSyBqq+dgjELMlabhpuQZXiwrrJf/RK4QDw6dtqbDmgycOvZpG8Doo7s99KWhNYE5hJC
3g4G5CNiyjERfNAtFvz9rpCWrdnEJLGYo8yzQkQyEgp7K3Ih2uH1JHLVjzGvohendQua3TJ9AuH2
yTJmKBojZXtSyYwvDUYlv0cpHwbaWcbhk/d93hCY4Qqz/ugh2dvHpZes5IrSGiZxpUaBBKVQnb/e
tTx+ze+ADa6Oxxr6iFo3RHP4bndSlft2YvO85lh2A6wUDYykVx4hARTLSLzF3CwcqOZ1xhFshRKT
YWKDBij3Hy3th4sOEzQN7c930wBC3JJ482FYNuWC4phOJ+5u184L8/bxWTMfkLJLZSiE4kE/MTLs
LnvAXMN8fe/3eB63QLGmRHVsKG1PeJYWc6Dm3ZFUvrGMQ5k4i77GNMw5rRgdSwAIQWEFWPi81/NH
TyN0cRDKdbG0Tv2EwXaK8fWs0AZBlESlTZoOtW6E06f5BhDWWC5SMkktj80Xe+R3zJGVL8ICaBhp
1dRz/be7O6vbqGVxzIzjldQSEVpIaAml79qZVefjo4klmj2QE6gHl9IFwfe+/w/Ne0x63hVy3aEG
jC9se4n8imZYhu35TMzlyk8J4snJmwYiPZmQEzfM3XOOrKtcRkUT/Z2gi/8aY444yo5rd5Fqg96F
0fwDed+5J4PMFS4nXZemKAyZpVMVtSvZkcFwrUvi0y98ZbxXg1j2B+jv6lYhRSxjqsPSVDzVD3BD
JXAs20n2vZWeJ1GrWN4wlagdcbaW2iWqzfjx4TepuVghrDorArI8M8s4spi5d/o1ajd75EB/SeMA
BnsVHzprmK763QHoXZKNq9ldcQ5u1k9g+JCI9sP9jxXe+Bkki++7Rri1Thm5XkCMZf0iSI1d2/f0
fNRxZH3573lvZbXCRel4s6gSCySaZ/uvASL5iQKUMUPYQSNrR4zhdWK0VS0WJWyGumWtHkkvLI1p
e6MUdx+o4UqJZgEtPP3btE8k/smQF79ZfxNAZO0qTNbo3PLww1s2JWPQd66ddFs2yra2jqxdzoSX
znBBkz84OvvjKLkHeeX4JFqyBjWAJCiUcNvxqN174jdoPab4JnxtMjnP0Xxvq8TuDi0IL8hxefq1
MWHaHp4a31gBK6c1oz32ERxFCEB9XxCEZ/1zmXzsrbvdrUkaXAAfBaJUAJ5VTnMYQ1m1gltHj2ns
1Um+vrAFFbENj9jiRxsB09X2IVLnhGHqqeqOcsrpCk54ehc+xCgjOxUURZjChlUbtHjs6Rq7fAIC
IMzp6zzZB8DcOokSV8aTMslKdiBpi+zW4tmZyHl4ETl8gBqe27DNUL+yNDPaFBV5ckuURGaXlU8s
7nDXvd3/Y1Ma3CWDVgnBDqhbxeGlD/f+7OWxsmNg3lEimJ3icRqkmHYn4M+mwvHcV9rkTLWcL+4J
6qb3yI0JGb7k8BSzIS/MLXSow6xUn0U7LyxnctZiH3nIG1EB1p3ActsIfmt/q3KmrGktpQxtACfx
FGOoGiFW+6z+etuXCa65F71GQawO6Zd1r2aPoKEjz03AiT8nm9ULLFR6LYm859gJpcc5D714L6sj
BQtMDXB3pHLymmarm/iHWOMmPmjoYqnFXpX3UGQfCyKkb8V+9fY+J+eJWCpmFu/O5OlZUk7EppLS
ZeqDW7QgwhTGVHFOd5iHL9GhB7x1MgfEX+rGEW2iybWDAplKpzN2/FKG2SuchOyYRZ/XBvYGLoWS
BysxNZyfGEdQ1ZDBShZUeSNYGmBYaPhErEn0SuN25T08UcS7dvFa1m+f+sD/w8VRXEwTcUcqv1Ia
G/PhdlBCaYXo3dI/BdoxuxNm00JXzAt6p1ln02BcyuUlgXjnibhAf6tgL0fpr5IC/W7uWP9OR3c9
Ero61cKRl1EMAW3xViisxkFdUO/zI++j5cvkw0FED3FV9/miqAidNFcUU67LNqcqM/D6z4FJcvVF
YGJwWw0iRDbvE2VM0k7JqvcZf+4XpJOjHJwXtAZAKWS/YVWtmeBXdXbgxRD6P95D6kn2p1+FdLq5
/1swMBY4045SuSDGU6sBnG812jw7jMTUa1TcSLTi8ycggOqPeFACVrdpWLDkjL23LZHc0sBYPlYN
EXcLtUkYoG28l3mWzTwOg+hugodhojbbBnaSvK/3C7Ixe47dn3KSonFeauvII8aacM0yOa+J+9Sz
ltds5hS9+4K1VX3jJoR6imHIUOOQwiDrSbUVAJxLvImi89vGFV/BYg4kVnZTnzr6IcLWfzRXR0d6
6EE1+QYHZTVzYdIi7VqXH2M50v8jV10wTT/Z4hP0UXdA3kIX3Z1o22b2reAsoJcaHGFCkqarhicc
8i2xkGMIfLNGu2RaUKWzUrTVa3qtK6Trzyg0uwAkUsK9ygd7ym+HSwsFpuR3yADN2TJV/i08Iu1u
VDCWqTm3ox32zOHziXnkz6KWfXHKCwJ1/Q1IM9tpSMp0wNbu67PfQtcN4GeU+BPDPmY6iW3Um+L7
nsXpCNMNTb6SukZzS7Hfs6LUNszgiy21o4ascHBNKIV9TVTtthRB5CzelFVRnXBB24mwZxClw3Fv
SfxMEEANmnYIC7ju1O6yNjK1vE6Hru7muaJKGvacUl8OuB1F8IpgI511rjdaMZnxGez8JYnW9X9k
UjwQTTJX/LVEyrQ+GyZuh/NW1L3KjMxD4Xv9RqcJJW3KdGlDnDjPHZlTT4PZUvr2nLI2o8XAJljq
1w8S7CxoxU9N6hVeOsthB7JQjPCSXspNGp4TmtVAyTQHP5LNiDXiuPqF4USL0bv/lXo/88DT6oFC
IzpbmtXX8fwojNkMvoj1swrt4+LqJe+7CCsR3Re0UQekHeIcXL2U/WZ7/W4AMY1CeLM+RWKhHuZG
dhkjWqQgpZzoBOCPvpBFWO37IMhhbo7aNHiWWSf49FRJlIDFnEf2VcdhQrPJpMcYbih8xm5ihQ0M
rtFm/3YzOJ6AzlxjF77SsT5LuyawD8/awYZlTOx8KbgvVl9h3Y4NhfuQWAAxMjQk2X+dvCWYHFAF
4PggJazVDAOHvW/ZRyQ/nz2vG32KLp9WSrmz7E2ono03vBMQSzu4uCYxJ/CMNPUZhdQhGJXSS/Er
LZTz2FhSnM2fdb51CPifh83PTZtIAk4j5QvasfyEbcIEIPd7ViTrw/7jtTgD4CvCUx5MMK6HuRd1
kdNNtb/qVjkvM47TDCl4bsF0CwefsexYTzL/IUxRnPZFzPt/YYbNj51t+M7zOEG98oFQYCnOndo3
iR7DtD9yl+2/+GX4358lZRraRx5oyeuMo3FMz/L5F5g6Ftf5dk/g/ZHAWRZEHGr9j5+KQGcObbvt
ZncPCU9LUhZPvufcX25lpDcEJRcF6oPRn16iFFrUftnHfsB+0KKJ7115vSJUrEFsWy7HxQwT0aVY
ud2BPTxMUExjMdZ35oXwlXIluLP40gQf1kbs83i+SwRmdQ4r5TnuluNcyMbXnS3H2VlPI2N8yh+U
RUNAm4xLgGn8hfs6YIu7IqMdILtdoVNfK05wFNlQFcbaoNfTjpLvZedrVJuJXiOL+dgNPKfTjnbo
2bBNdL96/GH/P2XIrhJp8FiAM1GROK71h8PDqt/WtA9lmJ6hC1PIUpoTSObfbwgDdMV21jQY8EB8
gkCtx4CwNYTee72X9+b2AcJ2MiCgh6rQK5XHvn/XlxnhpC+KsbUifibIEe6a5BQzJ4QCaVDjv+45
zfdRLq/RV27FNXYZVyyivZiPzDeLJvHNVBqKHKcIMwD6oCHU7M5XVIgIuX5jQvp1sIGorLTZxxhU
Rf+g+UsincTcV3tBwKt/fVrbRmZDpX1TaEkPkZCbSsjoAX0L33nchkX9OGaeQYHeMuOzv7kWlYG4
EKJI/f8tBNkT7ADiLK6sPSZuKBOSb5o8NCkIcBovCSxPo82jjui9Sks+dhUTG+eEmG2T4tnhYiId
o23o5G4XDRQYCHYwXLgu58ibIunxDahpx8WRm12MKpEpU7sspCwlW4Lcdl1suECAbGckBfLZYLhC
Rnl23zIDSze4iEC5x89Ev9jh++WGU+zmhjI4pAY2jJh/4JlvtklgVZ9NmVv0HCMzR1z0bx5Ni2hn
SEAXukOJT7585/DNK6fkLWCVH1VwRaJzcziWmSUgsSA0eAQpsr32mkhIVg+fgVk1cq66i1NnbP9A
fD3c6hF7PZgWz22rGc6ELU1Ds00diZJuNSZ7zuD9hIHHDiDZCFbEq5f/TlX9BiotzDQ4BH0D9R7+
QocrJl/c3sBHwNqaQiiTag6qLnHPMVKXGCxwhzBdceB1MpVJilxGNzN7BUxoIVRVyo/9YlqmizND
cUG9VoPi75w2QrEGlwNPy6LI7fUrhIgurG8HVQRQMYVFwMagrCuNOzWvepeOLaIjEv4urYb5FkrS
c08oFe3XTaZI8Tb+gzDJ1VmqhXmNfwrUEVKDDUwUicN5YONyDkufF2MDmO9z8Q0o2GN49P/lNgO7
K44YRAqam/4DJQvWM9RKFIndI90OiB90Wot1hTCoJiKqFxpkvLcKKPWsBINYc6Mo/zRDLIqhLt3+
o2ohYhV8OrXQena/Jd4YCxxDr++sQr4WWbkubBRspcolRidzmWK+JIZoexinoda1isw2Rz5Bf07u
RgaJE4NK5hZC9hDLOp6/mXOgpCgB81pDxEU+yQnQT6Z3jB5muxDr0B6aE8anoCgcemAOQUD5nHiH
W6gX65AgZurb5vwYQeEXnCZY1E/jUzeavTP8Mf12xtpAT8stK/Da1yxKeCJwvsF2eUFls8qQj3xa
Mbs2i2NWtlrCHdfNt1i1j79As+n6aY5gZKAUUopwEXk1BJIgdrsliSo+7wS4WoZdJh6Ccq9Slgk4
sb0PM9ulxgBy02Qjk4FQMR7Lls2r+bSYmyFunLk4EoVwVJWVcP0vwlNUHIlIn1IWJ0kGDGT5ui2Z
qJzVoKxPBMhF2G4d0I8Sus2UI8ZGJXvrZ+2M/LjbkAJL8PCKS3ARbT9fRBTCOJ33IIRT86XzJNB1
TseSmdMxtRtsBwLb7l2LB7vgxDoWFObP+0yUjz4YzImigmuBSTAf2Rf3dkBikLtS6oOpRGTKB2Ta
iSnOvFN18529+5U2kZyUw+A9qjJcfDyemrnDd6YCyCPlyCSsMIsbLhdboXai+YT+YzsHIrK4PVEG
Xqbo59HJvTfL+IheX91AreNuembqJkDgyYuwvp3MQPr8FPrFhjYENCxdXV68fiXtVXeKyZPvx2dj
WXeHmc7jVG42EkmEEDECWRpVLgpKGByzTGlbEkpCEv6Xd4K71eoSvh6q6V1zTy2XglqHrq/Ytgfx
WM4QlKVDrIZa8uhnmA7FpziB717G2wRl7NGJlCiyD2o23sbsJ0T/jYme23J1mwvzhydChM5hudK6
S25ui2BONQ51b8048IB0FsYWryq1ViX5rPQGUy0nos2AWtGSX/KpEdpXvRQm+7jmtfByqm3SOIeK
gvpeH9VSt8/rW5Q6Ojl4BkbYmnhFM1CztLtTwQH6XxKokG0BANXf+7JtsjPqXCwcf30WDJMQ+atk
SuFIcgsomzsBdCy+STGTwJlzAVKz4pLfyhR8XRppPbEYo0JAC752DjsiemvVn/s0lg/m4DQ3PiUc
V2WN0W+6zIZhD9/G1TFmMTOZRDbFPSbYR+798EOvDGL8Ksa5fD3UdePNF/P7xpuZS1DkCW8FdGJU
d7Cl9uqNL9XPrxd8AW5yqWiGmGM6+d9SKkhvdWCrLvSvbh5BdlpxyO6I3/7h5hSKYs4/xVccfOMq
E5qEt23NJt6kjGHoHnPYYhIOIrdanQtCrbp1bZqydfv2+4fZfcvMKPJpbFAe3mUgTM3d1KO7JOVB
IbzLvYOV8tmedM3DoEqBnKlJFyt3gIi0e8nbWfQNiJ5fGLJB6QxoIbjiD8nVz6N2yTU7s0bBfwYf
7X7yQTXvqNljtuhAzrAUS7B4PXFi/sFDs/oK3kmFHAaJ0+iWVhk+/N7j5nT1S7iSHM10Php5OaHR
yjn3SvcxyDE9L0y3b5JUgqHyq3rAsUJMQmyY+Qqo+De4X1N+rkyvbLbQcMcHr+ofaaeE7rxiQEl5
jO0+N01WGzLYkS32ZR8gAnIUK2lB2pREt46mZMppTVLNC8fM28ahORx8sAXYeTQEqldxFf0Rn2ZV
+wAq4K2VcR6YTHFU+/BopPA0LUSH9CIrYxEQqsznyRE8Wy/vA8Qvv03gg1MSwJUluLsBybb5PIG8
zJuXpIJR9vC5iEpJBUTfIv3qKTDGQ2TEOHIY/zCuOcYz3iWgLxlwEAKklS0HemzROE1L9vqZDGaG
Rc6n8pTXgaIGpffjUs0r23n31XQ3ZwbIE0zB9PKTKZjCrcorBN04zxTnzP8vxEMQbjs7BL2q1fsd
P12z4QvgzrwNWrV/WeiKiWpRj0nnaLvZJec+Ik5619bUTNxFY4K2fDLAb0KDEK3ybslficnbL2Gr
gs0qNfSz6D9py09mYO0KT/A7t6LSO3/9zWRWI8tiVN5i7ztxJqfU/pYlBC+ifxpc/WUAI2UjZvt9
z/002BMNg1px6HvML5eE6uutwQ+eAl1GS5YMuEs3h/ZJytY2aGX+zcrpMVDmW4yJTQfFQaMZzILE
zP6XAY94QzIe2S4akIE+exsnFHYTakwyd5H5/eGxx3hKbGdyJ9sl8CgIpINU7a8Cfes36C67VXBJ
/05L+itTNTRJZfggeJ8ZFtObZS8A+gLM51cOMlQUkf8K1RRsoSJwxGkybTd3HTgCtmqK3Eo9SdFr
nucK06WIkvos6+0QfL3Oc9rWXrl+fXc6EJ5oRQ9yQF8pwrGhqOCa0w4CuN1RPo8ezWoSo4yGGplW
AZO4bE2bRdhL3njLfq2jIWHboXpLDMjJns2DL235VH1zHbIAs4y0m92HOY/KFsg8+Z3/ZRbW3Jrf
52325sXzIvekDubnw9VepwqXA61ERrNahGc0KcG/KGAwNd4wcVgSAZeZEv3mE+Rt/HDcR/wa+iB0
/IVgBVyXRjoVSTl8Z7WLfmyT+kYu5FzjFDYQKI0eEYid5TV3f0N6KfHsq9UgFF0A6SZ6Lalg+kE+
tHAXQ3g3xUuktA5gE4hzndsU2DCXSQ9J3OqaVZZm1RxstWpjoyd0FnIaVfPfHxpFC0BAgX1wqEkZ
4LNPtWNurrbBXqbR8BCNDvjrfbtAUk7JVWgep52Yyw/rOE9OVLWgos58Rj/WqYWXqBgfu56UE7V9
zunerR18edg0bMmbWxbT30jAQU23LvJf+89OWNNJkAlVmfG28nig6EWxyQnq8kBQYTZdisDNPUoy
Wa0r6u/m3F+GKULBFdLOot2N6YWRPRJhcart11Lfp3jJbAXqIIYcOJmRMJKPmo2b/PoVWSP+7PWJ
8vQ+32L1F4ovRmp84R4ubnZSAK00BTIeq4EeKnNhs5Uz/MsjeUMDu13cetIMqbcu9+9g6ToOct5z
6O9NI0vxX9yT96Y++Dq4UsqCi+MELspYbAhSzyc2evCWlFwbbGu2RyvHGr64rGw1/Q632qOnzNqu
r7KJ6T3g3jFwHfE3tRTGHVZppaBppxwZ2903zUblkAhXbEC8azJse1Boq7HJDI4H9We6drA173a5
PzbAGmJWndj6wy7FlfrK76PmIbh/J+edNYmD5w9HZBga1JYl9ZW8EMdKbEQIsYKewCunRM8V/11A
86jhfkykVuDnds5qItZtpmvOt8KRNpminTO4hWQ+Dscj/FoKzTXy4xrrmAKngpyO6b80cl9SkXG9
to1ryECknE35/HsGCSmb+Ma+/7qCEqX38n51OUe82XHuQbPt+VzR2kU7Ha7GNgVKGMJY2zfYCC+1
eYm/wLJRDvXqPoNsur/OXEbgDuhEV7+keTFRwK0LItYTlxWD9fkVqGldm6G+V9dL/vRJbTcCAncC
CKMPLw/zlu/XH0NMPSOvdKHQQ3gsXoHsG9RVM1dMlOJSw/tF+Z3EyC9wUD6KezqTp+F+VWsIIyCM
tg/uazE/ePU6I6NsE5US3tdyhAeUygedlDaAh3WFtQxoq+8EqUhHKzdbp5rLQX3vVnKWtVGPV/0r
WWMAY5zvpPGqQaDP81RcHGdy23B9gN2WvhZoHH7tMMFq9nZH/BG8n2DIRPzNPwfxwfkDv57n5oAB
7nSkWv0Cfv0DJl0O0tafWgxIseqz1CbLNxxLvxJIhTm3hUcyklcR94pMRRW+5AmzTzPUVcIcjx4q
KZTmP93M71U+CrGw/RX8RbKO81Wfe96MsXfR74UVHhrOCfxvK/VruWGDtJaWxV/J/RO9g75CsAtx
1NMBuIFOaL6FwJ5mlIEj8yfRUAxulmwpOmVXfOlxiqReQg3Md7JdZC4UxPvC+psuQ5UfsoD6vSGe
n4pGdY/9s2nvq6xXLKBgG9Vym1zS9/c645yUpZTcURME1LpkeKRaFPnMA9xSXCNItJctGLhxUqfQ
FEatQr+SdKWe5VxQvpVDGupU6Gti52NkXta9diLZfBV2rApo77id9a7QCqd/XCHjr2rxFnECLtwE
AEO9TY6DSZNVDE3c5Lx83Ppa2jiRM4Ga3HCw3VLTTLme/T/JLat3CO2RNBeNrxbRnk/OBgPKYHjk
tJlSW7l9vVaFSoctr4mv4wktO6qQLs0EFlhGRLhMAX3BJQrk/OPLtvZo/yOuwqfFkQgExFh0ooTn
ozf1mqAR58nqXxeI7yheRWrfEiW1+hB215vbp4h+IYx1uu8xeKHtA66dnpF84/z4TspSz7Nyd5Mc
hJsAzZfWJk+q63fgBNUf865AnXtGyqQrMbDuZWeCiYSOA+6jW8sgSk52hCLPqjhQviLXakXG4BM+
pmRsLUwAT/qN1dK8Oz6h1rn5Rl37K0Q3Qlbu75voPF1T1DC3mvmXo/5+zNwzyMSQ+5wxlWp91RnU
oXlP1NOZ1zjZsA4oTWJZEaz2DORPgUr6AIgMZpO7iwszlYaF+mFHDlys9Higalsxflvp3DkC0yqe
WmYm74bWunNBj5ALdprHyLIRNYPgoZw6ySIVK6VChsMI/aXK5VZu2UpBWaKAO/aIa2MiU98LI5/k
AoHsaAg3ZwKfQ1P6VKJIiftvCznXqUXf6WQGQLrhL86iRF9eUFJVJ2oCfimCbimJaweY00y3Ftul
oGWstOSlly+Bc507QYFcKcsrICGcTHmpgBkxGM5L0D1RLMqX986SihjQrhhY4aCVD6uuUkmz7ItY
6Kbmp5FAZvHvmK5fdODbeEuK13F0br/u97otFAOoXlTmmkadjc70lJ+cEfqJ+CRYyf3BSB2teejr
r8zmCkhfcZKM5ERDhUmjlq0Mml1wyes/6M8ja5SQ71nBlt/mhp6sCriP1367arHoXoZiySZ5D0eR
0bwSc5eQCBaKbwSfDn4+gK77KpokJroJwwdje96p/+Rxv6ZtNiMjS9MGhQhE5FpmWdeNnQkqJNo5
ik9mSgtvZqEtYpPrgpR9RVr0nRiD8X++X0brL/vaXJwe9GpVlN/C2+8YvrWbRs+GQkC6Y2wyVqHl
+lICl2+I6laC+rDRk5S374UAQwkFKCJD9Jt2REsflxzsLH0FYmi+liR5Z6ddtrhqAmT8mMlEYhny
UsdUo9PIFq7xD1YxqBzEY/8yWk9psLhmBkkwpR6lN8A7jiu1+7nFcBiIo1fzf0po57vPMwYGAFax
GPWhkiA5eX/zFmsNRZr18lA1BjmEzYCFODDlN2Y/4sPh7i7tvYmr7Y6sYph3mNwbIUSGrOjLXlxK
2lNslrJ9/3HmLFbktkSR3/Yr8gnwDuCqYhcqG4CEgMjeL9rBfBokdjwE4wKayCUIRmLLqE1JigDf
+iIVBiiSJuapWhtjPHoLwmkUk802+kzn7BM7buQR+oHsTfSrqAbPsugy+KdL++3QDJmIOIeRuBzR
8hnB2Xvta52EDUNnPusfZy0pitiW61ULiY9UeQpsPB8nuD757ACD01QlJM6buZrzwRqpz6bIxo1l
RP5sypkLu7tKIr4x4RsPfuAVxoGpboC9bkGPOddbUl5I187KCk2otvA4EosdttSlrYeOxqcKcTLl
lnlfp3Uxr9h+oM5fxlT0+jGZe3JsWzErCyAmBZ7bg+tOPt+r+eJ5NNtaoDoyb/yFQ1GeUKhXFBfI
FUd+I7z2pl5+7En3DxGdi7iayGMuQd0KQm5TI93GGcLeB/bhQ7/3T1tWC156Y/xLf8uHEiPxypGy
IcZMc7Veg/MFUrm/1Kza7jGIH+lCVamAvQopAiSC+6rWgYTDrKoEcRUV9KMjP883pBUzj2qRcW4Q
NHfSdEFTinaLY8c768fx58sQi7VAhlQqJYKe7U4I6hTVFGpoxoPOyItcSkD8r6Sf0M+Ez4qqESUo
erK/SSMCpuT7xDI0E+ZFAhQYBj2xvfIZqhVS/w6vR20ZpAFuRHdhu4LB3N/NnWyKBlvhp2ARGLxx
oStTeYATaAFTzs5PRSvzV2FB4tG0rn/VFBF2AJ3QD3zTYCBiCxT8onykFWZ7gQAm++Q4HwmT8eC3
UZA6UE3TrBDEyfcePVTY1muM598AVyZw7bUUbmAqoVTQ75pH+MmPYDjGjMh9yoS5KmAqlNf1rzNg
u50jcfRncB5ZaLzKgrLTG/O1nd8jG9Ng6OexFPvlkbZ2JQ0VRDZ72uOQFcePNWcxoRI8lkvY+Cac
bPGqtXpc4s7k+0mSoOdjMLtspXIiqixcFgL98IaRraE2Az8UQLv/NQq4v0924dEesPf8uHYRoVWN
3ZWndkN9HLA0E2XCL/J625+mFUOxVpvty0EEr414yATyvoofiTa8/nT7d39pWaG7vfnRDU+pXAWQ
WuO3at2ZjPe0WRN/hJZfmZXA6omLglHHHIMfC69jSntbB9j8bbdWRZzVGetyxkuPgv+5dpPGAA0v
zQirSZFT5VOa2CLwyRVTz+ew+WVXslaQvGwpuMsSFMnvSJA3q1qA6ZIbZa+cFxXZjqZz3KYsrLcO
Ls5IABXAOcl5l3APrB6AaysF1Up1h6JXPCanKWdE/nHu2z6zZYu2ZpR6TaUJ6KfnOixavGV/QpMO
yUDDBcsWmihNx8vwGFn1rMktdClCsRqhblvVjCdC6v6mZLLf4kWC38SShXHaN3cJC0Amm5pRLzPE
v7KB5hfAHqy0adjD/9lwAoGaz3oyhP3MEaDBZeB7siNeNhuIkk93Lau4q0dBs1drjmkXaRTSxrKb
uhI3iufXHXuE2lltD27e6bMqmDN1B6u9jBLWS4fkHpuV2cTvQARLeV8TMUlrrJJNYVNXkbIgdJGu
8sm5G+6oPjL+jTHgC+D7ggiBKtbX/Ybpaic24w4USUBE2Qj0WMfiwFj/cthvQCnZ9Nvmh43CLd7z
okC0165KhK/zbzh6jETbBIGfxl0JqnTBpLoEUsMExz6tW4bUXqh1JlYy5i69cpkz8hKNN2Ky/Dnl
ycUJTbuPdSrkXKrg1tfTsfUxblLD8hc2Am858RIQhmyVHW4qwN2VDHRe0S4GIs70Ffnhsl74OxY1
ZxNQWV7vn8RSmvMSymN/BFm6WK4KHGlzt61Nvk6DuYiaOmTB5DCOl8c4KQj1LkMqfOCxXzz4cU8g
K5VpS+d35mNHFQP93nOI04cctCt1UYZBnPzU3jpOYC392/6VFTe+HSQsStYA4TJMdf/qIwDA4o/p
oPRI1st6VIxh1VyDe3Kjs0tk4UpMChZsnf2hlRlzkqRsybekDuyUrZ7hyCeY4QiGzaEBtIKnRb3Z
s29wuTEmvSGbCu2fjWSPD4K2BhJGQF6S3xtNIUViOmpZxNgs8swXOo99D4DRlmGnenndCd1ioVWA
EJjUH0XSBD1IFjMGoAwuwrDMyTrFRCQmKwu5jFo4fgYfm/Hjq7/zSzXyf4+RkXcv78N24hJq4GoV
rQDqhHiwq6qWpPFXG1SOJW5W1PDDzDDf9vAKPpuyWwbaYmxD1z4n+aGO7pKuC2Ipqs4TWbvqZ4ri
npNjFKjR0LMeo54n1QvkNhxLG0EXsitAnYOu184KKdBSeXe7JrPntWXVvmKto8VYYJ2QdxcktdvC
umKHlrP3kNr0PeAls+xsSw+vy/+bj4JNySqF4IFqn1DxSVCedQ/16XGEUfRvqAwtbzOeQB/wVKqv
tpy9FwXzVqnlamwhzHxn8v1uC63gT/DH8U0E3kqW6Q4BPoiDXlh64DTwoRiWL6COnkeTV+SmRVTC
qYz0lZ51jOUN7xvG+M5uQAIjFRz8a6boyPZG1Hu4FgTwiPSkZyojXWgusdhjA/Je54987/kZGFOQ
0zyX3LfwK1TLXkdk87AGRgDGJSofew8LERI4K4UmpOeVWq4LsL74fOgiYrLAU+T8DY2XLb5HgFe4
qQeek0JwgWREp7SzuQ0RuUNYCjpT5U04lUkpK3lLqi5QkfjJe+3WPPXYOEU2eRUppH8WQBf14rjZ
b6Z2SbvtPTb7CosOl+B/nkMQXIWjuayXIVaStG80kADNDNh/y0ooXQWNs5A1gLtWYdvG2yNhuTfq
1gtYYSrjVUC4hGG3pQpKcv5sbKKgQtqY6+4CdKTPaNqVbQ9MPjpsPz25gtyV0P9X68+hMwz4JbUH
JT8Xmr6H1mUtafCTOXRGGjYXM5cbmuBvgtYHOzL2KNrhvPtquPL433dWz+KAeCokAl/x2bLeGP+u
/VBa2StDL6YbcF8tBuIcoLf8KZFXg+Yq6jxzAODrFnfuQpLWuWRcRRmcG7Ak4TNLLD6shyFBkl1X
RihJreZCOOAA7k4cLzMqS/PLfyu5Ffu0ezknK6G0tHMvUucAhd2K7yC+IFJw62u9MVXRbcz3k5Ur
MPuvrDtAMsJ6ZC60GJ8TzdljrUZUbBOm1JW9KoIYoj2WQJN9SDg4uRNc8nRsAC7C2+blOFYlNCEC
UeTz7ukx0ddaB2lh06QgUa+C9Q1l+lHOJ2r+cPgRONcoo2nsKEF9M6uFK2w+7WFGcqPcvsRUCwjv
N+U8m/v85SZaFzSYumnWdEuVietj2iI6TaSicVBZKTNYDuSy9heuDyWoL6okTicXErvXq4vgzAYl
ptabIUtWUlw/PWcDOhxGGe2q5fMEmB/Bs2SIoO5zFTB4HXzJu+qHHx35igafagXNTHrDRqHqDthV
RLmPLssrzHK7+19mf8Fh+Fumq0cicnO6B9noqh550w38o1yNaxyJv/D7CphQyX9QXw3yb/LsIF+V
cajn/u/SKfrUn7pwvdwIAQB2kYkxoBfzv4xcrwFGlJ1R2kaW61KxNVlBFJBYZCofqvaFG+JM8LoS
OcB/ep88jIB7HD/v5r4aArAhjZ3RODdZYmzmx4GsGPqPlENrk8k44VG+WFW9XZI8mFjmQpEIWXGT
3mYGvzcFTAkzyFsfRpqMC7fhdDczrbC//L6UogA9JlVS+WWr+3RAHAlcngjUp/eG4HOtfxSXqKWR
CQiRk8IVPZSvVwBNBU6cI1DcBU0vAO0LvZaGISh5jj+Dj1kNuBcnKOA3754U3AFTvjamFOBAsJha
5zxF6JWo8J8HYAthlqYDKCn1wsfsFkcrAq/WoExKOVHfmnQzr3ZSuxgvKe69P/JQvb51QRHumrX7
Y3hLArJ/Mmu/jf6E1HAzvrIraz2Nei+wd0kLtlD6Gp6zyATe9yflUcEfLGPO7g+0Uo/jQS3PagIQ
uo49LxZwO+21C80Bo/I1rKLYsd9z/giaKrCknggQ740XGUrf/vri8QUrHdAq1bGBmOprd+nTjjoe
+fv7yng++nWK8xI+GM2YyrW0vC10K5VFu5C4PY36T9XsXgr1Rek4f1CV2X8pAK0a7hxx/TXxoj5w
W43GquL64C39FEEtkAXQ2DcOK89E7EzMUbiYuBHIaZ5bsJ97C23rr+uASgGw9wo+W5OkVtLbAxsI
3QVGzaJbTONo0DEJzrSfI5OY9xr6bjGo+nhgGvOOYZ82xoMzfGEzlJV24P+PHlg3nwidN6zIPi2+
wb5KAvIP+ojl7JWP72EQblcCZYeAvh8iiqVsMfhObuDg47JNlFV0gS8TCpuEXJXrIPDbbGEVDQ49
YkxMu1jPwi3Y9vBVCahohfks5G3BxELcA21Yn3lclnOhnnCsHG/U7XtyLawdyszv3UiuS6+1WxGp
Fkz71cEalIkvWNBR3pvtdvZxWkzELQwMBA7hfuomgLbfVCgn87cXYCCwc9E2b5OYiU0UtOl3QRcW
L/bdAmt6a51z5D70nYMhwR/VZDqG5p2khzZsN0XgodasgCLgm6IyZlyNRFtNF1ZNlNAGZWhYuI2c
+oSv1MJzcinRA737ikCP5tNG2Xrnh8zcx6/FVuU1uRFFNgtV97vI2Iz4ZH8gzZJ7VNU+PoRUT5Os
IJM7/Go+UCrLDhUXsq2oIiiEXFC1fTXYzoHBFT2MTlckI0kq0ojfWf52r+2NkePSo3YHR8G4DpNk
CP29uSh1zKN+BKSqr2Q77uU2Uxf6Fq0miSfIc4x6OSBhNzetWhX80yVJrsEQevFYhCPcGgIPfbQm
uB+sQ7SBhhek6+DJ/FSkPMx+Gg1ACGHmn9BO4SQyokhhkhzMpY/h4MR5yYpg/iDoTrxFFQQq1Zx8
8WjHr6nOpBMymbhR+qYElmhPlWcH5RkEm1dGnN4vcSKazVkixFHk6J5/p4pWN5OH54PUh9gZb5X9
HO/sl6vHFGw/W/9nEYCxXmWknz999fEGm+XpWK4Zuq7U2h/uuKD0a5WG3zzsZJ1paXct1gGqgfRm
He73kmVIcNGPzphzFev+vjQ8pQyX/04DL3YzEJXobhHrAA02SvCojg6M8YSpO95eTsYbXxfb2KlC
FhsKBYeAR9dwgVxfLAPCdeI6gcKCoOo22NVeifUAp1Fxvgf0kII9a+As9qP6YDqq3LPphwVhbwXI
PRixcJrY1fklH4q9lzhskbmCHuIAzL7mSkZX4SNEWretFtvY0qnTcHCIjqIhf68A0V3ezszIZqAW
EwDFu/4CtxQAOg+VxjU9n1tqoY6C0tYCzpsSTrF3lzDMBpxJan7alrHe2NWEKO7KekkxwD23Vo/q
tS9k8Amq9UMg82aBdaFBJhGlu0MHD37kbkK5nmrIUVetH8xFi5eE/UyeZXNJ7+oSmRekycGZ2bVI
sZQePc/zIM378ev4jqc2M/zLXQlGLw6N3BpXaPxCuxRwOKZKhFAA47VdzoluTo7zcJXyucea05EY
WG4BoLhNXkcyXJzBGHwlEtC/PqW/IjU5wdORwEXdoqZA7ilB2H6ngpMTdzusoFZJx8jfyplAlWjI
/Yw0D2VCI+gpdoQsmsZI0Z1Fe2NQ4/Gk2CTp4rbuZLalVDSwVa1vHShnMoa/epVd7jnU5Nyi5sgm
vqG0o3irt0r5aZv6Iq84dzp2uGvnhEIpkJojLvatLZdI+TwTNn+77TJAu3M1wFfpPgqDSE3/kPYl
8mwFGOS9dD1BM2UU2TSWTwlUj2/XnGa6MS8ACW6rOngh4cTx6lUQUrtDZxYItwVkhAn7XH0obNXq
buj7ciGrgcRlFF760Fe+1LbrK3lxdtwRoJ6KEm+EZGfzmultn6IehV5dKDx1ULnmnXJ/4B92cEfX
PizCfGI6xwxfqqyD0hSwFVitEhmupMUzdFwohvAavrdxEJOgXjKLW+Cc3OLwFBlcWMJF1SxlKQCN
Ya5VEuA11k6duM0WslojjnWp/prDxGw/sPtjKCXSkRxg9vbSqrkiju7asap6j6BhbgJTUFzKmcR5
gESBJRh9X+8KUKCcSICSGIZjgt1lZvOha9F/2KCGyJPH2aj/j1pAxBJzrouc3fTBsEBdPaGGoKSV
vgMTWbRetuRbZT0vdmfYzqOCs4GqJH6wS4okBm7uTp+G5XZGU0ZGNQquKjhMgBts+Ehh8+7EONUC
3W/LHUZHDOKbBe2O+YouAApPNRowSHnJ7qoWw/plpQTrNCi3JzaKv2Gdv6e18iwUxNj4mMc8OqGB
kmYjdEo+5D2ub7MfOQf5aL+kw1L1hlk2vIzlOtXmZCePP7UG8Glh41HejzhQNsh702aO9zTlgno/
gv8kFAhXOAStQmHUFEs/p5yHJGchKJn0F9hnBCjWLlusY6llOq0vsFr76GutnwMxMm4RUeWUDwc6
XwQbw13qVbBfmjcda4DAXPvFrmpiyZajW5Ebb06wDsxt9j3/BaXOQKXX0qX6nrpc/nDBugLqv4BR
1FAPbZLrmafC66jpmx/DXIzQi8yzZPuvDFaPnw/TgS1B2TAJDMHcjvpX1URu80kEh5AD7F/Bh/xJ
rWnXs/hgmv8xA19JfOANCSpVFCTLFK/wZTAQG/wIaeZIrPbixVyPFEQSHOKsTYRQ8KZZENOG8TBY
OohAScLFUuQ8idv6HhFbpmr/oCbSslxntlnEDIkwZVqsddFhk19md1LIAgglQXgqbrXFDBPUzkUk
G8puddHWBLbk0TXPgyyMUzoTrtOFb5/pLyfY7eFQJ9kyaSNxf7U5Lbh43QwLkUUfy92zQLb/fwwy
O9GZMdQ38xdQpXwYt1wsOh7hi7BDM/hDt3DWE8oW1IV++hQi18p7tqAqbaeB4bRdX23RYaUPV1fm
xKbi5Vf19fS9yunn9s7Q8sYPtRYFJfGpocmjwAjBN+JdS6cOBTjs0uENnnVXANqXK//BGBkYWrdO
i7IHm7UuhL4KZ3lPLTSCXFVLOR8PhmAjA78apKuBkNY00FFbD3WXdg9/gKt44bRlr4jXC+n6+E0U
NWaj8r8WBi4/h2O/6qxXNrySkURBVMo/SfaIRfZSjaG+/Pm7ua0xcQ+pWS7djY64I7RmrLgSlEwA
wSKa1jrpaTSm4xyhjtlF3xcDhVHDFeM49USH2HnRMEAuuBjxLz+bRVWz5qvNIpR0NL6BnjspHQiF
je2+Pcb2FvSl+Mnx24qXSrG7TfGdfOWlx2Qb92cAxjiN/h4R6dudRBiP27nOAKZALBqKtTC4SGBq
a9pJCE5Z/h7BehxAcu4Gq+/ltMAyccMZHymNni4kfa0aTHDo6PycmD2pvXlDCc2UxtFKjRoSdQ9P
5AEaq0XOUkwUp6b3RItF/YLB9MEg9ugGEXnuCCUAAT7bOB3K4Xqn6c3gUFsfyX07Ve9VQ1xnTW16
feDceWGcWkxuui0i8DtiuYouflR80r9t52SUxTlPxpgawYoXImI1UWHMy+9n8ebK4+Akc4NLgo4o
Um1uwD3csvEV56iw1FItR4qvZrGds2qrUZNqeF0of2fAVeQMGLn4JoR41HznFnLjXXC7C8wp/v/T
a71cjGCQfdyRM8+abk4YBvxXB0Se+HNNYAeigqkqmHFdpElqChABcVnmOXc/D3L2br/aFbS8b65O
1CiwFzUC2ABQMc7cDDsJz3wu19qDO25PUn57EPv5+7M9/XSVbe4V0CnaFVPpRcpZ+bNeSDrtZGp6
nbW6TaJBWRbAy9s6Cbe9kqlUSSu6coPH9L+VzNdvS1X5tHUvLl68Zr6iQ5WMbqgSODTbH+aeEdcW
NPuL5GL/UvdlZO5n+E+m4qVsDjj/TqZOhAzoNFje7j9fi4MxjjCv0JeEA4esg6Klehwlm3YgwyXq
DEx0kx4S9jc491avDFFTqK7BUAXizTJRgyazY98FydHXSv/BgHh+dafL+me22JRmoOIcz4uJC2Bv
6p88qCyICMsR9j4NqK3jks/PPTH4czeYSipOhSONsJAPRX1hgH9PZ1vsk1ioEcUfj3SWwa95K3GP
fvMtJcoqr84Ue6aCRm6vGx9/QiOGyWR+1L6ubNjYy6qKOiwP5ZaJn3uQXVxBrGVVGBjW0cHfQ1IR
qiC6pHn0hGMMgBVJU6u+1fZg5mBAQS2lt+pkirG3QWGThfJlrMITs9odMsnS41ws1pSFa16t0KKw
J3s+vVn53qZdG2vbK9PUowftCoLcchjcHqxHro9pV2/PeRWNjZj/Q0UIqeeuMei4efQ2t6tpekOZ
+DKESDTs5wPatObdz2RIHelicba8pSjH4dHz22C5bWf4aow4gx3AWvD53VNMJ4ODOaUT08mMe7Nd
ZmHXBHKOFVmjXbbX5BHJGll57KOhtSdKedQpq/g9djcvW5u4oi/ePg3yrw0mSeaGcql46QzwMVpC
s546TbBzXsBhftJ3uQH3oNu0QalQyiFqSLnV63XVJAyJnTRvhKRfXyQBkvjisGhNwg+yf6rmxYVa
iLEQ71g0ojaLgVUW8T/jOQRysOqvYpIisi3EJx5nkBAiJB55/fiA98mbL6b9rj3SNchYoHF31w7w
nvRlCMBzBFgwIOZIwBAbFMyhGfJxu/g7usx8jGh5il8sckE+7wI9q9yH6KS4XNgj5PqQ38L9A5K7
qAyfdCt/b+Tof8GnJrujZ8OeJrxn5TWOEvynxA6hWW7ZLp8UR+kHGrdWDus8dKSigTXZqvDnJXA+
LfAv6OeqpHnIx0eevLtPnUF4fuZ1LSXVkF8Fty+Avekft2devJ/f6p849kfKKOOBfgoCFYXl/WyX
b7HU3iCG6h2f8KJPNKom3smKSUBPNoOj5XjMB11fONIEXeSw+0E5/uOIL9iPPqEcTjtIV2JpzrN3
yEs1d1AtlQgsIToWS1E2ecHHiWGM/UAHqsMQu3W+fp/Ig22iLDwIbAPboqL7nDySzik0dFSk5jn4
YrMPhbPDm6UGuL1Fiwj4W4UM3nx06nHdc0oR1+JE14yEbYo0w+1O3X+ygZ5TBGXEuhTuUbNMylCn
SmNUcxEXxtUIOs4pazXV4yfWnDcK/b4/Zft+6lA1229tGFqibpWVFNkdP/AWnNk3w0eXsBSVMoiW
cWWg1E0a8pe3w3OCGKWyYGf7pgToEIezRD9+0jxTjlO55/jtvuLREXMdl2yKwFn35yE8k1j4EFpc
IBaVb/1qfCypbDCIJye20+FLDVMUeI+ml8SJWqgLjxT9eb1bFYvZQLDDc9UOyOCHJlZtOOwVRB+Z
mEI6987VuhyaODa/P2YR5VPDkAknpYAh0PypeTZY+T9oxZaMrUU5TmEguOUCZxKP/xp9NnNGDhR0
Fapaw9JI4OOUJtJLJzxiSs8FaZd7axvDGGGxjephmHshIr2rIZ/YNoEaHObOkxDX3KzZtzZnjN6o
xo4H0ZKvfPvoFcW4zp717cpTbzZQvcKOGMTtUIUc5J3b5vF6+sL1AJ0CxRbs+rFp6Ck5JIZ2rVIK
zt+JCZ/KXAvoRJyGzpyKCk/zzHcEThCSXwZCnIc42UKsQ7wUGUnUTWk8ux4ePqbflVLI0d9Ghsh7
Esg2nekLPbWOqFsb9N4fRTJhN52o1WocDhddjUrhbLbY7OpLypYGcpUm7/7aFVm1G6z/T/JEMgwi
V0NN1DxPe7YJvD6qgsyxsuGOzbYAlZGfoA1vPItBQyNVC+nezMRr458vYbWV78m6btOfHnAe4RGO
qi9I9R4fO8ZFPa/akUF3vYPVpLVjIMdlrU74OofjGqQzmwTQuaSor+oWggXWZNZlSNquLCvBndPx
8Ui8TLd6+YtyBEQ1yrgQgjFUtGgyPFV9HMrylJc0lg/LXz6Qdlc/3zTDvk3dZXg4UYXwCvfh9oNk
xsNi5pJi9JJBpF4uUscdPTay9h0XKx/mLBht7zm4X5I/tXuTCENrYT2VYyL+eB9e/mlbLnuuKI52
Dh94rd5noD3pIoqa/5OQYAva8zRQbqTHTGadu9YJSScQWND92pDjYnI9sZnS1XxTZYfog0X8lXzT
WI0Q8r5+P2R0Lgq7oThAD+tX1eTN9NiNkqoGKNt5l/u7GjivsEiZpoOm3BbYTjxLTAbYzYBwAYnd
8SW2eEviA0CiFU2xG9wjU9Kqbp7l8z0nGE36WehiAWiCmX5q7y/AIQOf0t+xu+vHNbisMiItHf9V
fsl+ChbY/Cy0/ydvUZzQoFZiVMY8C1/32dNwUsxtdotKWTGOMeOCG6yGnkrxbsYWAjgjVeaALWpJ
K36FFtECVZsVwuNEqV2NpjjYU4HDaWC9iJGyHR8NnFaeQ1RuOBusWcBVVEwpMFTQdnAucQcFz4ZD
q4WOYuibu9gVTP2oTBexMbyEIG9eFiRflKxA1IIK9BjSTI8OFu7FpyDtuELbg5QxbOIHMG5oYBFt
+hUp28THEZ0qCxOzzY9d7a17VdDRlNszQvqoxgU8F2au7HlTlYBMD5a/NJqEP4YBwP3EN7Q+kCq+
1EOmY1uTD49ybB5KXXz5dU+O/UN766QJAmHyR6JO5ruo8R8RvBEy6dHdel1PYMozYPAxAudwLZa3
Kc5k1MuHZ1ZrshK7+Z5IVWEH4pZWkQW0Up0spcZKbx9D1z5XlNAx/GsSe8rlgXeAYU27YlwhjuK1
GZLQDw3Tr8YnBmIwy3dzkBZe9cQpe4WLBPO12OGVDge6FKdju2Wb0eRRwlmLUpP0R5uj0cCdLvaJ
MA2wP4dK3ByIjeruQNVGCnB6LRaSnkJqjNPvdtoXphtqOARJTlAfmvhs22a7w2H33CskM1BhxcC+
qyr0ebknbaG63nj+tLGI+B40tsA7ulJSWNZ7bWIM7VvUG5v6y/JTzw0lcrqFJwsYuPHA6BI2h+6Y
uGXQfWklKlgEJ9wpRXFmKZAFvIxs10au18Bbtv02t7Jl3ilWPQlLWuOUWo4quOhDacgY8FIadneM
VN0jXqc9VE90I22/6EbKP1VTQgtF8Bol0tQJra88iq5W1l7Cuz9K/fkiJWzwFMoLbtidjX3MlK22
TOk7mVEBAwIaBPa6IP/FGghgprXxtVf/yuPik91vPDTgKc97j4HZfN7yKIpPGqqL/znx6kHPAOKu
rvF1w5Gh9s6Yi3osSAuhBJr2ALiU7vpjC6prxxCErtFpAyrzOgQwW48vvnqkQyrY4FfEr7X/awsG
K106PhS51jwqghck2pYlW8V3a9N0L7KqhRfJ/uwHKyDpJ3srpXmb26Zwj+sKVnd18DF2Q3dFotq+
4a633J6LHNunJFJXn4WDcmrWwjuY8usIcMMDFCqIdb98EEdjiXhh6az7kJ4CrQZtbFXtyoNdao8O
NUVp+voSSRin0QKtXLRxzYoaU627VGzWaDQ+jUo7hdJUYK0714trvHDT8f4G0U+v9kSojw4Vv1vz
8xZlpOZZF3RfXcxGYDcvNwguVdK5RazPfs+1DHd8qi9bV3W1e5CrSwFYZiNecA1SfDfbdfwb2kJf
dXESivP55j1/npuPC3Vh7E5y9kKfWYYnF3k7ZaEIxGAjc7BaSYsL8oooAtJC9mI1FNAavyp6ZO7m
6WdCWGjf7s0l1OLJz/8xNg42NGfl2qs2qeJB4atOlcDaPTbuY3L51AI3Ion0evkY1jsiAYxfbTIu
UxubqYsgveeFl7N99ja1wrnJxTQ3PmRmRY5nRENznwOc/0Um4OhYEIjkM5BUKygFLuNiE9sm4ZnE
NpxSBQGLRcg4MDJzYyZ4Um7VtIotGBxNF3ox25A703CflHI7aRir/YXIy0cTcBtFFRmMdsteWalC
gg3Z9BEpgNpzAWdyD//gY9d2rs/A6AOLWbx6X8vCRQRC1x0BCey2e9kUL1VwqAsZYSCBjvkSvalV
/ZgOASamhRoywiv9m+BQNLMdrq4RfoBcObRv+vFexMG3K3E9sAW3V/2IBCuE80q+dxwvLafxv22o
Enr2Cg+hJeRigv0Rjt0mJQYJAgZjv8wV5KG2rVXG/CZUf6zMU5iHOCru1zazYyUXQXYnvi9sRj1d
0AcW2H6P2F8lIOdXkbB9DmvWmOW+FqrDKpTNQLqI0HqjjP8z5lCNqCGGmtbPyhnbRMAvzuY65zCa
yMikQq5yBmddpkN5sMeI1OnU/fmCtQXNRlGvWX/xPA4SNYBVTJikUhyl2AeThPkHBO8KiIL9T2PJ
GXEkUIkvmAP/pG3zF7vEGVfaVZiuYNX2fhjJuL4AS9BliyPqjrIy++oXTMHko6bh8/Ei8jmOozhr
Fw/ufPKfb3YJtkjlLZtCv80xxFYYHGB656CXOVJPGNiJKZzmI9S/SkVU7y+P8M/qF5PRKlaVsyIg
jhm91qVWxGupeQfBoBPVYIj1XXzdtVz+FUm2+Ku+3tCA9Mc19XX3O4yr7mWqhs4MB/u0aQcaw3Be
T6t5WkQ6imsmcRNo6DbAuvsFKP7IpHOI/x2ccEl2uBjiGNh2eVy1134cam2Pb8T0QVrwXuU49f1j
ReEWs4vb/5kB/N1s7FOT7RJlLbQ6+2iPTANzOi0+hjRu0ua5hlxRqJ93LW4YM73Wpp0NmFdTIsJ0
yalXNzqSYuG5tbfU8cCV44BnvZ+KMBIfBW9okKCPf/0aB2l1hjR9gakmJJgla8YesU4H9+EHoRLf
Kh1Tcf7tdZRQvKhqP7Nlb9OY4rS8XGFv5f09hAIrIP+h5RFU1z4uDvRxy1+sKuTl2ju6EZjVL2hX
yTkDXQM1N/VUmPNcipFc3DT1rdPNNycJqB+Q995nUq8pP9CvWdYPu60vKPtxPwSV2Bbn9uc692Oz
m1zQm7umO/4SigQs1eRj8OynOn3rXWWGcPmCllf0xO765GT8iRIwERnSVMCIzmzTb5UxYwv3q4yx
31ifGVwZbtDaCa3GB0LaXmk68d4lq/EYNePwB09gWr3eDcRvPwIgr0xAbMiD890wmC376ck4OhtH
i/wUTsQ0RxUWvoEF+gnB/nhp6/YG4VORToP9+L+RSm7ftvD5dfgEf7Dcl+kIDUTB8RZB0LmLiXhu
NXIf3QWzvhhZkWo1KDj8xEzZ8XTMzQ5axAybxt2Hcke6lG/5S+VQsygBSanp2P7yi3R0trch9QH6
kqlWe++qrBmayHWkRG6b2SP2OUM1Jw5ZP/VmUBf88UjbQMR0jShAP+oVQkSv+Z1iqx5dtRtAxjol
mvpBG6I5qI19kDKnGJpV5t3x75+EKl3jxpkdB84d1gumyVz2ycIoY7QEfnfc8Si7SDq9kMohay4Z
hTC1mn1mXgklLoMg47ue2JLqlAuNvZeg4sXDSjEsDtglV3Jvs/L+QRmwqmW2vxGiSP0ZsMH7omwL
Wodeggk2l2A/IN4nuhNjuTfwRz+LyMvY+WWfn3ssA2yT/3ATD4WPFKRaxAcNoB5JWQd0bgfNGZVo
Ldd6e13w8poHTXBi+aRK/kydEB4nmlJwUE1Nuk+rWt2yDcFvN1x6kd1hwQBqw1L62XaPi+gb6xo6
D+kaEpl/ixYRoNuUSgyMBTr+LWMJP9acAKD69YRirbIh+oW/O5e9V2mIlKXjK3dUvsLhGszA8295
EhRFuT7WO6c13MEUB7x9uMfURGe71bDu3UYCZbmwD0WM4QP+Op8+daTu16F2AJ2t7Q6/cHdi/Etj
EBUd8/UlmfwdJp93JE9muZSPkJkx6mXpiX1VG+WlTzE3B9hj3yLbIAE7qnlqKaV7M2K0E2cMGCQY
vcxhcPihRWVTwEZlSR7FFBKfHHxWhO0OwWiXyyLbF4+WrkK53PCgoQ1yUl86tLoKETnRvquZB0a6
A1G8mIYSpCqip5GZnixn5ganeCzlyWjNQjZAGTJ0X3YTMsn7TTzM6UC7mipjdPRx2HSDgET3VAn4
rT/wEtZQVFw26FfB5eHhV9YGC8m4VzIo1S4HOBKpenIBC2vuDm/S4Us5RcSDhTsUY3ttGSQi7rC+
qy7WlW/OLh3/UBdW4DJl3jakz9HvHHLp7ATNltWUvuy+mLW8AFWa3CuyKu2y8A7robjURK+b+4mA
35sq8TjVJq2Tes65sdgvG5mky3LIpKZZwqXjj3QnsvbBa+5tZZTgQryAZfMJcSIu9f7RveFqmw7H
nQfvwHa3I8Hff6ZktPwcxVNCSwfuysGyALV9+0ViUjLj61X48JKJ2vKH65yzEhYGguGz6v8v7i1s
di5+GMdq2q1OPekhRtlooFEkxXoG+rI0cRiMVpZKo68TRuMSsFYrNEKeUPr+IijSnjTqhxxRRGDn
3R5UByRBQnrurMPYwbn45lyns7FcvdP/8XxUqYeDD8vo49kCDE2a6PFo+WAfLjaRfP2b8/s153dM
Q3kUOpvKS4BYtoSQnGbLUv1yPkVQDJr8dO4SPc3O7CwH1vhYYMcxnTsqdwso6WkUOscJx5rhQwQz
2draB7OrxYlr5O2wfh06rsG+9+aUv3Kz5G0GZgCD/VoOoHUFO2ct+nIMZJDO5/KlOXR6t1DF80Lb
VxQeoGci1oygtmB1/PslIPkx47BYiDM22KpryAWo+sU3KN8slwAkc7qNZRVuJ+XMDtChWxJ6NLeJ
mh0+Fg4HeCsSPrdq//pBWK+H8vRbTankSy4b+n+V4ogfdFqjyAnPd834tAGu2+1oDX9/cUgctf+G
ebponY9oBcphrhHNxXNgsXeBBQvWIFp1QZU7B/80HOMC2zWKe21Z8fYomVs83h6nq1s4rWIuczIP
w7Jt63GbpdIJgAN3nzZf7l9rbqwc5L9h3IIJCT+D7yovy/vDdJiLKFhuk/tXkuN1boLUVzEaayax
muocGswPPp6IoXjXLEeH99wglcRRnnfCoKy2cUdsuQIZeJUAFZ0RCk6tfiPvxnUHWNLM+dB5eZd9
5Ec3q/0KaR1sl+Lpz6EF0AoVYbnvZ0cyIC9c/JApGa/EKI5J3jdpDQT2ja1Q3yyMFz5VCuAFUAyH
P+ZaSRoHK4RUhRwPQOga6rM9PTy1XUdyQANrqXg853zkQE5u0JeH67Jg7DcxrryZDnz0oFnVdDbq
ynAXsBPP4N7s87Fs/mo1kSJIjtxu9oSGTf9rpvOaFTfTybe6AsmFtiGerkc6iTFBnSL9+SPKJsmw
Dm8f2Th+gGubzi3a1I9uSMOZtijZr7ulzjcFZE8G++Q0LwonmDUkF2cD1LFWZcFReWt5MmFXUT9t
eET3wWYNfn0QfAIkH2PYD4nJzwnvW0MqPwU3/rAOv/3Bdg+ZlnoL2bkmmidYHmcL4TR2nkPqA1nM
rUVQCXVhFEY7smHcDcKR4oE4Y/Kj6n9LBZUkO3tIzwzkKkpl/83UmXqvUYZii6Y/jhNeTbIUMCAt
P4aK/RTbJT2KnJaUOSqENvdU23Ls3k3HJjE4e51a3Dw+IA5epwXfQcl0zlA1eDC+vApPrrtv8Tyt
CI6hTR82r85+zLsrV0blKEsD2M2tje2SqjkkUktWnKqDO8TufTcWHxL037cuwwnvcfJnmjb92gLm
d++ibg6UR7oFujgdZLlxOsMeEBDQLkLL1f9O3+wWTa3i/QRGDg4Vs3AzPdbMP2BZdNV1magmM3Bh
AUpFV5dYcW9twpa4aT0yAmkVmc538lwBY8hY2Tj/M8cM9aCjbRpaCUN9cFxJWmDSDRXJUBpsN2ry
M8q+Y/e9xSwk5Q/OLDCCDIjZnXg6+Pq/dsU2C2FiwcXRx/cx8f3c/JoqPyFmoWukEdw/GB6tfxoq
AMJF7CwT8krVlYiECwR15L4tT7pLyyDdyHtHe/BlMWHn3SeDg27qe2PGy6oMus3IFr4HguXG/pox
DcxYNDtNxYDwziUngVDIQB/MgDDdafKIQDXMn1AUV0z9HVuvn3ElGk3bBTbmheEk3cZUf6LVLnNn
RL++1cd5fmxCWnWR+LY6zu+QhihNnTvKzA0flmR8sUipg1MZwiIbCKub3dbAQEiqsWQwZBYO4hR8
MdVxkJOv9w+G70NVTnpjQOjkOF8Bx8uONZXxm9wq7wc0S6/i36pMTYnT65jR6dIhzVr1xx8Mokc1
3xe1hcrTMd24y3bLQ2Xahwt1zRbzNGyYILiY3vZ4XD+k+T2BG1UBQMKZDDsHbNEHdA5G7uh96Aww
DQE7VKWI1q5NTbvi3k3+WedqbUPs1yo3NHE6gDfN/J53flZfmti5JSRFfo7aWAQZNWC5nIgNc4Ob
g6EBCB/wOzZqxvozADHHtCLB52u3cDCOjMzYKCjo3S18dl/gYzogjaO1/OAlZ1xe1LZu1VRGrPmN
otNJoraFrB16O3JguiEdCM3egs97uKG87SQ4SMiz0W3zxrHi+6+JRN+jqA7S/A6k568pLN2gZ+qn
tGdpOibot3xONVOHXhWIp/b/ZhgKr+qpJLPryvaRFsjYoamdEjP9Zr5OpLpUWDm9GrVpc1R19Vp7
1cwwBaSv/vFAZ0l6PqhpZFAJl7RtLZu9x/HmA5Gemgy2h5jpRlswrDku0ch20Iy4t9ka8laklsPc
8+aw06Oq93S4vwzmhF93pjWnfqFfppESX5HAcHP8HFcTmy1MSrNCSDPn4V1D1y3G/EbBwSTbUDev
n1amntcUT3jUi8qixp8t4A6MIjk9h4WaBaELswENTKFFMV0S0CWSN85B4fRr9mlsB1LWVMt62a97
USgUEln592ewygTWPeFHAHqTNMZDtD0LaW+jgKfCmjT/vE9GI10frPSkjVNblADE8bgTovcf1lFd
fqNyelhYL5AtQfEQ3UBYSIdq92UXfAXPGsOgnqEljsoJcy1lYRJKWh56/Ik1IXbfrlJpZGQ7OapX
l2FkuV/qFUs6N+fGpBh5pKpA+b88Pie0KHIvGgAUeITjepr06xY6yzzBx4zCsf/6v6QGmphIzjUC
P9MVipwW1dNoWaeSK2fBtfY1v+9/owG2K9JFbum6/9QE0ztQkU00PFnUVPC6oKQMwSYV3CR8hzSQ
xVU64WRGPO0U/Dwkc72kdX9u5/CkWyEKcWY57/f4tbT147dVwVDCM4ZxuZncbwepfm7rbSKlwEwm
PbF8czSdp9dfB7q+gsyuLkUjGKhbXu/F6Qfx9pIonMkYpxzyYaj0oiGAcAcpqBZUCJMSaq1FY5rg
6etYBk5uDqWYeq3fr0GTdClBLOAqKz2l6rHsUtxipbrjNWYxMv4d079y8nyd1QWRBXJgpzqPPhkq
CrbB9nda9L2XbK0mnwPgmRPCWUnWafP9m/+s2i46AtQN+7NcMtvulJEITTBv+WtdD91GwArTh3o7
KIMNj+yA7zGU5M7n14c5YVFzcnqKwOwHSU+2Ywb1T2x5W6yhTkI14PU1d9hVRaDsnqYPkVeTviNL
C4W5CcFE6b6v2fkpNLDUmu4zAwVVfdEVNHALqPO6XxFwmVb7g2QhewzFBqM1c6gm0s6gEzQDsXAQ
QE4vWmiv2dNrDG7+JeY9/JXy0Km85us3GCpwLFsvLF/QhdtpxGPgAZLeII3NfZ4MYNrLcrcKTEK8
0s7onYIYW8+Jk3lq9OBUzLIS5wl6CgkyFV6a13T0QeYuM5bhM7+lz1o/rMoax9Bmy4+/SwTiD7Zw
YjSQkDYkGoNs6D8dOvvIoU8vvYd8o1mc6+BhWzSFbz0xp0ilKspTbYqmLYlrIgFjShhSeRlXwIrE
940KO0HCihTShHVcqpyFuh7iCvWe5wNP36PtcikdCc82+3P6MfJvvntAw0S3tg5+gf5U9hkmG3Go
vaiKXxA0R/xIxWIcX89X1Qgp9PrMnoIpaMc14vz7EvK9LpOI02wgPvHs0mMmIoOAE5Et3JiRozUO
Dv+qII0xg1Ug0XA93DPr5PYxxI0DHEUgK3t08z9ivkc53BdFtZO1zwwaQ6pOgU5iSXwKALCRSYgr
wWdX48kYLuYCIP2+7wqIVG9ajaFw77hC516oTVDDaUAnyqZzKsJ5/vNCkFtKQj2liSpfQHo1BOe2
f/i1jYBCrl9HuHgGhgOoZuFdBQ4Na+8xq8JJNZBD7QD4H3s/h9Xjwm6qGLvGcazmIok0PoQrs8nV
pn3lKeKriEot0bfQvgnjjQ59HsgmerXGJGWwv0jRvS1lcpsLn++ArxQJNYwC8qJW380fOew19N+u
OCERGpmLOBZGYb6WuP0m15IxDuuDc0WjWc8ebQP2RMvHIHJNl8KfOyc9XUeabMutFS4ZelSTzSrP
4+imVeMvvnWlbyWf9KHLqcfckCGi1BYtaA2xHVt2P6phH7PsLW9KXs9iJvred+0pv/MfLVDkqa/A
AE9WhuDbOZrVjXkd8vctdc/x6n2eXk6aolsOWRLOQ6isw3uuRicgmgTHegYwKwmLQHbr7It+Y2fu
IenyM5FMDkNBgN2/NsDD8QJEiATiM4l0WHpP+V6EDkdppNQ4N+NuBrB/1mDRgbvUbGrwGxnV0bn2
HKvrIb2I6UXy2hMxpUznrszF86B3zLPQWJxgZqOv88H9vh511n4saRSbR6MOn00kgs+uX4pquoUr
jgxUalavm6FP3oRbd1vz1fklPJuqfEHRwy8ndTmIyrrKRJ98fJ+8s63f9vZ/xzVGuhTqlmaCYMGK
Ti/Ivjsg5WLvXGekzCvyeJKm0eaoKO/9nrD2G2orYhCsq+m/1A62DVStM1xBWh7RAXa2px6PwAGQ
3qDLOTmWZMfiaFx1hyyp6DwT8krHNUG97P0+qJKcOweSe7F+AN4h9rAeEfN/r290JtWlTi8PR6JB
gpCZE0xcX5j4jGiMWHn9ZR/NfH95BQGB1F+RL6FnGFPSssxuBNPYlzFxkkXNNBWfMEwuCBtMKzb5
6vdqVfZO7LvBhpWG658cSNmzlxxnzI/id1f++XSwMnY5G3xpUGHm7w7qNcxTqAbxqWDzwDR1QNIJ
zECiGRKNnHDStQwTWMkkxYBX1GiRIhMTvNQM0pb2ot6OlzvZ4UaHghksxEzlZDkWOMHD9GiZwtjh
amPt2HYxkICoxZdDZishIKinckBcYsBHOa4//3XI2LljuPEcDDUOn33b7MWAgYrl2EIkv8ECWMl+
W2q+TxHACYR42vi8d04ZMJrTiPp2yP1k/lFk+mVum/q+k3CTaThGX5YuZ4XG+BoB80Hlvep1GVMe
gcl4/FKGi8Fc6Da81EMECdLDyKJvfUUwzuehqFwUUPwgR69TsKxvryhcnRBjzoezDiZjLLhis3FT
ygUER18t2MPV+FxrwoIKfGWl2lDonuH8BUOj/NN+vN48MM+bIDbTHPI464D3lGq76zRgGT1skHJY
xDgaAnIWCyXQ9c1Ygm+Gu5ayDlzQ+eYglyTLI6jPrDA1NE3VAEPnsBd73skwHNnVbe4RgvqrXAGa
WDWH1xnYRBYGCfUqiFFW9aju0+JOSFX6sob0iKZlYiiyvfu01Ouyo0f96L2y2lARLGWUTPQqH/OS
J3fSNI4pTSF2H9GB1zO5kHvG99tyP5BdRqVCAjMafLeXEPSNpFTOabItvQHTXCbP9Cq4Q9vgS7Y/
+O2yP2mjOkNEkVH5SoeMu2JJOiAyV4DfwVW51bHt5wfrMXGskIk//gDFAw3kVD3fLGT0LUXU84E+
nTvni29InRkm6/xIYm+0WwlJPcKU5w+FNgMRhI5FbMmHRMYxbr+jca6Gn+tDgJUryyVKd2QoKOn7
7V2MWhrtdzgl7IFdCRUw8Lakjjv52UqtDl1jX007XWAHK/1TMgyroMcNMdgiLbMz0gom48TVnyCi
Y8tXh428Q2oqshjwflxSdfWnAe/zFcd6xWJPiHMCnYCrVv/V247f9uokB3EZ2LsVKZSOxVTRl75l
lHzctZTsLgu/JtGYg8pLtYH0LXPJsXEAQfcWC2HT2oqN/QMpztWAP4ct2LNDzA7gEP74bEpqjIUP
SWKMThNDSKDiU+0q88QFC1d9hFmmpfzJQSUCmN6vEB/hfmdS8+O2OxXbRJnj5wjTgEeY4f/9aeqD
GKvQOeLuBx4H4naWlNSIp8GzLceN2FBQE3SNxVP5AJ201y9KeEy7bXYEvSvcY/7zMu/RC7ZfMPtZ
LK7GS1XAP0YFZn7Hy/DZE0JeVFhi/eS95RnRMcc1jLj24JJNj5D3BTP7OMyLUqLFoXgjbQnyFd7A
J7zjv8jygZUOCnaMUBv3X/oMrku10TlNhJ7o0GnuZ+rGuslWrBUJonn4vnPHiRxHesIyDC8sli08
aY9xgMla2hgv6vbZlwXoYUt2ioXyLoCCc5OjHSP8bzbn+0iEHN7ca93l2NOv90LPCDZooZO4hgon
P/JQUgaS/m2t8ugHWyd78XlaSTtxIQgWlQhJr7IMXj1UDvGN0ZRug6ftX6CBrlsaiIAOiN9v6LGc
deArBeCRbEkfWQJDQXe4D4FPAAAOx229w6RBqCgK4EYQU3Uj/FQdBRMqZ7lLTMPmVVC6ZsOSABVQ
i6mkAGnr/EY8HGOfwWM+eTmeNtrORopIBY939Ei2YkYTp7FfR59y5IKOSzMHVHETIzHu462ogw6P
e4zedSKNlzdFRit7ZxFas0Wgt2QZwDvdWiiHgJNVjM6MWLTINCtQw22vKxRFsmx1b+ZhTDgpixbf
akAPiD+L1Upmubb55z3fwRpRvMiA+/JmrpBcL/qax9Vcw9qeid6olb35fW3Gn6zKVhDHLvvJjvHj
8QZfpUBNiXvQwxhXilXnTFpNPzfy0gnVSKtkyMKv3/L+Dxs5vHY8Rgm4pyPGmFKf0APWVl/GG0t9
3rTmctOSazw68kHMAQZWIE3Cr1HiEN8Y1yFmFJGW+oH6ptFM0eImKJTyPJ1UpNDM4PXU0Jo2CpI+
rRjtTlrbVXD3De3nRttOmp1vEdO6i42nnVw5FCAsc8SIzgjVj1erHUqT5ds4ALBY1oVPFoPfi6AK
zgFQgi1kArsLp/HW6qzMKbzcbl2WU1exqKgrimS/t7lMhtAM5+GxZhGi0p+8CyeEtE3u/bMCVzrZ
QoU5wwqbPYylHVg+5Lctah4ED5Z1vZE253t9wWa6IOYYuBMT75O0D/MscsYb7Be/duXyvfBs/EMD
gqsSkLzxbOQO3hqvPMUl61GJuRw+CxpYo4rllxQxFsfKeYan3u1Ff/F6GVUbAkvFv9R60t/Yq4tG
vvipTbKVznnivqRkno655qliW4sFKhshMoo050ieR11M5RZum+PHmvCJNGhMN0YFdb/6ounD8Hru
NYcSvjvjgbnmKj8t00UtWa1Xx5S/DBAX8Cip/xo0FcirHi9QTey0Utz2WVOwzwlW97nC6tVyInqX
qPVaiskgSUtCeGoaJ+YWSNkkJ6mO3WG2vkk7pdD14vAMSesKQ8dk165ZhZLHcbhz/uuz7WyG7J21
8dLCsMrlUAJHgkfao72dB3YKemZnycrOqfYnvSMAF4yjNwuCKuJtggntrjDj5UhZP16BKzU3trdA
WgqRQYdHb07civNqVwvsUNM+VmoIEl5whv9fAU2n8q3lgBYGRNDcyORkqCXeEsPdrH2APPEedI30
aaf+dvipOQhTXS3E8SBJE1AQjz6e8kLfz9+2ugSqTWV5UR/NpXQOrmvmqHBnlQF1MxYISRkOlR/0
0FeyhJQjQN8AFPJShzrhwpyDa/NG+Pm2srLrxXLxaqlJl2zNQ45FZYqYkey4qbXqLtoprv1zJN2b
szM0igtZiuYX4IcNxZTSeGO62N/9lafTcIg8u0npzhysrKWMqA3ZO+R8PVouZhDB0TPP74wvXjZ+
J/SnoP0JGemhTN3g4aL8fFZMwKUbrkE71a1elHcgjfW4fcPZ1AZewpNX8as5eWQ7iCcmnkxlvNH3
dSt5P7jnlUrv/Ec9nvHMcB2ikCwlAcQEkUxmNkYx8d2O77QmcrCBj9mlxSBXZrKZiCyKYEimBHvD
htIrQUpFWhR/cEAX8AkdpRNxBRdVHmH+fCHGsbC5tMi5wvz4FLAMcn95EItjMAzQylOwaI4L4q+x
pxNorT8loDDZdhsJFwp7yobFtj2UpljkhBag1msZtYjuaP8gWTjO77fQlc0mQVSWn/2P9HJjODUA
spqB2ZOwp4qOD7vW5FB4lJG+SI9mpzP+8UraB/BKgD3bryhLwHxIBt58JYiTCO1ku9T4ybTa7RA+
2TEQegn9j6zs0+OpHopWozdDzRvyAPRUleT0DoOTkvGyYMLPwf6LXWZ6MVIpLB1M6P0PjaSKarPt
KRRF7o6USLug8S70NRHi5hck4Qr/6OH+ebAFv1lml6Xum99vksSjjLkIn9Kv7ho28zsCOTbb55nY
pk7rjvgGgUU0scT0plTBi1RkYw8V8zNVflgYAbspSSuJtmE/M/24jpOGI+oEJlI9MwNYoRiwkGce
V7kxhYR8nyyTtTVACJtIkhBWscwhHUPUE0BCznrCSgcJU+iBP7bAkrrICMa4f5XMX/Rk4RJJqBJe
BacKBLPxw7gquqwpquCAkNSMLpsT/mMjAvrkI6QL5JnYtkW/5/Bh1pVNA3tTH0Jfshu90DEsqwTB
Lum5RVHw6fAhQZB/olPQGbKHEb0K18NZOvjmN4QbfwIrBuGXhDs2ex6+DK9tQ6uAC8XNmPfQGbdt
y8GaBpmfnaMmLK4YNC2lGzhIy/eoAVxpwbeHjY7gTRVSqWt4zeHR1HU8S9eH5GG/HHJkEZskQHSn
mzQv8/vHCXV1wvqGkna4fdFDBv7TkFXTM/B3XPJ+n1lojRizL3jdVT9FI+ZvvLLtfl4drJyMg+Q0
fIDiCwaj5I1JCBDCiC7mOjmYiKuZ99vlRAy7czKQgkhEAAZUmEJywab2TZ5ZO0KKn9BjCk64PfZ+
4NWqZJ/ythp6SgX7y3WlhsQABhIsXHxqK3bnBbGYLRLUZfNF5Em1V19tBknUCUNhgDoilfZ/Qrwa
8qKvt5OKG9X4+P84xzKQ0prqpybp80S3gW9KM+Jjd8dwf2FGlPoDIfsJFtyEi+Vp3CIVFXvvZ0vY
ENb1Ui8qi0NLmJM1Vi9aojozvIKlGUv7qaaPyzQJly+z41muk2gImLz2zAb0fugqOCKDHrRRMIEQ
4liB9Xc3eI75s5U0MeDLs4vBTX3RMXYp6tPHk5s4Lmqmb7yU7kc0cQA9NqYvdYg0fitnS+VD//+q
QhSSI3VsRTCJgBWWf3snEPQHERyLfRoBB+VUJyCzamr/XvEmODO1XoWFmvsUU4/IwUhoT8QQIvfc
l6D3ae8srMDMRF9FE/oVa3WLJfdV1sa1qbtV+NrKHiUmBBooU4PB27G+5/9WM01CJ1LoRtKHTzgB
emVlawK/sKJ/eE7QOglwFstPpFe5HUPldGI8TELfs3oxXfi6X6WeykpVehD8Cjr0sPMskeo3jbwm
V5pOnIoNhJ/sVuJe2nEpSqlFrYcbufZ6pqdQm6e3QssZUIGb+m7iyHlMI+TwbcMRhJO/fDnGjScm
GDTs/fLSrQfKgteTUPDW4QI/8pAVA5HaM9F8c8SnZ5S0yG92Nn2FmsJ7SKS3bytTiFmU2XUOTRrC
MYsCnQAxYmp+j2ghTTG+1D1KcPUob/qF8R3PZ+akkF3idMcHly48MMypiZqyHZh2tz5VGomAiYWW
fVWuCd/ssEl9N4bOO9Y8efu24JAsYV56QWmm33xJ7C5c3upakLmhRSJUrHXgPlGuOPm9AUz9v3xs
e3oA/bEMuvnNZ+vpoCFmtNm3VZO2LGYhgXx3CXPKj0rwU1Tw+vDxEML6kStEMX6kjMoPFH/gTKdB
1FfM7M4bXoaYP+bBhLweVG15KwUIv2TMj6us+A/O/3Db70wA8uOExMhIdwpKznqprrXAN50BJutx
d84TMeBd/Ri/FSWcVW0GzR9oKeJY9XDbTcAJih2sob5NeIUdjC+z1bXJWVhOkB11rFf1jjKYkliT
owN1e/sSxLfsdMF5ZwIqQgvRRWM6sRpRI3cGOdXDt8sef5oskD23jR1m8AjGLyXtcMEgXJsTWxCf
Z5akDWczraXLDnL1Gh7tGSdF/j/67JM3KsYAUuZYNycN6iSPvnlu0MtssKLNL53fPCPyArMIG4s8
ZdexaOJzy7c3tQlyiJmVho0ERJNdwf9Rk7id7jB2j/mKTugr2iaGf34QwVDCu2WpzOssBpuxLpLx
un7QlW3naezlVdsaWTZ/zBkSo6Z/43NbO9MRafEtBd2rv879jyl+ycO9R2b4YgbB1MHGUHGR0/nv
s258OWwFVTvNNN8K8S61vGNOVnHqkdWc0WDwG04Vj251K9kxPWOyVONEPOU7R3p+7+DB5dN/WcYM
lMdf2RGmNaaK1F24Oc8hjLdOvxsl4tas/hmFk5QWiNvTFnSwnY38iOMAKKpDGQ8wXAqmGZ+OcEam
tQGpxOoulVSJv4VR2N9a/VBGEQKMEUc+UxD6IiJedr9Ppv7zMIFnI8a/2JjGMpri26gNMd88Yfd3
2HdVc0jo7Tf9G4ezkPGQzTYOvCseA/3OMYUXOaqcVocvjC9OCJyCVdPbWr3m1l2cPi9VDxpXtY7t
kQ56jF16EX+SGAXLYq7WSG1cCez85wXQNZkalgdXcAZ/kGORth3ySiLwVTlA5HamgHCWb3UCTnxd
kFecrN24lCIXVI7x7Fn2DZFF0hsDKyjJvPxHFQ+wc4GED5GBu6wuqgrotypKy87TfYOorx27v0KJ
SRJU1G7xNh/BxH47eENQi862CmluX/WbXqQFjt/twNZUS9++b51Zhy7dWKJEWRNvZ+0/altiy+X2
3p0GKRRm3Mx/AHhXf4tCLvUQW6in2rmlKgtHKSgMrkjcCc5mEW+u3RrTGSLYPMWU7Jt0ssyJT+up
TDhm4a63z9Ch7LZU7pggS57u0Jmjwh8wwKEp2vfFpTWr4C/KUfvkMTTpLTP+kWSC73mCaYa778Up
XMUhSquCflRTvdR6ze4Y6uU3Zs8lvEUV26R9tOcislPQ3gHaqP6dYkPVd7PDz0DWmR0SDeVq8A81
/GAKUncIhSsrHZngwW8fM22V3vsr6Fg5Ci2B2/Tn35nYBzfG+aTOpGeb+m4cg2pmSQHl/BqQVzXv
hVkDxP59sWzC56QPSMjktuZOjl+98IJyw+XD1bThqnNzyExUNkPWbNr/SDLpO30Ly36Lk8li2jpS
qr/n0PEyg+MhfaCaPowx5kSmuWfKLpfZqvkEW0IfQV03q4f3MlMs4AHBwjma1gijD4G7ZkxU2tC+
8pJK428z4Epb2YEzAnNwqLGz2pZISySQF0JHUpkhLSQ8ZO/9RWKrpc+COZ8PjEpA1mMhsK4Ds1c4
rFa3a0m89nFgkzdPPcgU4Wsx19iKAyiDjRmjcTm5aHvvSO5lH0BQBhc5+eSat6On9ZlKYxV9LqVj
SfIbmR5pYKUZG94NIVFu0eHdwUaPrrwaUVJlRrPStJTCk/Ib6jUgtnTWq8M90+M5lSHJ95Z3hSzG
v3wAhWJ3RNmRQDiCMc5RLs69oKxKJfo+7G20KsVUVLE52yCkj0p06o3LIXky06Eu0KxBtPmpG0iu
0n77HkoJmFNhxGTB9UP3q6GMVjIw1nqFuM99D7pzGPvfruocph3s5fFK9uicG55UmGFwlDCaHmPJ
3qax++acwS5hZ7ycQ7nWHcbZl4ddWnuSYrCBgJiqm5t8w1pa69gpPlcLh91y2SvRmlHvy/+7Fq0l
AO21FiDHPTB/c7j8ALuyXV+csB/FcuN34TcaDU3Ur+lmwy+J5yMnTFbtEjBN9qNn0w++dYZck2/1
I0qclhk+5vTRfhGqsANR1fKSTD/0nWMtX1rNRhWV4t+VstApiMh4aQWWtRegqNqx6qwqPXzaDF4n
3y0nRrmK4Uvw1i1A5gixklKZ30ku/tb3pqdlKYjR5Q+t4wvJf8GsZJ6BELeTwBvGlljnbqyZqDqH
+YnAynr8ZKSzexWcucusLg+mrQcs8CIe9UJXNUjKnJqplmJes+Gc4LveNbok6oD6KKbDcKYJCvhF
MJnm/n4bZKdLlRHw4PyvagiLSixOObiAn9bzIrRgCNmK8ARYv79LfruYDzMAx2gZUO7AC1txQQoz
tIH8wan20N4fWYCtm3m9e2qhV+FXg3emRGTZIVRyFGaQcyYH8ERVDDzT9zN/iqFqHEG4jVTQlk6J
irEuW3n5KHxdT1tK6CQtu3B67pfA231xh1ZAhxrud7IvY3+kXkGm9TmaVI6SHCjh6mLzqPCz2Vls
InLTcr5seRDFYnxvFaLAqkhlsVeQiSw/a2MHRlxmz9plWtuJh/zrC0035MAp3NCyyJ7u5HulBone
3Lh80X1KPPJpwESpMItg/hwDotiFscW4MGo2+w1/E10NhJ+kLTm7LWLpqlL8LfiSpQy+WPaAZUPp
53KGQdw06hm9fzU5QHtWlr+xWeEEVxUyewOSWn+2bCiR3TycN3GmNElTkt0KpSoCqYzUJov3+lgr
8tMzgZ7TRsIxADPb3xPB72NGxzi7U4D7aXIXbIrpwXFH3s5XnvVhxJQ2vHQaTljgdli3YEVUa6fV
bOuRi/FbWY+seSsAjjysmuiVPLC0Mfekj51cI+TVRJZKElOnoVQ5DnZKap84KDzvV9r+epSC2eRb
jdBglsg1zQJyV0IVcO+NJyDAiXzIg8tOx5NcEFfjSCl7emQ3XYLOiRoBruTHuidrJzVJfxamcpq0
JX0aqsjjKSQkiMKe37zXSYvwQQC0LR2NahuieSdwegxiKf2YFegtXw60QdcdrJJ+ixk5AKgcw1oM
TrDdKLjVo22Rm9yRhQ/hb2WbFZMXMpTL4j49feRy3IjakKBG0yKA9BbeJsp1fGzaXK1vswsiT2/C
I6dhy0wbE/u/n/AvKkZBttLCScGomKHwhS2mkmGfruwaBH8sNUzSLHprupHRo0w+u+uQBOXhIujp
FNi8yiuBPOwoMdfF2xyLZqZGr2GW3YUAkulH3cHPo9eiuLR1Pq+QPIzeuleNQjCAcAiMpwpcNely
Ba/jVxRy1LHW3TZxp7mdh3WASkJhGx1OhuOS4b5rjt/ZbkXqUK6VUQ2vQPTELXd+iwlfJPaBF/C+
F4S1hna6hbWxVNRpmnRqLur6Pp+huC6slORfuV830+qk10sbwbHfmtBgIAsmCZ27lwJyJL4rqPWM
4WPCrsiy3sjjeSdKqRVtCho6O1DlbDFV/A8ZddwGPqldHtmYuHL66xzhWToeQlvcm2T+bJoLzyAh
GB5cEfgijCWP6N8mJJOBdj08KZ98GjUFozLwZpCqmr8drpMcu/M54IQfZ/83oO4dcbzi3YoCakwH
h/ffgvjjAUbxu9fOOBwnV74576yciIMlgkHW8QoV/9lTtDqJng21JL2aOcVMgfBxve6PDll6gRg6
7Wclghig6lgRjAmtsKJCvfSpWICLigMpwC2WA0F4WhRkJRrP2jPTYi/RER3ptXRZ4LpBSlELMbjV
H/i1magqiKz7lBuK55MHa3UdBOzC05Xabs2eR1JK1hGsJW4VQ3bABWVz3K/78JGjWTUt7YuR988C
wUJTZZLk66UHdCVKVfIdvFDt9fsODoLts4Kgp9IAq6pE7Epq89GJ/eghxAa+304P5IKqN80sIEi5
mfcCW9aHOetOmr5RJYu1yekv3h8ZCdIvYk8WqBgadiAKA2Eh2/zkNKMuxcPt7ihgc6vN/kZFpslF
zmbD84jDSY+z+40egMeUp3PKbRm/vYVJvCGlQSfXdTbIRCMleG7XGT2FPrUzy4ScgfYaDSbKYPWG
EF2QvAsxwxDCuXyVOyCZCq0llv4ERIUdfJiJujTzJfFSDXxfEhPqig54nD0CFPLAejbT9curz+NI
EYbDsR7EtlqL7OK08/ARssXpvd55l6JYyZDCNGtSHvWHXoVRvlCeUd9TAobLi9D39Xr2uiQXN3Dd
vXzPa2n5xr42NzcSnNJ6vKBfG9IxyhQWgV7gSKSSNbmZouHG+UdYGgGfUHrzDVug4RrIrfe5Tt/N
ad9j9yVF9CsvC4Mc5yGueBSB8kifYXR5DDBXd492y4xCOyzZt8s7Xx5R/yX5N0nu56DydU7N0wXn
mrZb7Azr2mNgWYVoGjda2aAZD6NfUWRwQ13tsazXCDX8tIICjppH0wzMzsrcX0hpnd2SZGnC+WjD
M0/qQ0yUdBcmVKlj8m1anysnV2f80uT2HAhNr92W8APn3YLzx2ZLbpHRQmW0EYbW5oMzYjwhg/Wm
sSCl8EfsvrId6klx8TBicoizD8y8rPR5Gu/TN0I2AXVe44+KwjdYEXBvdaDYrAbpqWZnBQhmOH+V
0RRBdYd7s57TlLZaAwHEgrmyT19lcJx1/WlhwyRfhwoCZPlf+CeRf/MLiCnp45Vb9VPzcsutszOE
frwiwnNa6FHy75oDDzJ59wHGrvbuVB1P5zICJqVMSPpUtT1f/YjndyQ9E/vnV5gxNUUwI039j5gT
2iNO8uob/bkVQLOAtgtd87MsX4q4Ug8zDz2igSi8xY+nMCOOnmqsgXoHG2xEFLm9Mm1yA8Np/fYh
I6DyLsK+3M3IVjcjwxw00x8ryEP0ZbngWfKjgAZjK5wBnvPt2lUhQ5DuYiBdOhGg06vBxxT3EIBi
v47+I1YCxpelfyv/nWkfZjRSC4O3wjb8Tz0FNQMCAG/0fzIRwm3BtSf+987rsZe8CsWKqKkF/+qU
7ZUAA0QpQ8QiudY5+ozaic8HPz0pUkzZ3igLulQXuIcOCJf5q61/utTw5IrE9CIA1bm4bAnmfoQ9
DnZOvXNJ0rzGpqCfHwVgABhJ0gDwWCSmanxRz2Yti30P4hJ8wQYxiyDAdqlZNqlaIGC/kBfjHnPi
xD9ns3v3GBa1f8FzS9VvLa9cNXLxy1mwd25S44khfS9bbuJjuZszbDfvLqs+PZ+Ui6JSTURa8aLL
fmlmrl9Crtp+MdI6rYC6Y1/QYzNP+zQ2k7qh09BqqN9LKrHGQxAD37inuDBANbZRPpQ9c7c/wn+S
cHqHz5CffytaDutmpdTZXNO1lT0ekkJcF8497skRexcCdvcggGpLPjgS9cgOD5wnJGkxpYku3Afj
Ckr1EwXxZToM30elFFWvHI5i5j/MJiGfT6V29AG1hyr3Wev2+EUHqh1DTk4/H0R3jV4uFyH7VCZe
xl5/Vp5iI1KfZgzQzehbdWW69t7p82NMzyyABi1hXcYFSnnFsXI+2Zzoep+Lbu6nhQjaGeGj5Ui0
JjPGuEFo/3p57nLeyx91wEi9yWTykr1uQQe7XPfRLospn1X0Fwy8tphOmwY7TpJGdr+QUWWK/Alh
vK82sEoyNr4gT07pQElv1bEZg7yGhWap/8Xwqk8jZn9sqm2V7zohKxUNmIWLcSeYatuAGnDNR/yp
qihMDu8M/KUAoIwVKtFObse0IhP57Bn8KXRCCknk+i8GkUaOzIBm0gIVbp+hOrEzayc56SeRl26c
l+3vghbyVtjRayl7Nt6XrqCCXBinv/BncIwFP2GW/TtfNbCC/A5qGMEoeOV/1PI6lddBn6otkzdS
oDXXMGo/BZnevyqIgK1VUx6qiNYFeCDO7rkdnLqYd/7FHDcohIaZWo9IR8OUkXQvCBvU63az369Y
YxCftWhBMxUGRRTaWqhWGA+Fg0F8wBSU5DAfXWHPrku8IHTLw+6iPUKWp84Afqq9eaQ2k1Icr6Jr
TenkEeWHPIoMh9ChaYTj9SxPmXSQ8QXcBLUhE+2GqeojzFh5VLN1W476qe0QPwXPq6p8PKm4sJpt
D+I3NxS9zeG6f3I1uSy/1rpnXZcqp35DEwbzPXx/Y2Qzgnkgd1H7ZwcNOtHwQjNVU0eB2QkcjT8N
y/D+efhuz+qJdx0IXEgFeg0LPdajo0HySgqsCkzAK5LE98mSVSvMvFgWIo7MFxv4YnrRUemt0GJW
X86c+cnzGLXpbkKyWWSGxHO3tjKCSfj7j817ijEqV4c5JK/UYneQVK/h/t1MwCDIgRd6wHxcLxuc
jlUGNpdujzPwJPWb7CccrJgaeDEkFpUluNplM8RbOK90jMibX3WaFVSjQIY+D7kWmms26YYvD8/6
pZMtchqmiqEnR81DUtKBR1lz95LkvetuzM7oWTHq5y2SNWWjFUEStYRqbv42wXLkfFiwFWvzLR33
Zo7pevJCCneRiLxNvk8WoLrpbKj2ggnl2ikXLSrkAhkqYfIXdx9mbNIedz77mRMX10cZAx/lTqcE
iNAhgBNc7iKqSGVoeDtGDS6YWr+GqAay0QwQb/yowfcV1yfXHlQi50Y7A570Dfs9OKazpY4J6iBV
ylLAm9t5g9x7AMqgweFEKzyT2V/W3GZbt53PzkTY9+k1SB/KAhvBeZbNuw9Jceafrw9GDsVKA/kr
mt6OASe19cTrUFjTPtGPuPqgxmwE0UTEP4meWNdFM+SKkTkDcPrcdyDPvlek5lX4pEWgxjCA754R
168MydZBTBU46KmMYFOOHCjQO6pgwuIoHkspR594WcJ0FkU/lkBpGa/IzED242byYYx/0JH1lVRB
Uh5/6fzhlodvvubNL29w5QDdbp/H1WdNH1CZ184PCN/kyeB0UnimW4RsPQ9FAMSwLUujMnBG1eIC
s9OHVBBqJcXV7Pne7d0rXLlf7i9LmA08aSvqQTW6c9bV5j8flIWxuUlVSGLBVqEqfhQmAxR46vFC
wynyO1GmSV8W9dhU/fgxRpL9OH7Wu/hjKZM/HDkVaja0mcq1EZRRCQkpXXhkup/mYQUHHema20pR
QQ4wtosPBTIOArFMWlENeXVLTh/5hzpToYSU6mL0NLW6dqm630J22zG0Zbu7gnWIH3QNTXkIbQA3
283GiP3Z28lVZqp4h2fqQ8/GpLzBoVUIwcAuc2QYzVz1dMs9B1NkKdVldOAQWHsCOQ0dgRhsE6Z5
oqULzwdt1f4AQ46tix89LoMJiat6vQfZC2cu9SVQFIbg4z+aHRgOcNcViXg4hUT6VmiHWgHs5B7j
xcxVtU17QsxU9dLV4lmaNrf08or8bhg2NUmC+/G+dl1YBUs+adKWqHyAyqMZLWvuUQ5yP4OlvKFv
PMr5N4J5xhDYQyGV9rd6CmWT/OZ/QBW+WYxRDsLOwPv6Ulw8vUMBr7f4oyvJWpyUz2VRRY20fN9x
iuBGQddSuZ6HBrG+5Ss0/PMtDPxAyjh+LQOCYAK+ZqM2aLzYKZMA4ZH+fD2IdydKroHuUUO4DU+E
47yzEAT1Sb0cbcorGHlGPziYao2o6Fj4xfD0r1pAjbR7VzJvk/FVDrWUUEZQ4OvBvXtvmmoW8dia
65PWsUcvz4rwwhckEj9woX3oA71GlJ1yo9d/EXRnM2B/eWNtitLhXddu65m150cEsudXcEup20vi
7ys3NRsrFKuKZ8iPvUw6AkEBS5DRDLF1SFXZ7q3KfiQmRtzy4sDvzm7zMosgqPz3nu9Yhoj0CtuN
Jecdlu7CmdeYWKvZXd0ZBXBNzJVRolCjYYsZ6VzDh9iH+opblnoTwDD8QXmzzV1vI2EXJ7uKwCjX
X3hDWI9QdSnjxTKhCKBflROsPg+f1FeMD/BXoR6bjtTV7LiwQGLhq+O16QFRwPPBFG1nc5vFzx2x
sEf6cOSYW8jLTuq5YQjJc2G8nwCEvNsgRcpbqcnq387jY0GCflBg9KIFuKiYz3lW3OsRayD98Eyh
USXUOW4hE8v7hkiHry/dTegYNQHh3NY4pIDGtDBR7IXlzalMJtrtj12WeUvzuyvw5WSxjzQurTXj
CpMbx6UP1zP02Tcv1s2qy1UAtdf+wtFFEIHrNQa4/i8KnKf9PDj/yOEz/soW8uOwLNaX6LEzNb5W
9Bj4Qr3QzJk0zcm0A0qA6zKb6YmDQu37ogTFQASSrHvoBRwT4H+c/mQUsKXd62ydL0bfiUVc4Nv+
KQjHKFOp0s48yvooxwWaUibYAJYGqhVOglexJh6n/ALOa45NUJO775ZXybuazFmzf+watBL7RIit
7ltaFHWJb+NMyawFumQprH+8kibivEfeZ6CljSu67e/mLxI+AxUccP8LD+JXGmS4IVDReZ90bbnm
Ts5wb46s6aafQQvFLR3EI703J3G1UZj1ay2lmvky3a9HoWqUM8KX/WorsYd5eoqXcYaBj2whWiCm
YNwJ2U8oteHnw7saDpdQT9OsYjeDSX7t1DRstzZ6T9ydVz8EWFg6wy2Fxrjvv5urNdrwesaV8rBG
68esCFl9eUm6CbzYEo/HLBZmkXLDSGYEBrRZY1wSKbWP1xqllPfQDuzSpt+fevn/rojqSD35wv1s
Fqn9vfgsmJGiuahfkXRwFNyxpqAMMUdLfQ9/yt0mgSMB+0ZvpJtEuDy3XFKoboH+Tkmux++gft8O
clR5gEQU0zwa37IJaL6A5Dxm0jTRVApkpAevvmRgiZ+Pa6ty5yL6eZkY9cC5SD9FCUmat0n1AJug
z1IlGmyKzKs4Ed2mpGG9AD9mLbGCyENxOh14m8Q9OwoGn0NPhf03Dd2hkTg8jsR1NBS4ZrkIplMi
ZGrTHzFVMpjrdRSrGc8VdY7STMLd6i9IBJ8avPQqx10dIzXL2ZSp0TdBcg5r6YnTHWKpZNltFpXE
6QsTy011O46TZl1PpOCGnZphAkoaYP5Pv9kbpJQAJ2Y9TLObcdb9jIOFQSskm5oDflQwoR0qtyMy
C7Xsl3Kr558bYYiU3TCsEG9DC2NHW5c7T3TzC0GvvJCq0yYIaXW13K2/gpVcDAsuAvdWPgdXTudx
4LQOiz8eff3n4D/FQy2lS3rhBxD4GHEyummC6iSEZm0ub4e0R2ZUxNhCgbviFiw90F+oh8Airv4p
cXxtzgjz7xAYeYDcZYO5GzGI+fCYVn5yVDcoGoHg0NdOLjybe8/CPIN08IZTzC+YQMR15gX+IrTm
8McLop9TMu//bya/afGB/j7djyhVgT1TQLDJFoyFxmbnJsrdsL9uVdr/b9xvB/yxoJBtylwe7FQI
RQ6iyPqfZvbZUyapvsGYIxP4d5KlX+TbIyV2SXl7m2vQAKNQNMBZQyX3djalPLIviSUU0NNhfgfs
3tkb/O3Gfyjh02a5DWamfH7JmOMrYyDgqf7CnExPYCLyqggvlWvQzwsLqdVzQdP7um05aed1O8Fo
yKrXShXTeoKboKQ5+zdW3h6PCs1whmNtekQb86OgOJnGQriBccxkgjG+MN2go4Cy2iZwIZD3iUUl
JrCTWftTLPABWipCyrGoALDTttibuEanwXNxxgjgiwxdw0UhHj1VqqItL2WiuBM7th7I2dgYKmZO
GAqTHQROX0ElmdAiPSR5PpUtOG4cJRRlpfon7goAbEWTcRWTPwR7n/cht69e92mSdaj9hhVyjJoj
+MLeLzLFXWpZJBoI8wd/NUQrSY9UqGYzYn5dwPzHDO31itEzT6ogQfd3uUQ+11+u46GKMh8F0yvf
Xeiv5fjOoQEONPXhpwiKLCNdqjidOBlmswTroFh3ijjkPmVNdJZplJBeIqhkCAtDyr8+bYhC3Zgp
zakBuFnBxpViYLo+4PKK3cH+f3F0aPzcEupAxbyxcVu3DHttRCZVC/1MMjkz9tSFyEPiHXeCtuCq
mzlspicqlyxUVeRZWnqceE0KYuiVPzgasVP97fXqhq1A0NNJVrZBgI57cauu/erCi4wLiMxvFlTu
Lgyk+ALWi6i8dO7x9UF2eV5HQ/72YiNZXgu/TDKD7Vwo5AuXAW7/ISMrZJwOe3h4SQDjJ1sXKTKB
YvbK31PAD1VeqLZyQKEdt35pQGh7GepfFPnDEEKH10LGfCdsIFcZkV0kZQiNfzXtb7Oa2ApxAiin
hHPg+jNDK6iXGBuYJH4GnCZA0vu+Lz4i2YZY31bflLypnF6kt1QT6cnHxAxiLZOUd6HcJi3wATzY
sE5IGm58L4v7sh0Rl/UnTYiUMwFWJFWurAxyTUHyGxoR0p2N2v7+QOWC2s1fB0tgAle0GV19LuXB
RRjF7/mGNcqt+z4DHv8N8q21PMH6ZUyayFizsVE1JV9BjDmpY2fth6X7+A9quWRXtLJ1blZaVUlp
3QNNrqlw5XdwjOQ30413AW+oDSPMuVkyafWyYwhs64G4DsthFpMqung5TPxQ9rUXFEq7yraiYB3Z
QCN9bH7Q9LYW/o7fOBawTvQWEIEa3Qtpa7s3YiDSNLVDU82iZkltw+l+0NPJZkwjJn5hvyi7BAmz
cqDJ25dYj5VrQHALFW5bEcg6rGAeVYrVEE1hmeXKopVDuA1qeyy9sU8GkscZpOQJkX5eCAietii0
jTZNVbZgB10LtS4/jUkE9+vHVHYyNZHxits3w7QKFHAk8PeniYUAU4ya7D8rAPihl4mMp+CaBSgn
yKG5LcJ6nFvRWjepFK2M0omx04t+z92lBQnsOp1yiQSpW9b8xHQ6t/m2PiQFVN/9SX154bh9CbmO
1gd55luFdKM25iUfcfI10sKmQ7tZaZm07lt0t293b/gop5Vh4HlHnoheI8cd7Gq0iocZ/6s5th0u
gcc0Lq9Uzmvr2gU3zryNVuBePOSzTXcyAvs+P03r0FfjLVTTWgi6p0TWUZrJNtubNrZNZuXbtMQL
+MMBafQQ9/VbPD2wMG7TxMP7QoaxH93yq+FvBwJvc9f9rSi8CnMVVSDLhNJJZlM6HQ2W32WWgZi3
bD0NNSdDGiSv/sjfeMzR8pZcPcHbpF5e8krpnAKY8OGXcK2hhPj30uE+/YIvuBSpsD41ujY9n+xj
3e3ns4b+5T9LDXp6T07g8a7QoED589/e0sBIVnhx6uNjzO5WX2beWAhLxSy2npSlFnw7VWq91Ndm
23oQg6Rdwdps5y7uqtD4JE3CKduea5qBtxhD3lna5nAeSlZlkcdPbDykmv3NmJgVr3O6/iO2xKBF
MZ1q/hnv9R2Mu4kTvexzycypUf0Ju6pVrzD2kAL+S/Bu4K6ypW6juYtUgXoM6hd8oqMSfvvkYpHK
fKPyst3P2cRmUO3BV9kKB4KY4rOTzBNuEhR5elLnVP7PJ4essPW8Cch39tMCrUOg6LvFx0f3QuoY
Cox4VxLUEjs2S9ZjNc6NeQ4Hc3SGJldXK5XJAYitwt93nn9PFXPgcadWR+tPm+FAPp4eLVKDTdCR
X9260VNHfayzrTGcsh1WeO7yr+FhGplIzCuzQdwXMpU173DNV5NvMjJjB1bulWhTy5JKO1dbhLl4
zOpM6cufJHYXes5Eq7IX5i9OT9sAi/8l7+qtg7n/msUZ1C4ObuUHfqmtjZJJnZdNZ+SjBeoSVIaV
Ir22MNAeXlwPOfb0y2zFYJvsL2pQCdcxkq1W0CuHbBJo3OtZMZJ3vlBuUk9il9xC2DcVQjmUR87b
ysCJFY60Bvu8pBFcS4to9yUtkX11cp5aSkffsCU4mMtuowr9kEEURhgatq1a1RTWmJMT74U0pILf
+TqoxFK2B4XcUj+b2f0EEl2swzSDowDlbVZl5NJT4IozwaxYQouT6FT6ARJTFdCvTfF9coKmnPx7
2hy4WcGiOy8cMfGSKp6BEbo/UtpibYsTKIMIS4uR151NsdDMuP4HRcyEEQAm09IZ3YmGNYDA5Vku
9ditzffbfwo6A1e+KfqncE0CrxRoN+XibJHkCVCiFrs+G20Dw3uVzwIvd4Fa8uKwCFkeYiDwbkzY
y1OIPAKxKGdjtwBqxgayknqGa89G3R6jyBZdyMPisnaxLkMRLiEpXRf2wBveBUdhbwe77AuGnpz7
QTI6rY/GcMpQSWfjHKfDADijId/CDzUjxNxmyefI8Yj/2mhciWjMBqkNAEHfCzoxkx7jrrzMfW1L
9IbU6UZnwTRLAjVVzCeIKpEJB7bq5Uk7ACIHNLBKhPqy+TvDGU89xPhpfb8NF+UHAjeBFJqQKbsE
Wp+9rUCkplnvwawoG1WzgDMmNObhihFJx9oD8pHn3N+3Hgz0Ty78ut2+JuhvmrfA9vHUGfXWqs4F
RnDW3JhU8/Dix4yPppLUv7IYlGOMO+GAHIx078NhcZZYaYXVaqNyACiULaprwQYb6ER9Ro5kJ1I4
FbuVsaNR/6zAQXKURMLauF0upTvZ03RWOQUnn999LkHVUYZZQAjGGzobGLPfQ8OqNV/3UHI83KWc
YRNaGU7fa0qGXQrPrzlRn9UiHDFxL7GBBxxdBKGn6bdVaawzUOMw75n2saFgZSeoZPbrNtmuMVWu
JHXS+ecfEL9wzVdE54R3jT8O4wDOC2UD7aJzCsWGvmhN5F5ATQc3vqxUE1A1vnCaBO27jYqfgMFl
XadXOfk+UQsX7i+auPBrIdORjfm3a4Oj9NLKUnMXzGIRMj2hZou45yJnAAPcKMQol+W64ssmO4XS
QIW53F4LOWQSxt1cQIkVlZw0TJLaRH1W+TNaXGPvo92jXjLpgsnfX/rmAs1dqINFcPbhWneVyjmO
iq4RrFNhvcwcMTXyR/Cmz6kvUsb+T6PwK85vFWUWHiYhNwcyIS+5CudlOgNmNrNd/Nsp9YPxBK91
ZJBKM0HDYGPbk8urcrDXDuLD5lMip14Bj7bpmzuYDsFalLaYaFWwc0Yh4COLCQNKiH3ufxqBT/bE
Tjj0hA0mpKED6/+JA23Tw8B6IJ6SGB6W7WHRo1hXY6TRsT+6KKarpJ9xKu9ejMBgoOMIGp747C1x
AQgvDauPG9SmEDVdclXAl3iJwcL/jUD+WGqoVcq5SlVSeiak2nXnEASB8ix3HUGZytRFarll7C3o
g0Hum9ySm85PRXT/B12IqZ51EZ6Fq/NzsUR2ssLRbAny+sDwEJfbCP4KJeXAJKlyqNi6bosPM0Td
0OpppHuhCkdULJsI4NjliRDx9PHgLDqx93Hu5TDaQ4hN5uyYeIu4XY7ElPJWycST92VsfabpXObj
DJl3LE66xWfkzI5aOoAKRyndB9gZSfS3Fi0SME1cJXfdYa7xhaZ2pmWWS7a/8SlE7cGXYVAUqJgk
OgKseVs8rS1X0DnxhEWE4nn5BX1vrntVRf1/IKd3hj/LupnRT0zRwhXMWzUbpKGUD1uxO0+MJAzz
PWqAsAcARa02uApjGaBpQ9iOfFASZkWHwJtE1j635MH2AkHEa4TN+2n8ZRwY4tCuLy8ZpkT4CKHS
fJVENeTCWlMVmO49vjOCBmPkq4mLds0HEI55/SxvoZFcUULxbP09jr/Yj1ISdmERF8xOZ5Swbu8o
4jH7JvbWVj4TzWw4BstVkTSfpBKPlexij9bLWMC7HB4xIOrJpEn5c5Py2XXWLNpxAHyfDIlMVzfL
UL4TSzSv3za6e+QUHkbocuWa/IPNPksVnYtwrnGrGPnlV036eLhsaCOTmt/mqJV8zglDflZrm2s+
/4lt+hmwmtELgpsgrzwND+dvaQ7L7C+83J5JGa2R7TjuQH46YSNrJ9IvtnYdqx3C9bRchAKvT4SW
H+4PJM6jDesumcZC7u0i+9TDQPT56TbRX4zxnShRqgWHdrRrTk1uU21s1Q3ma38DqaWVk32tYsS2
cKfRiDcB6RHi/vPG7Hy1fTdAeyeE/HtuaxhxHNHQJtFUq9oOCqqSu8nxfeugHekoTW2VqbotM6Gl
uha11N0AzSeE7ppnhDPV1KKRmIyMuGfT/KGY0Ie/Tcbk3P66pH6q/HhUPgXhmUAz9mJsMzywgWsO
T4bz3pLHgW9KU7i6Yo7vaga+eIhOJdY+OGzvxX/xFzBCKledYi+dVEHkE40VkAUH/KcAZfkxP7oU
ujGJRFCp2VWWyzQRLqWKTBJCMIX9T8vdwUjT16lKvtu03ck34hd7XrWHWrvPODCrPHQ5EkEeE3zj
4vXHDi8C1d1ISiloFk+4jnxT7KeXqFjUreul6hvXGBc13Tw+pRGY07R6PTg/9M5WahARKcxKPzXc
Npg6OLQj9X2bqp7Xa/ugRZi3rByfYCRo+eRZiKJfmKJ6k1yNBPaXMtQHezAu97k5MPb6LF/tLxgQ
ldbDRIiXmbUlPhSxTR1dY+A/k3Hc7BLRErOJQhp0CMWZV4BVeVScmK0mJEqWuFtpBHyBRCCY5i9Z
LcIIQ6gEp7TSN3gSimPIYhKZPl+q5Ikq+vRNUW50mJ5HztBwQhwgs0+sRVOnBrViQEznNPwAyem+
M/OOQVSYX3Oy2/JqxD7d3t9GWHmq0oNMxAW58O2ZAvAnul30sHer8rtZe6yxhnYzrCry+rhqEQm1
zw+3gSTNFIrlLqnZ6DSZxJQfAZlrild7Xk9bOTMsVBn3YWkXfncT34PfxqN2cCPTX/6FjIdx8hRi
DFBAZ4qzP4UVg2EkaupSrrLiWRNDjUP2lk/Kjwo4fASEEs+DmnhsROZ0erSjsG6NN9spgO/WdEGK
94+uWKqYiVGLgNwUt/D+ZUOk9x6Rv7U9jUrV3Zm7jnJPI6a2RlCrZSY/S6E1KjKZ5/uiClNS/Ipc
uwZnpRlk79vEwlK6p73/tNq9Twr4fZw9xDi0quCO3I39Prqg2WieCYd/lxL6/DmCU9usFOSha9Po
Bx1m4kvAtyI2VGsu3u/vq0r4Pg1HYLWvgHwXxI9Stw37YwuHqOyzKIT13lhGR0+kN+smENmqayoW
EALAXl3bJce7vofNvgLT2DDoi1OEXPKmemg0mUqOe278gKHWxpYfJIqt58SGsUILOmzVtAgFlUjQ
/crsH6lQQeA2vwMJI1ltDMmelQkyEYy6gbfVX1L+CPJauGLvaolvDUZoysxu7i03KwPxg3rdAqQS
KHYg4Akzdf0BRKLMJcTeTuK3yhNh/RaybjBbxVL6VLNZRB0XLHZhcMORnhnw40jpFlIcGx8Xuk07
Y81NFa/bnjiMuXHrahvYK3inM2pLo9lcUM9ztCi4l8rHeboQaGh5V0BvQMuTGdL0iGVZJbr/54BB
zoCpCcqjrzBFnqawO8ar3yivkGPpSsZAv88aCFNZfJ3+N/pglrFZY5ulEbuTr5kWeojE90A6uyVN
bJyGt6gV3w/f7MCCD7iBRRh9BOvkoF58ZKPBnFYq+gg52OgQnnrLLtLJr1aFyPl9hC/PF7BkwtEV
tR6OtCQgENk9AMdSTrM/iEylg7ht8a7RHJWsxFmJ8Gi/zCeYir+s/jb14G4XQpftCBZTca7Q12XA
DMBrbBviP3LGr4ya51fz9+AXOihF/JzZ/u/Aj6ZciT6c3UPBfZTAZCKQ5WV+USdWIoLEv7cABw07
7wGn5XPmu9cI9+5+HgD1WoOoHi0xmFGCHUmC1o7sjEVzEJkP5Gr15jx2eoe0g4iArxi4Z9Yi8CBz
SQWlB/ed23tpI4y3yAXF/4+8E9Nc/BPOqr4cZNPCajoA6r0yw99r/Y6GMIXmoGBiNrdtPi9KJzZP
bKbD5B8Se8FnU9MN7f3VkX5NtdHnKANxFoGqUKFP42GleLCEpfO7xCSXnwb6rTvaZw5ZQLcDhGmH
7kqa6f1e8DFC7Ev5Orfz9tmaUoroPJWjWgep4IS0yP3pnR6Noke20/OpiHXhd40CVs/SMKrENS/D
lID+qzMPNUdS3EcVuZROGnlhi9JxSvk5xb/A+V83xXFmKvBeg07Q2fqGxHGztme+MNpqKWaUgQFY
rhPHz5NO3fFMbu0W0IaoqDnMsDVnc7xJChFfM0kzgFNdrv4HFhn6p6fyMOMy6g20VVyXKLRcghG6
yBw7vlc+c+SwBqUebvUESccnMZqNY6FPG5X2H2YMXESIYQtzMiPYIv5SqeEM9OtR7njxmW0773gJ
t1sjaAivELYchRoJasJJ41jDs83ZmrWOVIQmeYwhxfiR9zFEv3M9kJt2XnzOpF4HZktHjx1Ml+eF
0l7/T/Nh4Godp0F1dbDZhouvJ9MtOxTU+WlHtf3+SUxGOrW15kDMlcbzEd02CLBhRzKSELpeXYDu
imocBGWxOixcmPI/Mwa3BnMErlGAzrlUIMBie74dd48NCdcSo8p9lTySchAKjWud0k7MvQprFzlD
SgE0GO1zkEWXTQRpTESh8mvSRJSXL+fFSVy9h70Ith11nJUPEqQaphJtmSp99hDcA+wBvP/akodS
XoW1ZHqzu3fzGkeGD7hk911KVL6vZITca7X77COlb4Czima47yU9E+LVPwEArp6WWtP0l74siK95
UwS5Yp84UywhHVdY0SL+Zj+LGd1tVUT9aq/tUF3xtXq+p50Y0vfVKBxD+ey2o97ZiqW2b5r6gP3j
jOhE54Rh3m3V6XxdVaO/EYgA75OMwoWO3nW4Zh5FFqahbwz1VVylBwIZVeqXcmkEVBECno1ue/xL
hcFIIn3qRlnw9Xa3f3bNEPyQn5fm+xvuoTkM/U/I7lZKdv3tHG+N8JNrB7dvoVhJOnNrLvbG0Npt
fRQPjJCynjPWlXn5Buku5QIr4iU/fkdLRHedAz1o5HpEVUd3BxulCoSTDDM61cb4Nnw51wPgl8t+
7m4Oklg+uWnHRvbTg4csnIgPHRH4MzMlMysKnCff97tQ2wOoeypz+TUG/1OenaFRa2VydQESBCDc
64+qQSQC4rmD4A07NoQ6uj35O+8GRVeK60t/FSPDPiQWxnSr+nDQIMqEG5kVUAubvmBDEF0LsRPq
6tFKvT+edPVCZfGjgtx6cHHbem9lCwonHyy8Pi6sfuXMja7ph4D2UCLS+zr6uSyAPJJKs3Ho3OTc
7Bh6s1dVRd/3fc/whYaciIrTEo3eyMdc2xhqxl3OfUZZGBaMIV0Mezwz1LNR19SA2Go/lwHfBDUY
9VaS5tBOU4p8qCX23cAPtjqFyqoQpHTN+FUyq0BMk3m+Ir/0qePGtpG/U0H+XHByy3VlmPFHLFV5
S/3tgfsUBwO2WwBUq2lOcdRDwIkrph+JdD3ki6/Lzwzx9FDZ4kEcQgUD5piN1Dqta990M3WbjdR0
R5I2oK/4B4agfs0xid4vpfdYQI2R1N4hXayIVNlSHhP/dq/itEv9l4iwPNWvfjkiBt3WdFwvalBj
efn2Sw+r4QSUxwWwBw7e5YRpFk6Ga7C55nhGkAsn/8wgTP/b9/3MsDcb8BTg+ocD8IyHurIjRlFb
uJVhjNRR0dGKu7ov9TEy6SheMrxlUH7WG6jV6vuYzG+m8fcflqoUeBLjGfSrOA5amZRg20Y8p1sQ
E2/uKgeGBQnzcD8hY4Tr0aTJayGpyNOwaQxn17SJ1X+knDghS2kknSy3AIfjEUlCkC7L0lJWebnf
5aknjWRVMULAoCAVIl+jp5rcLmt2FfFLYL+e3VnXN+FukO2XFA8Quw+PrmNjT4vGdzysg14/aD6I
9YKd8KN7eUdE3MqR58WFQg5n7NP31U7cMDfijOLad1O0AiPska15NIPjeNo/TLe0E4FNb0DiyJ0v
BacgTYHeFXxpfdbG4xGm6p8vSzCJWNHzTl24SzcDQk37QlUUaG3PKtauPqVI59TH/MayB67ye1sd
JqJvUWX5+A+I0RcVBrTkWN5wuLqx8kLO+6ITcKAd9JjCZbCTeXQzwc7eV66Sje0XfHMW22qI8zyO
aSV5yfttjXgYuQBcDyLmEbsr5tnUEWDsnmni7dcxgw41ZNuiUZfk51EoZv61mla8twewmjMAvR1o
sxMQ7TiXztu5HQFmtyYHVMFUjsbnNGvkfnGt74DpsJFOOpIhLb9QlL5B3lWR1kytuvg0xtTtBDi9
J/p+8RgQv7ykqapwepM1O37knWnpOwlWaQScwwcXoFTqAsgVqs1NHJb4XysTqtmEiXh4iCHrdtdl
17BV+iAZrfosbdQwGMtY487ifXCUjC+WJuuUBfvki4k67L0YUGJmjcQusbvRkgyt8zbFx5FQpcSW
XZNAhgQHOKrS8kuLZ2SoYDIKljuNm1WnNoppHKylq3MgdORsWej/AAtGClCkfGr2CSpugxuf8Uzj
YkkNcKZKspadPsr8T265Uz7n5VBESuIYIzv2o+pRweiCZr0k3pzAVJFE/rGniJS0j1jtFjkmL5ba
ZNA0+TfPNJwQkYYaQjUQnv9bo+jqJDDO1D+qcAtDvm9jOqUt4e8TilyKu9DpkQbTeds1yc/cwCjM
UebacHhno+7k1XXO3xQCh9LkFZJEHhxiuapl9vZVC8tEdtkY97wNvamO0qfxbowi/o4hR3Y1Vt8g
7/n0M3XcyVm9T2bmxcziaUnwEmPW/fSrcFOB2hGXmjiN1hdmQ0esIi+Uf97g0s9AlYsS5jTUZ4jB
GpXflbSRLkTGDJztIvMh+fopsDY29gMPUeZsLJwvw6fOP9PbesdRgwLlHe7G258qOWbO6zTWgIbR
gK6iCY4DlVWZLIgalxk1la9Qz6vCjXYWBxd35oNFn3VK0GMER875Ydh7sayEBoGhf6l1PRTfKP7V
Kdnwgb2v+kzWnEDvVBleHWlNABzjlJ/JRo1D5+QrGL99kfDA6sY4vDIXAJmXO573yJ+rJyQbzjS6
ydesq8485Xj5CbXwjin85WQs9yyqpgXBtxlN9z2GLAk0Cb05WAGVXReG2ubNqoX1hMmrMIDKCWRV
gdULcyLG2y2FS7zjQp/sA1dppx2iDp0VnmUqxLoCQgouzCk+rSTKAjXf9pJnpnBZyaV3RFiqPdzQ
TNQ4uPkpTLvJokNXpV7w6yQgriirH/8aFXyIeLXFuR6WZS1rs5MexHihtb40rBW5eWgNbRXTgDTp
Zv+kefYYsAe4+hdt/hQQWaCT9oVe+Gf3dOAK2N5zEHRxUSza5yBFGdXRLX8BqWDbWAfDaHizknVc
N6O3HhMqjAjq/7dhzhBip1kZjGG4mkFU91XrYxl04mKMNI+cu95B2OF5OEXdDPMIYtetm0OWxmD3
p2o3FdOgsQ29qLTwp+z2unszb8Yn/AuJUczNgxeRyI8C2gUnWCxEhJeoPGZbyxf7HG/PXuZNDJrd
cOpB9E44hi6ygYplFCA6W4IFzsHPiE8ta2GWg5yW6Ux6Um1fFk4nKN7SW8EgJmh6pqDSHEqE8cTx
i+w6swIZndWXFZ41MBpoiDflveXB+MGcEocTxCRjtUPU6lCXwu1vFD7oG0FI/NUAniDlJhhDKkg7
A6t93Tf4wfT4RQdAOnyRD/GP0teYeq1VR71WxYQqoHolThec/OdYb3fgRE9NN5XBQEZz57Ti5che
iOayN7Sk/jq39bUE+ZXt1cP9Bnz/w7rY6rxHCZc02AEu5V+37LDy7+n9P2faO471Y/UHOXnUAPGp
k0345xGyigzLFgezuSguXnYyAx3gxC+8qalyo4h9WzOYKSBZHa36kq/lVVoIZMjDKkGeOt79mEkg
LWX/06gc484wCq+w2xp+H8detP9aqbWwGP+6Ljx0MtT0l5IxVFaa2xXo9qATbTYFP3yh0yZuA6bO
YAMfiIfZGhCRlIHvFGruipyvjVJWRkYd4XTz5IUqXvnVHknjyl6h3M9BMSFLS2B9fq5+WdeIl8mr
DuAe9Vu5KjpMUULuzPgwD2lncjcjG/l12HyoR6wr+QcC4arUgAwdnA62eW6jbOiFb0B+nKZV9NaG
wg25Fb3r5lj3v9jikswy07XLQWijr7+YTXE3dVcKohxKLLonnuULzRn1GXagUpz0YJrdUi80rmMt
eUJ2pKy2uvVpwt1Z2792J9wdgWAtlBmR6f519hL29ZAOgOfFWzX7g+XU334xN1riqvJGBJ7AM8Jf
BLg8uxgCk5YuSYjkl8Jb6TzVY7lIp3rzAZXJ+Ca7Us36FuEudu1xaBpXTdAIhNXHgRrM4GoX/qCg
NLKYxqVVSIZu1E3iSoK978ljTbiAFvQBHruaB3GPXz7Qdlj9a6i9ylssLoiXgpjcSCvu/6ewZ7rO
SiMzc5edOOyXK1t+xHDqJxjmrm5ufiL6CNOfmwga3bylJo8jFpKGoYvwI7957vkr0F2AwlaNkqWa
n9KKATNTRx+RqIwp/MoFxdL0oF5S4fU/pZgg6pPij2+e0MNcIF5g1UdOxyUYqFr0bXTFcNbdUxYt
GraOFcOoIrWeMUuj8iQElsp05yzfKaKm0k4XWeTo9CKcF46o0Z/pnjMWeqkNfrLPNCqZXlWPUeJ/
Vffa0cfFJOKQh21l4JRMNa4mErF5pU887nyGGthFp2JSY2spBN2f8XsqnvmUx3FYAkfauj4pm7J2
KK2PqR6Cvkr7++KXiUzuHJwAEFmYRJKAWksDBsROqFblbVjf4/S2sWcb2WRQS5SlQMugBG9T12O5
PzpEr6fNawrCcXrqsH3uhcvQZA+KiYkHBjzX15ZzqaOT4He672r38Rj5E51IBgB6LZM3kfWaAE8s
aRLklyEY+QJNfSpOEEwLw7lmvX8TguWej29BVvOnm7kKrjA9mPOwz1Oo1rCmhytaF12WnnZMYbZy
GCRrAlgYG5hv3Z1MuGHKMctlguDqA9yTDQymmul+0FyYZBGIo3mDcEX4WcEjJJIRfw+vH0YbTtDF
r+cUnXDIfBxCKcTTevu3OCMxK8HAzkW9FOfFc9yChyY2xFPcOu2Ziye6EWthmjYXkT+iIAzKHkc1
R8nG53Du4C3c8xRzPXU/kmgdLUpKDZ4vx2VfzES6f6QKGbcVNhyf6G4VnrSsYmJK4M+MrOK5iHFl
MTty8IP1gL1YS2RnDVDoDFvvy/2GlQBB07lMa63xIvkKEQjQWCZvYZjEJisZe0ti3+f6p834MXA/
r+jtKByMBOAluGD4vFcm4OPB9/dJ+EkD8HWYg9RAAQkFfiLo4SlsRh4g+76jNBPTCOOKQmvIWBm9
vROZY+81+SXTXQIw1NVUedAtNShQvT0Th8ZwF+FvGcftfPxkvh6LPrJqfALR6gpc216yArLD7GwC
vsiv0TE1RSIHIBNcXd7BV2CIrGdXzwPy0dYVX52kGcGUmi1MYfj4GJGyTPNK7ScN4fNDvdTxS1N3
qOlevjlalliI/O5IZiVrAhVOo4v6jrQlmTewN9sJl9ewRKb+20GZuUSk3SB1icGg3HVDzk7K9MLW
mF04t8tVotJE2cGMWSgJ+qv1FiNRbhqGxWBYwUUjmpi8njqnuqmoxMmEMT2x7kLNSJl1sMEr4KEf
Pqh08vbSwp7DJIZC4cVGXgrQ8wBxUp00ygBD+HUj24mzj4/ouqcWGKrV8BzQmlhDRoHxGkXgImta
iarJnMt8s3VkuDeTL8lULGujTEz9t6BB0bHYUjXddFfKECH/lJOeq2cYRnR4pN1UIQ4obJdPwGTH
FKCaZbXzUFPIN9tMALVETKkbUaeKdZpD72Mwi7qduHgvxXvV+b0CHC6uYg/n7XNebq9MD4ye8U+5
0+Lel/a37Y4dkniIF02XUP/Ne+qQ9U3+5VOx3aLJ3YKi2zX0GGDlK/1+MlKfnuofcns0R6fy9Yo6
g9rQkWWXYnTtzFFY//0+MGasU/X3P6jQrOAxMjjszXcE+yflPHymUwxT31u/OhZ1m6Ohrdfw55OV
QqvsOm3zpXgHnIfMMS46TNeD20NPH+OYABFNGLcejD9u7wbDrnbUXZUVaZrJ7fPsz5OgTuEOABDs
QXm7t53f/kByAbXcaDdz/EvQ/woizk59GQOEzsPpYluw3opkhsG6KKmbeUOJSTfAHH54+lcill7+
8sHpFwN/cqLFpeCKIwfUZwgH25/Zmrg3BpVgh8ryKN1AG4InqrC2JtfwqFFa5W1t+91HeWhb1FMD
8otbrNUEmNEwoadCs9HI6F/r9TvBOzE58McgeVLFJAE8fiYomzvOVEIP7Nub9zGJH78PxKZMeSOz
B5w+uF9XpOWolSLzF0Dd/qKK/eCdUFg5E6Jpk847jv23GvPi6sygBQUazucV849xnkSsrqa31fT1
lDMwPgWIduDQqo+YHR6SW2OfvdqxP0A0j6p9syTWRjlKU6FabM3UDpOlMNYlBMOpNv+DVLsvZbSJ
cFEaCnAa5WuFeO4ItCguQ4HqVJ2p7bZfxeJsIQmUnr0SZvf56ps6VQGyjSo0qE0qRqNXpE13Qs/4
4IIbdlKJQbU+gEHuEYgerOy2aF0FzlX8S3VlQ/0qklPGzG3AGmyU8zyYEhVT3kcoV18KI+ewQRAp
+bGhNDnqHJGWwMyOaHKRHO4/aZfjo9Ok8vF6NROrwHSOLkCfrlYETuzmwEqi9Bj/u0PFA63DPfnv
nZoM9dkph5sTuJhrdRlA6Y3oy+mEy79cERqDiFEe17sv2Juk1b3x1YdbnvdQGl+NkUwOS0ataty2
LGcD1diSd6vXjfMPnrdpQRGy1oqilgJo5VsS3SN4N/KSlpM5HVpTKSy7i6FnZwtblVmKMVv3X8uZ
sG98llg6EVVDZn6PtXZCKiLWaKHi/5Dc9OzBg9wJhJNME/Ar3KwgjNsG5W6a0NJZuUORtP9QSEIN
wqXQIo5WNneQ2WtuKq8tOs8PzOY7euzk6phzD12Be62ZJBo2+eQSEiu3iAiSolWNmbFqtgzHXMR3
DdDKN/npZkUgm8QAAzZewMTkDHl8zX0LVE/ekOIlpNxPLL7QrPYwkGydCA3vbGyAPY9k6PvVKB3R
Xbpr4AHtgfokVWLf80beEoNzqg7EzzYovSBdJP0xKXSkdDEMMTE5wDI5tV73Bq1OOufnVlW7pim5
oo5/XhtpU8sOUu1UCt6levCpfUiETKH5/lMLUeD2BH0GMKOW+X96XqGeabY01xvei3S75po5ir2o
BXIWArMlV59WIVPXVDPVU7C3HuvnHL5OIn0520v/hCOwlsJ3Di7jtjFr/4IDQPx/Jqrb44wLIoa0
KAl7P/T+Fk0dZ+7ZZtlZm7Ti4gEF5t5Kq84Ne9wKmD8nytoUZJHrIzZ286zw9STnWdGZ2FMadSA9
jiSJgehnpaEyrhg4tziL20XMOV1OpFjeqLaQ9APVjo/GFVkj8brBIkF7I9vpJaPsgK1WHE6w0g4s
8NJpz/ve7KorE/y7XwszlSm/6mN3FqWJFE4hg52j+rY94MlytT5Im/Djg/vTwWGBVWTNAMlpgVB7
vbQRAaFZfYfxlXuLaDb5BY4DyBd7wv7/9FVebCGQJGoC3J9MMc0aHDUhWk2FGptd4m1mR3hndWFP
lSNZ5+jEqKWJfVSjLZtrZC3qimgJotYUZDsUHqvucbJrErqCAMZ37mQ65Tu8OpCvtWwqbvxlF5ia
UQ6FLyIfdMSB+ABGgpDdUgaXYOLX677Fs1LLve1i2AHVZAogk7eR6YdV1ON5gZes2uya/RFOXU7x
XGOVGl3njMdxL3mPP2n3TxSdteKcfQD5tphhP46nUxEJaaBdQW/TUfV1rIGDJGpp8aAG0ghXAX9q
DcCvqhQ9eBn85L4+09RYoLduIeGacMsvdfOVu8TQyTX7apUDwQKFV0BHiRTRTnvGaEndfMju0/qH
M8+7nbb9hklvIfD1NXE4USCo/ombRLX0MaybiDvVLMNWBL0OiQr56e+lPdG8cXqSDUbJYP++MXTN
2UEpxBtGaLyIK+beTJekpEjFyWUesReSCYdh2hTckBWM+VFb7oCelFj360l6Pw4H98BR3y+A7khx
SLU5+XTnM89pAvFySAxQF64lZbNGYFJGcT9Ll7Jmv8+Sr3piXc6qN+I/LmUywBO2X461Q/4Sy55y
6G/f/lQXsGVyKF03mLFbwrdGctQmQKlwBT5VPVprFQO7fYKg5+/9f15otcJjWDN9V9aeVRcv7v6c
oiOSyTp03gsesVDKTS9DE7JWOMHHnd1DwWMrNBi10KuHvRx7qSbdY5yNpklwWF/lztKhx8EXyXmd
o4uY9okGo0SKnLl9QaYUBxPNhOjWI5wiOT+QvRoOaBWgz3saV/J6W15zySMj+YXT7bVL74TXwG9v
74X+XCnR90D3Tu/hJYO7aGHK2ktCapqrvLnsEDpAoMriLcFqckOXmMbjkKmIpoS4/YdPo95nHWAC
2XmQSy2gljLcgsX+4CkVNEP4FkkEi/au5dXJ1YJ3Er4hfZHqqiRmy+5RA1Pz8Yb6AF8P3hDU4RM7
yW2s9vnfmFDruWU8UHuP5MuiyVdFIP5XBpTtQRcJ3LWqVL7CGD0ulMCkusNkdliG4HiL/c0oTBIY
SRnmlnNjbJUwwlRYHDiAMPJMJiqFeqqnwqbswazwPk4AxYzJ0tL7NL24b+hLVd/yzkH72BxwGVIL
m8PaGCFHikYPEEk99tKE4I10uKPEpoQJoK9a8M5sTg21WYS6cprVtii0KUsTqwT+6DFa8fMQvj3o
LUMyMw9zws5noOJY24yjD7Rplu5dl1MJeen13k6LsWwX6aREw7ELLp5U2sNqfHQD7qV0nyF7lQgy
sbG/SWGqDBm+FvY1HsZ8Uedy9c6Or3temOjQdHbx/s4eY8vvB+uyERONNQjg3P1WpgKS0XJk3zxg
28q+XmPmR+Y45pegx4KZP2OBDs60DwIo+JBYVVwKpoeoBXypNJuoDfmmHOYlbdb2dQ2U7k4Aq1Fm
PKA4J/4vJzqCzrpLXIrFG4MFCad1C2/OqxT3Kzd9us9pbiXgzfcper7CkgZVy0B/GySeu6PmZS1R
cI2Ec7Niw4Z9ZUnEXJZfG33mR2SISuHlwnkn7klW7hiB0+zzcFHNiT16eu2URdDbKyRSyw9sBzlL
DI59TMip/9agk4trv/syx4JjI5os8OdHlFUS8itY7Rm7jhVz0a/fSrEt+mjcNb2XoD5Ac9KOM2bE
j2TxlAKvhROTTlX4weNlyy+7DoQ07BYcXa+F0cf4RA8s+32xb22xzvQ8NsL2wvp9xwr+abwC57ms
SwwUE3AbggxFWbQ/2o86ERVjKAxKkVdqtiYf2uJAunt6gLr41MysLoUX6PbmDpGqWTUcb86KW6TC
gytzyX1UASeOFDs7b64R5cxsANM3Kfp7E98e+YSCPCC649fbpBex+X7rDOJPemegWFyjkkInUbzR
OlQX1HpfFFqIv8GBKKFLzpxJyt1IavGDdbmY1gODUBlZUJrQIa+MxQcSU9gII5YEBrCRrrMXT9/y
In71CfUUvRO1kEdWyDpRDjFpvti8mHx0xT4ko8laR9uvatTuRrqUFnfmVSpw6ShlwbmQUmo2/U/Z
vre7gjzL5A0RiQ49mwsO8gFnwnpqcBWsqts2fT3alobkU8uvvW+KjXaFT1If5mofznH3RTbS2M06
wmoXrQWZTRWibn6v8edZX0dQWnpsPSPcTVO++7earwbFoEv0wEiPan1bLmQmYXrhCjn9EA6DYv6o
GBqCvIJJypDIkSfkybIbBnH0oyHX/ve3CV83OJZl6wOkgBwQNA68Urgms38MLRd7EVcBVhavvrZk
gm1BANMLLCOIclipjo9DiEE6jnkHQBUvE+5z9ZhpVVHxzKBBiWehOq6fqIeEjLNBYw5+c2LKkzMu
d0vsKI2jxLWkmRTz2PeT+z5IaPUjuQZRVcQbInuUifmrGX0JvBRD9vYf4wgruT2KZ5dygFrsk7ff
c+N1F6QvWEBL5//xQhlX1CuGqhGl1mCKn0GZvbOOVzg4yZ5jZVGJv2LUkzdtUmpRcEFqMrkLV353
KUp4IaKPyqi5JB9OmXQm+lFgYlHXRpTPGtcNsQoynzuxjZS8Nh+X4nbje5T9xX4CjqFOY1ZPB7UM
jOQ3CsMge0kLailRhxqJAIFlv0mtCVwezw09qewOeewTeN/u/4gosYIArpbml+t7lBo0SaMZCxcM
9c2qalK83FV9uyDP0Q6CxIE3brf96JZN1adSPonbEBC/zzjuk6q8ijif02rz9Sx7f9Chmig9g+pG
Od6R+dFrx66YVureJBi3A3NBJ5ffA71v26pX2HxRhw6TLy4VVOdGg+WcatJZT7lI0MKNjv9+qm9O
dx3TiHOc+YBLA7djEDMYmOfAnyDu1jOzI8kkpi6llg9nC5ORWVFvw2H6FwiOapBzNYoJ0avsIedO
IYoe4xFO4Z1I5bpRoeGUb1MIHGIYBJ0sUgbiypsEiMX9qJm3RvtwnLJh2qlQ1TSrq7otDgR/stsD
vY+nRTheY5ibnzqRMHtZyYIBFoa+iAGOxffv9qHC5pxVKM+GDMe7KoU2QP7zgwJgmOEttmCY6+uB
NkBUungPGJgDskb/I/KuIaKxOYQowYGZPrXj/mKtSdOyuEqe0XQtFnlxoCAunq9YD+xI5Y67Vo+Q
2rZv2MoEkf4cGioXo1xwcH/f5AaYP5jhqz9E1316NLsRBF7kmeFQoYbeGWpBndNQBmuBPiiIqrNL
pkmWSR3H37gf8UQOZ2dx1sf3Y7IZZiLHofhQfy7OanM2gqJridGT9IGV5PpVGSa7DJBx7FalIVbR
zpwnYr/obJL/XTH/tC6zu//9Q+aCf1sTXV800nzsL14UvW7gSABHqVByWZ/FhM4vrcRbK/VkwIgK
4nUMAsWETnVAVgaFZcfqgXPqeFXXWx/2sb7b2WzzQW0XBKNgu6scFTpOu9JJ0Fk/21mpeCmva0Dc
1DlBEuwOef4zFiH+wddakECM1dCcAGxP6zMdSkirYazBq4PQFdB9sLcdEfFpI/3UZfH8xzytfL09
/SyhxcWbpacZLZgucH9XH3YuRPpyLsutgbx+wkJCkQ9TFJOoT1mH4W8Q2wXq/G/BLJVg3LfAc+OM
Ml14a5OtF9zHX7kMx1VIA0J6hh13u8+x8htzqaYmaY/aDbAr9kWQehqnPVeLVSP5wGEJRQqLSOwS
pTR2YqbUfdwvN8fbqk6htfqaq+yNXTba5r1r3BVDDhoGQ/6OYl5g1kI8AQjkhEiXyyD47kfpWzFu
HtHRTb6DEPM+LllHPJ7XipEK9uhd3eggga1oqGpRc5ePa388U/o0XdYqz+yWaE97rVGA/kvWI1pb
AJlF2Sac6anmY5hkrkFEJdK3rQP3bBzjECYDpUZsH1FHX2rxO10Q+pyI8UO0Uw8pvt65/Qv+onFS
BUq4Qst7eOZcD5R5EqAfAX2OSNfrp7KjhZqsY6nShvcFW/WNF8bj4Pe2VdbOCD428afCSM6DlxWe
EGAkV0kz5l+HrGSiwqcpr9dgbqtVQ9l2lqiuyvFE4uocL3YuXNMbKy2DY+ppkXSM83ozu4rhBp/3
49erFWRDNv3JGBjKoGnRu8Twqv2t/FGXqlzEXcYqPpP2077UEwPwq8M+po7uePAM9/QDlkJp4+q4
UyQOC2spaIww0PRV5V3c54nGvZtkjhUPqrFZohE9jwdBQUjW1aZCXymxorTNfU9htqMDUDz3CmP0
haMTdgWvLdgaqP+33jemiKj71lmChn49CWY+AU5DOpUctxM/aRZ2mdFYHpXCmNMqcQZg8a9tSIp8
z4XjVjrSjL73ldnMRvjbXhB3hlMJzHEwAUqjtN6M3NBsGHh6vnRI5FiKRQHYj6ZUkboSw99lTSOm
lsEpYb22T0s2dgHai9gT/htnjex+YH2G7jmsj0OTCMjDk/nJLTC9JUmfkoK1ef5/kOipkmTLILZL
fg08HllmancBZx62Tp0WAj+0Nk2BR7eSMhEfXBUAFfVTp9g4zcIdh3pIv+lXw4R1B8e1m4oKKSrF
tbfEsi9Bb5/Vs6XvSNx/WWFDmpa/3ngboZG38RW9c31j3atL7e1Y1twfHaYL5xLZLaRR9/4mnFuZ
3sTIBmMH3OqFQ7Mk5woEvcsbpUZkuq56gaYjGMzY9J5rCvlGiFV05r6X6j55japofwg07ZwQlh5C
NRVt4yD6KiAklBdpUCFPa+493jvuLjf3uj9MKvejlnYXZgYb2LSVnCa15ebjGbi3vzF3CFl2172W
jn/Tbv4h2zj9K2bZEbIr/lyjetuKNScSCvW7Slnk3GEffgsuIGtEXCWsQ877rgcOQHmGw8FI/SlN
BnGXWfu4G6Y7+LqWEPIQO0oNL9NtMbIUkoBSa2CSVmfywgRopiqDjLCRKIH0qX2Ru6Z+480QCNsR
q6FtgiA8Ap2e1eyzyWraNSME7TXZR26G+c7q22dDm4Pdn3AlgJ/WaHPib7F8joyBjEJu0Z0bBew4
k3fHu2HvEzxbgXLLVt42Rap2XkOGtqcW3JLtxTVEiPVHvXa7Ujsffbi2L5uXHxhp4DmJ33pn0PGx
UNQsxMTtTUQY0MbOVU0gbd975Lm7R4wJtRTb0xmqQdnyAqVME74PnQI4dh0fG0DT9dtK2Had7GzR
+s/hubw3xZdM1/F1+5Mv6kh+GBcWQPO+7a5gapoQKXNmEG87kC8guCA6/iNtgXnX1/vL5lTMCznY
zIKjMIPmKRQ69V4Cc5J0w/44BsTbVd/3XYqmR4uiL4+vKft68khg/o2jOIJ+N+exI3KqZn4+Cc+4
wRUerVMRsl25gwF+3RceyVI26hVOLh0pf3e2K/9IcYaNH1sfDCj/YMHOtRX1vUIgG/Mypg1wSdap
aLRY0zUBRwZe9nNdZULTjqujw1+dV0zCMzpbU9JZz6R8M12pikltqbmU3kSZnUQauNcT/ML/3fM/
XUYg2DdWhOQEtAr4fol9mlv07o12MBA46sZ/FAubbLumPv5ssoHzjF28vmBcbrmRmYQvHzFYBi9H
4uYPJiNS0ZZpfZA6TYECkssqy2hVWqmicc60jKtHJOVJq6wcsi3b5fjYPPXVS+0HgNrG6PTmHZtW
P9n+JqF6xrDupyI7iYZ6ZEbJhz8PRaUR+itXgeeGUF7MysmUK49N7akUlDrXO5fD+0lH1KwY+Pib
JTKKs4q8L8KiYK7kyhVW7rLv77Aovcwl4Mfqo3X2auAliMtaGh8bg4Pxjut6ZImkjZ24XUy7IXUQ
P5tyaFwhC83kTvK26UwAvidFnbn1hReA8ekBdTVrudNIkJgDIaiFbrVYVnVtmfQkyMzvsWaUi9Ri
ul6u1uH0uZjIrkwM6AFGG/qYSaP7fZaeaZW5w1877H1lYuISEGwEYRbvQX/7dVur48N8H4ae4K+h
zNfUwYy0pAm9nHuc+yuvKtWiomsxdE4DhMWFaBV9rpD5OZMDQJ+iExrx5D7qgIGIRrK7UtsGyawN
PbdO1TVcVW89wUF9iqmDieITRnvsNf3OD5P2U674Rkk30z/4QhCbtISJTmgoUqEOyNzIcVEr5PXW
OQr9u8slQWMfVxMVup/2PtnJNgTaMHc7iasN6/j8LQ6UUnO50X+5zC/gTYjv40eOMOLXFv4FqDwB
0CFl4EgQOMVp45axGWt4drfJlR2uIN7KoDYreVfjiwouY/CAY9J0jIHPHfDPmNLqwcwz8yM+hUQn
5nFv8qi6sLzf9HBMHGAidexCy9GADYk7pR6KilEgOYQEHt1s0X4ISila+63gFoU+GxZ2XXUmCsR2
EeIqQnRllcj7jxPrpB17JMsEB47HAYGAKue5gdEDk9ATpI7TodM29FQDKpaPyxnWmx/Ex3aJfE6c
bKRggtwIIFDheoOOSZ60E8jJKmOWKridWKMpHqS4CZsn7bWjpZ3hs+KwSJBp9OLBbOd+xDnY90sC
UN2ryKTa+gKvLsK22wPJOnWFAUc7bpInkAaNdhU+CkhM3lyFMl0TVk/BRF1sL9oCM6rJrpTQ2TKF
oyLguviAgX5o3Bb5CvFzrf0GWcnbH2EXkS+QY88do4hrDWpESxlKONCMHKxhK1aLdWWLcn0mbJ7I
ENR/U9LLv/2pJOy+prenJjfCAkWeVF3yaev4GSwnQJ8cXxWiQ/GvFoCFT1dYl0gNXrOpA51fWskk
ebQUkjqV+5n8KdBtAWqjis7/DAZtjC+MLqsaAFaRfxspL7iZCVkNj4MNl7bAp1kH2W7Uiiae2tpC
qoeZr8sa9CTNe42lRIObYgYDaZ+UWT2pk7T0UPbgIOUTjwkc8zZbvtQwpIoVfOrse8e9Z/yJSVYC
j7XzadGOfgvh9X+qGI+CkfE0BAgAVjHRqE/Th3WlYmaCSgxsBOFEQIhiHi4g2xGfyf7UpF8ffLmJ
5G61ytiahO2Vw4g+ZeeELP+jzW9nO/Y4GSfvPC5q83U3hWrAH22M82c5S9/ZjOWh2CHTsNbTE2H1
V+OBdCqRuRsWn+x8thayLvxYwEboMnwfwSrYXFIlVt/qh+MGwS2Gs0VJr0+U5uZZkPVgcrFSORAP
RAa6gIhBDNWDRW/f7hvxxEBbkrBbhE+EEy6hm0j3hW8/RpjcZoRJX8Bp3BWtm6Ote+OIk4NlrG5a
MqGROdyIE24kAiqtIhR11j8Q7S42Guqldcmf8A3fU0/l5sBHmUXBlNLnCXj6Z7JirueQxr7Ztp3v
C0oa4Jq1GsWSvihNmk9ri1oFniY5126tv5utP/va7Q1c7SleLje2jlXSL31STHnhVheVfnC2L1IU
J48mvIILhi7EkZ66dhNzW2Uog9fi/kUFLxVC9jdwCJhRv+D7j5wqO7l/AFBZIZ7xFXO0l+4gfGXE
wEglcYqwht+YfB6TuVzATiqeNnJ39PyxBlYYMKf/FDInEW9EY/fCZjrZhO8M8Wf5uOqa7e5RRAEW
MrZ0wLiiS79ZuERTlmCKop2UhdUuQxhu27Dop2j+CPDU7Y9ECdwsdDapA/IP8IO2siSrPuiP2KkG
BJYQfUafcOsID6dWQtBYcVgLDlZTz9teSMvcLSplzAGQwqGQXDC8/VHCtVylPOVqONZZNk0g7QnF
0HLe1fXx48EvxytApRWfcCtLTA1JSJMHiGsqCNF1GH2HV5CatczsofSYjECGc8vzGfsc4rTtFXJ7
tYphlWMhRHZPubLIUGaerljQ/OKB9Wdh+6ZNvOTwfbJhtoSPPOjkWKVaJA5PGBgtOJof1p+7FpHi
yGmkZlZHuCDQu4k+NvYgoLM1BtcZOFGtFYT5PLWjoz4Vbd+Khm+Z0yOfG+9Axn9K0viqPWxdrvRT
gwIcgDq+tYFHWQV/HVT/fKbyC6UvU+9wvcCbVojBEEPmUy8Fbfi5LaPnTctPXaAcxgHr9vwz3lWJ
k+0UW543KMr2Yo7P8yAa2sJi6o9kCic03uEyrYOGxbIu5V+cPKsUSKeTRzCDLudtGSZLDRJK69jD
5bxdAyCpZiElmcILudjXJk/J6EheQJ1EuXPOBBkemA4I7FbTP+cfJoLqI7p10GXOi8Ajyhzi27go
P+Ee4AHHL8H3piDtu52bjgf1s2tIbeujFRVMegbAp8GhpxWeJStgfrZJyyETzW/Jsibjn9tzcKdK
a5wnJWAYMoDoVREjTUGZQ0bK75jNGLREQ4aBbSObZdk4oogyQQX7pCBUlfRnnlz4GHH8cwMw2zPI
0Cpj1fHlxHjtB/mRrFSzvspNlkE/I5lXIxQbcAVTcoR5Ct5kLdbUPlkM4/76r7JbFcThPiAEElep
G8OQZ/9GCVhJBSq94saBU4F/V294DTaV3z2SFWvKcchWWV1EGvNllceAzui+7IyeY/HF+w7+Lhyo
VKMmboe7CTc+GI7otm5JbK7lo9z/c/623OFdyAHQb7kjZkZii0WKxQ/GFdRfLXZ31yQ3TMYdrhse
46AgDwb0pCCayYdD/XctjP8qQzOWr5db76Uwb/GgFfurpbVy/x8SDTQF6IpgziiMtGh+kOLkWdA7
I9f4qQyh4GhFo9OOD1/II7zXmkgjTGGEr/BKMPtp1FYJXs12PF2i8XWnUzTWFQ+IXra6Qu92KqLo
gdjIZcJoXAsjywQD89YhwtpO5tg7JqIqFNeF4Ecu2oKIBZHCzLBcufebQ2BEKJXEYUeU57gfqyae
EWpkqJCDIHUlhwQPGwEukU+Jv85+xxPr6XjnNp+hojRZh8uMYlwtyo/t0KemXyrRguSMkI3vreb/
onJwxHwsrBd1we9Tm7RCBiaPUF3Xp8ykToNTGrXeIhc6NL72DciJwSwhGkq8y2vpKEAO/aTASn4L
mIjwtID7rqH7+sARJpftbT6736BXSEr6YmOPrSkpyU3kYmCLEVgS/mxZKXIEQpOp17yJLH8Uggr0
XPJlNAS/MBHLgkjP8FwPWqAW2QW+femaQW0E1i+6xxC+jbVLVLkCaoSFQeGChtxovIq5T1bM5XoR
2Uf/C2X2bT48xCfmL7obaI+P9yTv8yjTTOoV0+l/bFJ73eC+j7tx57YS9AZTADKa9LFBrMp3HCgx
LRAKiR8721iapvVcnIK6qXPDtygBjBJ1oPFydRIWv/qPeesaila6EiQZEoyRQTMcuvE9gQj5goba
R+Bk6UuubL3x9MjndjnK16XXim4sAmPBmyOw6aFwpp+hUM7Q9w0q4XIce9nxqSQkRW6cFdp6P2tf
a1kqAnbNVInNfRz2YgFQlrzm78igPRb9dpiTv3szHxgnXcJD7864a4eJCWAiIZFtYWoVuGXrvUoV
7vkufhscvJ9+Y9NyaDSWoZ5Evq4RbI73TAUmymuu8rlgw6lev7C8UAYQiGLL1s1LnFJw9SV2a4xi
xH5Fg6gi6Ix1sa0aZdKIJY7EVT9ngK3waDH6CSv5tkbz0t81o2WowRYZtx5OOztT+QLv11dht4G2
QoYKPeueRxSrXlkg5NecqbUooR+UMiDKWjNpLdHq/YZKzhgwWrFo7/9AhNBeFlFlsuMPmh98A2rZ
WeE9G3vgsiEQyViAOcuyb409Y1uUr5iCANxEBV7xWyyXt9E/E0WPHZnJDbFwnTunA73hjttp0Fvi
76cLiYIcZK+Btb8L528/pDuzB7lCPwZjSrep64aTdoQDrrRvpLGnzWiaG9RAf5M8UX0LQC+2KLgE
uqXIT8wrY4Z4LJy8tEecGe2yhFoS7ekbdVxSNzUDTNCnM5uoDM56Rzokmp9XrZwkxur3H+j2fu/j
Y6uKGSzgGwjJsVSYapAsE/MRWX9uMeuRb/lpskGq7VpT0VWDzuUEKKEoy5jBKTbtrONOF+D+uHyK
DWmHqd/L/j/C0e7/3/7J4QbRYnzqfajjyPvvbMK+9hQbalr+oEW1qkTXuaa5e5r2HdbLAkl9DjTZ
QeC5NsbdVUz3zDfU6oJlt5fb7DrFgsRyA9NurRL1e+JKNWWSEBkHOndKdEHiJzh7i/S2TMps0fsg
ZJZ2FVDVe5Zgkw150byBaLNFzg79Fn3rGucqzknjXb9s9S1GpquSUFqjCY92UdzMqHWVyUV7+9GZ
OijCOS1zdnLNDs6BijpTFfeRVcsEbkM8WMHjfQbDceWtagxumcynwvSqdIRtN+E3W1mJF4zuI+bt
BxI3vtV7CAcJR3yLDLpX8M1RbS8q2F3X+J9hZJV1thNl5lEXdEWCSJSg4278MAssk7inSYSVNuUY
RnM65Qy6pUzVn1MG3gPzkSaJcQhf4lgGi4sB5+K3h32e5jf8cb+hTYLnM2xFvWwHgABlKuENvEDq
lFMfnHa7p1cXSo+kztxa7slgYcZPu4/A+uCr8UPIMptDOlJ9XjuBRUaGZ+edoIxoM7ysyu9UK+Tk
a3Fyt+7jPPHwLj7Jmcdi7FkltZsQSQJI+rjojVIVjnSyt3gOddsBvGPEGVLljPmlKctBQ6TltEyu
eQRdCvdUYB2NvQmE8DoYvI9i4e3tlAqLOSREVIR3Opf7Odbjp0xr838Icgs0z4Lss8S8WKKA3ufe
2BeT/kdYY4YQohzSXmFb3vgjBNUB+qfY58s/AcRVJXye+Je1KjEay26TCc979RQyFp6Ums4x3cu4
6LAOTjaCZp+SolFo+NVW6LuWDyh+hDSRLj4zjL32TpAB+C06LRfdPBv8VE07yqRvqOny+N0VXAQm
MOiAc5lcOUxiXzXCKJie2FrWUQRi04ro7rHNuiVVaDDls9GLtUNtzSgdcV1anO///amJ09Ia1MV5
wF+LN99tI7ivhucqNziX/0o/kbhfhsLpNm5ZZJIP4r1bMQZUj8vD54bYIuIk1hXrReXX12tKAPMQ
EXRv7k0BPdmSYE6xhVyb991EJ4Ug3lnthvv0jX3aDCJcko/XRgGEYNPIr2DQ0I4ZyVDGbX5IAA+Y
CL+rkC/HC3TaqLjZEmXw0Y42VG5oHBH56YzuS4aZ3FWRgavFmH48225zgyzATpQXz9M06t3bd3w+
VHdoIO4LlAuDgpvpO6opYxBhfJi4Vl4xXipxQ5mfVIdq8HadaReVL1meUi4j4vp3k4lbAZiXaJ28
fgvoZIpPGOmoF5AO6umiO/emKlqFUTpnqW4B1wYqzJDLpWSJPS4XA3I/wiyQYbl0D7IaUvdp0pVf
QrOsmg1xAc3xjkuNhrJR6zaatbbtNHLrtNAk9HftOMXd21HLuxgIOmUIWaJGjaTYkQOs1aj93ppy
J3fd5UVbIa75w7cqfNVWnuk1VXSdOibWqsdbCXS/GOdTxZJlh1+sS+uzoulBWUoyOmeREawDhhjy
isil8CpSHa/XkOaDBSiDlUdtpubSZLeNdLZL9Gi02NlgHl57TsoxkSindO2bY9BdhnfPJ5txa+y8
DmxUbv8lND+jbhYvytmasZwB5ZumpgFptwCSYEXL2uWCPtLYTYRT2RS9w2NkP/UG5vVrM3J8PYBB
+hKAAwBrzaGXsFcE2sHdANflWfVv/nvP3pXVsHqSzSfO7G8/YzWhLyi2XKfio76AntdMMJZTLUEx
CdrftB3YpvsijP3Yn66jGd5jbKIEw54vAxoCgEdLOyM3vP/Ht2R8LDrdx8n2tf0QxumyVg7fcvPH
hB82UJbeOr5+jKAveyw/4ENo2gdzbmQHdHYY4M833ltnqYi0qo4BJJts3fsZaBZoQSQkCXfbLk2R
BzxvWn+AnSTVg1N4qAlWe7hDvjaoe6TvinIA58RgvndhKoO3TCNdOPZsJLKGbattkBzZqPZxrCXv
J5VMf75Sw2Yu8JzbxrV36MYcNvg3wq/5WSMVW46Sjd4t3YrdsKKfgm7Rsdvj4u+s5weQP/ScFpMU
lC2BTwTc7Cd0E3Eh1HZ0CHJUJsJYNVkUhH8idxtlr3UqaGfXKa1KMTyOh9gxXXei2sOzyebWOngy
je1qmKYgDfxfFqcmpttG+4o0EShDrGQ5Ek8+WzFI0edUaBLIvzu6m5L5tiWsf6btMNgNjnSlWoo2
w8nxxIru4XoG2VkpISlotTNgoAYbI9Y9Qx24WvCbJRnvBhCXrSbd0S3FPpQCkd9E+F4zb9BwjlHn
zSlDVC8pX3S4GhIAPSO0SZ5iNqMA1kSkCBp7Z7rbCCcZiaOZSqBebqZNxmyfrr38qpwMrIOEricd
eZVsWQgn+5+8wNpmYhfpbxFO6Ssbipp7Ey9CK/Br+2cJRTO++KtlQkYWoNmFRk00MduO2/nIZFGh
lKUJ7zE9G5ZN0FBi8ZeTyaQ2ExpU6QEv7iQWC3c9AYjFb8hBYisCDSWWOAgOpmENNuq0aAdMsDc3
y8Ff6dSlwKosH8EZ1m/9KC7CaFvecM1CeQZW+8u/6i5OblRleTinNB09RYuUUFZL9GJHNBbrID3k
tkhf036Twmi4dVnWFp6RjQ2qgXCpXAmC6eAR2AWAvuJAiVGsYP24D1h5APuyTz4GnciJevZQiT9q
0HQoHb39E5CK1s4geO3nmiscs7S1Cp8GcpateH7ErgevcO0sYPMcDwk1mH2V8mYCYjsojY/kzUtA
3/O0/2EkR535BOLjz7Rz0IEIg0q7NupCkitDBmro+Wy08tbtVVl9ziciGY0mFbLkbyAy8Vh8ZA30
t7z+JKV8wU5jKiKAN4wW6tKbKJdrcWSDwxndQ0h7WGEYbTMJInviHlfFJAQUnujB7TxCJVtYcGyl
iRWjHZxxrRuNrG4l0S+qWXhHuyosItIKiVZJNzrwcpujmx7Ewmq/B+t59ZTxmaALhJX4TNJzkUbX
Nf9ABSD2pTAT1fPoyUYAVajUg04hd/vZBAgMh/l+VcMXtYuuIraQik7Xe1Rsntr1E8xMmKDGWwf3
Pc+XWL1Biad0Q6XPpiDs33AjPx1feFROny0mdbanTmc7ETKTcSgmjD53VbdhwQIQugXN5EVGEWuN
M6Q7/vwZ+sdXmY+F3qYQlZzkKEGfm9/y78fEKVRzcOdFRY70JQD/J5Mf12R8wtIVSIDaYrW5Mf87
vlejJgh3IvRhzzsoLS2hvsL4E0XsBaWaYVDKg1E/t5IHXPlnBOYvZTesoiF05JBJzkprY3Ebf4Dc
yKsVFqyxuHSCEV8opDa0lojCibLbPGh3ots+nrCnOw7fPyIoya3PxfYvhbhOIuKW0cV0uvVYsmHs
n8/OR+/vHixuj8weM6FgFz/4/WPKZxuaVC5OP0MF+mgALBliPAp7SOmypxN52LbN0YVqHi0wRbYF
v1VA0yfbJ8T5LtT3TtImIgeQHdwal7PmS9LJWKOO4AWlJNWEGScwPUCgpZ2fCBxN8YlnhoPsXUCz
4oKAlG3TqwB28vFQiEpfodUKgPdFx0spzlecSPpLtDwiukFr9PTx8HU0sBob0Da5vEEc5tQg6mWv
jdbsQmgS+SutbQ+CgsxxbfYXIqisqOu4md49OsoM9bTexUk9z54NHc0djWydy9SYyg6t0YGHdEDw
VC/JPbbLftpv1q1Xl3IRvHhyut9KVgHJQmYW170skBDLUHkydrBtdu5nPh5jBkhPNtJcPp5d4/tN
iNWzsA0/Q3YDD3WLv2L+wx/EVRG+UNH8LD+6Wi/MJsG6V3ks3WLLmUGoaclurio1Qnn4MGvd45zf
IOjUNKp/Lbgj1sg08TuVhjotZaTOPVZqyrjAk+ID0/+m90HLxX/dpYW+aRMkbOqhyQtye9Sk5yc8
u5hV+JucF8XAPXdrnzsIKV3iJ4P17vzE//WZbwDnGL0Z2+qJ8qlTQFS8ZT5V8uvfCXDR6vFRRMv+
1TH49L5HXH9vizCt7zdYrkNQTs8lcXKArRewHEKlX1V5MEaTe2EDS2CBT/xryYUsf26iMH8+fu1V
16Bc5CjYEhYR8bWyo5oz8TOF7uwckGDFNcHwrh8ZSvM9CN2IsrDC3q9g/Z9LbNPNdCJxf6v1oIN7
NzO7T2L3Spc/ocLuYXZWt5nJYcxBGs0otKSFLD5CWt0yfyn5Vu2XLZsA+cLbB947QoG9CXBYIEy9
PvtpOOfyW+yghudT1aIrN55eHVA3yOGKOFbiP89QusymU/0ezAtAfmvtrRTYjz9tASYYtRZjfdk7
xFyJbjszZyGeNP8BEf8eHT2+jhiodlC3ipghz3tuLqe2+3vscjzs1GZOzIyzIk0h9Yb2dOR6cnD8
qPQeHgUWI+lLSHq9hAMQ+rRt/D7pygWBokl3uwNrIKuXr31+ntdrY/n2ZdlQrSF2O3rntLWV4J6d
GyXwkmi044yu0iHI7v2kAdQLoMdIU23EzCVS2P9spwY2gAj4Vb6efqoyAN7Q4JLVsRpTB1WtEI8F
LtbtoRYYOSNOFSuTBX0PiFUgy4TV8kx7nKc3peRvHZen6lTH6ueEWsWXLb2VCZhesM8QFv/u7jni
0rNCwNYPv62CnMee86OFFqdKd/12jAv2pRMs2M8Hf+SWExZO3UgDZX4zZwttpNGzZTX4eSohpWD6
CUo0xSiQM3/dQuL7y4tVT/Z94f5TWQ3UBEdgH1Va0jjlOpa7lBuPhEGppAR/LMuqaeknWv9HWD8/
ky8suqbwzrEUWIlVnJyqfZtVDLXzQCVrvPGlpRfRz2lqb7IC7xne7etwKGKMRJrB8JzUC0P8q9Ja
kD89k4HDTnyCvYGIasqCPZOqybo3AikVRoXe2G1UZJ5rMTMY3y9kviexSwiSTVKyExjq3eGvfJj/
PGskOy9B2+ThtN6oW2MdwUfhAX2Z9CS0915UUEJH3GLpCtB91pUigXicfUClwtediaSvp2jqK5V4
mfMMF84XZgpx9NKVgTMI2cS8nnnee9Dng4SL/nvh9PwWqTEkuzt9cPG3ESsFC/0OrkPCPl3mgw6s
hH+clmfiPcX6gXGRKql2/24C8Eor+gWdGk+6QL0FenK3+Bb0RmA8zPJ4sVVGxbgWGhSqyfR4h6/4
7iti6OS9aFGZo/E4Z42S4xDTeUZisE5jlEoj2I4lw+jHdpDW2CSo9PIbOg/1DaIS+UguSW3FptQJ
/ch8V04eTONrnySe+pHH5JpGLEoUqj2uifOWMWJ63/n71OZa/VrwEL05eFdo/e9GA31Mr2qvaL0A
gMidy+aJktfA73O56pw3a4tdwiY+XIXv5nsgN7t3XmXmo76jbPryuid6G7Lw0JrISYejIe1ZbSes
E01JIZ0XdXsnnkz/MzdflTgPYBMJn/BTEs7Kdju1k2cKgF4kKwwIM+3xXNZfxjHyYEfcW3HB8rBu
JUZx2h6yUZauTqQyOXosg4zPNyNaHPFRLZm6LWup59r7WbC00/VQTgIyN7qwGXOOpMsE6IzNzM1U
pmIfcyMO41Nkf5Mp7eD3SzKjoNtDWvTdkH8Y5cCkNU7i5OsR+YIFsoMhgcE1SP7KwzmHmbfgYMbx
af3KwFOvTUiVLR/flMm5NVfgQ/JsbxBv4IFOAV9Lr9ucurqYi4NjkmDQFQ9r8cysS/lky2zotUQR
axnDMznFO7xWmdhARM5m4bXCaqVXeYJUq4Obhs5Kk/COgjOVj5e2vmu13xzFI/w9MBloFew3IIDT
OmgWp87kf2IVQh6IcCik8WkietuPdH5p4reYEP/GpGf4BCD8xAZJxrje0PWDaQY76JR1hg62KwK9
Aqo+1VJduEAsx91wkxC+qS7tZID00DcLFHaZFtFWP79s0Wc4f71JJMBwnzTERFZsuQqTADZ0olZB
H6Z639rGuN9NIHdbIp7kiNTFsStqtA7GFiTp4VzZh5k05Jit6fogOJ8n9z1l98gvh8DKFgEzqdMZ
CHR9PjN7Rar5Gx5rQvQi3UAQ3UFZqeC1Mls/Vb3JZ6lyQ/zle2ME3ehb+xKZKtaQyqbmixb1CzYW
Qrw1zcpD/MMgN7UXY3jBP8S467JKrGALjxYFSAxIqS40D+yYtxJ+LOsYSuLbzZteWFbyqTQZk7Km
2UC9wyGJm2lvKkixN1yGGYkfvgwEVmd9i+qOT1DbzxO+43Z1pnhrz+KTJYMHs4r34BngO9T6BMqS
FBso15lSsjQZrXFCN0XxnvBLnZvYcHyS72AR8JdtnsBI/KzwHzmBtkSaof6RhFLrz9LiPuSKaXMY
RD0NBBYkZd3SHk057zcuq7aXOq03oDUOB1AbcvqJeuqO5qjq1oC8dVV6qsVYmqy/1ZDBfAaBNYai
eM4yurGpMk3Tixto/sZjkl8diBA4lpACta54zS8u+KVr4GIk530HxmcosJlXNHkMW3mszmJUolFV
bNxqZTi+wmoIFrlxF9ahR6LLrLpa+zSWLvlIekebuoNbZa3I8ygL49orpLBzPvzJ7r5N4xDA0zgb
jZaBTLHn1Q/qRA7ExHcHOoIBaViHFEZd28byYHt7aBpBGyR2tWcUiBAS4fI2s60oldnGGgDyUAx0
p7Y0SRBNtzN7IylgQ0nDnjjbIloVAWrwPrPxcbw8ySwOy6AVodu/Z4jySyTAv5D4WRfnzNf3hGRq
nvj21+PejYQMtxtWCpYnJP1uz6wgxkSaBGnpDPLWmqwaEOO8lGfQ2fiOoa+TdWg097RkJEGeqku3
4B++NM4KnrH59WS4e9BBBJtBcGGKtaOIbWaEkCENYMboL/OhTa/twkVy7c1JrDKN8e8bSmrKqrtc
Mojywf82m/cfJqmZw4KrW5uA3JYhrXiuZ0f26B7+EDaD3XlCuchceluSJW27a2rL6dl/Bifw3rg3
+hSiHa2cllm8W82ECJGXIVn8ShXvDcJgft6lz2IPdQrvGX8V3lmWg7U82PtvOHfDXhWaQZDM4i8D
s+MCdifxHsEuvHmP5la5/O+UbdjN9mO1ca/Ub8c6al8a8M81I7tkdtnvpk9IYKAGk7aDxCYyLQ1w
zZqt+wLPJtC08SIcEegAGCQgCUXpgSgBlfkGztodFvjYDh5RYWWhl6jBE9lpv0SXCjF/fiHKnh7O
cOuhjHmy7WAQL8ymXIn1U8Akiyjq8hhJz8oUW+j1B0ry/Zifkjk1YAYUIXLh00wpN2ljvX90K7iP
mu+VU0am+j0tAloV1ObRX30vDD8oUm6hs9th4VQx8VjNr2i0PYlEDpz94+ulvng77qeVrFWpdBHz
ZkY/hCELt+dOYihuKlOw2RoSM5YTqUQNjrJAplXb22IxQ9IUj86CgOGTk9dc1rAwpEFfXLGwKxuz
TnvuFPMOqcUQzAN4d3il6+KjRtwS8xE+ZyhcjcuwDVik9fZfSzyii14ULTGop8hPIfokJktD6xPG
UljTBWui5d48NulH/5swBBy3dcudNTH7y3u0oWmzGB+PERAMHbKEz9mT+4hcUTboH9OcUf1iDnPe
PAkBFoSpb+1aCODT88hXJPDsTA/hs2hBDhDnTeI1iVIqyOmFftouSbOaRZdK/Zs1zFX0pRRke5fY
nHMmyNc2iHw2wAF4jXpcqEa9S5WZN1lwYcJrPv7gp6N/ZogDl0jK/NDz5Je6Q8ppsALau+OFzT2Z
erbJa88rTUIZzQG5TMn8KxsPQuhC6JgIvcxO5kIFs4EX6WV4DsjRHSb9vlP/HrnrVEp7JvR7p9bb
ZYLKdn0K7YD14w/T8BxTIFRQhiBRsGzx7cSrLLqhFD15cpqgq7CgANzVaY4s/0jkVRH0Lw6oLtil
WsjtZ8NGdTjwfYdDe80a7p0AnRDDNDWKZT8OyUOlHf1B0VTJN2eUEueZAjIy06mmo1RKebGgNLtP
5yixRlkcH27pnLgle/Fqy3B6qrELT0onD19LiQEIrymUNrfVcdJgoibZ13kcjef3nUIXm1GgyO0X
`protect end_protected
