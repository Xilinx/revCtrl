`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8032)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9TaBM/i2ZgCPEH+TSdpehCfjbUj
/XmKL45eczCMcKYnyQPFoB2fnevdjFZowlTVLk35CMBd/vPpJZg36EztmnMalx6gwFxB4DvZWaM/
L2uFdKUbPyI9+VKZhbEX7L5/72E25VLkyTPl1sws0CuKv6vAeurfB5IAD68Jm+9ZU8ef2WUfPezc
A4eGc5GvuVrvW0koImwYlSoNQkiiX6aH0y6KbCvsKeg1eSBUGUNB7wNDSZ/gGr7hlmfERutyMrM4
WSW4QvFXK/MBI966y4UNeuXCoya7+0YSHlQoWwHEab4TWYRe5DRC9duQY8WJDQNUUOUquhdzSdbX
xxDnJCmZWco4MbnFufX6ID7WHEqowaxID7B79RIY4+BUWoqkYvNowK1fKMw8Gi8iYxW9Jjql74Ph
NnMTpKvcTBDE4W65BJDWHqk2B4mKAtb17Z4KNZdNA3MQEH30YV66hXrwrA7Bdl4ezqni/YyqgnbE
ofSxrt8uedCgDCxajAjhcig2Z/W7WkUTnqaxOuZyNukG45qb/DosvapE/KltAdNjJoZxiP9FEEoz
a1Y5uh+5BU3e0RwfmgNYK7rM0JG3x4seXvSogcb4sijIrEpnBnj2L1jFFSicYt4w9IP1CqlHCgMU
xdnEhNDPlcWm01dFhWjGgpVCh46837B5CNFYZ1KjubfFm6LxKbeZJgGKxZS8Ah65KbiaEy08NjAZ
N0Q9poFVBO+ulq6zh7BHaaHKqpYXy1Lm2BLw6um+MaNjrF6tl7duIfJ0BRmqasophTaB7wjEsGld
hdi7yLNlbbZuHroonpr/f5QBJX67qPEujp3kfLX4kGNGN7xe2dTehwTQJo+EbbKRQ36fp39LDwhY
LX89sjnE46L+yTcGhyc6LVLwiXiqtroWIWDFceXPRzfry78RqDw6dp9SXJcWsSsqcxl8TUEYbnyy
FldNxQnqmo48HM/JcKCv53QICVjOZUAs48EBJS3pryK5AGx1R+puo+Q5ggrbo0DBbZwu48Tr432H
MU6hjKbbf/5O/6ihZ0p5jLkkoudJaYIdDz2rFTUMM0U/bYtjXLFRZhbq8IwdTHRh5n1gNmwE49R2
8/jT5JwNV2Rnz112wViUnGKIUK0rnWnyy4cFXtsOAkj/mIb/BU5O0ypjgGHSlAnjuIOl6XzhiFKu
mYJCBvN6NxzBZQz+HK6XoUEmb4zMvXpFKFgzgtxOAgZkZAGMLCsoJl3qw0NlGdeKOYbCbFITYN8l
1r7GEN8gvp9RVPfmKPpjrTZdn0VnudqAWUS1IRPnIojI5HgQ13vdSeBbt/bWzFpA5xoyAUxvK92B
QgpZrvLrlviG8IEtKPw8LQRTVFhfoE8fApHgwv7IF+8Z/Hok9HDwOjWRKsUewPi9n1qAjWqExEm9
hFcanK3hjaDfRbm1Fk6o1TkvnaB9d4fZJ/bq7ECXHoYHYYMNVvUh2pfNPAneqAtyLooiNKLr8UDV
ohK+TE3pbtQqA7OwjLUf7Z0wQHKTLk1le3nMG89rD9RTeDIHySrsn4+G6n/8pYKG/yAH5aMwLQbZ
5Slf5Mr49ZNprKaywAubM0s5x32Cux9mEuBoOqZxXfgBCKoOhThxZw5j8Px/8d/h8zILoRTiXuZu
rFO5syHqRibE/THiaox55E8k8z8D14Tv2O/677axbpB/CSlakACm+UWkPzkk2l19Mb2z4oGtwmUv
wFYhYVho62R6D5fwCm3BjKBLm4hK1Ij+0zx/o/8cgDFnWh6M9v57ZT/2gJI8GQRy9bxjX0TLCaVT
R3llKL+D7iMUFJuuWKFw8RE/xdvHh6a6F3LlYjSfiARZmOMLPlb1qsrcKq52wUDRNr+X84byK5YK
KWN+W3OVXYjAVVJ+pFRIj402CXvYeeW1q2D2qm1TISdjzUsRp04v+gYMSKFMOZcRBeJsgM868Wa9
dJUgQo4lWK1AkcNaMWwWndxMWBdu5vLBQimVzE/1NuA0h/YHhjLaJPnONrKWjcxUl5Hd1NdOP+p+
OP9nnioV4N5zw40CjIKjA/CSxB6dlVKB74H/AKptDicLbsCbOLfOcD3X3e2cOFRwm2BqZY39izfh
7uWC/qX1zcycRHEWwiu+6WmXR81/8CCP2G6F81LMeikB5P4E9bRT+KdvyGgFdWJ5Yt+H91102uEu
uZM+zWlwG0fcrHFFs0N77/3ugxrHlHFt59Ky0RFMs2SZiCAxB5d1AD6ZZHzsbqaLfUM0BnUKrG6B
kmF4Qryan+JZWIHCzU/XBt0KjmDxdOea+a23t3bEH5iUYrcBHvTsE9DVPjeo0+LQDi6B/84NJ0VD
5T7A9CeXHrIrJWWRia8Os4BMXljSG/T4eG1DfrqrW0J+liPdvF2aycXuyzuva6aF9WseYE/uI0Dz
QHUa5gNr6F8AhUpPGGhkaFz6InEZC1d0+LpdRrvt0YYljbq9NvZDUgizbNEZkcD8cOGUenKeJDVf
62S1TCxyfeZeplwkqiv1odNo2nik5n5mET798xBIdp9K/qMfMTG06mitiZB+1cC81+P1EDtgK/zv
NAM0VglVUcHbcQOxPG8TONhY5OOPjCFMwATQfeURhberQmt+s4MNSaFhdPtV/sAQvlaiJtSWxDPL
jmyQSlx/u6UeGzMkZg2RFLTgOfHHl/EcKp72Bl6GXc+uczOwXWTces3MdiBGpNDrgRXtLmpj6W/I
4YlbXQnFM3u1mGKHJxHOMxgyXnjcIg/W68dt3474JQwvVSrqkwxY7NUGyXEj1tqGt/9wGubMyZQD
0H0MYgjFkGCKZfEqHC85/p7OwKCJDULbgUbJrqehoZWS4ucrY793z/LKSkgQfLcUj0w4dQL9h1kJ
3wpHmr7zZD0b6iajFoDjdMsYnQSmiia4viAfLV+b7/yLXGuNR4NinCo0CrbpDFiEzZaL0aTZgbLR
sw0Hb8xiviOQdQgZlrGHv7b2GFsKNDKl3dvpB8HPw1GP/I3rvysY7767hrBZHji0QzWW7UjWiehc
ogjWFht7qxvfgYCGx9NN2MjxAdGXRe6ODrwRqKPkHAlQhVc/VIk5hYghTknZDIymddzoDiS5o949
hE3ZwIMunSnxXFC2nD/rR5JMoiNfg5rztSczsQBsJKvAWpTOHKj8suHwx6v3Aa/v+4G1EcIYN26E
fdauanzyjcNkKnGWsVFXRE5sS1TnI0Jx8K1XClqeBp1j+3phFkzUiGI108WBmXWWB8gcbu/HSK2K
hd6i1o7snDPkH3ceByFs6dB6qfNGaWh/QGn7kyWY+PEKoqh1UJ9SzjVfTd+IuRo1Nqdw8q21/gGJ
uXxA8OYEuzoKlveL0SOmtvdcCbunUi74Dj8Qqp4flKZUT6NB3sBUEcGoPsH4fqwj+kkdTCCJ0Ptm
DJnx6ghM593ZDX5ctbkZMajuMgLVhTKEhAEHiSTYzdPW/pzGPjSPZtmrer5YcVPhijz0inyaCB3U
wS4hFaja9kqym96FPFceU3iLeRUPVjl2cR0n3et8Zws6ucF++P1m+KArqvf09pnHCqRUhUQ0xa0a
MkMIQqqP7+V0GVDIMkIL0fVGo2aBbly8KvyFYEF3jcCM0oqwO3TAs8mh2xR+G7qo7dlCRH2ert6A
3jX9oHVLNxGmod0+0R3Bc567XjGi+NKcKnTw9KC9risvGuDDK5Xx5/nMwRgEqD8wy8M3HHQ+Tzbq
inkU9reXFQquZxkHoD6kgi64FCOxTEgsO7vF5CnI43ufH1km4sflGhlgqQSYs75X8ciyFyh13R1T
Bxv/iYE5QMi9YCrhXu93/el6DT/FJW7yGYh5LicjfRIOzZhqRGZLkelq8MSxtnSFARTZANDgP4go
hhssexRAKzz7GVDVkZdg2jufqF9MWCJ86bfNNwh3iwz6Bfu/w0P4uTt3BAM1ei745D70RIhkK96X
r2HgsNFAiRr0xPNiDSaSscwEDK/wvAD6GcoTspzQO5fUyhN7NRd1dTL0ni5T/YuuiJRR7x4DpV5L
H6TeGnwRZrZaw8LDe9d8GX0g3cAn4CG1QM0oWXXDO0A756ZEOe2E65YSpwHlHo5U9jDnV1lKyuws
Td9IaQA+dOAir57Pq8tb0ovQVkf5SQhUp0fyhhPtIjk4rilCl32vDbE4xjJgzwcQSFjk/DRpWhJR
E9HUF3SOJ7otS6QCYRMNaFtY94RW+oEmQRufZjyvKzJw172XCWFAcjRzyGxr5Eet4IB3vyA9qSqH
uQlK+5O0jPbhzhuiHgTOilGcvg6ZWVLdDos6zeV+UhC1SCzqNnDxtD4/HkEdDTvNAvC2xlCD57hz
nA9HxsD9iwnQKUIKx/2p92XYtipHrl9Z15sY27QTWV5Ya8YJNC1CDY3OGmBArfOyjYXXJ6udhDrB
C3jJsxHjS0hxDuN5UZ3GhGHjSDWicX78hnK9jLyHVndxUJ7vC8tOwJQALlUwENbbZfVujMYYXkgS
//s/8NZzZq2xF8pqOPdbU7c7Q9bwLpX9NnGoFBQaNjbTdMJlNx0/1Y3AgiAcm/rNSSuCF/79eY3J
ionDh3A36Ey3n49i3B63Md+OCRr9ZPWFLAz2mQ1to1uiBBzgJLXPv+v0BjdUsDAokZiab9Fjv4uI
wteGAygry35cfm64Ww5fs/yZ1C7qvl+VHYtd8LQzbeQAwuuAHTcRa1zshTxNofgOrIKhoDTumVRU
pBwBmnpeiLNWnMaZbbOl6rfIHhh/aIsvLFPWVDE3q4GRtnARj7JXqhyS2Na4whNp9XdidlxfLYkF
4n2nlwQT4gOGY1k5HEZGm9feO8r7v9lR3dIcrIC4hgCaRKcEXvtUsgViX7hDltwqeqLo1laIk6De
yNY38GWc8GheqWteN+g/iWl2aRwyvDYqj8jbwwURZ3nao/d178EFvysIIQyEGQJ39plzaYQajRLb
BwI6Yr8Ye+CuDgQhbx9m6kxLfsDTkNjY9Pfzt5dqyKXeWrEUlneNFuCIL24OTiG+/6VcBr2xmopC
AyksYXp4J9dIDzmjfsTuC3BoL54qGMAqoaM34J0OHn0ZIhvykBsl//PNZ7uauAidbke5l/0zFwrM
MtpD6dm0NkcQYl+cEnwtp2Ft84mdVcGcMKvslKROUCKlcwpWcsXe4BX1F/nM3xwSm89EO1pGZ757
gZ6WwvEGQfwwcAr38KoN2r0+KHElKlhsp8S3W/bQE4UBzrP3fzct8EXGXNbEH3GLMmZp6/nIskcH
EzGAqJSKG8GPzN+vOTWvQNAmBetpG6dp6pjor+g3L4oputBkHHa796dBiFNpV5JFazVcwrijeuv2
Zjmq5Tm7NVSDOg11gnbQa7SnhsfnBBkBzgCmUVqp7SIOytxeJM8wbIR4YMPBINNXxLpqHl4+xg7S
1R5ETBt/fcP2WjgvsGQNBYWGZ0zYLUbRspS4cOrl3fT9IF/YsV74yATaKjDDnbS0KPhhD6sUPilG
vXGR+tYM17Oxs/GqociEGl7DiPtGU3dk13t5hPOxVSSQRhNa0ympfc6HdoV66y7apO4gNOQWwP9O
qfhwgKb1iQKvTGJ6OkSJB585G1J+CdAWLyygFHJYPBhwSZ5zdWUabtQ47xlWmHBDTa/zUfDg3O6o
yXaFcSjCrmMeDD9Z9M7nFHChINnbcMqlyrR+uHEZj4gVLwkJhpo4FybVYjJHxyJKN7izKrbHs0oU
auWZ8rfNkoSsz+CywffkWxM8NbJpOULdtWARuKQD88iwwr+gFeFswAVWjVURWaxIDYnKIkaVfCzh
J3wICra2aAPXc1AYRVtXwsT7lm3m1SBrXhjDZmpiH+QB6Y92nKmhd0Qw5hZNLMz5xCKAqLIHxeso
oHh7IYEupU/7UvJC29LrVMxL/iPyjiofPtr83/6PGPA9oaGeih5Qw3UXLwlE9UoKaelDUh0eR+hD
rAYkZJHmP8putPSfoc6QPSxLTb2ftNxfToLV87N2K/G5cEbjqS+/1BT648/CRdXDRkMCYOpQrqWk
K1EAeu5ZlBfnS+WGXNO/Ew+lO6HwMxWIuc6dBvDfQX+1U6PDa22qUTwU5n2HXvOvZjRhgbmFKjGo
n6Ht5tM+vRLbU+lOVuXrYiSVFUsSLTVP5K3/cVWfniv2o4Ft4twzwr+3t5HrfEzjBaJJpnvvRDgE
kW3MXYcz/wfJV5tIgqROCiz0H4E6hj4lg6hJPHBF1X5NsaAaZ06DuD2S2aJiB5sM3vk3sksbKTbR
d0drBkyRIEfENxdytIRHoAYn0dwciD1dSHk7ZYZQQbrqiP2E1muxN4eJ6eD/a1kK67akOetaA66C
A+P43YoihzdQb/WBmhQ4c4Z4zhX9lHwelFDmCI2540NCzjaoXjMAztP3howSDLOJcscLZW0/72gG
sWnsteqDotzej/NJmVrDcW0sUBS8q2dHOTEsdINIuOxfkU0M7Z6gCckrpG9iy8S54qajQ7W9jWAB
JF70vQO8WUmkhRizzqKRKgwVFe3KUIHsvYFtM6vJrlQ3yhK/erEwSNUDi28T7MsperelUF6VFCOJ
uViPtTue1IPWI7rDAhHdvUK3eTyr7NZ/29pCfh9PhVhuS872Ej4PzhJtBNU/bi9Sgi7lJp7Mr88+
0JOwKGnwbK5XPSIRNGZUlxdiKCHt9xBtQmLohB0IoU82u4Dfu7czL6UWYk9efsGUkk+jEiJCH/L0
dvO37jSEXU2rho9mxH2p85m9CrphyfsQg4FOVm36xvoAgJ6qxCBoLr1H96rTk0+/wODWwjqTqY8o
fvcK5cbXlzcwa454TVgdk1VgZDhJmYLdPIr3fCgaemWKGsX05DjMlP34rnpkOXsiOJS6j8BhyORT
Wxj4WX7DWnA5eHEKHfCu1n+z4dEI6MAmi2CBnari+FatXtDdfkB4VKxmO2aJXnerT/PJGUUrorrG
Y6kytKNx8EJk8E0vxHbGeQVPRUBIVgQHdxLAfX2QuQg1UmP6fmia541dCi9flapjd2JVVmGF6ggX
jE5UsonqP3/85YnOyUROE3yXYaamrAWLq+eRpTLQjG50X3sYgbu3ESbvwjtAD7v38yCHI+CF/9Xf
sEhqnx79EPKBtXdfhyroXTx7KOrkWPWVboa79ae3ZHljls2tgMzgQPJbdsJdndQXVMNBuRj+EGiY
plSsPcMi7ZfIXm4Z/WmyplpbS9hFqBBEY0HEtEjZzqYqkzEn49vPiwNcLhNVYS0WzAVEq1uAEatY
zEi6NKlfv07r7fMQxgIroNTsBhC5DbBucLeLFAn4oA8OlarYDCKKlz8n9Iu9vCkhRlEkXgcUxnXY
SpjKIWG078ZeU3d7NbJ8aTsVLiotF1V3b68WJF2dDLBFAzPgevDIr1l3ew61qlJFxMQkANiAMp6x
mG4kcwdDUUq5FhLW1yONfrDv6FbSphzjYmpjuY7uUTaNw2kwvYrcnZztwJFknA8gIQkPaXPoj66b
3Kov1VEPgOwWeIK+7qL9bu/5fBtKGY7Psh73fiupx24U/QuyIVdhFTEEB4pDq4aNIeoM1w==
`protect end_protected
