`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21472)
`protect data_block
td5QFuuLITbKOtkE3oI0mGg81uxEpl4OzFN3dx3S1ftkr1FB28AsEjJ1JzlMER3jugQ0XxNHpZ6B
MQSg9LCC2ub5LNwlhvbYEAYYqCK6ZgIfuBIOXcuFFCv38YT5eHX9DfFv82XjsC1Pwn/wMP5pa47z
RkUFjUxny26VVLkcvVGgbXqytVTR0La1xotifeEjVydMrmZYXl4iOFvRKQR/0EgKCt57YTzbnIky
JLh6DJGnFSWystzWEN9m+rQ9crfQxmwyJpBFPQ1QII2LokmEvRvosXL5x6beIuBaCOKFsx0OiJz9
Fg4/beWAucsxlrFBfY/gzEkeEt5K/rjVYPngc4Ri0EFvyyEvbMTir4tc8QjEOnn9jRDkcf/RS36Y
ET0rvaIgmsWQK48R53jYh0rnb4crHhyLle/Ld6omDaWj/Xc5XOaz7Yz+sXCm0nrOX+sXMiBfcHEx
TEO1mvpCCwn5Ok+cna2VCI713hpjMb15nBwhM+WoRwyBnqoe5vDKSrQjaVTuWrY2fmHYY68kaTt4
xpCVojqKrWy7a+Wamu1mLLgiwdDsDUp6PYRObD8mJ8yNnRXCxYEDjTYwzNvwRyrh01T5LLpJqoAU
sbw/DUe18Jk8+2esJjmEp5zF9PntzGnMXA9+Fvu/mFahWHYm3bdAKTbe5ela8KxKQPqUHsgyQM15
EnhwMs8hnDjruyhXcCN2lHx3DukmuLXdqsrZICknWiaqWHUu99PPdhun03ATDEtu++uKQzw0sW09
64H6tdsC94v7nsQDL5JTFQqvsJCDcgqSS0n8mtSh0BeDXUI5mQe9umSEdBYNNA6BxUtHk9iTOOq5
nBkxTVY74Q6qr9lYZb94esrUFHy7pAYNw6r9uqSAWHq+oUwopvBh+pGHDI06L2Oj/Jtap+BUfHsU
GqdxBdAo1DfPL3XcZlxzJnc8uywtdTILhafZn/UwT8nK+LeSCbCmzTn0oRagUB7RgwZOmpOWvV6l
BwrNUBDfWk1f/ME8J5g+j4FPYi13d5gGlNil4ZE0mKQE1W5dHoe4+h/JYQxBwYHw4ovf3J6NwZYm
fpdzNj7YR7ClMGtgHhVngXMdbXuI2RTgvpJEUcazZzUaBmtq1o4HDItWBAZSHE0cVJ245qMiB4BW
/3BFsKtO324KIUVUgJiRDgMOI/4ZuqtQJRNrI5bPkv4u2Ot7nKBrYaXsZ83Zcyc2Ia+MZQfGNyCV
xeVhpStbJLmk/1gpRMqA0tJ1BDg+7KBCYdbqIT/g7PaIXk0x5eHwv86wdj4cMn0b5eGMF0whx57h
Ofkg1KV+Y8Z1GfYG0v668LTF9lOIRxP6w8+kfVBYM4vBL2b7cMiRYknhjD0x2PUx6iGZL7yL5d2D
PkIhLbsNMJV9eNZHNUjeUP7jEVQNLjfqdBhmivvB/lpv9bhgPvTfDyxXO8gsI93LHdC7QKaULDZg
IvbptKSnk+7ZZFBpRQR14KgoB8KtZZ1WYVDQaTOG/JNW1aKr76M6wgqTJjdsR4S5xu2fZoddBIge
xDLtAloZ2bLorOMs0WRXHe0/H+jER0cA+zouuV9x2PUF5VeDVeaCloQ4vpT9UOo4wwVmGoJD89VD
iPWQsLEjyWhiobmwvic+xZZu2HAwFDYhsbplu156fr/tvRbxOpaRHyUp7aGO2hT5o9ozgIH92AAx
ujHnIgCzONa1i5y6WmhDPjc5c74YRxJe1c6E2l1obKOXvrfdVpmnXazOiqiloEP6lU7VBEoSK7sg
1GBH8m4zZaLT3wrUOCZit9bA1gLJYRRC6GIOzJMlqsVEW37m9bGoEZI2yRjt26UJak74AmZvzNPG
lZinFl+r552cMJptP2oiVF+CYiR2Z06PNX/+ylaLN0Kdl3mylfcqSrKGhYn+w6HdoSLh7UmJH5Lx
z4FA2bZF1wjsKRYP+8j2MUPu4suN2OZ/idT7ORCiG0L8dyZVniCTeKioH7FN5NNk+R7infm5RUIv
+YPBkd5pxTYqrbWfBxG3AYDg8tzlrAUletO0pKL8sA8TA+Tg4GcOLI+u3NJ6vXoevXrVEdGIhwL0
nJZquKUPzHPSWaYlrOiTGHtp6bu4cvcfNJa5Gx82YDV3mHX1UIPsy68odnhhzHf+5AxVclQO2TDo
JON/knNhKALNy8aHdNJV1Pl5GwY4U49xY3+Z3AoAwxn9z3GwLJbGgSLUEFFFb9AKnE8QEGy76OSf
3YohxSpvLynF7FADJXIbXOjfR8NCqXHlmZ/FCLvUFRT8BG+QtGDAQR3Kv9XGECWw31lmhtE1ch96
gSoz2rnFpee3G7OslLRAQsfIHrzOJ9hqA4Nuih445q3DlQhEQ0EfbdYcmwTbMVR47lsjZHt6WzF/
M7DZD5Qo5kMAzrCgpfTfJHGIGXEOhjk9108zSckoDBgDSyFyzneHjxZvLD+g8i34s4muAMnexZKv
S3vb9sIfjhYCbVjHoF8eRwikZoYvtZl48DsPqnZ/Vc/q0EPFGUt5Pe4ZUJAe9BsPJRXWOFhceR4t
QauH4t/phDuuFzvexGNJ2DPcZmn9d/9tKk/H/JyfNiQwjg+rfXdknqzdkdyNCuMjTZ9esKiPTCQO
y73apM+iWRHHD4+FHaRuTZf9fiahWaz8O68wG+dqOOuLqbbQPux7c7ZR1iFR8Os9CiY1lPfkk3Ia
+CoZW0ThoXMJFowQrFHFdhOqSpJE+1hceQ18kQE6Gtu8OgL/iuArj+2ebqEwT8d0XRYUDr0Evi16
A9fzcb0WPmHHnNYzvB3X4aIlYVeNnej620gFYFsJKmzFK0oO7duGZjkQHisSzgQjcpzeApJEDD3M
TzzTMXG5X16IavxWzZ7N22nCPsnqXVOEhFrRPAJgEdqiiBd91M4ImsDMDdgzG07+syrbdkjyAKRH
sNBj6tBUMj61rbZl3J1ei0UaB58LcV7yywxqICg77PuSYOT4DoJNMjLX++dRVIZKOwwniIHBIj90
5MaZ/mxZiLECrHzZ1FmivVZ764O3/Xx0EKBfpnScjuUBnCmWoVTIesUp7BFhZ3du1I1wl9TTAyrc
khww4z0ZzsFigGvyXQuyusG614X7uAgq4BoqF+xhEm52GQx9yD9WCsYV8nmlgBKCSep+be4N8xfC
4y84hStLX2kC1p/DTOFpN+bcxJqCTwVpCQjYomp4JenTcXtqnV9DCex61yhQl9agW7NWcvS+0ccs
tdZN20eqMssptd51kMPs+80SiqSjQ5Ry1RjYNxRmM89dmVtV2qRhhjFrjo1m7qfPUBBPwJWw//Q6
NSlOiMKSn1Bvp5MYEB10rSmNBaeQSA2vek8hbelZv88HilLAH3jyKKZgEY93SqZdlwPJx2zBk0cD
rqH6hNKMIhJMEYRA+XzrBEbjo7Dg3ZbOXD8Oa4P/oTw8rLWc4ux33AS8mp4au5HvSETYoPQiryaU
zNkMMA46IWH6Dgll0Yb9PIS2A939B3/fqlh1NZC6TUD1pByldTVFxgQdm0EAZTh0p9X1pXFpiweT
nnsio46quR5HNQ1mHFo9Qyhe8TNZWnPMphrvbQOxSb/S0aryUPmyZ4EGN0UvUxu/6wdKr9P9/eyw
jygMn25Kk/az9xqlLFgjDQM3zAw4KRAAOgvegld9xsglZELhQLyhREEBDL42Ea6CFPmw2HYb7YLc
z6sobtIGdfg0FqcxvoDc1mVgtYJaJH4ZwYwYt+/M0FJfZpuHVAopv3N92IJ0SgT8tZ7mBo8MJ4xl
R8rGR5lGaOSxz3HizMyDI+Bhn/EcE6/+HrKt7e9zDKZd9n7S6zlCkEkFoa0vDCJszVH0xbjI2IGz
vgkMKsrbCJ473wkrZbBCteI3ZI9ng8qejm4F0vbk4XuhC+Yq3+TJcBWikqkp4iuU03VoDveffmhU
+wylefTQHMkZvZ8ov6u6M9iKULlXXmw8XUv0cz+IFaU15a1yaHgvYVKpI0aNslGH0HwwkIvWhO1t
y/pr/sR5kRWUaBKRGIwjnPL3wRjL4MvypOd3usEv46AB2vVfI1/V8t0oZvCmM+pXGKlyT+JaD2DW
lUw2Db9+dgR8VnNXVqeslwxxzLepcjwMrALpOgsxcsUTwJ6QDttTquglkwYpU1MCL5IGIs93GW4G
2sqPQqodIHtkfx6D5qG8LriMwmNDeLYzMzR6IlHt2b0SAnYFQNDb6Xg8cszk1hNRrX+wOGFleohD
KT+akCLxKkWvZpo1OKXxTM0Ta9d7GEfOiXjiGS56q4E/uxB25IVI6aowllXGybQG5oq2kySr8UB9
eGFv+wBlN9Des5U2SV2zEVAjYpbwHnvbYzMQolWkDomG7qc8Fo/Z7/BJxC6OhkfuSMFMJGGqk0CV
v8clO5n/EQXjnRPIGzRZB/RysG9Jt+mB+s3Acs+r+uPjrARNvMvv+rKy9dTIgFDiKbWw7bXRhGUM
SdvAmqKj8pAXkB5bj7pzhrm2uJ1/Q0GlIqTc56xnrNuQPHrB/Kr1zDavwz3gAbLikrbgkMqtBR6X
0+y9m+fE8A4LlSLVNu9xbOseeBEu2k+C3Sz82LW8A0Rk7A4p1rF7EGsm+GVYIF3ZN6NXsrHjpApJ
FFebhcpwbUAt+SXHSEIGUgXqhUfmuoe2Z7cpPEGV3IAzNjPH1TzxXFZ02AjsN5QntN/4EOeIIjvG
UCGAS4uz1AcmNK842DvPxLa2SHl55LvYQ/0ch/TRPwGdMjSPF0lNp00vUR0ZYCiLXohMEKORtjWf
9BysfSewxCg1D9b7qnSx023WMSd5oFRZefUN7tL7oy6dKdEvoBDeBWkLmCajs4bTFSqJGdQw5lsk
63N9oH94czC99rMQRMCy/BLVK0ABb1qNcEzxYQ6tVTWhYAG8IqdDOvloi0Xf7p6a3PRILVKHFjFB
u5jyq7iRl+kODaKt88gLFxxntxall2HxzmRRskd5ZX5v9Th4cKycaaA4/6WAPNNBOfvtsImSCURR
vWK4gRp7X40JoIXdTiJZdWfELHQlNhZLaczkhY8qIvc56NWnnzOa2kRAnnT1y5tu6ojr27bXTBk2
V7jnXeSODyCNwUZn2L/dI/BLd0Dwe3aHJBaWTax/6KyXJrY+OTfBpTq99UsGQhmw5uUnczqRPVIA
jpoD6Zt1+iu6ztE82a7YVghHbtFhym/b5Y8IaAwRSqld45iuJqIsl+Y0UArCjZmNSwKk83gP4X3v
ROHYJ1KYYZlqrYe7yJYAuM1t3lkxVlGviZvnMEYalPh2l5cMTUygjM1qOYNlMboXrDU7vFcx6LYl
ryYRMH5JOou+iNZjmixDzxdL2JE/+rS+db/L45wLNl+mW9ARNn1V/tuaeQSlOJa0v7y8NiegCJ4K
GmAi51nWwo6I9UflQb7mwg2Gx8GWpTu+QoWHtCqx3kzHP3q7awX+4ioMLrNqyXM0TiyqDv2ASGke
NEyCLLjVNO8qzigbWKb7zeNuMf0u1DDjOiNsw8H5Dbdxsi78YzXsSh7nrKCgSKEBruORMpOWrYCz
Egq6Koq7zOXX+fZRtCEL4Zsn/P0Wn/AzYx8FZMFHDVFoC0sE8ukgbaL0r9IGwC9wwcqHBkm+8HRD
shXoh6KZ2owH00xd+tyRMdypRDYN0/DIftWM3wAxk6lkE0iwKEtL7giSTcVOeE+cyW0BfZK7V97p
4U1eflzrk/ZSCwE76cD7VZtRoxr0LHpSQw9ZhE58K/MtUPEoeoS4nG8fwYX+Pu1UtHxCtulCfcO6
WQX62uTl/+Iq7oCtwTbbDSyqW+cwDGHyyt/jMR/7JEyhKn+XcRhu9QHELQI9t5vpZHR2RtuZVEmZ
Imrqm6U5Str4KbiWXAEt/1pv16nhBTld10in3Pgaf2wrRUndgG1QSoyaKde195Ks0gWLG92YVKIZ
O7Up/P3A9d7gvV8QpdcMK6ePc2Senqqq6FTIH/RnfEsyvms4kahMCammr92erDZr76H0MJLM7pKY
AVzfWDCqBf9uDIq3fmRkqSYmerWcyTnjeoj3BJaQqWP1rEoXNH48u7TWbTW8RbV2GTVMRrqgvEsE
FVQEPlLEicpwWeYhNur8W07diUxuTIEiqaORDs6dPArNbZVaqqCOPnbDn4ZBKYK5gsrJw2G1+0a0
Gls8NVbOdSrN0XVneoB3HADsN/2XaOXqIUtoqi0FXHuhUCXWkWQ6d05oXNGUE1At0lb45jT7Pf6u
DNhiRtgngPutXhOLtUPquHF323dGH56ZCLEFTq8KYZx2YSo/xAc4dz9CICTAoQTTwev23gRnhw7p
pt0+qnOvG+reT9LB75iK/MeK7Z6J9ZwiaPJog520/1vt1ibaPwLw0x1CIqVs+jA7UR4riYHhKMP+
0sylgg1V/f+y1Q7Tq9SmiBsGUku//pJfDY2Wk1bJSw6oD8o/rJjtB2MJYeNf4UlbXZiz0YCSEGlg
PMMKDqjUVfdWQ/5mjGvFSbS4e6yaC3yr48E3t9CKZ/ltZyYmbreudNK1m42gSnSbKvVU8hWAFzEy
9EmxVJrbf2pQGM1K9Zb6aoQcjwcZk4XPqAMOnpgKiBVSUCvvEtkQZRHv+gGa83MCjV8QUkgw5l3m
SFX7fBE3E2K6iva53X7KenLNqy3Qbttg3E3GqlZO6o3BKlRvDPlAkDJ7eswhuksVBhiG4P+vFw29
y06UnFhJDMRrlzSlSvBB194rGLC+IVCQV6HTqhrx+tb6at4fUYNgWX+Gao9cVQLdB+cm8hwTSkhE
QmrBdIy7z1zpOrU1aZeJBWF8WKyocxBQ4NSCA2LWc/xLzvHS7gkEIOfiUI6KxCI6ZI2Ay7LJ/Guc
pDWU9yAuxRMYoQCUKidueWaEO3cq0rp/Xs8MDGC2vLhILhdZJ2F+ka7q0kiYFsLWCTmZxtmA6QFw
A5g5JPIsW8/0jUqaTHPsKFS68P5DyPvXhA77PjNN3Wg4H1tB4wwlt9CJiVcH5C1xiD2yvamMcfJU
RT/Qe2N3SBKYpKn55Rt8j6Pw/VIAFw+N0r3fTsnFnsk1jcIi/bl7zcmX9zoRfyVRyxawPkXA56jU
fNj9hjBRFv2pHxJKLtozIL8x7TDKpJZj41xstkOIMHWYr2HneWlFlBPBxcjrhKaHXqBAHZ9ybPzK
OBcREIBxSs/a2ce8ozXM+mj4Q8vRMW9bIgko4IAl3gl0s2qrm3irqpl3sfPnNF2fzwsLf+cPy7+V
0fqHWw9g4sOwnT0sThjgZw+MPDaI+nRrIV05B0/2Mgo+a7bs5EmybEwS3SMI0fU6U+c2nCVsLDbY
k2SnkzWlawDYR0Xmjp2jjd/kYgjyGk0LU1XgQgMU/sMyjecZRnQ2LVkZ4PPF/i7NaxJOZfdqgR0j
rAgz07YdMXn6DefvyRRFotkRgTJ1yAVhNzcZDpazSVIGzWwqxtrzFvofe60mACD6PtCsBXXEhSPm
GKJElENIh5t4fEgY1sU1K95H6ec6XY2tN5jAXxMAzM/rpENyPWswi0PhOjietuHXhF6yb1ZOBWYp
QexF7XIat1GHrKYqe/qwzv9o4uiQ2RBjFWqbgamtWpL6KxGq10Zk74HNd66/JbZYf90TWhd9aBnk
0h5mQlIuKJtyKvJP7wEiPjUMvwa/uqTBv0JX8fcKK4yDVjulWQnbpyl34CVp/wSqXEZhyNuBEUW5
eCreXe4Uw8OKaiWbBj7GTnm+NlWvFPuT+a/K7sxXy4QgQhGvJo8QRyh1DQAX82HsyVJVWU+N0cFk
UxD3EPc225h0Zi7zc3w1GYKG2i1GA2XK9eXbWHtnfmzHBcqeLUIs65LlwncziL3vb5ebPYDQqcD4
chlU4rQBx+6IZfJ+39H3pigU/sLRO9nWTVWOHeZ7b87zkZoNUK/blvwQyzAk1XPThKuFFTM04BZf
WMt/je+RJm3uRoUXXCsbFDQf20Qa+C6/cbrFnKj9K52M72TE4K+zXDnZ4PhRVScPz+G6WpVArBTx
D5LQjBCUCkJRU1koNZpqz5jJbpExxiG7b6kKECv4wx6MSYLKAbo33EUzFxdYRbAHYEszDEP9OpYm
2VhKueLzSmQH7/LjwYuNFe0iHEg8EclvX/6Z+sBjfTt7WXPZ6407/0AIVB65uyEenfY8SGGFRJBy
l1R9d3hHJgA+vjk3rN8sQSx4MyeRO/PcJdnwMSp1yGkh37DpyaCAEdZEUqi7SjgtcdxxS2T3c9gb
NdCzwxq6VTUZShzTULGmKvKEzuL4EWlvIF2zUnbiigsnHf/OOt2SEQGBSKOjuCeQwKuCRWAi1vUC
7twFDXracC55Yc+RLLtGGqrnZj+H7em2o0ULme69yhHGolTHNYyOmZpHms32onVFcHXdXtlozSHg
31fD/BFEZblLFlgpVvT+fc4wDCn6UgNlBpfTISS41FliztxIOsigb117VSlSZfF149GoQd77VjFz
NEfW37JvWi5KxffUBog8lIp5d1QNCQiN5HLlOJXjIEyJmQO0BAeURdHV4V3BbnfhhDpaCfAx420V
49MH3OX/+OjnFr9Ifkl+dJidwiP1P5ow6/SNtSLscAEIbGzM10onvr9IcMdrLuXAtfG1S33g5eMz
Pj+WiAxHMkHpjtQfD5LZfz9ua0rDCuGTbhU3SlcbwukzyEBk3C/BlTo3zfWTdU+4Mv1H9rhY1AsO
BgsaYGM1KpSUq0dS/G2w600vIXmQYE+gtkYFrdsit95PhcdVvJ4zZRgdUqW4eAsVEhqTmhUCuTO9
vDBww5+qeb8Y2+rCJ5uRVhTld1v5c7yaLFSdkiO9vrpHu4go/ypDZCrGG7F1xa6/rXL57KMht1I/
H6CnMHw4uhpzKy1n7NorPs3+UmmedZPZVy2L7VCa97abJ8qLJhC2+5r9Y4jvZhuIyRqKi2DjsJ4e
YVyikdEvpUR0EelEX//KCA4YnGqan3ldiFxgwH0OIfSyZfBrdgsR89LFZIzplbqVRSsft3x8JyFe
j8v5A0A4hQN48TprLs5ht4GE4Fs1TflRrh542RvmD2seXhpAgbFufxUhZSLI2VlsNzO3RLROi1Qi
NhAq6CDCEt4KR/tkGPsxARKlLzzVpakCKI20sZa9QZkgMRtJMqnURzgS4t+2OhcRxMp9UKTYKjB2
gKjxgGRuiDupmvtrH22Y/5QvIFwV/b9g2bIFCkEGFyqFA349Jqw5r5X1o9YnqLPk37Y0wAsJejge
08krWcszraNEj7Ilp9ZrCc5NXj8KC/+oNVhRIFzApV8G8YfdBK9gixzLonnYIru1jMOrzoM2k1a2
/1q8ir0/CsPTsWR+Jc3oS6WmnyLzhHJmo0GJQULzcL39Cp4yuE1QoAIhLPO7AgwTfWw1Tq3cJ+3A
qrIVqPMRVEG/Kr81hfz8v/1T1kvPQJOTx45OGwjXEVRBBsF0LBVf5G5yOLuJr8P6AfKDir00U9Hp
n5ECxyoT7BlTkSNjeagBTSRZuYS6q/gT1qKGxjtZaJGx/mVS6f1bxnQoJqpoTFKdsMhl+xEGsDgr
BTvReP3kOEoCvN4Y5g6BgUEqr5eoWmy1r+vF0VfshrENy4D2zR6sPQIHjojchhpF9N6YsIy3kDE/
CPTHpriYDbjVvxQdzS96aMz3bLz6w1hfLZemIlJkKQYuhUHl68OuMnkHhqcFjuVj5Fgzju49NO5X
P9cuWyRl4EDgYGyUfgQYUqmTQEDCwwPrXgGeNy9mcNdi25JFC7jOaEta5iYumJ91NyM7p/FKIItb
f0hf/2CWvuE8pAW38EM9bQi4NSOdz+tbxaKYH/+QdgZLUHoD0+2wqNrWGX4v5gNYqU3hDYKBaWc6
Kfrsanz0BHzlQti2PMiRfUNGV7yPVGd8owNm2reWL4CZqLRhQs6v1ds7Cqbzg4OOYk9/oqBynv5o
nIIwFQ81U8KfBktcClfbAs9CVJUf4OER1So25CLw+Z/0FP4mtbHNFt/KG2lkPRep+/69/lx0KNjq
OosqMuvBaPxr1z0WnHAXC+FtyMXGouuE3mApED/5OqpV+QJV2gj3KaCaq6WhYk0fDCDL76JsccNj
nPt/XMcrGML6+8vPC1nUsAWgg1SZk6kO0/zimODo5ZhpRysfI0auSVCvMt34C5FB5XjZQkKyj5Ti
984nr2TcPwkTmv2eQEP+Pdllc/rNPy/B68+g4l9ky/Ea04x7CWbclTukkOPD3EP7RefZq30N+tmQ
yXAVlwH2qdvA56s2VEZ+/CvKFRWVRJxlAEln4n6Jf1Qu0aIZMz+dFynuaqdvrgcLZbOcHRtOr4nc
9pX6u7NxvPU8Ws3O84GGM8nasRQivg1UfYX4uYv/LkcGMVMBKg7REd3eQr+XnOX7A3LlIrvZjuN4
kt1Q18fyj6uVDEv+GwE7MUutkLskneghinEj04F4tWIOtMidurHFLX+R2wntVbz75qsS/LR+lCgA
CmnmsEXHhfSzsvcQK/9K82mcHtTHDEwEYi8sV2pgwSixNhjNMNJASlt+sfFXommDLQ6gXwIRexj/
s38H+McnV9CVzo+XpxH0lzhMjLX17hWtPst7YKQ7AYzJpI1vKq6QSFuQfPT2MiAW6pfpUPy13yFf
A3xAfSbAPMqBOylaOueDH9Ks9FCWe+n8jvYmkRi4tFt+SFe+z36zCIbUApYhODbCyhJQxPz4miAj
RyopKdxLDJOdRxTrFoFcGOPpd+rPdwx4Ll0dwpryI4UPdapM67aKiqaCx/lTWQz2mwtC+acyHQvd
94GV6Pvcqdz4njYV/qLYA7c8F45UUZpymoTVHFV7SBstFrjyG1zS+n6dHjl0xEKwNiXGcJu+ixIp
9Sn8nyxWjvFoRzLYYo0oMf3n4Xe4Tn54IHjgj5WIq1XxvIy3V4uyCyyjOKf2m90bvUV7coslupkS
hzPc+irKrLk/0r+XhAV0QE16p4zFroXeKWDsonbY0Lz2k74KnVzO33TMqXzJI9PWqxP8kuZRLNH4
aJDGnQNKlcnZm2n8EPqb0n/ctavTPa8X9k/7FuyteUobe7FzxWKw3SNmpltZUZX/CRpBD6Otpknm
QPqcD3JpjLzzKr8Z9v+n+6b9cyCgu5yxuIWouM2v7QRcOTaynvS/CCU2+2B7tZjYUlWp9IGGy/Wy
msg+KR+b5tLYdADJWAlFH5IvyucQEBjjgmtg8fegsMqgH8sk68YxNXTk1nSb3hrpfTt4I3grnusn
5gdJrBAA2eMYsmUlVOlcs1cs7AvaXnj7cTIPYo6ONYD/Vej6XD3AMtpRUw/AZGomYG+T70xGtJua
ItjZQ7N8WQLA2R8ECrx5kWDwRx2Ha+spDvz7kEfcGFJjBTiK9LiG+/M5lst4yf0UaFHgwgBQOYbM
+QMTN943Fj/joQkJE4l9tRBv4/40C7woEQhc4AOvocA9P8PuPOKw+zkZU9HIUnrVm4cXgoJtmHI4
yV+D0tGVMn6rZi5Fkv1w/xlZekl+7JeFlOR/11JVx1KB68Zen9lgywvLMAEk2d9jn6NZzqiwZMtn
A6uv08K7Sz4xSzPBsHp4PdgInhI9sm2ltHNWiCJ0GJioUS0Dn5d9bd962ajGelkbdC8guoMZBEOj
13xLEyObFs8oVkvjiEc/Jkk1HohZLSeHmPBcrmF8vNdC/EXG37dAWBJVBRxWiD6ynvtm0fMUE5rX
1kK4DaADeNkd/DTWZxRUyMMjBQR4hBhXtl+lJf2RnqA057KuYMTptT2njx/Ih1hJTzestwPESXxn
0u96eTvWxAVFwk9emBJWrEQiIAuz5OlMyEcO8GPOp+lqRYL9m2t2UT+HuhvXD6v7ZJDEX4chIq5z
w2HgxSCyHH1mJ73jxHg88acuFxMEgqja3jXD1IcJqMt8MHliWsyCf8YUX4god1xKuMovVHFRE0Hv
2+x4Aaf1SkvAVKM2FfpmT7ddOMnX6I+mjlreg3AwV+f/u8KE0Z8wa7oLY1EIcsNQqcNElg9Sbn+y
sH/91FjxEELKyiLgBBAGs0JxP94DKiMdBAcqwwqHMf3zxtGkGOQI58r+EUuhtCIIUOaDALSmtDC+
CQUBo6HSBJ+0hNrt23XKwp7E3XaIbYPcJEMPAFzXrlg1qLoHrb/TzMLr7SdaB2+Xv3R9YSBWDmhc
Ca0iSXp+MTrSC8VAGwbK54jH5Dg+L3/HjLEqXGzxbxUN+TPXPkv9qqVHjrF7kMIHoQwW3i0L5JsJ
QFVNh8QuqjyVGtUF6zki7x1TFM0Z8LWcw0Jfl8UP1ZB+v7Z9cgSJoOb7YgFi4pavNQPAacI4fRby
C8juJNlVqbYFzXh4ciQcdqcLAmT6lvLC+YD8UROxsNtl0EIsakUEv+4R2WgSY7aZnZItHqUm2GI0
FEhXSiwYFJ2mlomvFg/VsagBYCibdomSD6/U4fcth4OJEzgJu2wAjtwDXlL45xMlgbniIkMjk1Q+
K24etMwd+ghabGpe6mUYHLEcJOqtrTWd1xAS+DOaW4Ot0Jt49Kp+kmzYfuskGZgYsnB1T3zqvRna
bOstpcF+K45ddes3Mr85Kz2JQfIU0fL3THMaH7f+nhrT3rF8/UBMdFw8pzjOiHafjSqE6Uh1DqOk
1Woeg8tgf/cr3ZUfVr6Bm/v812jIyGCneVXshgD7OoasdECJx37fGnfIZ2GTdWaN9Ccx6CLOHcE5
yDv2Kgqgqlm5XVLvQ7W8inKFovAV1G2/sXLzoT490+KJr475s7EwnKy72vxDEd7Ce5/dcY655l1H
iuWuQF/hhLDjw0zPvtxJiJ4oc7aot/iVH4vLSASYeySHL0MorZSt/FUdWUKS9xlwWHyGum4btSva
HoMvrwrNMv5zMVc4o0Ano1Byjn//nmMdF+Qdanp7ZIKFZfK8IRkiz/OBN+L+00bjiikE2gf8qzMc
PgUfZWpBb3SxpbPZ/Tuz38hdsnpZdfZsa9AdeQkeBxRI4g3X6/m1//c+T0ESSQ+Gxw9SjuWzRBz8
RcVjjArhNKcLN8nVzuwFSRDFLOXgAYG7VTxj4JlM8SClA5w422Ww2Bx7+1Blq30wFD3aVxBMufzx
HzQ04vof2Xo0y7K4dRvy6RFjr+KmEb++hCAPVojElL9K2JMf+MhcCwJ/pb8YB5JdVU4xtUzsjCPK
TQK6/amm9ilsFUJEgux+EL1/S/z3GnHTViTlgoXFHCi5J7qqkkxCwLdUpmsAj5QCZwn/aWcPpbo8
ctkZDYfUMVpSDCNR096SWvyUV1P3Ure78FJWG9211uMF8vmJEZNAJC+t1O98bog/PTMKMy/+XWM1
nVCKvdiW25Ses175fIQ6il8hEEPlrtZm16nuLxJgHro+y396qk1EECl3BGILGW2dlqElSzkOFJLJ
rDMn+b+BM71ajTkWrRs1u3jawgVWx+K6J2Nj/tnssJ6kjixyKs1bNj0Jdybr+mC8QC+urBgi0bZb
f9d0S7SD/1pHgDljSsB8g6CitpQRxwAzT/8P9uUlSR/m16p/eMHcbIoYA1hjtYHJZUAUqPi88dG/
sYZiQ2aTRx8HBqOFG40bt6qX/REyUBFEacVlDRaDT8OiNNiKb8mLBNNfOtRXaD8MKU4uTmTFWWQy
zDtIZUPR+5omag+4ulxxP7JLmZIZyNuoWd85iISMf1aKF78kIs9wllKEkYUW/1IpDlj4e4keNAbL
N5H3LWK+/q/SMWH5IzeubIYtUBgS6I5y0il5mGB+K+JDm7taSX6+neexeTWJLbBgRj3bZoalaDbP
bBdg+sLFquSOgKdOlUGevwx+W78fwLFMUp2B9MY6SY5ONtGM+zRQU9IiP31kKKCJC7b6gfGbMNRB
k61NaB3nLiWKxEkLeL58hvP6Ekt1KDUvTinjgoCCHroafmQkmRrnt4VidLSJHfpaQmBgCSHRXgdf
/3OvAViwiWqxlIXlQHS+U6oRFroCM866L+fdODbao4lieikj+d120StBTYQZX5pCOWghqfeaTWQH
z7Ep9YXqqUNEMh6ix1aYYd2LGw52F+K+A8lmTClmcO8ScJzHLSCkxEu/+PesfB1x89ZekSs/c5R8
PbsxHeAUmbQ8yTP18m4zi/5qCIeSMA2fwKwupqH7J+mqx5aAgxqhpBkTxf/ProlhT0p6hjy9aiCG
Z2+Vml4lEtoEb531hm6Q5KjGSTWBuzD2V3dFQm0k2t2b8heFVnv6djq8ymecEPgJZGDIAWMsufxC
CWtaaZ0z6LqBddsmrQn4Qyoq5m91eLeGJZjypF/R1bLReiB4EBmKz1mFIUJ0YrdevsuwfO6kVR65
qmdZUwZlaLLmqgT8v4A4amdop+lAD+z0qCnR+fUc3VXWDzz6SJnJBSyc/PZ1J6pPBweQIH7pN0eQ
KAeKe2Ypcdl/HKUFyOg2TXhsZl8zbzNmSW8ktOuhmQ61eWyf4O9p8aTmeoUi/Adb72BukXzHzo7x
QVOyPy3PXOgR6RcftDYUctiThnoxisge5/GhWbXmc+WGayXbRHomkD56Le9DSWraYKuzCo0Qcx3f
wBmvB5nt1j3dz9jKXD4ejGifXhToTsgp+fsiB1qczh5XFt1A13mowfxLWLhHy9QCazQodMvqXM9K
cWnmhchsnCjfHghno++oRf40GvHCdgDVtj1qBIexIEsrSE5t7r6G2gv0h3BUbBNOSWYOpuPuChKY
YNuzATfSJPzE3F5NbvtQzoi0p2dxUwgbQGwXcQOSVMArp++Us/h/HsMtMMYcY4SM2H+jwtgd9/Qi
RxiaPuRItzk5p5yY+GqinWTv+Ic5WZRgflZelWGkNaox7iYIL78/O3CnAqy2Uf8p5z47WZKaVmuX
JKEYbpGTFaejONMTutTCZaj1PjmuNlHmI7/QKHG+34wxIyGWT5Mcx6wBUJcLJBZoUCdwjAX+Mwb4
WWFbicSgLPHbm7pFU3Um3oryBD5VMf/YoWz0+4fuHcqsfQDhRF0LnpMMw/iNxoh2YJIKcWR3vnlI
tCDfxnqbxhxIR51bQtu2p5qf1nktegq/vwlogGxfGFqYc92i+KAvwimbdIHQzhRdPyqpY97BwJvP
8ox7tIvMkkMkbbwG1bbohAxhjRq9WslYh3/G7d+FOngqC/IGFC+L24B2k7imYuPIkjXU6lPaQyuI
JJImbcvVmVkSKH4oOwFKgPTy+yWmAX6NFUvvDaDH92F6uTWRWvLN7pSSor/lzSIA7i192AX8Xqq0
iYJzd2fjwjsz+6F+6bt/jwPWTTmGte0DHxLmoDRrPg4oj7VwaAL1JuFqIu6wElhBiOwEo0GtYoj9
aE3ThMR94D92ppPMJOK4qGdFy/dGZimEnvEitKZE1jBCkTilZricJPQ/z1WJ/1dNRLvRq68bPd7M
0afJhXgnKDNJn1XxPDeDWWJvKIPjntIVsOAKApT59oj8cEHugm6VSKH4Z0VZO2PSHhnpXhSd6EYV
Q1eXYr1GlK12EviAPSDdGdDQ0CxWhSUfc2BaF45M6BSwvbCyN5XkYPaZZ02XZ0CuqIje89pzmeRa
Jf4TyQqNbuiz0p55A6bsY4Ji/o5ijIwUtx9p99/LS1vvtSp6SNtm0THzp4zQl/yAcVm2TfV28i1K
14f08H6xMJ3R1z0gu2Bum79feoFC4O0nnVvvhSmq2nB7JA5ln5syhJQCIIsoCsH2KOKKa34AbQSg
x7aA/zownWD8ZA8GzqK5onFw2uV6ZD670WpaZY1GDPntrJ+wH6SoG6QmDcW9gG48ZKIlkrsjwRQ0
rVOeqyPJ6UXW8BF4LVRzFlX/ZUbJ28b3sB2ATH3QrYgya2GPvY9Z9AZ+L7cIrKzXqWjUg6qCA9J8
9Xxz8KQRi3AlE3hD+7cxQbmn3X/gv1K7OtHkURKLCniMNzBV7zYEndkL0mbYHf8gp406hHrMQgMj
zB+4lLyhEQ3D+zv5HMHNMxCF416tMM1rRpyTalyim4rjm/Jg8RA+AJP7vr5zOgWNAsj006T4CKEk
KVtxoM1B7VTESly1hWR4vKgSPkeopFXli8vlWrBKNAyIrrcD40Suk/RD+Jxo/rLRHTxI8eptRISI
jHn1Jcxr4tANZA7KijaRxmE0bocCcWTJM+RbUq4/Jw+TyOII/phvlqCU2qHxAu2fWgfWwztjohzD
CXuZxkG9gNvugPz+kMOsGe6qigNC6c5xsm42eB72uKhIc4EmFvkyYW8r8qeTIjbxpDghwH5FRs1p
9UgXOrnNoAMUFQVLtE2VeebtLIfM/7lMRz04BUOqgxHlnLygaOC8arxklxEptokNZzmH/Im4jTnA
txSueKJr3rH42vXNwRDlHErPgR0rPFplI70FRRb88I4v+z03nLrK9scagNXADTW8yJ9MGOX60mEj
fBl7wk5LwUhs52LTENczPe05onnhxx7HCvK+37H9zfdoyWzul5kqACH9aRdJ0gjvpgH85hlxxk0l
vIzJSgRKgW7R1R8G9nJ8ezaBUe9kGMe4ztWL0lpvHMs0WeMA37ckPL1ajlNZJQCQTDwVKQbazWwT
eNZhvRYHHyji7zZpxMsGGsZF8C1BYs9PDbskrn3V/KeDjEK7pzn70ArXcAO8pUhsR30LbCdvyW1u
xbrX7h2sSjvng0eTL9iwEWNJYzrra46Abv+i9OjFK0HjPQFCowh0qmL0M71KSGVj0gj9mcxnnjeg
N20aEyO9aPw6Bc24wB3EhZ74fmmz5oXiLvLwFhvSZUDjHQ034En+g89X0D8L7E8CBhMr68eTQCn8
oix5A/+tVqTzpxZXXC9LspxQNp4GiAv76h2JYJ2pSyg9XEEmY2DkVI0UBSY0WdFWJz2NuF/hcw/q
wxGYkc4SiFQQx1jkqryalECzuGEphvjrzobctGYAvnQH6h4ncjE7u7E/1ZTtRjoB3IZve+YN4rkp
VcHVAq645mPElCZkqeQyr6fDy+Np58N1cFBO2o1J7ueESLFFyOxU2Gky/ALrxPRooLIc5jZRYAwK
54CPwLfKqNTq8LTbQ8WIkowBceUoCeauEUUcXZjNq/zAwYq/KD412OFZg2KnD6oxF6E8EPnAD63s
eQODtsTmt9d/uBsnTAovhhBhKBAhSYezt+oMoQlgFjG02GWybsDa6pqugeEzjGBTGIzuRCHf+1SB
FlHxML8+SOwTmJHNO12SqCBnFkvWg8h709LY7gwrRBof8k0cR0rS/mUrZwAFpCfzk7p27+fDNp4X
s26njnifkQai0tSOG6LQ/FiD4/v/sJNOEG7GEovcdciNhh+4Vldz83TGtc39qBWlT5HdRCecb+ax
WSvbFiZhdrbuvF9E63yxJMQNxanU/DHxadfpA+QgBtI6LcxnS5Pv1gFYTQe3kFR6bTbfYoSC9HHu
v9bBDl1ZODTI9bVJmax94kpGkH3lz+907ss9+rTf9uvUrRHeWe83jFSJ6DgFOqL0ETHXzVGe4i3f
uKgwGBkiCytnNwUq0/Dyg869fvfbADtjcY8pkfSoD+zGS/IsrGViNNawhAXNUJdPmd+DxOj07dPO
VcCsxBfzi2yeqMpk9jUgboU6RIyQ+pJLq/bsV3jONfj003wu3DhqKmEMwKfZqwxvh6wrk/lLkiVq
XtG39bymbsh1quFRy9h4dbbw2zUCyGlopWalcZlQcMQv4/LGJ7TOJCO5CoTOm5QcQlVMz/Oq1o6T
7PwohSbqDIXCRUtq1EiqNjTufUdRZ0zouauz7KwDMvw89iDr5ud9hi/koGcPm3N7iMINpxtLhLFc
qjg3ifXLKTEQZp3+ej7KqyN1UEwP7XrkflYpUdJEkWlrDaT1xFuTvhHIgYhb+dBCE0ODrFaOy8vf
DnJczyaiZ+sbelIIQf6gjOh7GwFzwkUMW+8vixhaCBcSkduyK1ELC7kNgPDvVhVANEppbuVaYdMR
LUIzKrga2c0JaxwJMb42JdbqpbLp0wjgql3bd4UBqRoCdbLwG68HcSiHqxEas7W3z8xr2XUt82CS
xVbtcKP0qzo1YWnuYHS9k7SA3khEqqpNPhKK13WDcaEYBbJ5xnpRnF3ZqRB2O9C9JwX0CMjgOS7o
XyLilQQZbHFKMkol2xNuPfOcYDDLinwXv3KFAhxYeOqUipOB8rW8LK/qLrKA84mKoJIPcOJGHkcc
TuPuF9beqZlriNCSdKdMIyR01OcyMatsbFDcVvH/xaWMvjyE4LJ3EdPqLS4oowPpymwVyopoJCNb
+lmCmrgYbUpcmGIFBLPRGsBD6scpksOaIVuwR5Rf6ktt1P+7Yx97P2hMPDFUkJ1BsMmwEii0rz/r
sAkfTRNEHkpZlcyCqNW2FQ1AX/Vg+9lsKoAP65r8p0CsrgDT3SZshOvS9BKSAhxM9mV81UadFZ0k
eJPfqdZk9tdnmFmYaXu4ecTqV1meICWdxylgXZ3yo+1r5o8iAY3wW4/FMhHlhECqHLuhu49EtJVR
gpfZrmbs8tikTsS9c1AGsajwys7zlaId5w7BTlxX2OV7Z9KOYLgE4JJKBzWzpU/GTIxNYJN2W1TW
cj5kdirhWnESzpqILRyFYKzXCRC8AzoGa1qGH5lJQxs41iC78zG2t8ty8q6D09QMV2dU3II/B9hV
1yJlPr1rRdrCVg7L2aZ7aR/VAAhXT9Jr0TpsJZQP7/5h7P4YUzDsxPsU1IVYhvdqsabVY5bNLW5p
Q+afSHdW1PaQH7FZDjhQ4OzXFYoNZtFrSXNsVIgToLr4nkcLAwl7kuaBPeQu0HKEO61SeCuK4FLz
fSN4RKncl8wIUHhpHQg/wED/uUCRdmk/WHfj047pL1H1fZhsT2JHAfCpdKF2KrJnqN/QzxDQsbZb
mblHeIy5nWG5dpYa8i24nI2YR5gORz+bhV9sxYDI9T2Ypteijq2U9KFOfnTapv1z5GSm+YezxHll
loHRgB2V4M6KyEhGWdTGj6dXseGCVZ69Dm6FaIYOkCgquPQr8LUyRiq0zH4HyL3Eq2LdSGxKeY00
CDGvJ2xncNvlvW7abEIH42pSZ/QKRFVsrw41H+X/lc2GKiIjlfLbYblsvLcR2M8HT80iJ9pjf0qg
ZUuUGDkEGtxXLGUpVPdu0so9mZMJcOLmjKMI0xC5vv4rR2r/NOQlAQ620GwwJ9Xy+0cIDbBdxyjo
dwpSRhI5ARIrcF2l9T31x06TQTSvvOVTW1g+WazClNx0uvj532gybj3G1jDUjakwQ4awtwFGT3mz
XHCodg3t/w6xea4QScu31klTYELpBIyfQXnKvq557XUeTkMPSNJux2qn6FHDtCSHcnTgkgnnOybI
lg0VCnvV6UZH1tb1Oa0Rq3EXa9QqLAMevik5vsXomk6Y9FGAU8/WwY0Gmp3qePus/+jkAhf/zrof
GsdPTnw9WbERvj6ViryYteiRFZ1PBGdH78CZfNFOrZUj5ORkw7FBkatB7sAcqQqSuMNRzvtYFxOJ
T4CfAP95mmpK48/Fe08fRTbOkPW8ecx8FnWtctA+jjlQkTErubq72qAaEohq2E/rO/Ud8dQNMYCh
P+dpyoVw9/8QQZQLxTUCvwiEbR+Q5YpMeJn+cMb2GnAvfz8msB6yxCYDXIKonmfy8s1l/pTOEefN
pqCAYhWZ9nQuXUFh4mdh/qcfR/hZThOwICWAzBkn2JK6BVutpoRndzksuQcwbd2+wIGLwWiZVuzN
kYcKc8b9XvERpMefhx0khZthb7NcTDicCIFElh5zwXnPeTDItRowUXWYf5RlV+SGDsNgproB2yqj
8l4/ZG0wf+s2gW8+5v1UPcL0QjqpCJp3iMSpes7rj702pBdBp/MqZZd43RebPzsD8TNTc/rgLqtH
A0fkj/RuC0NtkFZFax65/ba/kOzXQUoMphTRTy5Yl4YfM3PtB4GR+H/KfKfXMqPJqyzvHTiOuE5Z
TdTH8N4XODUS0djJrYoitAcs+bd9WGsClsvE/n+SZozLd9ocYbdDke/mzvlKVQN0F8wuH/fVoy8G
b8zYS5CYcLdFbwVHigYX1pHOsiDquETWpFW2TnBtwS5A8velzCXDW5A6eatFwIgGC9rhgNlcr2Ja
XP/fHicXc5IEhgw8C5Lg9Hg0qjO28J6rpfcDwHdiXlo8y+D9ecpztJgarZL15wKwI3bjW3vpC+/o
UM03cnNxamMSwi7P1eD4cAgfd38TN8KVE8a+/gVPsunl83jxirVkLftLdKIzofTvJkOy/P4I7N7/
lOAw+o9rhryxggDHe/bsphRtgByCRyQrnE/L7uDcAmQOvlMQAtP9mPRsuwKJkaBbAXTFi3gLU1Bs
fPc3byB9TAgdj9xQKGdf5hmfZSKNYA66MhhGltC4ecJBQqeiPJrKvuEuCEfDerYs2JUNwO46QFqr
UiD1EADdr3ATvBXZbNdoFgwswidC/CyO+VdFj1W5M9p8t2BoIXVc9xYNIx4iUo5taS5uWcXufuQS
cGhMT8wWNlqpxNff4q71TfbyNOTOmZMktYj58uqN3XyTQDVkAcdDUeuUjyRGVIKnnBswle2v7hY4
cwQv5d0tDNbXHvrecQA6cOy3dnfRJnkFmcVALd52yoDfmCwqX+wnaFaVrbG9tHGkY2z8qv36J5Fp
S7v96NQ5U9t9Ths2Sv2/T8JQgU+sVEuwZ4JXPp2JyGkNoi9maIF4DROxJrkVoAtTuxjrmtXkT4Za
8ecqy8OpnsvI3Eb2wznAZkNcFgR4MVGjoD5AH8sXebxIiDHmz2188b2l722l/JV38r/wpDiM90eD
c2soCyY8APH/0IuBb3TUpSvS1TNaX4/O3ejZZP5fhloGwf25NruAop45cTeg9MRha4Ra7kFsnHMl
9CK6RWgloaZad+6cuU4jMu9dGhyt3N3qJ0S1b/tsNT49yhheo7GT9u1iJjjyIPpmJy2Y+NY3botN
oQhLJNQEeOQzOqLc20oC2IbvVbFowS9IuN+3EGYYmt5h65dk0yCipAvqQ4fTID+UI9lmL8Mmqwvi
wfD2/w4MXB1EwmPel7Y13KgUXakQYH4YRPHBUI3YRjAAB6PX9TNvX1Rh77NfIvOtL5eIo5ncBVLs
7papg0KZCgYKkH82HcXQi62+Ht9mQD3sQRGLX/QuwjNxFYVQEBpe+VPzOqFyHBbHwF5C/xW07QVc
rKSEEgY1jnIlTazNIr/sME/Ifp41K5XJtmw/heVgi6I7z7alSt7/b6iRIfhBYC/WEnzTERcbjRlj
+UyN6Ha/dbOdOTn2+gZRyA9IIU3QdTfd8NBY+1i9KJ9CfT6dM2/pfK+/IfVQQtuvo4gyCkL8wmrS
7zLLQqATmXYth+0ZEHXkahFwof4BxJ7zXVeynYZYncAwz4KaS4rTpxMz5hiFlF/K8o8JClPJk5Vj
5wF0hC3OD30YplRxQy0jzJEGBKReacSe3PT7Q2PNKNQ0NHXUU2+8mnHRzeS9QS3GLGY+9NTznAIC
cLLJTv7NO5L6FRj1ZPOhUOkebMbtNB+WfSZHnaZt3fTnLFJOmZx2lPpGfLPe8A4UBw5oLJEVcLu6
XVcCGqd1Sn5kLmKmcaYVnubG8Lrtb0ftUyDUIwwRa4KCQRPQFljrBDBH8dC0+Q/tlma2J+qULU0s
2vabg1/uDzVCsmdqkOyXGvqn9ZLtzXVIaSIaSKWsEN1uKm+zLnNYuB+QWOjEkdrxVC/pebs/6T+k
Hb8gLcu6brjoW3ki71ZpBWiBFXuu49wUsFrbsoZv/rZrVTEgqWYhQytL0v8M8VIf89XkaRT5mXSS
Ojh9z49lmhtIwDgJuVDFQD3LVgpNKXGr036TSddg/UJbiLhTwDGjaN89RqJbpT+8C8CSlSMh7PW3
s46LuRik8+rMBBj9I2j7MmL5qrzyqHx0i1ckdShQ+NTD4AyqhqD0/c6d2wbUcxgP/IHweI0PR1Wl
/xyETgSCJFFlmFCrSaZhlc2UdfO/vtyRxnjo2ii5snxuwHG0zUARRFxd0u1F4xbbG/BvyZhnSPQf
tMgPL4gHc13hqBDcWu3TRfSSpgVfC9/6ZbOkxWSbgHDkLuHm2pKgnAe5d4cB3zb/OGZ9orJo/gF+
heJh9TEOXYAaZ+SoFVLRL+AsDf7AkKu5pf3c1Jafxbc0w7KRXvpuIMQgrIJ74NweSzaky1MmTifI
EcdP3MixIECWOhoKcICxe443AOaV6tgOv9GEK1cBCvxg31bEUdw4pIuY+D9TswCH4TZ7xx/n6r5j
/VomUO7Re9iAkeOGR4o+eQ0IWcETehf7JwAbVTBxIvWp92MYWXrgH7n8wCwGGRvnqqhupQeqff+2
iBI7A2yK1EcE7Tx8NNnifprbNdHPvz88FAFx+ZAQT/nuEnrmDQIKqeOqY8ubhDxK0gVUwoXgCseO
42ZvtVkvsaNnHcfGUeOXjOfudWdm2DDjKx54eOf8BsTmwJjWdAhFrFlFi+/6GwtAzxS81Y+Ci4DS
sptf3cSgml7+EeimXefodtPIGyjJsZc5DKttQFlQqAy2P81C78iTafye+Kiv3+TUDgOBe0YBkNAd
/S9o+T+vT64xgObSg0JvWcuZ+PQeGY9mQDBcMsMJxgUFdGig8z49v7o0JCy7NZmN17cIOt6wEgqP
32yruOa5UI79AD2DzzsMlyEJjgIPPPHjuNSJB4Bw7ubVbe6RkJ3GXSuOp4T25CmBOFQ8jF6A4jnP
r00UmZxduguYAEQ+W14V0DcCsodwYnqmL6Yc97H0nkBkXsLlx/8j1TP5y0DPoPUXDg4LlZPW+Sr0
ZJJKj/4eGGCycgWNBWYnKNj+l2nmLDlo4CimYiIQcNbaNgkOsW3T7uqga6a3RSRl1pSah+y7N4Zv
4zNrZQeaad7Ha31TQiAVFF4Tkaduj/98UpicNFeywVbOWRP0FcSPUOqEF5Y6zgGgoPQIDYtNbSsP
YZpCSFn9qooTsURahyFvq7OJDgUtnwHX/R8ISCKlzjAiQMiqYetqEhKap5IE3wWl4yDfqUxSY53F
q3nWJUeLm17NbfH4dUQSRREu7Bh5utZedb3tIar2OeZNZqjpR6+uDm2bVLmqGVuoORpnqa5Z9+c9
6I5Yfq8PUjFZhl24fcL6TLQ9XFtGFQjeZagrV/LpURezQDcnj+ZC+8CsR3sUVRau6zKWBSElXVRh
mNJc7J/p5CEXHDgE6TsMPVpWh1NmhSOgAiWWPF3+DGh5p8aVoREWvMjOqkxZg2tI9zOBPKAFjhqp
nmbEF3yGeq1pDtwKVIiq7y/8mAaqhjnqejRpnwkUlDS4TZq74K8PT4hh+facU9OKHzZ7XS0kORp6
NxAJPbEn6nFHRkaYRoCu8Haw+6qm0kwEwAYn6F2X5LuGziHQG1dMHNLPfeIYOkoyb1UwglALx+0R
Qv6h7R8jP/Qfnwvu5+UZnf95Rh8LCvrkcFJpHhbCuNmNb198BdYePkPSahopM9QbDIuqGGb6htgk
Q2wVLdsgFW+40FtiC3gLthVLZ7z8tQg+jTz6VxGlYRveiUoBIsA0JNqi5GHKApu0yQ/V0A5UII/+
fhk/IF+g+laxpklR+C/S5qPe2oL51/y3YC9in8V+MzCvSwlfuHYrD6vYYgeyRkwOdd8+eFRvTJ7c
lwH+Vv4O9LhD+nyhuiCBX0+JLDbXgPRZ1cwu7vYajxeTGZePFc8L+WW4CRUJvC6AQ3LBBDa5R2Df
wVSLH2ICKA7o7AVtNSw+DmKc6wUGoSH6E9m4Bwly9RoJCSd077FhbTD42EdisxjQT3fUBaq0bZ/s
C4szdSKwesVWp5vdVU3qT8vit5XEc74Hpg7jfg4PO9hL19+eBl/8oB3Yd1bzaXQ5GTNC0Or0PH0l
zHnOsMaNLcnS6jEEuGEWv2X0+zm6z0mpoFCNxygN2TeNd7lySpf2MTQcT0oBCGZR/DJli6nQUm4j
kR24+kwqoa35o6WcxLU5hTjfTpl7NTbHUrEhrElho2MZaKSHDwMJvcuV/IvW2O9LQz1F132IJLBW
hMVLE28Q5Hpa+KaShl8WtqHTNRBSM3tjI7mZuYBwNuQQd0ZaIH07kafDndbSDyNj7bZ8qEAQozgr
NWxszp2JO4s3EdUq3odB+R62uOCcC6EMlp7UYt34fUpnn/SSpwRdutIw+tBCGY9tzCzkxKs5ZHHO
Re2+e9V96S+PPcXTyC3Qfk1+R5jc4ZZn3gS4roVBsKf42+hTUALXBiUQ0LkyOWjxZTFHqwKSFiz6
hIS6jdRGgdPd4W03iGcZ4NMj+m/nnSwAq1RrWVI4XK8FRIgFz6vjEZK7NBxveuH4GhbMvpVPtY8U
RdOR7Hc+eHqoot15RAR8TqzL73TNKrToHH1eia1pXHhUSYqx3CWqEWkO/2DLPzMeM2t+6O4nxHrr
7zIuzK77RkG1f4lm2jMhEdm+UvmMO65ITP2ZvKLNIDht53SJHUGuWrfEEXtdea/1gYPM5chJAv1s
XShpJj5JIuWw85ZC6WTaSeAqM0i2C/tUBeuNNbngC7CHoaiLePlV7mtcN0SDrTNxwfXlGUj0/Re3
uuJR9F4dJblJf4Hl9nHTmEmx6ZgYcIglJJaXirPkTym6GGwDPHSnJ/xbjjcqAEjTi6nEqYjcM0tv
Nf+H58q1uWHMTe9KnPlQZNeSGKokQ7RRezvBHod9EP2z3ibQjH0kzictcsGs4uRp917nK2Zm8eF9
8sOeNWEFugmvOHM1ekUWpkSLtx+DVBzGknnafCkLbCCXqLqRir6BV+/bSoo5dx878Eh8nkFs5OgK
sZ1kJWIlevfENHXswli4i4ZxU0KGZk/XZ54lr3tYjFGAGyPOQpWHS53Z3yq4o1hOfTG4n2ya82Yh
FPNQ64JK78hw4sRkG/9SdlqfcizzeIHXd18ex1cHRaV+4OS6gAT58Z+wVQ5TeYes4OEq87p8pqy3
ErknTQh4pRWnpWTHZd7UDB77pNPxVwa5ivEk7Ntx6L0/8upGlpdh4jBn8TfV5Bk1MtA/xZsJ5rkz
L8jZG1c0aIneTXhoJpZMlSFOhd+zlInt2rXPZwdiAhSNlRQPCXq58I4YCYGdYghAynzH24cFSIub
N+NCqmllto7jgEjv6djoiUDQCQm0sny9cEvONEzQw/23mVyFf2chRq+2EAT8kvumlO7U7dUwGclJ
J420HmvhTuFQAM5j/Lc5FSNf4nFnxNeCTwj6kh+cdx0kLz7lBbjQ85OEDrtsrGWzsfVRhRr7qsvV
O3ZmUPsG2jW3C51Wnb8CvC0CObJxP2XDEsMl6VWsDFI4qP3hGVzTIPJ2g0O5hM1pkLKzzlfiPJRN
J+hgZbAm1RLR0FxOcogt1Ua5sy3CsiqsxiDDoE/RuKyE5s3c/eVbcKlmrjPAREpfgusRNeeBRZcw
IGFROQiRgVlvcSDY5znLsuNUZP37CsE2BdfpNvX7TS2TDsFRPuw3hD4omkp1AlTDK7QW+TImaTbv
MCEqkLNDz/tv8AOqDpTK0NK5peBy5uGn1O0onac6BgkzLfEX6QW8G2RCnDjy3xRA1iDVZdH4qWcR
XcRpcusl1pxuYFXjz03/PK37QJfD4PYBfEX0gLlrS+vy4gYPBuVV2GJsJwN8tnTCa/eZLku1JLFU
OudSt908gwlvgJUGzmQDQOC7+L4QQX9zTl0uq1ksRw3W9mQ0eo9Jyu9jbMBHIyTdzlmvfDgUfmY2
c24Vlh5tNuDKpOQicsbLGzXaSUqAOLCm0q9SLfJepeF5K30qvVrVjDPezm9itcyW02hmfkT+QHgA
zCadHh2UG3vf5mA24YAuQQ8dboVuHa9q+9+2arc7asr2l5NTEykaSbesPeOSY/WHK9Mm4yx5uWFb
pbOcsNpF30viKFMEnFXTxU0i+9pFMpM7glk/5nKuNhAgaAAo15dTimZNmfTX0+8n1s0m9lH1vGDt
VrG3mYl3VegFKm+JwJdY6PSxYx2juiQPdK0xqZNjzB6B52+w8Fqpz6G9KTKHotSKfe3DlcRTLjUI
TogNAne99hxYRc3/E8AJg3FsY7jdqY/cDyIaTl1hZdHJVkTIeVPW1ilv2dVeyFY63cwDrNO0R3/2
5EiYmC27ZcIkQqbbfTi7DRko9mgjVuaRfIMNeqCcAvr2n+tMMdhmZuOEBLd9FypUKU9iCkTLkJoq
yMBlJ07v2nJHFWXRln6+tbscBko6UiqllpM9XKogClPO0TwLPh82CqIgAUuYycCApyJFoit0qW5M
sVWgO03kPFobN//BnKss2YZimK6obzqQTt+gqfv3tcTgGIKMB7ufnR/+qahdSaCerOYHfr4TGsKD
5pH1kLJU0CXJxLvQSkeFmbigh3S0ixafuQty+bJ+pQ8WypvuEp8YFBplXZiuvsGggkje2xgTNe0m
XIkgYN5Hjz2h122rM05wy/MYw/kgv+3SyTnO/PZZM0wWlOM9fTqYwF6rV6fS1leQyJv+5nRnUOl+
HEqs4vJ/Dbaaea+WzCuLxAIGUM8m+AvFrjh/3cjKNPptYr0vlnEsMhfz7j/w5hqkCZpCYF7xDMiM
kRycHCr///X0/YlegdcjouIRNyEWP/tdIxDWKG+htZ7zCz+35owF5azjPg2hmrutxmmgSdRsf1yS
XDl+P7zAAfjBIxPdKR2pC20UCwCQiqhtr6LzxlTHqItf2FKDoO7RHJnyL2UbFUXB9Q51q8ETxmq7
nm1H3RMk++iHSaQGS9UJwBDLrkK8iMCLeY1WmZ6UF3u4tqjKWPZsgtje4PP6rNP8Rn/SmMSVSnBE
873+3TNqDQEezqz9grsS3HhIHh90JE2HJbE5YarUbO3qiqam1uPi5+/LwRIph9EZlsCiNKkILYMa
de7B8iy61yZY0cmbAqdAuDBzVk7OOGSZC53BDr4hEn1+w9joXUef5q8fRkqCBfkz8u8zPMInpJPx
ditTImk/aO5pJaFBx7eRWfOnZ5tELDIGa+6BPqPVsLfNkPK7HOHTdKVhNFrYCKIDwv8S+d5eW9Xf
CXWcvmf/koBfOeEIFGHxUPgeI07i8IU3QuAjTcY9GVTBMePtGtDuB8Q2T5MarGe7MeGfvvt/nmmO
ASObNkZT8Voe43oMCQrsfC3QjVVciN2T69wJEiXvDkeP45IsqMXIDfMowqvOSHk7EW21BMMsHvmO
imb81WkSynG0VxIUUdCZGBBnYoPZT9Ku5kkNZt69ll82LDeJqGrC/UGs9HOApBCUyltBmnKtovIl
yoWh6Yt4zgg8OfG7HuG37zYnNfBlgabAf9xOa8f889IJ4xlyh7R7ynU88oDil43l2RDB0CU1BEYF
EPQRW23/TGu6w7yIpbvz3PwRSCViYP39QfhLv7o7+UOGbbnCr4fi7lqp1vxnY/S62IxHs2N0QnwV
fmC1JHS4rqVo6Ye/NxCzPur8rFlpWrqZiTFd3o+cjhkaQhFmn+i7KFfrT2mWSD87m0sG7vklhn4r
PotoZRy1gcQRWOmxl+UsULlTXY3OrscS13Qb+hKJ+mk7P7bsbiGtePAA+KBHntaQoq+SHMT9qUva
jG3wgDy2/i7YTCHWKdkw9PzdS1hSIr9+ApnSnYS3dUpQs25/CdqLQgHqV1KLdGZ0589UCixkq5Es
kEHexS0q1bsDcbBCZ4Vd/v6lSASwan1U+5B3s8gEQZMeoa5lQ85ABgQl1ykYUL4GYyazRiAYDxP+
Nw9PxWUnWvJITIEtkaMLCRwn/KNWrQHmikA9gjJ5HRP0lBKkP0TFMPbAyj0h1xROgKOEsX5Nyf60
2SpIRsHEXwGvssvDUEkBYzvHO8akpSUPg+VbnRVxWplICHSWKoa5940j/Dw/JMkg5JllmPFOvamf
XyDn0zl5NZKo9i2LLfv4bi+JV4IuBwunwvuX/QYlP9R69vCG4b7cuS7iS9aM6IB5TbHmtU7CEQJk
bbx40RwjKlqprx3AXRgn7mR8QhMdzS0gLvbbI3j6V5oeaw1UfkcTwvCRCSJKqqU0z0OVrx3R1wJ8
u8HHkYjC90Wu3HiWwOqeMfVp3uT8CfdIggAXBurZe9LHvGGLf4HNuTKegURfbdKQir+L0FjvHbi4
idOiiFSA3ZF0uSGycaWgcyy4IURSFiHNtHxvvAVRBVijQQM6kWO5Zy2d8dIeX3H2uRxTzjyq6No8
Ez9BKe/mo0Js7etM7slv1V8xwtcYxGgmB7b7fiSuENevo+5ieW4UQhL0nkVU1YiREE/Z2P5b0blF
IgePXOnKBSvD6+mcPa6rvby7p2p/oAl41k5Tv79EtQzr0duRTFHp++I0atkHNgIukr6taQRFG/wn
PHi8jpkJXxBXRxHQHO673v4HsAkDzoXXiHS/anOl4aWp2wdRb6RalU4WFmwv6Ve3nnfGFiBKD0Wm
tvnoIhQrAm3k9M5/fV6WvG7TOJeiKhT9+Ll34RO8KHfXpzRPufYMRIjAMnnJh68cpcHyDBkSiJWy
x8wsEILf2n8eRTT1w/3UDZMhtrE7W4N5P5FZhxqj4SP5atwaSecL+Q2PsVEFORmxDNm7gJgC+G1L
D/RwZ+9nIEb/b5BQxGcp9ij9sEQPsvy9MKNMt/heQscbn2xvHYIPl8NRFwdTdWPaM5xK1SbT3m0h
xLpJfa/DHlLRczuY6blx3d9xipLaT+arrtMJaU3BeHGSRHY1LlUpJY6KWMD2YH7ru4z3YOWZsx4P
rDG5jHj1rJ0iJZKsUbttIbEvs38rOeSQQo9PMFJKbKw/tW1xK7fWwghov+ASEAufF6dH3fUR37LK
uJ7sriFosRw4FOWRkWcHwGwd/BTGo67Sj626XN4LQHRfxRGZCpBi7FU0UxzlA6SwZZnW/SkCDgkk
SGjV8InAYouzE2tlH0ak2GY7wHFxSDkMfq5aemqVOevangCk/O1CF+SH97Wl5RgxdaeMK9FUW6BU
TbvKJKMcyfKJTJH8VVLsQ79CJrvN4ftTIzFezztfm+XB3GHKiY8+6g==
`protect end_protected
