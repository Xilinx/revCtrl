`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jNvGKMNtWEUNKagzcg2Z6WIUWv9gWJV7my4RvssH/ux/cX8RktigUyw+RYrzrXJGrNW7g1x/nBwF
74yzP41Y4A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cve4pj2EfLuhqfhnGnOz5iUJuIGWUldTY5TKWZtU1S3TPZ4r9ymlKXit4YnjR9S0JtAX1GoFuudL
h/jZOj05rTC9CmxzpO6a4qp621eKZhXdyOHyWMf8jPXE24P9V+aRttTL8nXifMfo/UFfsvRfUHHL
a0V7II16UbNY0z/aQ74=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FK+UvGaeunWTo0SP2EhgyPGTZaNb+A6fyrB0Pb4mabhgLBujusE/NHHToooQsIrVtG+iA4L6uoFa
xZk2qbFfIXLgeHkE73Jf9tkvOVSfNHKkwE4Tk/zJ3hux51whzpeHeM/jgYHXV/AGxAjK7wYmqNEp
cavJsaWgLnwe3yjG331MbcwzkmgERAfcBrC1i6iTT7oe42Z8bgt2QuADWtJa6+y6yzc95b43/J72
7JqV+DovmhlKbNR1biVaDlEMoR8wVeDr0xj6PecXn0O/DCkFw3POXJoaMT+xrRj1LksGsCY+qMlG
IfvdA3kKCxIRZxGcAPvET4wf6cGXK4CAVBa7IA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
z2wDansBNwtedB12HDIWNrI0jJ9Of4AnAAv+qKssr7e7NujivlJDkMFVu15DOLNgNtFvyO0niOHn
/kdDAjIwQtt+ugBkFsRzbHtzg25iwcWgxIDasTP9xLaasNHS5B2OfeSNk+sAZRujgTnv16OLLpuj
xCVg+ocyScQyJTN2fY0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dHaEE44368Lqz+gkjyTg7OMF1sLix1urvVlzCGNFKkIp5zxC5Hb5ei+82XYKqaRz661xkzrxnXIz
CLpQVXEZh1wM12r8fA1f5G/ZuHgSsoz7RWoNbHd4G2GQJUG7WVKCnogPJmbAQZpXthW3KW14NIsi
E34leEwjyTjx/frRrPczvVKGoZSH0tKOZiCD2ER5SRLpYvlTJUkcUEXx3CipAjm/wVGV6SSyQJeO
CTF45Rt8GOFQIMhL/GO7xMB3lpMvQg6M9+8i4GbdQOAk3MmCg7nCiIL/ptz2eDE+txQ7xQlXt4Cv
Iz7BX+6KUqHhfTCrqRi9bRB7HwJgifi1MzfmqA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4048)
`protect data_block
dBSVDAWiIsOQDtztSiCUKV2dJjLLY1u9cgJNvfNDnv1h86vDqn8lVoOz+Vo9VeiO/U6bUH5BVLiM
I+s+Dn1Hi1GqUglU1a58QdP4aVSm/Em06R56xFVG+YWqGCmMLF67zSg6tySpnQsHJgH24U9TiZRY
+251BVYlX+Br7+BffoBkqhwRliAI0HHcDHuxuHdrh0hWx+pYY/t5ghmqL0SR9MVWnklQMu+9s8Me
uhNmy7rQ1GbWeOboHREgfl8WNEUvtLV6Jl9HQESh5VH0kpdtsj5mGXYRAt6xHY6CLzle1m6g93N5
sTgW+TKh9k/yT7srN7f6LuWqWPeE9wMDwchlAcGN9+tH36F0RogjnvdlOp6k5WZmSiiIkleFcNF9
9j+d4aydVnz5Oqiks1gSZPEpuOPXA7WSaEMhPb+OyThFGBhF52RsUzzygLpWLf32yL0hD72pbzFj
YeFH8T+gWozZmS5RzA7o6+4E5WDep6HG0yCkGNwSRFeoEPAqYgaIvcXNh3ZzPxMZOR5Lqyn0uQLG
8GqOI8e3J8yNwmek/a9nPRc1ITebCeBFaeOgxlLvct0h/WO2IgYRPqijQKLIfExQn294RwfXapLp
FeL520ypq1TeR9T+R6iCwawSL5WawPFraw2LjUZkVVzVpoB04uxR/oPuaY1V3OIPC09VUUtDX6zS
HzLbS6HlJlc+cPon5U6edz+f+C1mFN6HJMBGYcqHVX3xGvvEOBYUG9g+lFHlj+T7I4L/32qC9fa9
5XTBmtZxdIQJnTMEEjCGMFa3By4Ju4hpMFIo+kh+3d9exi3hYBOrnIHZH8Nw8pZnoCE6k/7eyype
OkUc61M4P0JAcYjCGrGnHDEOwUC2iUpuCmbXNglIO33BUb0hbzHQY8MD1V4ZOBnJhZqj14RddIKn
AXnwYX+hM921NAcplLl8MMLJvoq5vrNhwHU8qFWOnd6iwYWRHkfL5RJ7AUqH6cSzWQmkgVIFV0WS
k/B77XlE2CBcYiA30QMQMi9GY1m7c3HjhfgA8ZLlX677nVhvDEmDZWjLP5FqS1uq0tXlei4Qsaja
cJZ5OrtLC4jjFxQD8tYVQQSas3diLD2J2ZL9VR7VTHRPnxtM7aE31o6sFkTDR+la1pKJeW8uRXlD
c8RjCV+l5pW0eFt45bIb9HQkEN2ShuANTiEz/VxgrQ1nYaAlnwBsKuzdUhLEzpdyjg6IyQnXLaAx
YL5aRxnyi6DGB1WhMFQdFLiCn3Tm3b2/cmyGZCESp5lf3vbgsUu7FJtiEbl9XwZGByftOUXaP994
ohFydNzvGK431WPcAlNRRgm1mPEyY2kSkzcqLAhaJft7+JCcwlmY+urWWPo29ns99uCGxReYpmDM
25jlNIqAl3nOfNTiYZwKxBGyhgPfxfD67ghqOLB7EAQqyfCp8Bt/7DU0/8Eyxzce4KVSuNmP97ur
iSs7hsx1oKa6gMuKXP7hKDIdq7oP5327zm/T/UElkdfHsAhOF412FBgPQIECRj+R7KIeRroR783p
mQHR+j/UuzptAdQ9aUjLtfdTGPpoU6xfRZL+o0I0XzXF7ckMmVBFHAhMahzKSFMtRx3dEYBlYO8i
Tt3q7+9ZDP9feQo12V2JXjTHw1WtNlonp6dPod3RK+lFsadre7yUel1I0J/M6SRwanxwALDZB+EW
Jh4IJl0BOA+8e1nPulK0SF6KB/IwYXvPiKQCjj8EXQEvOa53ZwyCQW6UcixJQDGaV8DZ6yDtStaj
b/+HB1XGj53XHqvhNbAugDGm1BhtFJfV1hDdiUXJ2s9o3flhLi/bhKKaOCO6zmM9ik9XG/TvUy0+
54HBrGyDNptxj4pdZG18WRapZ88BbweOx+YBb4eXZvqQItU8qY05VzG2jvTu5Hk6n2rm8LF7KO4N
Zh7iHeE0yB0TUpmgY8PNfWAKc8mSwZtk3f1bGtTtsygFsbyr3un9O3zHl0iCXAUbZPZUxercO9et
8Kna0LPBQKA/KXV8qejrOTbM6ajTn2lvSfG6gZpOZlPCrGuAuzToJQyTdlUZiJJrot1DALVyGZ3I
J7ocBwWPusI+hWBlTWHk1IaBzrfUTyiAU3QsWW6AHkF6P1+kWHQO1zfCSEEV2WIEu/M8S/aeRRCg
+JsaUeRzv6upWJE+L6pJ7qjtF2cT38HXh451tYpyvoUlkMdWOPoiLzc2/WVotQ/im5pC6KEwGGqZ
iUWrMYrvmR6jQXitmav1y20i7IxOeW1cKYbfo/7trc8lgkIF8NbwvMmG5J2U/JRh9Ubcs9TtVu6q
wFWtL8vZlgoUcdwFEr0IqURotqPQNC3Ksiq1ysC6Z7ru8LFQgcF9Et8BtSwNTKgLP64LdnrJwPuK
l0QJT3Pfb8dqRovikzq1h0VXRM+QD5xu/6XHkFUYvoem8KrHMUPYHjF01f7JYxLbGhCsfxk5NFD+
kPYxyh0ALimB6ePRR/K3l2XP1EIhrjkdMrYWmuRYqLjcIvXTqXX2oif4d6cMpHL3Uo/5SXa0Vmq6
1eBR+OdauV3fRdMOLUmb7Zm3I76gv8Bk02pm97f+FV88eFuJ3rjR580VlMjmDYzj6qbIlRGljBng
Spa8m9H2J68uOCJ4c21Ja/PWaJWjOvOTj5MkMu3JH7xYUsBH5LPt7oqcu0z1LMQ86jv5NQZiIJut
RInRLMaKBLWiCIXmClX1jFGuRagtaaKEKBrRzAdoc3WuKsAf7uAVN2MioUGV0LRnjRXSdn+8221r
9xvJ7uwnePfOlSkF88GMfc29CNl5vF0jBw6ebYunRfIcKhIRaih3MQ2lsntWga1fM8jNlwn2tS70
ZtqIwhRJ8kBL1DrvwCwFDHPeLr7R/QRDoFxkohUBvn1B3EMKzfDfBNl0oWI9ER7PL88zCUN8rV/W
G0XpW0N2CqeOwiI8YLWWUP+Gdi1YT29vlxg4Q5BqF13wswh2IYwLSwiPDT6pRFpuxaPCSp/h9pwo
ALBiL6P+YjUlIqnWKpqy8PPoohU1z+8c4AMK20qNgkVkYBnlosvp/S2Vumo+AYZPSim5v/fChQkQ
a+/8AxPIk79Gb11BnlHDRxN8DagDWmvNFBANXGL3zZ+C92niw3H2R7JEs80+1vHBEkXi4dlGmyg+
3Z8GZAg92g61X2ahlT9H9reRYFwYU7cPxjOWZUQO3K4abo+4UtGDWyTNPj64x85NrrZzU6HR7hBf
VDPCOqGyKJ/mEiJrGxT/1ufeiBbndsx2T/US7Tf/YwYaA1bSrzM9zd7uoIWGuimUn7nxq/I0nA+K
NMRdHKoPuM2/r3/Ut76kemPpsVNHe2SA8Q9ySGWXqhIV/moFwwIWcI4I2cQm+VmkIU2N38bU5o0j
6ys/JNkEp4y2VI5Q5urdQ+cfpP4qHUVfvpsaahYowZFHJdm0E8vdxtuvPwSxjlTWKJ/knRpLVK0Z
zLhkyRSNT+OdHBOeRDrRJdwrl4JP1CQRVdUqnjPjNSFIYtNBkETJ72LXbJ08hEBmS+v9bXwgaA68
kyNYsvXCjE68WphOb/JHqzT1uKEFFR4HI55b0aUkNA8/HzzpduyvhHd2GVBchExxZ78sO27wx7mQ
4zlYJgyOUPPElGczKqK3IzCVjXgenh+ZcP00+osMxcLjVRvvaEComEIIYu82xk3k38sFotiFTNPO
6bfarYM3gn8oWYrrlreJ/K7bPHijnmMJ2ZgfatqS69VpWCifGkUQN20ZI01bAYVzNMVY79rd39K8
lgymFeO4ePOjDsGriS1doZDtJeAce0lUb54B35//+yR0fPDoOJxxWEsAmCP9IeNTty1lFdkb1Yft
ibsftUw872vnBdkrTTYvRyc03DUMBehL/9cyqdcpVPWUWctY0UPVTotUeMZDgXyBfN83HxdUwgaA
sL02mzn3FekER9NscNJJ9h4snqwAEKV7uhXELOLHuBzaC7T8qJHHbHm205NvixiQwBf8zGZmcpCV
jqz+qlU3vHM3kj0I6X5sHCDsTi4LTiKuYkgtTZQOb1kL9kGwxm7afwoK6uAWr8t5NVcyXJ5tju+l
hIcbKF0tXFiyJqLXDs2jKwy+AgaNUpw3zaT3RZr5g0/Vpb8L18kUe8/nyPAWm2JyfUxAhGbK2P7r
UzO56b/WkvryZ8lF2loMiM3I4iw2lSKixRFZYpO2WIexKWjS++zg6o/v62VqUdhfEfafvfBdgq5X
rOvDtLbY2yp1HxJmWEN/EmzvUf9RRVLI8RZh08u0brKhrL99M39S6h0J6T+8DxhQLn5+5FPuW8X9
AZngW0lweP0tAcdCnSetSzvb4GLgwbZb34VJqD69XYPTeH1nefsRqqGVWwVouuXy7dI3LnHhketv
NZBynCEVNiIuHLwNNeM29J8hDdvy3iNEugUF6bAX9M+D/Yv+Sjps4CNkbRGC+S4uHHqUIYjGUMDS
kFPmRmfLOwLAXUwSgePhfmuclE3ZmIm7jBKf8FuTmcG5s5bj4GRHBYqjaJkOe5vz/v9UDTyHazEj
hAvlgkpeuvFzo1mHAqJ6FOpiDNccBWtuesIVhS1q6b0MqHu1UJyxNsH+wW7zWIbt3yCmhuEqxOyR
6nwlX2mDuLLzicUCkvSBhFGgz0rRnBZqfZ53tQ5dC1rufZtuOaZLIsW5diS+H77SWxqg10MUfdq5
n7WxZ+ty5COD+f9xuqMtH6GPRbZZZF1bZE9WCmgf1/hM0C599Y8vKf7l1G8qie05GKXKwKbaU0hY
R8G1S9o4cIYoXe7DtpKVZoUhfmmuxsmSFpYfWARfwGDpUiqa6VVfaKwOEvro6twRdjxnXH7YSosM
VUbKIpZFb8i64oV5BP/QCoXtKhum6bk8TEO3oy5f8kPDNivrK59ZxvkQI+HV+TxPj+MjGW64+qut
cwNkoKigcJl1SH3wWg8mxOG9UQQejxDQ80sBn23Gq3fO7LvNG6p4kscvVkFH1vt/JiwKioi0n5Mg
nZR0xZHULMDMsbJ7o20ohHcv7bRUBxEhK5V+aAHQrwMwHfWFErtI0M6rx7m5HGt7EcNoUGkq8mdb
SobXBvyOOTJEhx+OOVjJnB+jHg4Ysf1dgyoQmJiOQsZnJhd7hxXT8O0v15tKz+i6f1SRpHHZKPqD
r6eTpHPgjr6S9zMHqwGeWn5ftyyep1tqz7lzPzt7ntt8ioum4oSVqu0sxx7VddXqbiqpprbSoR1i
N8+d4pA+8dEsPGKSlDPOS78xaPi2Y3+nVo2C8g+OWFq1xL5UbPO/qXK5lrN+lx6Dcmv29FQvHMrh
hVO7Yn7Fay99YynoNeGRjIcVQFxjGCDbGzJtbYu0dNbh98ur+ELM/XpZGv8tYYpjsOYoNZHba17L
GJXDsyDI1ocw287b7kOZPp2GHw/RqVWKVviLxVDVz+s178B+LsghKCMTFmW6i3Ra4oP525wJVqqD
FA==
`protect end_protected
