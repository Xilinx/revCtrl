`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
crsuNbGKr2+HGjsnrWAO3ApjaENLE5lmTkmDpqy6wXOqFQIJnrktoh4R9l/TVlY/BEwSOhFtvEbq
RKvf5np1ZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfoL36fNI5DjzIQX15YYPTK98uQI+Z0aMjl+hiAVWq0lzClrfpDjXWaPyQGiPvnYkkUnnCNmSyGP
qGrNm7GOsjezCGzMgQVr0792OKktWuV2kt0zVP1RUZuHk/37eznwh8N2o5rw+1YzW4dGzl1QbJom
tmB1UpBcp868gDBGaIo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nZKDyxkYA9uy2Xb3FwpEri9edMFM6SqsP4Aed0tRsVeeX445M1QANBu8GOl8sJ4QNxr6T3VU33/s
FK93SNbe96iXZq7rd0ZTftDGFn/wlb+m7r0WSjfp5pkNrLXaYMROFr5Y+cSF68dabG3s3COIhufS
z6LjxtxffkVZFl10/p5NYIyhVlCgj28/qTLowb5EYe1tZ0WPUAxBFuTyFKtX6X8Ha+x+nETiYK6i
PAhbV564AhzWOG1ohxDJJcn/sq1JfdeuDFdYSbNKycH1TqhYGY4rODz7EB10q4+UCVziUOr4Tv4R
NCotWnw5vu+fF2mIxu+vVyyYTSX+rhEfPs2iXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZ2XWhB75BM0Dt/9VMCHTjvBqUtECoyfIkFt8UyDN1IrerieLUkQavGMJnAyOgfgB2F9GkPnzVQV
7H9tsdZ87Y+A3ybRmsawN7gt2tqx/GGsvZlikuuSepi3sHN1vWxch8VpcI/SFn7CnlCh0jupM6VR
707+yLDj5AJkQVyH1LA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S4eCKuneguafnmn96ntdnponlGVTmyJu6zrxyF34ICbqsowM9Vhvgm6poU8XDQ/BrjS+RNPc37Fg
G4CZX64FNy0IB8M93ARmuOVvrGN2bYMf3jNRnVO/z1hOqr23u4iXXLcNjJcX+q+ntygTqDn+dkJa
tNf5JDJd7KcZbafDC5iOu1RcjafQnwlpqyaxuvNRdQkJM7f5tDyB/fmqWMaeSiYSf6cbwC2Jk6x0
7wUP2rAkEzcYQjkJqSGT74QQ9ZxpJuO1xNUbfsJDlmWbSmEyg55J46Q3XRBw9O4UV1TNB2XnSxvt
0rRnDIzS8sn75CDPR31VCmG8K+PwSCayofA3ZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12128)
`protect data_block
HGwVbJA7sypyD5yh/+WUmYczAUp9Ilw63ul2foAahIAqxWWNlG860q1IJCvcDi+ST5/TvxcuzPir
qt27wGW80Ur84JcU1ohvXeBLj7wUxE4SSH0YZIS2OeLGptmd6Woi/81U8unCKXYvaMQPcML2PbCK
1eHC1m0mAw6MVGLk5Z42s72GjDdmV6hti5evWU+/CY1OBTVp+AqaZC1aYiUAW3PSNH3hY2wA6RDF
cs8eggDwyf/bgRCCicfm56kjrb0jXfM8Y+t+uTF8cmBa1Xr/Li2UsxkFw4tyTL21LEN3rjPGcl7O
uopWN4QsSquJktHagfDjMwgNre/nvTDCjB+O0v9AniBJzkVrEIUo9ywzYvj7G5BrqjKVf31OAQvt
PMHzIlmxTUBlNg99Fy5VxvexNSr9Ebq2F1tlmykUWFpS1SgYsRnIMs9VuFtzALOVUkf6Mhmszvxi
OnAluGjddVvI6Yx4gBK4l0pa8g2XNjqneRN6W1fvhK9xtE+uchDketyTzpCt7dXNBSkRQ3Wc2p27
mlfXqIUxOvOtilV1vX/sRSH3ajGsEo3yzl6aJFQ+thavccJuNEuRrv6j0s8I/i/0s0+iB/Hvo+u3
46j6aWVNF6B4QNqCEfpSDx9U52IoS8A5U4Ogruxw5haVjsm/EuHknfjLeEOYGu7owgDd+s7PwCHW
mjC9+Zrsqz1T7i1K1CaVYaEFmvzUG45zLDOFg/m5jiXDaRMeYnqSM69ObmXMk6jdIi3Wclw8Sd3/
XJoWCaB8aDudmv8PwPpdmjKb3SZj3hWqE4Q1OAUckRJf74uyzvl5uyJnKBr6Iwq1TJIB7VeXqWVX
LXVnvecsoWOnfmizzE4iFj+dvK4LzNIptb6s0DIlr8N7OeBONnyHCuR41EoA29rYVDX9hF88/k1w
YHJOrY89dzo8BIXUbWq8C+9WpA6E3Z+rBt06tSXdhrrfLcaKPnrzy/fyUSLJRcwxYSb/Nrfso3o1
KAwuPnY1ecvnmmIbdTD3qt2/JF3chUfzFQQl3MJeopXta4QZGus1BVRudgcEutHK1RP/15/8WJ8I
MiOGk8+NepRdwIpdxgZf+slfZhGmXnQ7Jpxzp6OMHySj9FOrcMaPJqKM0T14DjC1MIyriaMLBF+x
5NG7dSwJ8Kz/hXLjMG2xkrwv2NuQanpSGSgYWb+bx3KuPUhc6P6bKGy48A5VhoKnXe8xS6gMyH++
g/WpbeA7EvoK59Gu/9jifdjMAGD4KkniNy6z6rzhZhTApRjNY9CoFq7SkmgyGzxoIz1HbNKOpPxT
mxJRiffnv7g3EckwbO4NZN14gHJtcCvE1iRqCkjMCzrU1pYyz1ca7HYDbTG8Uz2R4kxfuOsBX8RC
905yLdYQ+G0B8+42blj0kpLZP6nc/EX+ubb91/89gZ/Ujx3SNfih2dN5HzFZZZTZ1ilcHcKg7myr
t8vBgWShj7Nzmi9apVwuadlty7vp2uxFgvloG0LH0F3sIDo9mwc8w2Zym9LOys3BgTDNSfVnaTQs
G7E4K4a7VVIxHCyFMDBJJERoEXJsdJiZOdfridTpriXnH4LTuuZhllYwDrDUpELI+/6oCd+zmgnn
FdjviwIzImfuZ4PD6KWZ5CiZrhmfR7HdQwEx2VHtM8BRVKEyNXMRZtJurSlVkUcWhdISsAOz6u3k
jDSEdwQ1jaRwHXDlS2jj1+TrLjRoBDWrlpeKblOXaddj+ID/QPtYk//DhTYjfMTLeJIFEfy2uJqB
S510/Asz4F70bgv+M9oXdDuP4TOX38c+ycTHBDRZblVEJnKYHel3I7Yc7d/QFqBbrRN7yBQaIoG+
wRMkaoteiYGGtth5WxmbN4ArydUbU5VAPUBdxdj6TcTpy7QQirEGqYnkL9Lwl3PrqOg+YFK+0eRP
unENPUNO5+gKssjUXKusuOm6/6Qtb7UNdOvNt1vy7BMQ0KKt2S0y0Ugqa+CXbjfmbImG4GiSDvJD
daUqU0h7oEH8h8I64M3qNdVCsOfoNKas8tAOI3JXKXaDcsm9j8X734t8hgMVPFbHyT1zaBENpPGK
avvlhkZKB/DXOE5pPd985HvpXnJb8PiqHK984ZDuq68cmbYgygm8GbyyX/V0Uc+iEEqbbrQi93/z
YVBziDIlXkv+CJZj7RBNtaR7bGr917G3rgD8dXhyNbrZpzEFVvSCNTI48ZDLnCmPd+9F+44v52N6
Xrt0+vM163mDQv4nT8CdKGbWnhDO9kiR70B2sOKC/3dkaS2v10Uv02Wj0A5CP48blpldH/aD/+1f
bhTDnFfeuGbsebalwt53ctBF43vnFz+jzViIaSYaDO9/PSC6DnclWSd17YMh33KkS6OaJktDktE/
uS6MTq7hwydKWDByIQHrNvxyBMcZiwexS+onyqK88NW8XPf58KlggHs2Nn+vruEN2EM6PwWRHIEU
IraNe05amzKjo1nl7U5nnnorm/E4GxNsAtbwuUoGIAFtmh0xZjci0REJOKE92gdFkimAOcYiXg5w
Nd8fxJO1hG0l8FOz/am9RQRDDDtw/66ne9fg4uJJbfl5qso79Li/+7XnJqhfcyvoDoGUrHVLnmfr
mwU14rV94YHvoeh9+ivlwuVKFwZpTvXkeKAK1CohdeKGzd9za4CDYqjSlVnE7/KpunB/Yw3SSilI
oVrh6Defo4DIfaLDt2bONpIv/deNeGJ017m2cFdYiG6Fgi2oPyxLYSAtXK9zTUboRNsSgvKcWCl2
LgME+YO5FiBqbpV6jV6BWmbVMMztcHEAJmIZK+m1t4ShVl/d89f+l30tO8mEktI8zNeWtgJh9lpi
dThr0VaJkYLw0LtbUikPeID84avRd+s1kO2CnY1q68gXYEvve+JvohnCWTOLQ3/mLKkHrD7wm1XZ
FhVBmANleZkw5NNO4tCFzRsGSnjeLWhots7/SHyzyrujUJowgPPlZep5mflnn6I1W1Wskce9jLjD
mYPaw+XTl72DRhMvgI+gyxj3iVOBiaVMa/OaoU/DMMO5Hf4kqozBHUanUw4DNHhqZcHnqGht5mTP
ZIOMK2AUWfLQFXa2SA8nZflpMOCK+mGoth8v/wNEiJzKj+4jpM3r8q92Q/AI71NQqPS2CVw0NelE
yfPEqwLUAuwKe+QlTKInKSqLdhX1o83YDM9IRhDnnfHAkM8wWfSsWxKf3hKYL1BYmTDvaCFF6PPN
kMV+tWSJ5zpTWP70ekh7rVXd5hux8IurTrhxF06oCgF6lunm5jQGzWIFh/Dd2R+zvy/9cy1g5Bmt
5sqp8Pq9Kt2jn9pz8pjv6j/FLfuRCaCKEJWQ+lnvTbZJmnMKsdkG4qVsumdYk2NF5n51AOuMs1fz
RLYEfcyY171S6QG0WKDgyks1b6e/o+VqHwh5dhVHZDsvA9zIu3brnkjUqzwfP50oASw9av1MVCAr
B8besMpufehHOpW622z8ne98nVAVRmSTjLgYk1X/Jm0fhp9v2HjqRHCVSidBQuZp4Z+2AZF7QzVl
GSr1LFDe9guawDLuqilighr52wMTBS+KXqiWWy/IxLrx3rNG63Fnzd2gLZihpyw7t1i9TJjwHEHE
nZLMFEnJ5XnHESJwG+Sx0pt1g8RS//tbr6/UdDa7MmvoITli95MNpo+QwYH4yn2ID13nXe57ReJR
BY9pSeOhpl2Bbfn2szgjyASKdeCiyKTbJiw5xagS3rD4XNOjhuR46RbzukAQfJJ0Eb5GcPHrvkvw
Tv8QbXXaOVA/+DG8sXcBEqA4Lke1S3ISI/FFHUPhLMBlW/KldEnLE90F8jKlVD0Fd6LfkULh+qk1
CWnAYsyEEoQQ9Vz3x3o9AHkEvr44wLXNDs91A5byO5YO5HnmX1JWjS7c0glVOzf8f/P+wTiz6Weq
6umCyxX94a22yXg5bmu6mzoU2a41IMMbg4L35cqeMLdB56muvFYr1AZYhRwWpceVaTbG+4FLLL+d
euflDF3LGpNuOQRs0KMeFYrk65bLQhIG/DgE5qt+iZoJN20NRqJCorUY8d8WucPiDKyJ1d87AjmT
cBOj/PpxVa9+UkEjYqANXXFUbCaaTjcXp0z3FlVBZPtvWAcRLMPY8gFl2bF/RHBnO1iqgsZVn6WN
Xhr/bVAcYRmTQQbu4ynvfCNDUnT4SkWUNFpHlxdOsu2NmuNBpD4LAEEvcXlN9KcR0ZtiGeujqrqb
obXBCW9Nx1Ivwp3/Fb5LnW8i5Z5Tgc0tt7RQ48gVbOlzGix0Asg+GxAy4dzf2OberciQk/1zj4s9
4MhhcGWTwcXE6/A6mH/wJP6sMgoNQSZakDpdj62bwdmNe6DiXEgWxxw/AFm+jqWkNFq66TkiZiu5
DwiW4ecxDGhu+DW9qOM2Q43A9MiHydCZ2x7yN8B6sk9SvN5vG0CX0W38yIU1ReCJE0QzgWFhbwIG
Rc3upmJPNtazAwZzs5p6SCdAVlh3ms+1/7l53bD+7knclwAv2jNk3VzlGD4hhGMfQ9Vl1i78UXOv
BXAFwbZr6UNN4/XYPJAqtenvZ3LwYIRSVkB30ox8BIvnmS5tAQnRnTmHRGz2VKQ1avA/E+C/SQrx
2UhnR+R3P26VJ+wO+YVU8yFjQn4NsgwHpJo4ASgwYiJn0yvo+VslLwe+4anN0wAjY9mI6J79GkIe
IM3uYXQ7PGE/ND+roynPp60vKa3aqWOuh2OZsrM8TWpzRyndldsfeYswNHmha4+qqFzFpUS10PTg
9wekWXQXKcp70dZHthdQE7ZU2ETWkBj9uJIb9h1DuNB4M6ZX+ZixuJABDjavYhHkSJWw61HEaQ5+
noShX4MOueoulwa8YZbFrKusd8KHvnLxB4Q4eQQDLDl2J4Zg7Idet+6AHhUM5wOQ3856wncF4Mav
eH4uxxHX6xAxEOz/gI9Z5d08Jl3lu7kTM8fGeSeDXVThC35PJMf0jROkKw2W/39NxlFB7pTNvJ4p
Rl3NfUhtw9uW5Ng23pQwkHsSswCCLwC60ZWnJ8Cq+UQL9QPwjqMNkxa6b7lA+InxlMzol1dEKuqf
XsNt++ALHRABFj+fOiKruFJlofhNNrZA5I6SYBBiz8cyWu1Z9oOGHx9wEvW1C9ykxncKUbxQWZUL
CSpAtojr+2xKpOVxHGAqClhVdgpAlcikNVoA7+jaSVSyn2rtcn1p9wPXrLAo1KDRwE9OmJT+ZsAM
cqRduoWBmHk9CKRYACAlIOIIfrpceEMkUhsrv7nhSWh3uOjFzxvSbZcYO4AX2boV8iq4JSrcdzy6
TOCCdVhBFbptujL+60uT8bk8thSUwJyuzQH70IhYW63XULst+YJ63UUvLmABWIR6yANTHdA0NCB3
Q6yPQsycWsFaDTpac3+cymE3krsr4ZmvxhE1qBouZNNjtFePwkCWqct0Tn6/VvzjHg9cC8z7JiHV
fLGKu4j+CcqFY8QRFfoSxlWzaf51cniqkBcWQyPXdt/v75iO8kM+TA/MC1rCpf0rZ/6UL1aVy8pi
lI5we/selXg3m2v2i2q2d/x/BHCILrl/qn4xboDRoJsqreNfLKA6KAdiCXbOQ4ZFMwYdieTNXC5q
Lrl6Cu+b2KchLBrGvaB5PKfnNQdz2Rw4gkLV48awSxRRdrt7AK7/a61pxK5NOL+S9Zkhkk0jcDru
U59/7Xj0uA7s9qPnpwbjWj9too1TqZa/PTGDO6uIQ4JX+aCVM4R/0R0fjAyPeDubOJmgsNbLl2fS
IuHx6YLgqmOaCPpsYYErTKHcebrkbL1XilSzVw2mwyWx+FESaLIUchePR14bUT1T/8iQFeFT3eMs
YZnoi4D7TuIvAdhwM/3IC3cgVAA+yHDHX/d3j3JQLiwLBVNN6RLyahiEIavtK1a3jLoJVE+yIRgA
QhsXR2dgB14Vq0lywNC+a+IlMkP7tL4rsvm/Ze1vU8x3Ne2uQ2VURtG9Q7VoHsFPW8zMWeqL4Sk2
+GHgJIHPWEz2g1rwWuX5kGM3sTWgfe2VrZyJe9QT51+mZjkzRwKiIC4Qv0Yy7Ntgbi4Zh5qpMT+2
R+4yGprcIHaZxaTK5CfYMABr+rp7faxZyRGsVMKZPERh322AzDj79SLI3FDkpg3x1FT9PvqvBQY9
yGUjN9QFilHlCVR0T5aKt4/Y+cdp8n2Gwi5vfRu7DIjFxUim1FnhG9pFDed7mwFht2yS5gXA8rus
BZirvYcesGn5wXbjKUBhAzVD+pkgSBuk93y4KXrHahqJTt9ng6WnFCt3Yk4/Wk+D6yakWTBLp456
F3UzSIS5NLo0ag/OzGS0uvjYUoh+F/rfNg29+XvIkVqHjYMMq51fX+hbUICb+CnMBNCS5LMSv8fr
oXE1N6RJQaHsAbxwZi3i5g1d+Yq/R3V/YXiNcRxpzusoBp+0D6iEcBdh6y0ZcNlfbMfHalhmb9Xv
bE4Z6/NNp7s56C26T2qxMjehJuMl1RBwMWrkE/J5BUUE6KsY1YeYZNX0djtU3WHzlkNF2NGiezFi
dheQx4v0fOkcXZZPh5ZasvPFLrzYNDoX+m/8jdMKs0PkWTtc16MVAPKCAjVA2NmWvrzaM3vViH0V
judih9hirX6d0/IYiKZ+NoynByLjTUYLNARVIXCIRUQRN4ZVOjwSeM0YgpaVc93kNqMiC8q4arHZ
uQbTFFWK4EJMuy9K2xR0K2BIJQalByx4rOe9ThIN3sl7+0VDEullDS4091Ly9yMInRquwQJxiUUX
c4jcxYSp/B4BkLa4926ikW3GDJk8WwF3mb8nEd6uH0AlopLOYnICgI4McNFFXCo3YtbKWxZD/tep
W/ez5C30nQmrtZNDPQK2lDLN5UvwxOkefDZC/SmaMA84GOvHFKRMqkqiBoKMDfG0oCHC98e3TdzB
64fRYyXlUE03zFcTLe9Zk45N1MieA1Vs8P5jQoMtuX9auHO//i/PrwNEMz5C2FFYn0b8XGALoyeJ
ZIzw6bvXzR8PKU5qynMoJ23fb7WXC5CpKBZyXl88iEKwPojNUcOHLlVErs63t4OsQKC6ngTnapOy
c3VNeH8mIg+svd/Zvhca01dBdrBmFPMSNugL5ck4MsXUKeuyxzuPIW+JAE5hlIF/FD4ERtJ77JRq
BO6lv9u9Bzem2C9oeI5r3KjNzhv8wEBu7HRVbMyYWJsOltfrXUXwtMV9079UhgJ1qiOgxrMv/SgN
UZncqO1OkKFe9NNgoEQPtmpFxsLKPmSkXxOz/oanYrp5sv1y8y2vCfEM8ehQllRz/1vFlw5A9hau
TgFK+GafoHxqCKX1t4hz8Qm7wk0R8w/vK7fxV088tkP/NwZGuLrS/ECAyRRjm3o+OXTFWURFCSVd
kiilWYQyWi2nPF7uTLLzDoB/F3wBLYWdwcJhd+y2JHxF92WONeQJIU0Qb/7rqmmCvjAzELlFxeJs
d4BNy0i+ke13+x0Z2Nm+S74zfZFWtYO8LBLnbQB/0BJvszT40ifX+RIeRlltKM8bGHWXlqzaZSq5
RH/ND1Lq7YjyL8r/5s0Eobiwer+1EhhnESmr4CsoFrh4eIVSYSr5i0UQ+B5YcYC4g1aZhpgV6wuU
mHE5fGafFOFOYDGpY6cFTq2ijUP91a/tdtJAIuYEJiV/V6C5rKllwsHuavR5y0spy2Mgz095IYiF
s3NzpddQRYE6d4YwD5QB/a9lZwzORt2NLLSPSS0tYB6uvbE81GJnZRF59ywFQupI+i69goS7cMYh
dayMxPzrPKiDPwsdoSuO15TnIyWyIg/UpeZJ4uBSeOcJXsgDk2cnefQ+wWrsmMq2IArDap+xv7wB
Fv0m2tXZFDXxZToCTsEtb33f01U87kv0V/4QgVPpm4G99pILEXdhvt+sPn7dGF7Jw2ur9jd/8/cl
wyI7Ii/JqbbUYdhB2zWW+wy/HrgSR+MerSyKYkOgJxXnPEdKi3SLgkdqzPwVcDocOn2uTgiU8Lww
Y7os6SzIg6s9wHc5mwPn57SwuNIQ7fvXmo7+W3pjI4K+h37AsoBa41ad3HYUK8HSROeue3dwa05U
0eTSHjUueNb44tYTZNSF+KycmR9Kq0P7m8K33Bmu01nFFrArMYN4+uq/8ttRcwlgEwtmhrBUSm22
RIZEidZK7mnlu5Vys2bGafteNp50AeT9rD3Uzp9bC8BTg2t89L0k9DI0v9rE99IrxHKJZtMAkJsX
yXcGlS7JMJ5qucBOoP9crim2eKdB1L4S7zPivROD7gfxMIG9k24ti9ttvRAy3xujBJWWQw5o5Z9L
jcNiBDUzTCwAxecYjo2v2gvt5yBl6KEeS70WBoUzer8FzywJeo81e5TRPac2md1vhyKlGQCkEFZs
YafMwbpMheT4FALPE+6RbWLBXQ8RAoJ8buoj+ipLmqTvv7wC1PUierl5FZuVoiTZsbGI7rbehj/M
uwOuqwy4KMVL4QO1TGigpW0X8SGo9bbipZK0NbUsAcFnvbr5y73jivXL0A3hwnn8KZNtuTjvTDvE
jITKNvWKu7IHvyOzwZTcC01vUuEwDYgNsvermaq8KtYEKOm4915ey8IJjzTUBkDfIY7ahAm9odgg
/fX/W+xEq0n7JBk0XptqKkSnntjaNbqMqCTe9qym5U0MLi1PVdGlHW/4NQ8a74iJwq4DsvYylE6p
dXwUd6chmacOlPWCIVibI5x+PcKlU7WtV5qHukRG6pgnX6gheVpf5M0u5hyzMcSoKbTRen3Hi+LL
jwL3/908lBsGg4cKST3/rUtsgyMYXIiAXYcAiwvgqXqMebK6pFRe8c+Ec6fQAKkZo+r+/7e26KdO
gSPfvyN/EPU2duLw7w6wR6M12Gm7PaY0YfdouNeJ9mMyFDcrYL5RgH5Xf3S7wNZgwnx/piQ3LcqT
hqbWYdc+QllS6W+hnzA1sqCrnzbCQC2edaMFC+vGiWV2lomfWMtn0CrsYiSxRUinDCLMKEfG5D77
+fU8+nktZLFeM3ZjnYgEPlBno+3BfkqDvXEWt6w1iC2UvI1o80ROzrfrsuNbnq0IzUkz6GStNJFQ
Wt+m7yCMWLDgvHCO21MrfFFGuJ8gHeWe9z4DmKo6IN9wQGqHvhS4LRT2sf6ntNLvZbK7oKDbaal2
/54h6in7YTADRoBdYizOSzeG+sccG+bmYQ633foRxV75TMvhvlsHa/xEwgSDA3l2vFxV55xK7n25
eTcyp6iTptirIot80xRCSytXS8u70Ra6grOZ+EuZM7MxCMkXTTvKlhlwolJH2lmMYs3FrCPwHR/p
tktRsEnNv31t4SAcWxGiAlOjh9mRJ7BBgi8094dJI1qVQo8e6tAxdJnM9qKWLMCvjgwFKgYybNZ5
aIJamYW9VN9149Ih5K3RFL0wx1vp7ydSuhWB1oNo3uvn+yzb0qFzAjgQnwTeMZO6hGd6LC06AZ5Q
Fe0FL8785IBgisrNVIwAlG9nry5/+2pwxECZFTJxqhxY/Yn3oBkMlsIOoF9XjeabBkD0QyFvyT1a
Dtp6y1Y7RHfHKOJAkPX0QiLz1Y63HAlBNbYN/olWgg7h2hLLEnU5m7uQNjFYQHeC/L4mlu2I1PWB
8rT4uXycAJAzLz5P851bbBItVY0JAOT//Qa9hHZHZsG48WUlKldBezG5zWdiMTuclMQ6b//JnDzV
JtGySxjdKO1R+NocyQ3qFgRfw52zRKwacqOFfaenVVPygiaInQkWGs9+oO4zToCGcyuQpLHV++O4
8ptEXITxKNE04g8/ajmDiYxFAa6peydJXtQb1HupyUa2dnLcH5EymRAFKru10E/zRVOLVeNzxXQS
E+ZpAdO4zU8dNv1Do7PiB/tSaZvV3rghkzvAGO7U5qj5GXJRSokPXIX2VOkiozBgj1SBq+5rOYTp
ppxc9+D7sx2PGxK6GrwsjCBBlMu/5j7nnJ4mHRgmRO4hgp3S2QEzwPGEzZqpLwjrFwv2FAKPhdYa
0bVDCmGXJUe9mDuzS163PcMAPKuLSRP7/X6mCqLeqYZky9Owd/8HuPK1o2PEv5GuMHpQ8puk8oWY
AcN02NaCq40p8OZvl6bZSgVOzgkLLL9TgwAVyE8tMF7/Z0AZWusGw+/CMVJzYF4FbEF2TR968FJy
n9PtEJFX49DJAo/IrxG4scAhcwVqj2y8JpzfLNxhL1QIjRKowHW/FrVBlOz81Kab2jJb7HhKvdmg
Gs1RoEbxMf3zioek411cGZm0ZR4eu57zKC3mMdavUzGESE1WjyHspjknRbVRp4XC1JcViLx/GeIa
D4FnFYKdKcRZdXeHWka2wWnBStbBxgK8j1p/QF3W9KQgyoipnrgeOoBcICyfaE5UdPmO0Yhdyu9T
hze/rEkjJIr6TeLbyo+tXLHq19+1tNWrWPedBxaeyZ4sLJOLn+L1iYAsshH3PuNr0dVrAI20EdBH
M5bJzoZhLpc4mr4bF02xgILMzeT1TVVlpavmmEFzticCJ+ybdtlO9s0uSIQ6XJ52YlE4Yq9R29vI
HVaTIwEwJuIQu0sSzKvPblj/YXM9izG42UMJo52bskWywUf5jTpZTkM/d6n1vRIYsbVaO6k3ESbw
sD5wh7gZ5DmhTsZDxw7dhINlXC1mRXAone2KaQ8QAxat78B64pjNz8BlkXwiYsXwY3v1wIlHcgFb
HbEY10FNDEz000fExTWzbBL9TnIEentc/pRektIP70uUO3oRQAS2p54QxWalAR8pKNz1uk2HzM/e
5NLUw3BwNhgqsfn76cCK71J9c7zVKlvRoYSlAkhejNi92+cpwAjph2bPLBNkLtwkhAcPWPgrZSc0
4Mfmn/q3wnkIzWgtVBogrGyz8FZpgfBQR7RXNnij3LsHUj1lJ1rLv9nr4cXOYT8sRVkcKQ4jYqDI
aDxh4aNIkvKr8F6uIx3xfwCyKZ5gF+wkJvNWIYNNik19vD+r45fNawpoGe1JiYfEs/K+O2AmVqlL
LsJx46vJn7r2ybAG5BWgV2/Q9tq3CeVhu9SZ63ypJB2276JalI1geW3ePu/o9avZ/uvl+i7CM2h0
kfnZFaDPHwvIQ8hXqZrZd2qh5Z76x4Fn1QBGLObI99V/p6v5H0c45RWInZDX6qZuvVX8PLxQYJG0
a4EuEW0FwO3HPEo0Bkm1ve8SSb1z8jrCFHVP41HdCKrChuo0rxxPoGXFtsbngw5fBngBKmsbdXWm
OQX8ijaQ/xkkgj24oEfZYyNb13vC240B5I0GNrFt/lNc+6SqQlOMKAtdjbVUPNqTvf5SYj8bvEYK
Ge7XaSrwEj+LwcDUYuQ6RoeWepTlSLWdakVULg9l1TGPtZrBckgxV6rgGI1TiQd+/v5JQg0+7aY9
ASz2z4yuKQhDWwHdd2nDd/kuU2Uhj/KYPZF1js6xk+WQVx/6lNJSAKljp4ed/PozqmUqYXCpXDkM
amifWIUq1ChqhZ+uta7ObYi1eC87nSQ/NLnWrzCrvBTGBK2atzoAsjOABbWLxT8dxDb4QsvXN+Zm
uaun/Gyp41R8+QrXqwqhQkrw2dxROy88VgXBPQVWh9uyWAqOoBqjFQUIp2aj7JhDNadtO34IF9Fs
+uydSFkw54aylC3Hg+s3F6ELD+sot4DWu+dkQB8YriYcMbyEVHow5Vp+3KhdMLpa4vC644PbFwKJ
mNU3tNWywAtw9WQBpL0uOwPJI4RDfRav6S8INEJL0nuuvKPwyWKBzjpmZngZPu84E1XkO2DQm3PY
NcKShV4RnOdE9uUGY4qyQsmMfoskgVXHhFr+nAf4B5+T1CLrup6VDUhFfnRL/T5GdB0cAjMRu+I/
btn6CoescNpv6Eu5tdOW+ilaCHokIcCN3g4DhvgihQNoTS8o9oDOsBhcLSCZTNDVMEM8+fbFLHvd
VXs+C7P14z1CCB+KUsRXwLNmN2B7cmSisqRD6BSw9ZjxeSe8RugwJ2m+qlVNZ/+LBG3KKO1sCWTq
5P45uSJQBrHeQzBsiPZHC2AeLlTrUH29BLOHlZNZZODkjyu6A9JkFxzbOKHCQWP/gz60CKvyEVFO
amOPuNH0mZ0lgZNnJ8by3t43rlAN9LW793d7ruo2pGle5Kht2szp9eKHQJkXaIJeLr6LlJdtwrYt
RYGGzs5a4LAurmfsCVkaSgQdWRCYglgQ6lYfWCiQPZS1yixu93CIpjX3MHlTQkdo1Gwt6hY+4oon
q1CYmrlozu3yyhRuyRwFRNTV2vl0APzgu+OsxbzhZFFspr41EnTqTa//JK1DhKVmdILrfy7WwRsZ
Mqzm/XkyB4FzOgc+cBOsyQJp4+iDnIX1VwCIbrXTkxLuim2zFhBIIrHeuJLROn2vosZQ8J3qiFsi
dCeaKBMc9aYpfos42yx+w7dqwmYzZWYcYwy7if41cJImRwJT6ZoMi7bk0L6kt1lkvyLA051kq0o7
n/UcQIo01Icmy12T3Byp5zzFMf+FfNKb9KwO4c5G02YQKQqTzAklAFgpce/2UrhQexnX048HNbQv
j/CTnJZ232sAToF/O/q3kKDoY+YpQ7bqyeUf9nAVF58NNy4FM0EBxN0ganNHs3AMK4a3QDw9CJat
5htKmJfZjftYrT4WPrQbKcHFXxR7rt5+K7FhKtKwVf4lrTGoSiYBsZ1wsh4rxQLKDvAgbIFWgE32
7EDE9ILjE9T/pOfYn/nrTEaTmoaJamwcpkAFHLkazG90iGrDC0XiBT/CWINA/C0RF8Aputn1uJ8J
qeskc3g7ZlnpcrfQGlnO00Z3N9E756jQfWysd9SstR57D1ndJFtc7Tma6XAYI1Uirk+BW/gpcbgt
Y3jQsahXCx0t7lDsl54UR0jkohJqozMtcRm/lqPFWZAo2VcczJ4BeLUoPjf1P46DMnU4IR/0Kqoc
Xr4PQqtdfX0ZTu9bj3Cm9OSkb8tCDmSk+EZS567pMgdlquYIXqGCjCQNyDi0FEsaN104ZsSloT2U
s8kyxoQLqSm6Brqt9guxRg1BjodAwJ1rrG5JzCksSto+V0erRFWPJodc8KjOoT+9S1FqMIdh1KsN
BcSrbARlv/7ywMM8HZkjfMUQ+KxfjNsnc5ltBGmAJkePOtjNnEQTfnGJ+LAee2F0p38qGzBlH+0k
P/t9/paxzpVO5x105vVSSqG/LSmj7Q+BSp0psey8nXIHa85IiZZTrqHxxce26LibyZfml0dHG6j0
Se0ROXz4OXMC+1cNYhMI/EFq8UQGcDubPsCTUqk/W/C6JbI7nhPKxTGKQ7GN65eOGYgngIHqmXDf
Oryu4oj2CFErDs6H60H8zDtZa+SerxuQ3hGst8OBKikzWieEI0+lqNqS+QWtvvYRGlarxNElxDp9
00ELKl3pOqJW2/oh5SVjOjlL1tATQ5WGBMkq7uwKcTq7+ZyTEeqepznnChdjIiNONL0Mtxyg+XfY
Qs5R4kFzekBGK15PPsaE85FX19QuwpLmKf+WHtqvfYulhmNOVVXCd+D8IkbiVAQlB3TI62XDzcwv
NeuGdQL25mFmwXtJ4hMlrOpfkqN45d7trFWE6HF/0RzkPchRLxQNCgqYZjPXhB6invTfdKkBrR40
+w3EyfSn9d7ufgTNN95tFMyX/bCi/IoT3xAyqdBrI2g1iOlzBXhNvO0HsubYKCfhw2R8kM9feNR7
7t97w20mAYWmz1vv1PdXADqfNO4Yo2BYYzXdnP4e7MXeGUH30E/b7tgHf5EOLUKHghf/dE04cMI5
17d+1FlrlFj2Lkj3218akPGpHUR6zJv/8kk+bMgy/tr81alUldv2cFwfMbCF5+/goObbF9/e9uou
glAJTv2ipl7RB6VKwms4sHvGuhddVjPqxbhQ3FeoktvFDuwGsH2DjxvZ42wf2Och1UJE0Z4WfQk0
24ZR797NqnHW13hfgMnC+SndN301fjngNmnMpFob4SOd/BfdjmbpkhkGUszU9CIPHbtEPi8ORcDF
NGO2sq1S69MCHVt141VreyzieNo2wZMDZX+ePiXX1QD7HpdyZ9o0EmSm4/K98qHOBXp7qhGquua4
hmutUYNwXBvtLtKgbjDMuNq2p8j8IfChiZfjApryiPL7YZMKIrdJb40ZaF+3G25JlsrjNrMEbAOF
qfuPQKVaE0Zkn+76CsBi27jEVZsu4AL7doQwzCJZsoi+w1cKOozhYLDuMFs/cFlpxsc473jJBE4k
s0ceioBXwGB9+MV98gaOFb68z6ohq/kDl+Mb7ivbXgZkDoEjWXMyHP6xflSBmgN7Gy/4GLWem/jX
o17x05smhbzknED8D1hIJXzKW3qxMannLRvi+XdCTY/0HNPlm9WEar4H+xihJ2rjelEN07QOrr63
lSsPRD634voMQUZzFe6q+3G4GQESG9mTMzr1MnDVf57GzvYLKv+G7YcTifRGnqbRq5db7Pj5PUKM
DruqPuaGQx3ZvZ+YR0ZCeSHhl2Ia9XOEm/SeSZUPtBQSAt+yRu1lX6fgG2QHqzgi74gupzuk8nNC
WwNoxfrdFLGtC5SGfdNA3tN6tl8ZusvUyAW+JsMvUdkr1/PVBKF+L2ewH/I9IywjqbQxhOvrOUVA
4xNYz1Im/IEyBioY/I4apc0IDSHk3vKmSRBONZc8wwL7XJPPBYgk8WrkCJ5YxpdIh5ngeWN6PXJF
JwGJzTWgXrX9QWTUDYt+lvk5T2MgrVgifT0CbNEiv8WzzeXSOsNTXBKWjumeOMi9UIHgOYqzwYXH
CvYEztIOBrUwqc9o876EY4eGzOVBZZyvYgLMANfEDnKbtLIqMdhLznKtzRt53Ovd9+9VraYVaO2t
KuWyW7HK/WXVqSSyKWEq2HASHNawFaN2J42xUlWCWIoL+f9hg+AFyoX4Wyt9YdwiU8QSWebh5DxY
76xgJMM2zL/8xbJ0J9w5jVHIACG0Ea1K3aTMF9eGINah/vPPT5LQw6onkyECP44+K3Kr0Ghzalil
CcY3x3TZ4RuoeFjR3T/VPPUdZQcxpkv4zxPZFdocTi7/YsFbpBqMGCkhfAFnMpmCiA7msC0Wto3/
c+kVZABt8GfEopcUwjD8dEqILzvx+cIWs5Fa3cdbHcnOMszo+F0i09keBe/c//Osdi/35YXAFojJ
ZIkmlGfVjIJ6f9L8jrASYB8O6PSAZHbxIrGiinSKprmYJFJpSwbfKxmTjyWGisFqQe4Fc80XZH8a
eGEIe9oBs5dHyREX0IOEKYuwAZ71Tg0Pr6TE8poIbNUyr1yaJIFCjDBS+dnQU7WR66kDuMm9vvyn
dYyZQ8Cb7rS0ePjsxu9YQxUjABnXHPB8whkWXR4qgCz6lCO5Vfdamm/Ix54FfmpIasd30IUOIeeu
h/s1UKq5oK+AFwB4RWgJCvgXJBMcFg6lHz6D9U3NFigVQSrikM6d1lDn2bUOkON4l62YdOskqWpB
WpBYp1sEjo/FneOKqQyfLKR0v4aytQvCePIo95KCnEMLys3tHngO96rE8E9V9+2G3Yy7+kGFI1eI
NUHGaNTlSaNwnFW/rBAesm4pI8yZLp/4t5r5lEaazo5BKq0FEZiWqQqQBiUIlTtavyiUnLGlfUph
QzzHD/ZtU2mNIn+glUiRCxEYz1js/F5sY9QHAD6hwKmHUbasrohL7GNREqam6vIvLoZuCXYMwIpd
SzqVhrbA0mVoZ7j59SQvEAriBo4mL2yzoWVvrNKdbf4TIPx1J08+dWHiD8QX1S2Pl0SYLB4vDQiy
a8QzEqiesapivh2PiwpVTCNaspS9LGJTHtt9EuI7JZf275gKCer/3E/MqEtJ5OP+gCHM+ZA+KRkB
3Lo2GBkCvOZEMHce2BsafbXX0z9H/uSzWlK/yKRnE1iEv5u3p+cCjCd3mW4HvElik42FEWNuKILp
uHgc8x2K+WfdDVEAwk6eCz6mORpo5eahsXJDC+m6FRA4YmeEmXzuUftNl3Z3Uo7ymXgQGrSpyEFI
lKHUBrc+eD8cresLSVEBDw1xUVXb/ED6X2qaz76DYntrmOtC1JjGTKx4SJu88I8UXCWD2+dxTiNF
8hCXnonpahZla4ssiJncH85izMawZza6Jq2zWFq38NLHxkyF48TNilfU7BXwtNu0UMAI4VUo/VBT
zhm053/D1St6PtyBEczCcjBVKZDPTeK05jw/fgTDDvQ7mIhOuFkh0i9qA4iMHVeAtVkS3BTkkhAn
UPnxF1rCsjy8Vew+oSxYQdHODbtiTsLmtuZ38XvB7qO+7gs2Ukq8g2qybpUl3KxWvD9VeiTTqS6K
FTJg4gqlx/E2FRtKu0SEUYQ8W9oWJgu4otzIEILkR/vC+DCvMq/A2g7PcaY=
`protect end_protected
