`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6336)
`protect data_block
wrovcHZ5qwQL2M/nAHkX4bSVoUptwBOsC3KrcEauQpvfqtSQ9szJpHNcg9eRdwOOzbYZn9UXWEc4
P4H9HrDsM01KV/qrnwKrORL0Yv0jebDqFfiCW/atAJHmadKpvFJwG1XK3ciLl1Eor0LIO+TGPsnD
brw/DsSO4Rappgf5WYxQZpVplRq4LMXfNJv9WDEUr59jiXTEqrlkUJRdLjlR/1KOPlL3I1ZlNh3C
P8b2mhoFpzbYNdfAjerAOOtTLZENmsnyPKltbMCWUX83YRWudR7Cco4Q5POszkQboaVR+q8cN7IJ
YEb/fl4QQVD3gywZvrocCK8Pt6CGHvcqHbkKhmhljkpFGmwQVj6mv8Kzhqvb7ItEYMQL85XLWpSD
VgItDYGswSn9FvTjJszgqgiMCRtPkaz6W6wg53koESufXqodtnSF75AKlpeoHsn/9f5DdF5qDGhZ
eW8eirnaxmDdknencD7cq6/otLBTJIz1zpxpXb1gkAhpsFw4MKEerfFJp2z1qnakWWY2qj68JDo6
eBbHpGBnWfS8uulkhoq/bNu0GKv9Tv69Wve3E+oi25TwwUSQm+2NcVEgQ44qI/EI0ozJWnh7j+yP
1kLlK49Vo3eDOYf4pyilOyAuZF1Ixu0kYeBr6VU2G+ptreugvWGGebnUtspfBatEhpiasmTTKqVT
qWllctTPOzVUcRl5ZkjfPS0+3qk9mNmicEYaRyk5lt3THY4aQpv9qEkpvBOYcnXl4N3WLwCHqd2z
ML7wsDMQmGrM084rNPfQYTwA/Zzy1i6STFaQvq7dcc015DFkISlxF4y1IW6AaGH3pe4GZrxCdxd2
KLMx8vWLqAFQnmSIldOWU0pPi7nrQdeOV4pB+ks0hIoYjZNGQzHkp7oOHFTmefD5xS9gDMRVwH85
1t6NX3qO1lQqgZi0Ow9qnC8I/C3PfDJS+nvxvOs1uoB51+/0fb1W6rLC5Z9XUwycGPOMmmKlSN1t
cGVTtS5WsrXlHkTy3eODi8ah2devtu652EA7iqkxjIghUeaHiecxqlyKdGhhlqkR4ARtbRFgcPZb
BjcVtJsKYzI7JqlnXmqCfH5XLmJoUJykHrFhV/zK+XIUMAfkNFgRB3YN7V4S/nCMUfcQoU7jItty
rSns1abHHjpDTizLE+8g9R6qTTRJEMA9AVI5HDGGJret2T10j90p6j1OT/gaEU+hyNfvajVACz41
fVAEvKavPSC3UwvUvxHVonIfc0ttaxL1y4v76b1f2a5RD3A+L3ANowy60dubITaQAfvAd4L5G3uL
Nr4zEkDS6pcGZ6oLbECAYaN24z0EmvmY4aA7bcj0UehB8KM4Z6DKId2RPJ6SczrTkdbxkvtQVLe0
lOvJXIVmJ1abhVM/uEkszg3BIeKjablL6LrQ4tsZhj3uQJfG+uUUSRPThZCRdOHTgzPNdWkrlHK3
vQHPUOsA4cp4kSZCrkAdQVfmKhbzo31Dqtl8hQ9Qe2Vw4JBr2V5aojJR2xW46UnKQRgXEVt5APDA
w6AUD7j5d68vHFYK5LycUsn/1DfigyHbPCfoIKppmRqvY1JYZtU6xeA2trCb7Qejmvi23h441PLx
ok1ODHOqKPIgT7MgTfXI754+SqDjwfh8DzbjoItNs4vIhnDgCB5riXrFvIxGr5tBm6BNmS41PV5e
8OoHf74QABGnV/oLkhxIQPsEQSZ7zTmtB+l6DjuqGTAEUVcf2evoHvsAZ2Jg+VwnFtuklIKwoTfu
XNW+36at+fikeOf6KNlcNyarTDZxtLzj9NMEyrZwrWajoMMxVHRBJ0SPARnLIik0lyUNdVPY+YLo
R5btjQQnQ0FWnXdbu3g62GY4KecMR+g2GPyWo+9ha9aLnlmoMgIfXluUXo1mng5Pp/wtwBpiK95Q
hIE2ydQmae9eaLKkedywn0TSHyV5Bh+4da3RfY7sbDFgYoiP7NezLd1mIzl+RjpqpGGQ6YJ3+MZO
AkisfMvUeWMSdpG1PMf1tu3CGzUgc0l+jMUuQF9F3eftnphawXI0t6mJ3YGeMjrr5vWWCzIKopKY
tI1o5kOtsZuj5+vDNFxI1WV9HzVo35jUIU13L3+K6TTned4k5NJ92uC6k94kGGYHm9/wBLWSHhVg
AV8Sr2TY+MtiIicrKCNDy2yWQpHTvN1sWs6jW0Qs4ThCY/WBJK4UTJ1onFw+ZAyVgJZBEBMZRQcV
WPgUQax/o5eyhJMymSmYTN4JojXwvpEov23guEoSR2rwbp7nflhB3chEPZRIzbUnTsGAMZ3l0uPK
pRWABgyrbdRAbSsLOtE/ey2399oOHv9jLc4HwIej6HvBkacPQhRmzNsjbvuYBPYX6EQufEQzQHjR
j8miLnGqIuM8wNqmkJ1mTBgdwbqmKVPSeUTxlG+QlrdvJCX36QBH2nF2W483qu5WRDVr6xpYLgYu
Jk63BRFUct67tpBFxByDaN4b+PjQKYd7iCc31ARU6C9GFhH432XrsKgtWxWnRNM0QTFnsm1olgbF
F+mzcyAwWZ0T7ZPDKcRpkmAe7We5YNIDv/UqBPN9o5DEjoGsJH/GK6T58BzlJUAFawVHih3RwRuD
SjN3FNUFhFHKCKUljEX9O2TiAxAqGejFOJ8zAWtJA+qgwQFty045FWLErPj2Gb/S/JKkDXtNsK7q
7gKzvihYsFdD0wrjFObY4dvGGOOVYuQ39QegpDA6OT+UV/t4HZPY8g0eZ7SuF3LmbMG40SrGILPs
TYlOvdvaibMDssgqi5zM2Lc06B9Ih0CBn5uXmzmU+T/fnQFxJ6IFzVezJKtDYX/5kzexz1mVBJEk
d9NoCBNdhWtJthPoNs8KoQyHOJpER3+8DoZcvhv6Ho873QCPSufxztkNOYL0T9B6X4ZvrrznCVB9
wSRFrmMT3SN5yBaJsrxLtwTZ31TBEuOk7XPye2aXw5WbeHT8SZcH2Yhw/NqMO06oJJbOv4IWo2Uv
YLFZzIJe1DvNzmgoNpNF3j70t1397A1VPNrJyglhsoyfZl9qbCzgxGGvpwPIdXq9SU/E5txn38Kn
+cEOuw6yaSlqoF1dKEa3fn27qHTXG8yJNUBrUuW7tGwyO63/69AxGqlPZvodS5NsTv2xGkqh8DaM
AiA9BzQlu8rPZb+MNzVNdOvjvO9JtVJpP6CiQX23V3ZE9GBNvvyhAGQqDC449TjbGjw5bX8fpjFO
PwUBxTahj5aIjYGC/3gtjULPAfOF+cDbdJNBu+SoEfU6B2VPGUd043TTozF0XafmG6pk0NdcKz42
hcmBLoI0igCy4y+on+rNT6ivK4f8Z2+ipj4Z2YUeeykp3QrzauDuAsnJB0XU815h5niSMm2u4ZAR
/lbIdDLMM4g/2eLgNU60Frmyy+ddpElqkpCefzuC5AwUTyFJAxWRMjGMb26562PbIi0Dn73J1cnL
lMMH6cBHoE23D92150tpCmkLv9cULRY9pd5BcSomDgenHX337wFl6kNRJzvg5rLAi8J2vcn7+9c5
XP5d8bF8OdILSFUtaMv60UlyRW/2djyBrmQjJb+nDryUu3KBd7XpTaoFKI9t+/8vhGYEfSMJdOif
XgGXmmni6MAnVsySme9+u7WzrJyS6sRbN6nkw3AX3fVg0IB/ud5QULp+Vm8XUTsBuAueWIohMz23
nQH/WwzCL3JrOMTRT95cJXx25V5mHBBxsipQHcjufnAjYhqrIZiMthOkz66altlSrUR7w10tMg8X
5nVEHd7+Actnx6UOyIPtQnMKSv7Ym2yL6mB7oV3AlgvJdg4Uj6aIw9JRX8pCs02RO+aZgnO61bYN
8uXoHFYuoKNQgEoLhMNayk0qri5jDgd+/601RgFEQyBieRqUAEmF7a2Kw5jNTeBCdcIX/ISicCQq
ge3FEdJ/EtvnA+NrrVqjE3j1OO+vhfeyg1fu5bGSuKxc5FTvcqRWVGXdreEvp6rHKsBmmwOS2RKj
fPfToueN6A5KlnYcml9yzrgPd3QzPVwtDXQRsiQ2i7fZGEGItQXYauI2/GyyCXa5y+bF8EKQoP3c
M0iFS6I2bzis0esKnuZjLsqCAB/nlvbnFkpWaxhOsKF3MlHf6AWlg+4pwtXpjZj0g3lmdX+FJdBE
ytAo5+ZSmh79FhDxRIe36ym8WfgMk+dFYR2DnhNf1b3bM50650nmAM4nUGtO1nLpIXaeYVcuTawi
CJXhn3BdF+remeGPs2CNBZlzz31/61mZR+TN/ej1n2RigPFvKzHrPIh057JHl/ty3QA7Ff0VU48i
B3PdxF+CSxs25p41M+XEP0XG+WT2rn5qZukXmTPoHghqMcgav5Fxdoc0DDyMHkQbZnryyUR6EuqB
ZzeLzw6QiiItKqOzNeGFjwjM6+2ZUAjNMPzDCuDzNFarB+VfnOSJ1F4sO4g6JIQVYvoem/j8YruF
ErY2U+u9UAaSD4yPOI14xs2Y73WTLsosKrfoDu16u+nj9ebtlzuV/y/pbIVtqqyyTlLUU//WnBzU
Wrwu2yJmEXvWM2yNOxU1wng2Sti1dPjX/6x8+tc6F4Vd4l0lyUE+R3YkA08drsLSyQD4GD7e+7qh
+9JoBG+HVCTBkTb9BqULfAdwkH/cT3QPGXNgFeW+Cu2NfXymaBfJHyrIF2FPYoS0V3S1UOWNV/WQ
dQJvL+vVphaRXYkOjtb0yObAkU298FYz28y8rV2Ru965FWesNcjknM5n4Aa661AO2lngMG60P4nb
V69o0+jKm1vJCzR4DBGNrgKoDNLmq2OXU4m2yoq6QxVKeEljRFOd9BCIXsVe0TteYDFKdmJgV786
nCddfk3ZMPX+BqUIxmcqBZmIgmLJD/gfA8J/r4Bi1V13BzBLGY+gE0GuW4+y0qoM9NMWDKaJfrCu
2J51eZYJWMuYLaTG0zDYwFBaK6TbZN0b14qBvpSyn2PHcjxkD+af4M84E0Lz2ehj9hCi9vW0OBYH
epsS5E043FvbwRxtNEN3ZvTzksO4z1gLmhAI2lIF/JwkSdGY2OokvbLX+6M1kAeNfOGO35mkUuKd
wKzKjHbQuK6mpLoAHUEahqrCEdmG7m/2+A5ItANdfvYYbtTL0UPffQhpGaGmp1Ax4QFglFwUWgba
x9L1D7L4FlTBYrGAEp6vXaOspg4LbvL3nWQysNYBvroxbXzahgySXrSC4G9XB1l2T784bc/spsd3
oUR/LZKPlWuClat8qIAMJ6Gwn+e2aucbRgZ1xy7pCSAqgl5Iva2AlTq31T/QwgIfZATM9MrO+v7Z
yQqk6J9XDRkMsHzevkjp63rVt9Yw+Fi8hQaRNtM4NGicaNLjrFr5PxK2P67V27IMwoIHA6ODu5Pm
x+Tlazckzsg9V0SB9xaiGfZIx/TzpV+Ofk7oRrlQ1z1bSVAM8fne3cEzKMYFuscORHZwqqiB5eo1
7H8vt3DGvtUtTryn6lhApWkdVDRYvBpqPBg2XKMrLAxH5TtvknkzPKSOSGxwBK1P2pPHRh4pcSaP
VRYhh3UGC+8ZoYwLKxl7rYUCTAZqif/9CPyoqg8Jv1Q7VZJtB9NrAcDgGalX5PPGqvR37weJ6MoN
e9eo9SjxzOWp5LoMV9geblr0WkqwcLKDzk5g9NdNVw+iZurAoZ+lqE5vJGDsnrcwI5NSQjyRZ123
r3RgFr4OdWWRZU8l2xApoi5OX3Pi63qvgnJmN6bHqwR7abX77v9GrqiqZWahpv71mvO/ZwUI1uRJ
8/IlKS8guxFhH+Qe9T8Wyl2nLNT0PZMBoYrLl52OgdWrxS95895pQASzRfsv85umtM4ZPBXp5vtV
20iiYezO8IhbhQdChYYPxhQdkwupqrntCadcIIJfSEFms3Br2tuG8M9v5OuXhe/4Se4ZRKXvm4Qo
jhxfLkum3prH1XDOeNy5dh6hHJXebUdmgYY51eoBPa1zeXbxBYJVntQ/MY1vyU8FHIiTx2qMcCjA
VKEqKi4U/XpS+Gp+dBBzyMths/x/uaCoyv2nCpdMiDOEG6gcTU2KP+9eZIa5STi8Z6skw2NVj8ml
PyriDMUS8kKEaa76mwnLCh7qSgudNfZK4zDE0wx7DRXvLaRsEoftreetPupjCL91RZfWZtI8onKX
6HDFZe1Ji+M27LF20NDoTatS7mhmgp+9YDa8b3/Rb8NZjJ1nO93ostQEfr+8ZZT+3suPzpgLN8br
eqcfqHABBGcLIgdPhQk28rfvQmxFMDscQE0bzZS8dXsOYn323SBwK50JmQcmGrVFzu9ohO8uBMpE
Lzz53yRgz7lR+z9eHeCwOh0WFBILPqxSp/B5cxVn30p/afao1Gth621gPLdalrTWX09+XbLeoQ9X
eWGgyl+5hPhXednJ3rhBHJdweT4Bhpj4I65qaLGnSR/J/LemL6m56h/BOJl4JhtJ0n4nCW4CCoUC
c79hzLXh1QPn8Chdrj6K58LGxT4oGDIjFVglSG+OdmQ9WW7K4lP3b/ZRzJ5M9PmRTk/IFme5eQyV
UA1Tdv5Hln0w6pQCPQftAlI3NMch4Mil8VPdc9FdGHumrG9LJ1PA4djnlhnj/0VXP8uJu7zgyMVi
lRFWnWh4W/T+5jEEE7Fj4QEtJYkRMf02QaLbAZojjD9PgHaJJE8rJdFF3Ur0O2x8kek+/rBAqTrj
kERi1AcK06bMuGX1KFBlhPm4bu+x1Zy6uI/vSwEACU9R26oK6EkNeeD9A2ilun/AOUn9UrqGJMjE
1NhWbgDCclDqHH/fCdwQCq6Np7B56JNazgerJby0D/9++1+UGNtkvoVtceb88E3lDeQ0yvY5n32S
ko8EBp8xatfK9NuVVkE/y35UyUr11JJ5CBeTEJ55TqZ+hfFb0m5DenVMCHvPmE2nnnUmozdS6rsc
r4T8gsUJ0Uyi7cl5JBcjun+MbDZoZ9LmQsxIPKStA73j0QQMPE4LYtn8K65ewE1k1A2Rdxn/odVA
c2UKN7sqUB7tLVl9+atLwZ9PGNgZteakT5H4A3mh3ZSgOUF8Ifx/wAgB6mLndCXvjBf+XwS312hH
u4t2Km0jE4wcSZHT5I3w48Y1Utg/dB18CWJbse8nyHfxeK0Ak21xJQ9zEPExD/Kmj9YDB/Xbselw
U4rWUFZIGvxhrfUSEU3AiIhYRYUwi7VHDxhf3c1L4mWqhdMHE0HGceDL9yqSm175qXOWp9MnfiSj
pwwJB0oizYF8I8QC+kZjHoU7Ri3uZ4RAhs7+IVWuJCbmVoOi7re9sOl/T4dcsAi2Vt2atC1BUsqx
rPH15fR3tlj3sycHaC9fAcrtyblhMd/vaYt9Gq4Jhb/hnR3LSY8y+EEcE/PWThdAhrTE7DNOx7JE
l9ZDKTF5ASOU6AKbiKw2OIDxbEozA9LK1p5hmZJSNkzcIa8XA3lHKLWJfrtXeePMZWbFKrDzvjEu
LQ8jVeyR6FPga8hRGsM78SHgw0UrKu7JInhwUU4oTcobZxTN/KFrl5zGCIhAl+p5nlrjgjVeIe/x
5CVPLOQfyLo0thCVq7ivbwiriIGnFsocKn/PTbX/yKH0ZrvW8DqfVH/vls8bv973f0Jny4pqnuZt
2T0aarNcr9uooE/Ax8hrzHHfp1yqpEz/9z090biUl80B0pS+IWPrL2VY/UiCBnN2r0k7rsawKDNp
FsBuSgghZTeecnlaX/ySoKaaEbkaKdVUDmmPB1wTESX87e71WUd9jU3ADrsakF76jr+X+VP9dH2k
kdYgvyRw0YGLnikuvKFqd4JzBJtmnY3nyYzQg1Z8+oVZ2fPI/hpdvkugTTwdpQIfRs5AyW5Up2yE
9C49RPIyvt63Mm/K69Q78NioB+kstUKbYodK46g2+5Q+06R3asGpT7Efp8kFbUcaTNHV+mCTICeZ
MEygSf2RV8fEFPdqHM9ZZiLJXb5/UCcck+70wC1f5bUC7xtEfR1iYZERbWvgaevX48dJDUjAtOAX
IHirNaiqyZ7w7JyhPckt9jO383+DN71uuav3GuQkSEmrmldmduue95TShJk1WMxepsP2eSXc7/UH
FzYZ9lwN9A6tM6MetLfUl7zWwfNnmHi3I/PEVcM2Ua6EqnbkQU13Pj9wtvzQ6HI5QxJL+XtiLhzV
Ph/honLyErwiNX/G3JVaL4mAxR7oPs5XG8oWlgdQqt22LIgAKC35HAb7WIYzonU6wJk7qZ4bETF3
iytyXjtoBw5QtKICuOpFpce3vOtE5AtSSF7NqV1kA1L9tI98cUfwpUlC/PXZEq9BGE6UAeasdmXA
rjzJ+X9bLebac51N/DDm2uQBnGXcNu5xLrkDZgQIL/SH71g00bmiU/33/XrRZQAvRygzg910EGdy
Uxy95ux8Mq63VcJEv5HrW2B8wD4jiO4i22slavg+o/Vmm8mU2K9NB6jhu55TZgiVYRILcazomEGg
m67jSI56Z/T3CoYTiehglR/uqUgz2RU/xdk7uI37HQd61CPS9S56B4t3gycPu4gBCr7JhVx1Dc3a
BaFxGAmuQ8Lr
`protect end_protected
