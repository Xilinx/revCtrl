`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8192)
`protect data_block
0eB40Voek3XE4QOCP93RnVPhUSFs7gsuZImk0NukmPcJTMD8K/9fx04PBknLIgTxGJzxdx5dk9mG
3UaXP8sAn8MbkbpLuki8LXZVKbQTOs4uaRDPEqLZbU4FWMpamBYeqWX67Q0tQfFedUfXEybUeVVz
OdSpbYa5GLEe3y7hDoau7Y4W4UmKK9n1NlsYpxuW1zzO6nozHZGpUoadeWd0emq6Tom6WnCsnvZL
Dt2SLFVBEy2pU5ZnFMv+4b7Phqbv+LFtvD/IWv0/1OPIRX9P8KONKvhl49mFDuW1kQi9Irewojjl
Wl9BabJtisT5ljEBq4AX1WEDGy+b7wmY2vgw2ALfqQvsl/Dm6fKz1p4Sx2WQCe3BryJTk8H4uVFM
NFc2JoXylTMK3pBbnO+DbPCi1oxavpqOZENXXFhv/uWNHzqkY1fZA4KJEwmqSJCP+YckvvttzkfS
Per7kCZSV1yqtA7rUHVkReC78EmSsWHVjhnpD3J/xB1YrPGIT8RPxyR1sDVoIelAmDsmtMUix0b3
yNSyn10NhRF4ZOe9acl6y0ePRP9Sx6PEnKnW8+pIIqeXjr/AS/au9ShKGvwrdQMheasZIY5vLtWr
n9pi9KqHrhhGfJ0QXjPmj2D1OWwjMfCnoqQaaz8Tb0f3+rA0avh1uwAI2sYBpY3iHh3PQBMIK2G9
Guj72N4j5BeGcuO5HWAmHwGZYocdo3bvclzOBr7t75Ng9s6hS4QWDCCY2j77C29ad0/nTd43giaY
wx9NUdkiIy3heIwaMNAvuHF6IilgcsWub0Y4UNBtlabEQTWx4QvP/fHzPYI22ghR6PFQy/froEKL
Dnz56sV8AgpGlEeE7zfQAvwqLeN2sGW4JMx2kOCJPa2OQqvZ1UEqSEp9O1KKbS7w365W9ee03KnO
4cpjdm1BOXQcNzFqpedexQ8n3zHm7XmugodTSlSIZPlTc0i9zLrxSVl0/PFglyViD/brMV/4nrmJ
TVWzxy4aBGRSkBYc1Nsmsn4bslk6HNPj6S6vCjLqezfffAv+/YVT24zW8zEhT9t1HmnCLgZYlfDh
SiPJzWpW+6IJ7kPhFgl7N8KDIEH1Qflcal+8WVSN9ia+5NdQZXafoR4GHkYTytochKiJ3C/oSyI1
QCih5OsuaJUQewHL4jHn1aW0g9ZLGTRAgTHcrbhTcph73S/qwrDsl1T+dIyH/yIXUt9jccdSy5Ad
itv34DNbUz9Fubbbv1Ncd8S5GchMjsuqPcOrZkILy1BFK7+Ww36jsRN/aBpLIee/pl0VblgP8arE
MxJrvW6fJiyx2KSxUSZxnNrrNv9O2bqX46wmDi75CcJoXxTz1v7gEHsGCHOtgCltHxrZ3AiY5vpo
RvRhQNvSbonm1/LL0Q+ka1UU7k7JvdFfy/gCz5busNb8H2XK26DAq9CmC2zuF/EJ+k0ZJ70czHjM
j/eUt2/BxM6q24DWxmemjQgj71ItYWcOzUNDQchJOVRs3FJ7l4K596VU2WX+7W4FZSazX/ucbflz
JwQRrOZNapqUkqjt8wZWiP/QDGdQbnmBWfXVhytpz8AGuAVYxLmYCcHZSn13LVwjYWPWZRvr0KXR
OH0I6pixDumB1HyVJdDweu9iV/kkBJq4aZ4pn0YVp073OV/JR+sNorh3+MNKk8NotjTGigXrhPxV
p4+a0KcuZRzDd2p8aB7uKCsemnyhZiWw7beHyZAqOdEaIIHGUscEbcAqFBbLtEvKynn00J/G68ip
LzzBTQ5yZeCD0mxrQl2a960xjBR6vec5m4OVVBn8HjJIxvx9VP8VdJ8YXcMVfggv5YCfqXrYX9rA
PpuNd7Scm7eZ6O+6xJTix2xjM3nyNds2ph3j3LfxRmr+Vx5Qs1uXaER2qPJwUXp2X4GuLXbOK1h6
cEdvb020d6DQWa8vgbemzQcftzYnp0kAWWZ8t/i6mU4GLhezmgjtxRf+SR/En2HVu+qFWJNtP4G1
T4f91o62FxmglmgBcUl0mho3DG9AF5x5GekvXbNWypZv/EOJHV0qFEQojyXK/7sFTLiAoxX75OXL
xot8k1okuQQPTfI6jZIzE3Z/J1QjtsiBx4MoElsZbMuG1bROy59eMRllGxeCymY88+PlrAk53SOm
krFVlVljc5bT4yOC0dVF+G7/U4LzBqPqyYdIOuYEE/wmihbIDmCkLqbki5Lt3cNVvyit5vixtm9A
89JfZPyxKhkDDJP7K0F3JA2pWPvoLFoP5iFpDfnvg40JOFzhbz5Y6WJmMAXJvC43/XdGOESXjZkA
WfEd1R6/LAzymQFoN8VrWj8OCvJ6xMzzuoUQbN2Rl1CC4EoJtUFIiR6NggvzlYkGfaiZnMmscpHk
J/XArS1lqamNsMJcm1T8CKDfYGKdnokQSh3iu5z9qckR0RXcQnzFxIri4NjrefTy+HYq966n5X0j
R5W1uI6GK44Nv+oJ5FvYuACU79hE6ORnfg+KAF5S9as6FdocPM+o0AEbEGrYjg3eeQBVPDCmkI0J
mqUWTo0lX/ojC2nJ9S/zZPdixoLLetRv2LGzBZNXmzMXMRSjvjHOXc+9gn8OvX2upP0nKSedgaez
9dKNLD9xHqOKsTtgun33ONNE2b6wNUe1areDw+KJQ2EEliPHAI5WzjMUawv8Ou3gnvlDztIYI1IK
uRpK95+mhCi3eYXawWYjA0IJx+vKP4Rvw0OYhibOWScgDTlAtlf8Awc8bFaTZX5JolUb4vy1X3DQ
ImwrNllnyP4XNDT6gvl0kZBzsmrC35gtXkr7FbLcMqg6gk1XPaBqDY4tg1p0JwfzwwqO16IFR3vw
wdSMPLuP+MxA0zjgnHsVpkv4NlwYU48GPJr3tyjwNN6OeK0KRudCmm5wSM9wr/rfOeerScXG3qgW
jhO8iNHaqKot5tf30iVAXdsishtewW2yssnRWZB2PvaNUKNCm5UQPdwSx+avP0I3jHCRgHmdkUFF
jBxLaemsI0b5DcuRfjhKyJvsLcuFxY9AsJQ6gA2cc+JeArFMRg4kWTGBsNzohcEoxT0pU/wxx1/i
EEhIhnHtbCfFtvEPLxStm1PqK8ivq6Ra48csEhw7nw33KFBKEu+fT4cPOoQ9G4/0bo8xSL+uV1+7
t5uIhkGqJ2WZgOAekuc+qnrWdJzvtgV+DrJUx+TEvj5xVaGrtGGnHGc8M4rCewHO2BPnoMsXDQFW
Ilt5vvyAi/punuMlqUwGsn7crmx8NSSoAEoZxavDr0j8ohaKM4wQaJI/G9ppTKS8hFcLyWSVuTOl
73NpARKWvyMGW1zS9xZRS5XYxo9kWc/aivWFjLmuoXn756D0HsR4sMXBzS77PARZD2197gGjT4sb
nt+9lvDqajuqNZ2m7SZZcmlaRxcV/SztNlor4I1o6qUfRvEaGObP2P6mPy/4QiohBZq8atKyOsRz
Sd+Vk83TJCc0OnMJBtplcTS/jfMCRBfh2UI6Li8IpBEM4KfBjfFKXSJRHNvbW/TEXWVnU3wOC8qg
IixxbvDR0jli/5pJJLhkLq8vVvqwaSdRMuca1r5laoBTz0x6TAmF+1R+IPaLxlTTC81lrnWV2Yf6
PJovcnAzjnAWyDiJ3IfpwicgvPI+75vIgxQgoPjKHsNeGTt/jOHllpEGGU0icb8Et8uIQqBgwR1Y
x26+AL3Ky8vCw0YUnmN61WtI2ejI3gjfx1SK3MiV8bFpldM+bmQESG2G8oVDLi0ONHh7uI6lrR+Y
DDTIszOYSf6uRf0cv83XzhoJYsrG97XNG62H/SB0PE+3BeQxcPB0T79MbELm8QIqT6KNrTZfEM3i
CNwsuR3znviz+InBgJRVgaPIqMw2hROa0SDPyP/HeM4uwSE2eW8LRsoEUC/IQ4V9L30AL6LdRErr
61BguTn/RKDfQDMS/y1A5yzTixohYtqtb4ibFpVXcoa0UuGFQO+IVHcGVGQ9aWLGmX40119R4Ywy
vCmiMlBFiO+nGNv/6rNMRwCIWylnRpz35s28XmjYQkVateJuxTCqR8a/41xwml/tc9AulUJRlB3C
KhVRqxY411IfxWbzezKeEJegGACm/nFYc09FbCEnhs81QTXI3jDoWx//mY1EoKP2K3PJ6BRMAlBI
Fz/elHqR0ZWYa1sl7olmwaO89uZAU1f4R69NByfowJ2TtypX7aSvkQlCCuOQSBaxXOmQCX123KJx
4PEKGLHcXnnlZjfBP7/vOCFdEZ+uhdQG3GnrIruVuDZUMlzSQ/97D9D+0pU9QSD8bdhhIs/QavEk
EG/epT8Hj52BosfvHlOPjKwgS+y+hyiOxUwa6sqU2yTbO+SIOPO8Rr2fSsubJBRWXnDWrPiR+Zke
bH7YUSIWtiZmubsvtrD+FOybDbeKtLQN14KU6RctxOE9fHLrVpmKqA7l5B77nRACvu5xcUqkLdSI
lzhVGqEAwR4MAVs/uwp2wQhwKyV2+7dt8NQsEvhHnuApZfiXuGniJjZW4TUjdfNH85z1GC2EyB6h
QWQNLXA8SBh8EiDWhY8LA75vkCwZCWzMCUMs3iWFy4KrAO2zBLpsreG6oWjG2+TAzgdY8gyq0EM0
OPyZ6XHDfPrIx2KjitF9fObEKlVc/jwiKbYLGdO7MmojL6LLsawgsyaYLOnOf+BdzrU61UZkmSlo
3aKMzXzivIz7A3b+2TaTGN++G2b22rGHXVajBzOVmX1+87w7FYc5vNzGzvJ0so6L/EokmaYANH1O
lziJALPtlhMt6FQbhGJq17tMsfLfNnpHmiG7Qu14GvlUUVvih/2tavM+PxrRh0JRm3YZhM5QABSO
QBf31K/2lmKJ65PbU+N53cqWm7Z5SQoGoYQQOMZeP7MHtGkRayn5uaiBltMkYh7NAVvGunvdYP5r
fDETx8JmN0DIsVUVCuK7wx8BBvLUfVngGw2/3/JZcYqmzf/+KJ22kr6bfQn30eu1RwqHfMwfchS9
FhgD0q4IiGYqgBV5NgeFWQH+bhclgHqpglAVZ9zvR6ZiwELnuR6IQkrWKo0EOLgS9Q+ixajQyz5B
nIwTUUNKpbI0qstdYMNTNNrONgyfExmmkeR/BoLRRZVhBMFtzlISYVmrfzIhNIHF2AwhD6MXX9pH
+jwXFpJWDg0QY7DZAQH6SGU/gvhzTayU9hxiGO0o94ocpRlWRyBwctisYg9046Z10FeeaU/ssWgj
Xye7HsIrJiROe9Jws7dkbRkNzgOpkdMqW05riSt15fp3s4U/JhhXWEOBBsxZoxQGVFOnxa3N1seC
Gzg/xCNTWpwI9tk2A9wZxjBw/mlPeFbAWndDhe3K17bR4ToCzO00+n8o4xJpxFCEmtkopXmEqHJI
seUFCq+o4SaB+R7L+lDXrRmgAT5xqGf6jjY2x+34reR6SKtHZ6cEnoeqHPHoeDEnU4K1pqFEdiF5
ZL5ugvP6K+JIUl1QfVPPnEXapsyuC3hP2fd3hjU/IYJbXTSFhdYlN0Ek/87fF5eMIdOwFmjXW+gQ
LuPN0Jgr18auhwD6UAL2zJQJCtl8qya3f0hPanswJEQg6t1LfPdG68Hctm3oAPWEMmlbOxwMX9uA
P3Uy/Nu94SexTOEMVTSmOETy4hF5cgsUiU8Js2VF6qlwNbF2Kx0NECPWD3d2KXG8RbkNjTR29wUn
rp54ki2R1DgCraia66RhjDauZn5/bk5At7e0C7cPUtyoRPeocg4GwMR72T07bAWqpWy561VKor9m
taxM6o0V6606SlYJfQRlesp1aRpGYLScjdzw9x8TnIpG/bQ48FquAcwve/7nEl9BjZRn18R7DhBR
fm97N3ro5XIewAOsIY5glXlKnZYmONaLvdSl1i5UpXKUXZhkgMLYa7k9k4uSjjT5smGLMNCVg5xM
RnLL2ixyqkv4/A/7U7+cHxpVy1eZ1d/XeLMSasG53U1iUtbOtVjk71P/PSXVTJWU2zTLwOg2zRGd
nI0PFuZ5e/DcOCQkhWrqZ2Klj9ZyzO+6j1MEI9Bl+mQI2hdYyfGF7o9fYl+d/1r2dBt9Q60VQcp2
zSLxerF9kJ3BPt3k39yAEHRXtjJXqysVRd3Yfoeq/kKEdr3L6UbP1sUW47gJ/p2F6lnr1oK4eeDu
p1m+r/3A4rZkVRxgjPEgvZ4KbB6iN/5Fh3nT5ZpnF1TkLmLpQIUZ62uTrTFFP2JlquXI5dr3Wtkz
v4xMJGYh4gZkeRzDKoy6pAJM9YJPqsC8kkYNobpi71UtnR5lk7vOPlTjvy0PiUwx0IoYih7fyksj
XlF5XTwj5lvEt7ASr9at8JHTdmVCtHziq9UTrm4V8brTjYim3NSmxdis1hJuDkGSJzzkzAGpHNTD
P+ifjS8Mh6HdKtIeeRBXfjGeCfGKTpcwlJixqmNWZo3dgjXFxsAAW6zoQjg3XvwpKWGj0jXVRlZL
nNAbC/z8/stRCYmw9J/6fIJIoFAhC7hcrtbLzgPSq9CUMS8EqB6XbCwH9FC2l++SzMPXl5vve80y
laMph4VK7BgNhg7znQsIAISFfNVcSArLCBDDbs/Cc8DzJG9bcA5YVleiXpQBqPERfxzbXjK/S0/q
9KucqSN0WtTWj2Yaqic4tE7YOlBP5m+xijXOngLrlCqrPVpTe0BGpFZaR7QvegAIjRhiYscGcmIj
zpqkeVYl8Tvl9o8pNXfY61a0sauj+AbGWTJu8hJVnlBOIdIlUnIYYJvlWrHNTiM3U5660lSWjKZN
MSNcJG6VVNxbINs3wEKJgDdo2drb75esVyhf7RMU3zfRKnYStCe3QidARo0IOcOiN3DVwlxFjKB0
BgilkS4rzjYvUnDPZjxG6wtAa5UG9/TMavQ73i6x3CV1/ZnK9wjv6RIXOwrOqpO2Bk2FML8GiujQ
zh5QdTO+oSVP8gsEXMaUxwykPg5TVH9l3nzbK1bZVdMinY93WMiwqDy1GZpVp/BTgxDNEldemp+X
zql3osxHSDid+y3iYIEhhHa903tSG7hkFQSdo9HgK1/8HNZiT5AgZsLGSVOO0ZgoA7r/FsMwhb1H
DbF0XQHlx//ahujRfvajwrJGbQw91r28Z+RwDINTmIEj87TrCFAQpCtWNcF3MIMOdMVY2wkKEI56
9XDApl6mftZmZ0k8Ij4Y7+4pvbdeM/tmiOcj5sgZIl2RVPFfZGP5q8OUMU9uCDNa82BOOF5nFogc
toBUy9cj2FHFx735R6L1O5ftSk/nkHefScca8wm1K46DXb920dbX1UJ4EFsJ3SgoRSvR4pusJP2G
jKUM4jmVydj4u5ReBdcMLU9AHNB4d8M2z9wv7FCP7bwvk6BetwPUcw5my+GMnldY1QhbAM8ozmZa
ZTOLXd6b2Ai2Lc0MfT7PUOmg94wNB/5x9KaFPQE+GONxT55Y9dJhfYA12xYinHtGvu/l2JMBnf2t
cZCse3F2ql7esnJpRLyy+6rOjyVUd7dLAYBnqS6N1HhZK1AAFe6DVAsGiDJE9cz6S/fjO9i0sKG9
aDbWAGP/ecpW37Zs3+V0juWG0tpyhYDywo3i2Gt7pk9iiccm2Jc1M2T37RRbSjfMEwYpy/1dRFoj
qFyDOBbuEO3Nw/RYAGePhaPM2i9iRcuig6iRRMYZv9ihV23/6sHQQH3R9myVNwcPsgE9zeGaD3FX
sOjQuc0gLNcSiQ8sK6t9afIFOBUzg6M5h0nsBwDWVJpd6CguOwXrsdE6gIVABG7cJ6pc5RdmYud4
OCITAE+s4PBka5HtwOnffO0ZZmCLXBrUuvpmD2T6PzTJ599217pmeu76xIWPlUwK5KAh+bUvQ0EY
3REyNOrS1jskz5stJUX14CPyLkRLU2G/8vpY/wJVl99L3U924+EwVaQZlVhjNoEF1j3SgCcBvfyR
GpE1fGht+K76CKTIOnWkyL7iPjV9MMmI5KEwvhRV3ZzkWpInXb4qLSD/0jkTwcA0R3y266itW31+
VRpgcFuaerKs1SMGo1JvP2ci5SMWHODma/wGb97mVtCT0eSRSaD+hiQMrMc+9OMyTj7u3/BHbKZM
rCnryRqR6ONUCqQDz7swzh7khCipjX9+faTF+xY57DjkmaUMxTGbUHEdsvjZqfjeEsfTnxkTf7/Y
f0lQewXmrD9PMyirrVW9uAEcg0MaGxX+4dPx6ZZoOF1rzAgNrCz0SLK99m59VuiLLEub7xcwHXI0
RvTHuM2AZ+vYjnfSeqMcPd7Kwmzn4QHBKXphpyYwiL5zSZ+YfCs5r9IXPQLVtGgV5jv7ynNe5/Kn
1d+WdJ1E8Xi6JRM0LzZjgUnMZXYUFQEq6NPAH+GsgCtA+wsO745QHKMlgA4aVcinhs65A77Mlr/x
RC8Pc4U/k1rXf6gJBBaEP7IjT3oGWXg+EPzlDFsFCujKblFSVoHXpdjOdpcVV45BGZjAfmzFxAS0
tUneFko/YRmCQwyo8AilqGKF4sI45F78arV1W8Ru9G0m9313ao7McGVOYwVOZ5tJdeS5ViYNhAO0
MSfGReeesIOEKF95UOl+QkBVqCuTw3kVf9KuFlZNqh75MjVvbaKr9FGiWl9poEzmw1Z5YQ+nkOOL
YD4o2cPTmNWtBkr5MKGE4RjhURcHVLL1LDwi9C+9QwUyIJ5zBcYG6VcxZpWX6+xmYntBS8ROehaO
FkVLZGEh+qCB8B/7cG3PrhtIgf1xxCHf498nt16ZaKOEpFB1Xg6rV2aUskhhjfFfvasNBHfAVfA1
Z6LNv/y0749WlA84cipzsviK6EkB0ShPtlTtHBlORJvv6pHg1oN2xta9fBfQJC4fxeg/wP0YAnoZ
vxri6a7E47g0GdNMBRSkKVdr93HNc2QAZESXjut96s4z9lVs05IuWj1l/jLYDJFY1vPs33FLaxT/
VvdAGi8eg2IzXaDeG0WP2d7J2MHXbCYTDx8MFrDjZ5JmJ6W1fu0okksPYRHR4RQgUjKH8GQpnOID
q+z3rKC45EkVmj2XVcDm30NRbHbeL1TwQV8Tw/U5qe4u/MUkkvMv4c2ralmViBz5SOjbDQXSBZXE
TQKyLqjA848crWcbgDiHtCyVHYy9qU0fouiFMF0nyFaU/ZxRGRltEVyIlIG728BnRwcEcQSAq88Q
Z42U/PfsK/YzzLR2mIE/Z2d/jlNdUgRqcWLcKwbrHeZyKaKc0GomAWqndB5c5jq6UC5/1RrZ2/qz
io64TujnVvyGmSX+Q5v4DGTQhtVJ4AMbmY+GyYutlQ09iCg+8zen3S6h6ldLCWKpL5Gs/HYkTl2L
tZVMJOlyq1+f54epuqrCoV77rZnEPU6G1mPIqyQex+6nGsV0U1N9pRn/T/lixoPANvYvKwzVP196
LIAS1auFZI8AVnGpcGyB5ODsfjueKJ5VP5tzy+TCaLYKmE+6b7bbfIpuA32PvTCX9MbXgTuoJ1eo
n/sThNOsZhlsdLFEUaSVgXcjIkFMUAllkI417wy7Qqg7YYUNol+5DyB0AfS0oaZ8k5Zs7wC8vjAj
FO9hgWLgg8ihR3iyQ3FiWpt+aS7A5t7azYwumTCUP6t5G0J9vfUoZiBgqPE5eS+ti2jJCdjFIEDH
i8W6VcTwUMLBFtM7NyeOUDrVLTdNvWiVjFoD9LZsuYOzGUaX9Wdj7iKlfouDowblCKbu18DFZe+a
2tiXuWd7Qy7JmKYUwnIZtsWWIaLXO9p9UtZFHnwLSozvHmfxJxoHTtN/HFb+eAwuJeiuf9xxCsoW
rZi8YtFDgN78QYxNLSIbEMVWG9Jcx1zfYzYkNw8U5W73iCPEqVvT8iWzqBHP1Gp3mI8RC5zEZlKj
RimGXPS+3d/Dl9MfMiE2c7gYeaS+A3EtHNHnSrSea/Url3Xcde170GeKIucaJuHRY8Mjpo2m4KAB
tBaC2im5ScGWYNaUFHVQkxyaASZ3Um5GRtquzX0+n3YAcd75AAY0u89o+bMX62CQo5mErdBN7ZOv
L0eAx3N0BHISqI4zb1dcopymatShvZ6YhbdX7AYS9byG6dYQOx8fC/nw6jNNovgdpntgXygThskq
ZPP4mnTDs0axjZER3ldaK6LI7imzkf+Wfgm65ljevss/yEMnqt/kApvG3SUfZJvDsNj6hY5kesNd
4SHQlfUA3abT1KUp/+3I7Ktv4cbEXbm8RQ3+QQOfO6Wd8FmP6zyZy8LvVVozpixCB+CpBoni3L9N
rsPSMm2jitfTncDE3bF3dEPy4QnhedtjO7VX1nBdriw456t5mJ4DcIESJ+w2m2NxD561q+/Cnm8K
/hjsPeGepQI0XrQNMztY5gkaQlWXe3gRA0hh13Ue6m48EiIQmbCtifYZLHiFEB+9C7L+KOEHuUBX
nLqPDtLk2s8AlnplqBVaB19BZZZPzEsHm2a00BsIZfS/hawVhbxQE29KoMp+TK90Rqgg+KUSAoxW
ewQ+/iRuARNc4i2eFMQF2u9G6+UwCsrBRGC+dCAn3RKbuFPJsIv0TITgUqEtreCuLkQzuzLYOLlp
FnBHwegiSfKSt6splQ0XecprLHQXeC/1kY9d6H/D/r6ya6XbxhqzzsK1+CMOIrrPYLSajJn7jX2N
YgyD/D6/qUmAXXjSY72nQi92BcfDqupQURFFdAgk6GrJLj41JYj5E4BRB1qU631uxBWBzqurH+aP
q2e+b0VfJG8knQzr4L4czC5RHvUJ63TbZJIpi0bo1WbcT6GQehf4JKjBnXKcVgVctgjT/RgQhLI8
2BaWtyOmtaQ2e6RSONBrgR6nvSnNmzJnSDulLSjiojAsPCaUiXeNI4w2tRnIVfReXjSdHWiafwdO
26x1pRJphdGXRS/bubrIsG1y5axNriiKn/rMNUXiNMAy5HUYxI8L0Rr6YwefKZnAs+8nbltRdWAI
Ufhcrwhob06eX+ymEwHUOmRmyyP65arqgaTWvPyyKscRKGYfN4k+eMuQQLkhB495t2Pqzc+L7dnM
om+mCmpT1Fj5ZqwrC0m2G0ugdIUBrmRew1pu4jof2v+/WSkCYmAkjgg=
`protect end_protected
