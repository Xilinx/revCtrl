`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAM4ZaB6gj7rLX26j3rNRVyvmaIAVcS6itKZRSj0uY7WnDNt7ObtoEjMe
XnZlGxxRFXJaWkK4r6Qw98G538NUJ68nBjCaKyCnLZVy0pWVoY8/4Ki1bFJzot5YjUnqkcZ2Sc46
iRvv8irdsZ5VoOXyKamj/w6aELMyycwfJFpZNbYDk9llDety76Wh51tNCfwD/OyH8LD/nXygqNGK
c5nGLcyJA0znoewPvBazwiYxswIvntQ9ApD/Cgu8cHiiACI81cKmVjsI1OjXHO7erwwX2Sep0vHo
kDQQciJrVUri2V4XMuRRo2GJm424nqoKbZcG0K6srb91nBk0EJ5xRVLZXymS3TY05m767+gH8eAs
pZAasgOFWtZiqUEblan6DZW8Zp3E32C45II/Ff42vjv0I+ShuyLnfKw0UC1pdQ1ZOKqABOlNDXV8
TAgMveR2uJFFosx1ETtcnHq9YI0kKmgNo2u4cWFE0Vj/jM8gzn3RVWK6eHIXG2xoOHrSC4lHI+Ff
k67X+jgha/ArTMLSXtZsDMdqAFXiy+DbMkaa5Cx4fEiXdbrVbO3AFh3L+bZrLJ863Z6dSzPOwW79
gRPX7//1G5hyKloSyCV983eLGYAdF3AIkTrj0RudJ/ss/OYr+waSJmy20EcA4jJT7I7H3wRTrulr
GZ8B2hUYIXkmsigwOfl1LXOhoVm7057ZL4iOOVYH4W8QVuVQcb/4xFInLQvrPkce4XK5ZMwvh7Vv
rwfmlwjWQqjlklpLLG5ayzTCbQV0h5CTfD/6pZHtL3qyU4NnGEVdtmB9jQCbnxQ3Y+pYDbrq5+vI
YWIFg0xoWgzUW0EHorcOL1BzwA1tGUcGJ8arrxX7gj5on+I7EbxxYC9yZQkr+/3lpHJeUg3OAkjO
J7VluwSbMjNirYvGh/3Q7AETKUb6mp4A3Y408I+5etSFqnrQE95j0ymoecoGzkbg8W/6spyFDKBy
03lVBiNew2plE8FtMQ3C9NLt2ycixTWeRNdA/9D/d5t8NSQQ/wrvQE3Ne6L2hyc/Y+EfXagu640L
oQAX7xQwst+BLBKqSKGKPerX2NUwdNQUBZQDBh9oXruVSoIzimF2F8y8rWCz1bD5pzGe+HO7Dr0y
81ml+oqm/poBgWT+cjmnF30XiKofRsnoCWlIzpjirOm7oPINjgg1CuvRbWGqkKyEsa6Xz6IM5ryq
/S1SzJWMjLRAvkWQK34MqDV9q50GrpLpruZDyoDhvnMHLrOaX0JoeRU2NUjnglsMjeo4LkuBjgIi
OABHghPrIK6SIlrQm1IeAJ98iuPxLo5TOdSxLwwlK5GZ7xeMeV/hP1uwQkdl1ugooyEajXGdsyuE
oUIaJTG1vMiZUORDdbnIkLGpxcXteeKjdPO9FpYYvYfQ54seo0FbkOB5jnl6SlcfQtkteSQG4Fmn
LPoi0VS9rEg2jjpwLp80gTEIoR2V49Qbxrb8pIhDmNU0Z6pyMXx8d8Ed/6YTfbLzLT7TREtTISiv
B1OFTCu9QDQxnSZOBONSZkc30X+DusrP1lHJicrf4DwpkgrDWu7vW63OMuWjepF9DmDcKY6/rzek
c0tCyRswkXUhcnpJblQ6HRh+H5oj+lja9Vyqg8bXeUDHSxZd2NwOCXtdOqHYdqOtjyFNFvjIe8pt
3yZaTn/tgk0eHLXuifA2pbRY7EWKfRzM9XK5ry5rNM0wIbgl78qAq5yBQo4zLW2iHhOrFkqg4dfU
e/wx7jWdjyM1vgh5W6vSc8i5+0LD4roGL5bBF9Q1Y214984OZG0HHYtLE7sHbLx9OBxqIUciY1Oa
lMJyIPMx+4LS9EXKCJ0Xa6tir2JIBLqhPDEdwAz4+HIZ4xO5JEDffSWogOpPbsqhsAimcESljGry
xeghZLpA9fuVG0el/B40sR0YyozNsIb/rMKha4M4QBsBsKjoSNnQBLSW+dbYXOtLA0v5M827uITg
TIrq1H0ZsQNsVZd0Nmy5JJFgMx6Upc+sf3MutNMr9seGzbeNhwH2826UjXTCBfLPyrewY1ZQcA2L
kqXJzJJGmVIZPxIQ/RbQ4j+PLtR0+SE0SWyrfncr/c2bcfKNagYMaDxYVybWBh/6M8Av0uSpb/Ru
P6c6FCactYkKbfpr41QdZftJgrcRcwYfxfRB4hkeY8ZrN5v5E3MqFhs2sTDdFjA4vTpiAckfWJr8
Uckr9McR1M4dM0I6ess0up1lhzAkNH7AAb/1jXhTkBiBwOmvIGQ2PouOyOTIJo6S52OIGJqHb3sb
GwpGrv3R0IArr225UsVKcEXq46yXzzyK/m89bmtck76NnRHQERK3yzfPK7XxLyL/hK/xUHWmCbc1
W8Bq2OQJP4m1qOhZ08aMCf3sEV1QNxt4symgawLa2i9Dlh/tWvueNnHYD9gpuKnnjSvFzYDodRNJ
reO8BbSQSXgbOXGb8MzEwCyeTuv0Jj313acI5ZgKfThw0331jgNywRvl5sQjfn50mFwYu4kwmp3G
5WXhqRNP9UOr0nZbold8dlix3Nz4kP8xWQoH4q1wBljqY18arH/MHFfgYufHjVtOO1zHBZ4+zsZJ
371upeSZ66xivwn8jLaD4auG9C+Y//WSvaUBLXJ4wQCDPuNnmEJ3GzIxogHf4YQZHHAOazXZHQLH
1oZBo8nV3Uixt0Qm7XlpKK7A6B2wgDNCVvgVOyGhTHTddODwwadkQ6/HIN+ZvX+TVDD+2x0GfFBi
AaUppykEpTILsOvz0e1Bs0byE/GeP0vZvoTBSL42dKk5cT7tUg/B9FOPGhaHkCNZUzfd7SUv0/D3
VBJRSznCFwvrU85KpL3N+ZLcQ9X4zplU+H5Xi7qTiinxJCGs48LJxGy5GaLkvy4ciQgxTBDsDK2f
nrBNRyStICgF7X/Fh8gpxhZG9LPfsyhvIlJp8FDkzG8Ad8xpDg6gP55okGapYCREs99wiH1kZwmv
dpFc5k/MKpMDZ7XrbZAEVYtM8Afp3UrxTZQnUgvoNQAFaMQSVbWokopSwm7dkeAyGia5rJWlQbcb
qou/OOG1POusuIgTqzw5cZi1/F0VtNAfMJqruEBAOsl+93mmYPPzvCRxFtE0kBhPUp1n99fltpZB
LoEDUK8A0EbevBq68yQP9uhrGbtN6/LUDPhoY5ig8DxxvksRTlh/+fWIa8PiZiS8QouZvyLFx+3y
RxPuqYNsFZe+ZyJheVZ8B35UEYDya4XVm8/Wa7gR/mUGpxgjEOpdkoqzHzdrZNTYsNW576FKAJXr
RJbRXv651da3xRrWnf0T9ujhdI7+zajI3lx/jD82Z5F6OnbpC8LymSBSK5MTE8dZjesJ7To+bL8Q
OILxU2IgIjMhvfgnYcXJ4CEwQjYvac/K8HjwfL4kLPrRdGElfUoxTqPg0/eqdZ5ObCQHrcyYg7SK
1862z8aq0+ar2bcRm/ttU7ab+X3Y/gzhfj1XT6OlhYM8zXFOCeqyo3Q2OeeKo+2be/8TYo35vDi1
kBN0/MXzBaQUHUc85PcV44NuJt7snbNE1HgSXkwYdKt3FeOx0oL0iwRXvVwbA998FrP6qnTzyjpq
FgHV2qxYVCJHNto4FZwBY4VALFOMFxM16sDF6oufm9C0/h6YhKpqqh38buq135iIXlg5vsugQow+
4fwk2mO1z31zRQjuKMbb5T8HFWwauPnc5F+NtmvQ+wZTPyqyzhh9H57kLp/p64glxT+Nhbohpfjf
L/hlbNDe8rIZiBAFxKgCTRnefAc6mvjvAyaV8F/JcCJnXIUcVMgAj7cQxb3AvR1qdCBBMtRhq/Rj
Lmoa8mBsxq+crQH2JqPBnhHV2ww/3TgfX4nJzFrhANoNcBPFtdzUuAe3IYDTBYbETO+QC46CctQh
w0drrf8RJuHVkQ94PCMq1ij2pQC7O0IkVGqSaJyLQLKip+YHJTivxZD8RVxNOfTVPnh+Wklj+FiA
jFNJESq9nHcHdRfODurGa0EUJc8V+fMX1H6NR4i1Eejgtbnfr5dcJUNbMxoQKRnlZgfnBMKeNXEZ
LN2uAhUZ2k2EhklnOZwxpLdYE4T8Y7/Ibx2SKg+GFdGx9wEiFfKeR+gjaYE1/HnGUihD3TWRt2XR
RA0IbgassIVYvrz5pA1oimIeMwi6gXO2As1r4qwWitx1NH5wTHfU/YTIMAKlC+jBRA+bFXeZJQ+T
tKn8x1+2iG3fvdOw0+zLNCtPwlRvs/9JIYMOZT6XlDjYr5pE/BLRhNlFhyRLlUPZExHGMhjunlbD
ER+N3Ipla+AUcMVKb/aA9kPRA1rM0+In/loJT89Rk2K5E0EHA8CPvJWZDNZaTx5iSQX96oKWnotz
FHL+OFhy4/R6RzFIUH178erZ2ECX9/RUTkrAWZ6Jx2KVWxLpsnV0eZNTTCcWFao9PaBiR41TD3Ii
NCUZlKglCrVTTGf4OgXzTICvxlX0fPeEweTPXwi8L1YXWp8Y1DG3HJhg9OSHT5WNe5icosIDwvQa
SaIOOTlYWx2SMA4wjvSuvoLq9CKt84+Nu5MrICT7Wu1SC9c9wRmh2YNchd8JhXYDFuLyN2oyRTc7
1AKKKe+scO+hYITNWxgNDUXp+1vmm7cVh9MxPlWz09cNq8Kd3ikDyMEtSj2YnoPysc+M91vWX9VC
TqOBrbYoxaHV/a2Y0L3E2GagEWyi9oCQx0twt4wwz13sppF4DSxaiJnBMgSvl5Ep7bF2zDYM64IA
H2jwomX4uNMITw7Ms4LIv8n+UcNIJv/f/gydlocPxu5D+SZDyAxgZK0peM71Ud8Luh4Y8EeOiP+3
s80LxCfc33pXRMZH0P9pteMoOYNPUJVm2YX7FjDLRo384IYZX8Xo/2+YxxwnCytqSt4P2jZsh6CD
zMPnWcUST7vXarZZ4/EBYpMuXKavvijw1hhvsdqH2RaJNxKZSLyFF/ogKhvuYx5W57UPvQEQ5tsM
+SHXZINajvSyZmM2nZn4iKLX+c78yWxaaQQZNgJ1Zkbkvk1VqeIYAWlDe0oZo1+0wrlxrmEc39O1
e+6jlNjIUVHoN5QM1f57PENQH4+kUUetHILGes4eYe+DGwhnPExqhJkx/GIlC/PrSxMvIjijHOpw
6WHXn3zSD6V1ZUGwpH2Dvp3mWlPUhBAFJILa15vN+AVnWxu5M3xMhAZIfPU8E5av2mHogvDKCexL
mDeOR4RZFGiCuB+y5k0KmIRbDmu/gHJQLkqRZivFtUKHMKuZkO1ProH7eiQant6XojVZvfhIEGUm
gUjMAVo6DQWg+0OF9CQMDsOtsO8d1I7Cz4JTu93+KKS9HHpaN0GrXnsVS7Ttg9+lqxZ75nID3eqX
MC8sr/cBgywfVIb0ACieoxn0ny2o80xmAIDCF8fI7ldXWh9S9I/L6SwGgCrJEem6sQWU2SANyPaS
SeFUs4wk/3ueVs4Qai3PWk9mMIcVJNAHUWbELkfbV+A0jExj5yzrel9QvwrP4M1agBl6WlUIO24v
16Jt+Uo/YI5pumDxmxg/lPudmX7OLk5N4/ORBAAvCdSwf+pjEJfvWu9P6y8rxhRJ2Lq4ep1UWpoD
4mEuofw+Aoli6elDnNsVxEJv7sPuBeVxcjwrTjlVYYzPHy9yZ3gaEpuSgFXj38VFdThFbFrO9IbA
AGzZ5/di4qK0Nje7qpUwrqQ/EJ5Dw6WaI/2yc9kVVNxC9z/l8/w=
`protect end_protected
