`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6704)
`protect data_block
wrovcHZ5qwQL2M/nAAAAABEDKcEgBUJmN7bEkSveRawYiynkYmXJ9wjpvTqiEgbRHFMMlu6tkRhf
Np40Ht0TN2uVBlS9KJhlS0mv0fN35qMRpYlLhVTO3PmEjwLhbsIGdgrnSyE27S5tLh7PAs/zBUAW
kefg4OnpeVUbYshM2GmLF8di0LzshZBVMjdvv4uHIoNnlESGdL1XJxY3eL4vixqUHKNTVEncwF+/
KdW5pi8is1wwyg46kkxKZvfF96nI09KINEW182yiYnA1e4qNyIwMA1bAu+ZjDa1ta4v5mUgaXz6x
NRr6SI7/8lorBPuqdTNxRq7GhaxkHvcaUcdLyUjSS0aX3s3cjp3X4hqqy1fmHEoY6a8zveKG0z9u
bu3417MHcJUtWgzt7Nhu6NVY3PWhjzZpVCwdJZIzna6KCpqafEVlIE5PlStpQk6yHjSWamlN27sW
CvMBFKMuJOZzlG6z94SCVZfa17GBFQ109Xe9emeBfw8jdwQ/2RScWQ2TOiME5KsjAwtL7TvBaYOF
qeTNzjGlpl6C2MzV1VWAJE4QDaDOgg76hv+K8bXvwW8dPTzXeda/Q97t+u0ZVkXrl0tEnR3lWzNK
fMA3J4P9ZEH9QmDBXTE5+9/3jzh55B7g5TaF+dBM6kwQsczBGT2xDd40fDZUNkEJSplrbRwSktJX
mMqZKzFjMsgeVnwKZzTzdglplDZNKg8Vm/Mn6eI/Z2kWKDwLA7DRuGXDh7DrZi/xffIlhXeznJY5
0zmT5w1gIm+SI6ijisYk7K304JK4b0G8GvdqWdFrNHkD0jx71JJS/T5wL/ZiBd9gdL+uHpqHi99h
XNs3MH8DdtnO0uutc7g5xht4ECfh8H+HRibYacu7WY8dOTgWhF4vYe4O3VISWf4WuvWcPArZWdqT
NH4aojYbsWOl59CSMARcHifb3J1nqw8dSwfcJdvSPGeAHGlDZKBirxwZ5piL9K/1hdQWurYDOci6
al0pnoJ31qV6YZK/PdcjlXQw8f4I6fy7xFzzfLDDDTa6pUySDvs1XIDSmxMgdswM3ZPgh6CvD4SQ
HH5yBEuPBq0L+gZDcflpNBTTK3EO6HlMXlZGNlGklACcktyZFwufuc8iZQF3qxB04u46xaoytypO
JsX6pU8Wo1Y824AHB+tFk4+E/sIx0Vzb14wkK6xlAZ5GEhL3cNj72tT2b8AgGmyiAmnwh55x3c1c
5KIA40nGbCYx/mjk7UTA1b1jEs/nBzwfyV+CzV5OC8XxeocaEOC0VISIKCU1CgztDNaoNgELvX5i
SZVdDYMKUJcGU5F7QHa+ir1670+WxAeryr7nbZ0feKIIX5PVi7yGNDgUqf0DdPkMs4pJau2z2Uyq
8KJqBJNOyOKlrlnxal55TRLN4OmZNW2srXk5j8aKOVN+vj8BUkXN6Duf0Sxb5W+ldrCmi6CIgzGW
GMhKVFBPnxRT8pOZ/Zar1eD15r+Ot5qCAtLu0EQOlt2TG3VhNeLozcmPI8yvaOJKYb4Pn/jFmM+Y
foXyQF9XIrU27a/9vlz6wIx7Ygb5mQsVmUhqOlUF1B+0Qigm4Vw6pAGiqw7vYnJB+r5hgRgOAfpM
Kyzg25QTvzO1X9Sdc1XqYkIHP0188HPMwXmbZp6IlsDpxv5vNcPdxs/siPLhqWHsJbHe8SIlh8mG
wrvX1pLGKB3Bvj2RJ8N+H03vM8CkF3pWRNHqiA+1l38Jdg0m8k8gu6FSvSvd3JwrMdw4h54ccvru
G8/YTYJamTUubgXmDFeHywGtrGrW/jko9INntcdXbPEcbkCnK0RVOjCa3gagFEXZFwH9fwEldjm2
wAmTHBOgC5ColaONCRSfumIoLAchPygfStxiRv9U8DYQ/wD9azTEw0nU7pRIBB/pDIxIXqfN6fMH
meHmvedH1BxCcRWZICLgQ50p9v5gmhaK20lSIyozGqDgrhdJ4yUkMoM3Kz4DOf38nfDifxJIZFnZ
cU1sI9imqC146e075312huva86gJxpS5uH29eBcz4Mbksj/fVXQBTsnJVSbR95L+hAZI5KbjKmdD
sA+PYRcSof4ZphY69Zn8rFefmO+haeM2fKTkWIdt5DBRi5cs78Nyj0U4twXOBAKcju5gia0D8FRo
Y4b14RlX6kza7hLWWoP0Ot1BpqILIeQLWYfx7RXz+go2p13E1x+M77IlqWlkwCo1hA9x2aY0/2zS
g9m3e66QVkvWGlVU2pOH5VNtg8VWZQ2pwi2d2sONMgLg7qOcYJKTdHbBITwO32hqzqhnJHkSlpWx
rzNYvHv+Kk+NWLu0LC/2aT5yejYYFLnIrn9ytzL/bOlFhL983phl7XadA5cMKNzOQXvPsgk6mcb8
1EolgbuNzfV+2sasm8FiFTcmqzIyndDp/UZURz/alNePZYifENJjbvDOI3yvKds9EgxoTkr25N2b
Q8DFQTBosJLXMbFVTBKRdfqWrsrwRvOc8tDwmUquzKIN5qZV6hLpPpHv7kzuOV+8GvovxEMsTTyM
1qDCnB2A5s53qGBnICvL0UFwnwIlH0N8kZiRrwZ1Q0bBgoYPQKwaRDPMLk2hWg59h6p99ME6pfKS
7V2Q7Tdz4tKQ8HT/fwEnRp5owIhNWbXkG8OLwBy7ic7Mr9q7Ul8BVXA+9qTx/kG1LrpHjR6Aksio
v4eX2EMPO9YdcELr3Et+pzU9PhyeDmToEih8GE/i7Dv3F6tiCQAuimZc5MxlDtdofjlZLyqHYDFQ
iHtXIbZSWgaNZpIqkhArGKi6bOWNBWYLeeIDy2522Z5D6pXi86EwNkv2g4TTJQoM6pkRnSj4Dv0Y
1JcArGjqiBV/A6+Z0Xpl5qAy5KcLYoEUeNHC1jWIYlJNwccpnkodT3V+NvtY9fnkqzDrEaBnZDhw
s3MSeAfevzl1GhSCCiizrBYm5lkUcSTM5n1yXvHh2F4RE0HocuMrfCco3XJvK1bwy5iFuTIts45h
djfrJSe0bIj9+bA/xDMZ1EjMysTLDUbONtddZ941f//nPPyk4+kiwO2zK4DNxjQhdlGaLWjQoNOO
dosbZIM+lSYaR0jOhwFbgJGqxLG8V2n3fhXxNX4EkWAmmvyLHcjeRCH/hIhVetSUL1LkzKEyWbMc
pMsaGJDTpsso19WmeZOKCKxtp0S1kJ4TbRQk2Mo5kVP4QvRIsz1PIcDGNs4OpltZbC/4HNfllT1V
J1j1CxA0etA5hGYtBAmnXtu034tr3K2GVqI87oS7pJOs9YEsYv2LPCUpJ16zY/Le6upoLcPjGgIN
tA9NNnETug+aU3CxSZI5c+PRtWX5GKkwzg3XXzWbDcIgXrvHe+bc5SAEcGQvOcMgSiu2s/08bSip
uNdZn2KLZYIpy9zp7Xksjs0TOQxVLIbq7IfXjAnOe06X5+nLmIHFqwyAIAYEqhQYvO46YdX+wyKY
C9LD4jMzSUco5Rwg5cG4HKTIOzw7wwrs6zebEHv2KitqMPRc2pUhvDYq3XWfaNZUz8/VXL6VdDoq
zQnnmg8q429PEwkCuUt1FPww3kbHdRyxhNpP7uNggTRquKHiH2Jod3XvYLNggFHIkXkgsh2Qm3+U
1AlU3gfKiGj3Hmaarl+/EeZZClaY1zOazK6cNmRyU9iINmD3o7X07HvGT/+EehrWVZ1Yj7cUafjf
ITAuJphK1IQBFm+lBSGon/C8j3j6F5GTeEFYxuIgiwfoBGLgRJDZWLNbRHpJaN1wnGPrtpPSxoiV
jBpVqjcj9ePEgPbrT78SIlq10o9Ul3qHgsBRz8qj5Mg3gAVZQsHTQRwZY+bCS+DPwMM/BvCPcoOT
QYA5rtyB42VFt/Y8ozeDWS0AjXJoInsbIwC89d2nc6Pewmlfx9SRxOjHijSdEVKlL7t/1x/cFM1Y
3H1jx79G0nApBBpZB/0NxqKsXvPf+OHAfMCsp9UsMRzqGnYoGvAIzl59P4sQlAUfyEVEC+cZqSNz
jGIkcZU17LpZgPZloRbsIHzdSDQwVHOGha0LsrSZVI1rHiqkAwIjFPP3kh2bbUt3gEWGjzMpev7O
yi0vqaMrJOOENzOC9TJODjA0tXEdbprY1CeRV+r1OsUeWJXsYA+aiYIcXLfrogzPf/zkzmTtfqWT
Pqk9K6hXvQINyLpVysk8jqeEuEZRcJ2ZY3tNFZXzUGDKsJ0gK2LLGQPbMecUNF7Q4rFOUW9XlLiO
vPm+pf6PlmetrjxcxvPgv7mr9vVoD1nPnOPnfJ5acIvESUCfy2zZ46ULAu1HpJmorzfR2MjW5nyc
HcRsolktCDCa7WkjP2YNAF2Rm2XVGLFHKoLskhAwyhcg9QgoGhD1XvmlwObe9yi7ZQy6SV1Io5Ct
/qz7O519QloFJAw8N/3+O5o5m9PH5IdYXcAUbzFNXzoB19B+Tgy4ApXYrBtcTxRgjtBjmDyqkH++
LQgULsG9kH9PQkvBvOj8r42Ywomc1PF39ZZs9gwqWycKKzwC/XnJFqjIxG0RN6b9clbPwKWDMLQ9
yfvb189fnc+oxm5ZG+1NfB8m0I57yoiA7kNxsKTtY1nNddSUqbJT6+5TEgy8iYuL895dSsBw3fIp
OTDFCv/G+vqw2yBHAsJU+pUYNKIrC5szF1Zc02v+TtixGCepRspxMuiY4sbK0DLcmreBsFJCOdG0
/B2cN+hWGvok5k34gW8f2hjFVPlb0MdygYn66xjyuNyfBejK2UhmFoyueDnPuCCGqoP/TJ3W5bBy
IH3E0jWq6ZyKQjgds1AXg4Q9KeZGJef19pe7ud9tTMtaKS3lUqyGbIviffp0bdSV30QA9xoOlzO7
GqDjazfX6jmKnh1/+Y3XDOx2meYwVBISHdfOP/pJLUNX7f4F7+tOPBcFECIE4eJTjClSgpXCcNhh
Z95ZC0czWW3GGJH0IgSkOnp5n4xmaLpXHatdwaRL60yNXJfTlf3P/m2KPQHSI2AU8Uwd+e7xwMd9
Ge/AGzxcXw6Ny05nQd2blMDqFvSwkB18aEylnnCLJ+msRk6gvuTV+rGjNTFJE3vlwB0u1PRsMnxg
W0+0hQqSgYABkzayGS5ks7f43Hz0jXioJbFDwzlsFFLh2tBK1n72TpA+vrIMPNfO3oaYa7Qg1aUa
DTgtF6ZdjuTFXvUW7R8xd/zXj7QgNcMYjrnflDG2GMroVPXBg8ppTjtn824V+XeD9S7Jm89FYhtd
COql72vgjb15t6TkIsCw/U7l3cymUbA4ih8Esfeh+104NXToXx544zi/UeuW+SgaXQnvfRm38DAR
wRRPSrSP/dFScntUUD88qt+HesNqGxd/ypkJUIfb0+atAYx3LWJ48HBzqX71g6bmTkOq+3jBAcrm
N1TLwJbPJ6uXqtI1JwLx890Xj2iTrWkC8PqG3PBLbDB/ESV6S+R9biIkBDtqZzdNGRXSEQzINFbc
mDAZIpWBqXXzGwmAsg/IGSu0bX4QaitAXe8U4qe+EwtLXVlCqdsBSxm4Co236psBvTxH93kggz37
Ql195oc0zwvNJfS4mXvZHTpkGC8vC0EpPucSsCK/kn+OB2IuuwA9B48DmYToxP9O79QK9sF1l2Zz
LdBS7AEwRZXeQb5eFTrNOCZ6yzzjVKgKLYhkZMSyQDlEQm3zlqhdQRDpiQhWvlquETtQpmPJibDs
LHRmOj3yQss5tFf94BGke63gEIldKpeiNylZKo1ZM/GK9cWP2o3roBQXPH8tCZUwmUFkFDa96RXb
EAnjZv2Dwmo3PqxEqw6E5S/lJPerNu1cVbH8CJ9vvuM7SytHQ4YZS91pjxy96jfif4qkwuwyakWg
9dtGciISSqxZLB5xIqzf5VxDCvZ2TpYyGpudfCTXRe1L2CgNLmAS1568+zshgV4zdbryOX1YSWEs
QZg48Bx7rn5bmIp3UsHr7QbvTTgE0Vp5E/CZbJjskQhH/8hxht/xHGJxXb4J+61OXl6gIV4tUnu9
IXThkWmAQ0Oe4Mr018ibdN1HjgnfeOV0m5vBUeKT1fqLWoo3PnYlaaKKIXtpffR0QSqHUqiXbxPU
RCw11Z5zZoM/aNbEllLJPcK6iQJ8TU6RReEfL9lgEWnWGmYIB/a3dDaFmDYftyzy5/RjsE2FDO6j
6Z1xCPteZlaKw9uiNrAmpQKQcXoZEOnMigCRuyH77LUj5A+a8TYl40n5jbkpXBIAgTAV2hq2veVL
vwBj4aQUmo/I/MEfJ6h6ok1ctuOOh0QH8wlQxYRAhw59TbgX8IvE6YchSkc8fzaQEV/AXn4+W06d
AVyNNNfzVgUDRU63EnPNPcnrDCsD4tnzzvfKaIpj+sPD7bnSqLK9VJIUVFKPiiSTez+Z7dANB0vy
jOpsbHNPmX8qQ6gXFOYWdoelZiI7Hd0vMxHB7vm6BilVkLnlsU7ySYXmbgUJnCXK5LwrhHN/vsX4
UAARA9Vtq082YimhP7nrEdYRwP9PG/W7ir3nIASJO14kgsBWYl5f3Fn2vNymv/SQBPLMmajXmfjr
tf1ib9tR0uCnfq09xyCmm9Z9xer5tbC+dPF9uuWO3FZVxxb2P6eY6NCjPhOVbB8DDWip3C++eU8c
VLJAJQXtlr0DDIQ52WXvWFVZgFr0jcQd04mXkw3AliluZVQNdS6MBkJnjBaHg3Ml//60W2ddd8nO
caYYQgSNqvN+vSM7P14tNM+FvKxcbPLEzQ+cfi6SnY3Oc5r7YKQUKMvbtEuZQnalAa3IzdStOCXb
hrGY1SeNYLlEJJkvoI0SQTZ4ll9hFKnMVwKKC/6lJrTrt5NFH8tDb9EpU5CLvm46sJgesgnaZ6w+
IztbVjTFqA8WTIrQMKoeFn2T6R2W1sXsm59DTEO9UVcSZbdJB53QMG0mBUyCp1QHW4LlxDDuw4eK
ttwSMYXQ6I0hMRRoewcyeO7Tu6t2CRGJzLEThBNx+v+uePjeKAX7+LX3+CKn5o8S+2Wy66ZGB1qE
IH1YThYvBSow7dlVfC97PRvr5u6RMd8vIAd+2U86XSRPZoMxdvAmCW+KECViVOiJd1YCCwxh+tkO
6Lq80dM8mbQgc/c6x1gWpNqaIwhc8eHf7a1FVMp7Reo4P46tkEE+44OowVELX5uxidFtNMdGnOXX
HDowsnV6PnNw1ZslAu9zuAEr016XcTIIfTEMgIxmio8UV8ReQi2xVaLnNWgYaq2N0yFBJDHAwtda
4vH2J60lmUBNZvdBeGf9V11BkjBLseY0pw/hautZxwyCEAFNBP8PK2ECAuXPx7ypUfVPHMGH2kn+
EFJ8cWS5z/TW74Hl8P2ZlwZI4VHslycfGyRiNLotcbhxjklmsdQQykOvZ+aiM9iLUNrpgzJpCYZb
0IXSjunkO1kGi4WeUgPN/ZYQ9oFjGx9vehT6DOV75orNj+E7PGV3t4g8htz2shEf0hnPGcTToDj/
gNdzsQX8Ka/CNCEbeh9uN5FxGsnt9yeKKCf5O7F4x7MEdo8UpbLRhDI5MdzWvJ4ZLSghjbUm/f0Q
KgbdKxl/jqcBb3Pgn6kBEIBAqrVDwzPiioULCK6fxoaqDPYotpHFlpfieXBPLf6EUMl1gPtM7hCd
2z7plXjxhvr//+4gwPn/3cYEhYj63b8lUpaXv0rVcD0MzToatcNII87HBJ7OcRhjaS3qWQhpmZXI
jRw7HEWwyjKCxqtHUIYfqV8oSCvaZue1WUnHxn7k0xSRpM0hZ4weGDd65JT0nK6n4YiOJg7dxPGU
oB9l4FizapGV70gEhx1AKhk5geFLNFWOSjdvoTHBG5m/Z+VAqVHPntOWxReertrqR5CuMHwQoscS
Pif1/x2iBFZ7e2cYHV2nUr2Ckv7VYzNROOnyVTmIDCBnCi7HVU/j/v77sj8TujLOCw2SHHDd8t8V
C0oa8So8WVyygMV3zRT1xK3cDp1Q1SkqDR3MhRLu4560hTxmJry5IMJlhSYEheyujo8cMCSvwp9Z
twPyUvoj+wAYknORKjueuFx091Sn9n/JDfkOnbC9jGMqx+IdXhH8DvS7DQgc/pvsoKENEr4d+pPO
f8W+2QO67Teiy3AT4PhzGvCMuOg/vIbPsI+cagfDldMtv5UaQnbeuC2FyJiCq0briQ1qvrGdPYK9
AZ9VN1/yam/q3GxK4952sXJ047W0UgYKASvmTEgF/CSoSVVouwbMuquGUrnpVUJGc0C/gC8GwYHq
GXxZCZM3hSiFUCYiZCPuxqGQ2vDs4Pg6F4U0i5j4MOhoYHoNWdCWDluyvqBqgKq23CosN+HgVkmP
7VbZEWTO1fyMEERsF5WKF95z3Qo7KRHihzjO1mKjp9gU17zndYT6siG2Wa799u8pzaSsRweHIFqu
vGaGCSahL97691gcnlxCdPusZ40gbgtxmsoPkkjmryC6ZOs6c4LdfM0G1uiJFpm6oTybfeStXRhE
Wn3R8no1QOtL50PbS14t9jUmkGEL2FXhIn/Owt/72qgFmkZ4zfMxVSR+PQB9lQgjGnApW2BmTDfn
W829xQ1P1chylZ4wXAXM/Hs668Ra2KxFbyjA4fe20lpp4mNuNBuyOgn2T8RD32OyQOyvB1B8f5rK
L233Q+X2yT6zy0GULKvOC06H9bmUXUj+82jFGcPugwMaF4wOoymi9R1jacovzQHyrY1/VUDFK1et
q2w/SV7likqwfiirEVatxaT+WlXFwAPXFCdlYf4cNvHKZQnwufUHov1Cs2XlZW5St4OL2VTuvz8m
x2QZi+EJrm8p5bfNsZnpbWR4ElNipiBIsY1TsEylPCbKwblgeAh72P6MFQQRjwzMuTZkYBSF53j9
9MHs2sxTu/740HIhoxphfMe9e+vitub5hkgOHRTti7dgSwtwYsJMKrTF0vrVkxZ8IjnCt+MA0+9J
jDaP2Bvr8U7xSbjV447S4YM9sVt9ENWUb6f2fP0FVcgt++AuFaAh0hSMdYdgajFLnJjbvj4E65YJ
ZBLl9rU4j8DvoKLbMjKjEzDMN5TPSgfan5Do1fqWkWckfkU=
`protect end_protected
