`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9216)
`protect data_block
wrovcHZ5qwQL2M/nAAAAACcrQk6gQ5cRWKUSYsfWY3JSbGuqK0BUPAmWkkq8yWantsYtB5iyuVFE
dVbC9HbpLV/L+TDHICNczrZwQ7ScvmIJdEDkgrI/lhrm/m370fvL848Zt2D9CNzjzwNcdJdu5jum
NMD3j2U3S3/3RKdVY2mOO/xN1wtwfjk2DGa3OsXgGwW0vguaVmFQSswiXqXte6R3YjIfmsHQifZB
N8L4dT7JbugvnATV1ekDU0HdHVsD8BNAWOuBBzcDSMs7TfWffpK7WHPtp7jVRdAHuofKUuGDfbms
bHeUl+9t+pV81lRXgIukIk95fNXY0yGNnyp8rz/U0aT3rqRCDIXHfeIensBUeQUxUm3xrfg1uK6v
axQvysDkSAoNVS2FGMVuQEDkhezUu+Hi7h/lxIJg46ZGFxzJqTdHGOmxCSFAfdK4XeBYE5lW3cXQ
xDk6q6odGimV/IPQRjUzHR7JvRYXgjwkr5O7JpGYeITcAcHroDaE5jhSXm16XGd3PUtlED6Z5zQx
26y1vyN7/fdTzn5NQvsvVvbUVzDGVNjTleIOcyT8wJNmH+KyX8BbEjeNJeZS1Q5+k/dWI22cSFQ+
7DCYuWCC5biM6Nm/+LEbtTAduBj7USjkTIPH5PxXwuE6oWLDqZkznxPUu+sUY5KTSNuAgbOwMWKV
wxApF6LH91Pq+0uULtqtGszApM72F5BpVko0gkTwqfCbfXA+3xrIZZ8njwnl2YXaXoJlzuB2VC3g
gOaONkycCnDKUfZ6wKpgvgT0u8Q/pVabiowmZANnPiazJJ+hwFMyngLb2zOn1VFxF3J6/Xef4pFK
ChE4XjhDNrCSBzxW9kYPJrywa+sIahhBHBdmYe5rBnFnzTuAfJz28y0wIzlJsmj+GHXlPM2iWQ+R
1rCz8rMGIfmyTEEL/8VTEsumJPLtXwHmcvxBi3Mq8pRUoubMsokxAR5rMWsOzvQLek9IdWucgmMn
srrNO5u9iDodyKV9tZNlopzQOVg6S6l9eqyDvVUShUsVaTgjeBlKwzjJ1GBx9BgZR+8asEyn5Xq0
/hZKKa+gPQS4papfNRYNJzz89iAZ6jip0B8+5RcsGuXIntNoMIjb9ce81ElORtzBLWlMNbgg1SUi
EovCE3VsdEK2JWjuC5/X2wzcveKu7K5scyZFU/yHT0gv5bArJBIEVzQudLuUuChJZD6Ku4a14jB3
a8652BXvChntJaqhvWSTKNoby2oS3dp8xzFECwNHUx3xLSc+90leW02f0ssqfTbeRFKPfv1hiHXS
zKzowCJlPqrCsw/olOLM4wwZXJfd5B2HWuDrL+BsB7vXy9+P99/oOM+Nc+v8DpIrU4r55O8Pyd4i
igdyQbwdfJi9Wp1c8flkMswozpg33W5i143wYf50SpeaSzg1E0bfXpuJFXijHYRQeDUTfuRNoRgZ
5eOnC5rJ6aNfKu+iJ9IaYiR4mAxmWIrEGeM4zvE1uKqu9LxgqfQr0SHm19zUClx8NubczcpJ6DHu
0c3yhzQZUolRmleaY1hNhUiTsHVE1VJ5JYEyGMfa3EP/fUgkZaDnlaQTMrRSrflKv43HOe37oETE
5WDhBU0h0PAyCS0hsDiguqoqYZaduOT7znNcr2/4BCjwxaCoolSQcLqm3DZJAVkzTmAMrmdLYGoQ
jb9LC7KF73Y65LQzfyjRMEnh+/Gcw3h/mQhjnZ6uejb1ej/hPy+onAJUG/RvEHlLZAN/x6ij6dL6
r/tkCwuVVZg6MIhy7T5BhB4vRuMdet5s3vLP8PZ1d9S9ZpqES46jra9lX4aeamWMP8zj8mtRS0ub
YQMXnPuViuKxh0XytIdv4Gya6RVsSCdqlwD/H52PN3iIAMpbZIBVIYQ1xXvhrb1qvoy3mwdCGfs9
08M1iboMi/0tAEKjDtusfpu/nOXutzcRTqJLM8cKv6+Jr3yUDfajqJc5uUPv7j2eMoewOweTDOla
CA38qZYVQFphkLorZzmTr+c260FnJHiOkWXuVX8LVHezPEARNncyDRbdZvMNXip13l2ep/Jt7NlL
72fgueHmfl+wqbPLzqicXRqw/xIXvPVHdg5eLhatyy3VvH79J6+AaHxM6eQJDJA702pqT1xnXy0n
ytOjBipFxPF91jiUy7Az6pA6SiywoKmKumkIlCPAhMgREMIdKbQ/KeCe3Ob1esbFhho688vqw7i9
icF+ptu+1C3+3d4FqWD0eIirMSImV1GLs3hC1GDUcMOis24eTtB8PbbOkAGemKV2LpUuMgcpELJQ
HxTzfN9DrGvvCo1qlo9BqN5phJf3NCMlH+p/XZagN0oAv2H82Ld+Xji+KpoagjxXNgjUtsmP3Z7W
VXb1+gOMCJAd2H88pTxgAiA8bu7q9cOHh5CsRQUkd0rIburKMkWCj23UBhzILhttk8zpL/4RaPy6
tRVuRIqhDRG5SwVBGdJPjCExs8cUuHSvYASPnoLO6WfADIX2uYjoBys4H4PnGXRbJV8O1PbApN2W
Geeij6YEOzkNz5TzrcM9oHwUTSDYu4VLPSd/23AuNisa9n/xhys5Eebc0TpGresu6XP8x9Xn3mGf
ZnYNtxLdDYlodYGh2twS+VwPiE1iTbyON90FMR3Bh8We68c5ApCaUQDm2+cAn7m8GSJskqJbjzUZ
M8sww6jRhWaT7EF60BIoRzouyQzsLJEGb51m5KnZMs2Xej18msQAo6fhC/VzZiPa+YOmlPAtMUHW
S6EDPG8NkoyNavOsN+xPFa+R9UCKJCGQnyFoB79mAPPZpFd2ewIl79vSXsaA9XsucZhB5nq7uFJb
VuCF+mQLujt+4Y6eoambzfqNmrW/uZarJBeCMWzMvhjv+El/3wtIOXFZDMX3dgJUG5Yw1tex+CYi
qxorG+iC0Ja+CRoenth843i5dt1Dm/UWOSnj10rGWgwYDwwLPEd3xkT/qTGc+PJLlRh3ZytXqok7
tHC+n0ZVZbRpGK8pihTrCsG7JUmzCbUAKhDcjfCGUycLpHNYWDGcksQIjGPOdgZ5N5dSQCoGlDhm
IvwlNUN5MQHzcPT8RZfUyCSGTlDNUP2h7zAhFPStOh5UNdTNk3NU9FqG0Z+3QQxvu0uPVmvQOqNi
TJJinqJ9cho5wH13hJKLUYmh+6IkhaLXNz/FTVWvi2UoyL97iJk/Nz5O6TNYAtJpnn2QmM2fqK4f
Kmk1pipTzjhZO2Zh3/8uNr0sGbbupReUomgpBERbvAqohpRr+aPkbowmLWAS0MSd2SWKFTNZVwSB
DrihKkXKEkfCQtJ09KZzxYjpWWN8cqnffloBoZxWaI61rIanqu+g77D7TnSXlcnbiN9a372gWez4
WAo2pzGQvTeW9uEo7tTPoDOI+CLAsRt2ZXaXbyiMs2gWF4vbXqvWiubI5IuZ3nF4dSzx+IXihw0Z
9BCVqggnM6IHDMsx6jhsQVWVDaMh6UROXjy5tTxhrbc6+TgSjQuSrGaiYRtDXhPTkMvs1CzWBexC
dCTlU2RDBqoq1gdhkTPLPvbiN8yBBTJU+hM/KgfjvJrlmTbFs4YQ2URBzmkX1EQ1JasEOCBIHAHE
9GDoMmATdYUBbZABg9ZfriO62Zkbt0oENwiJq4AqWEqE6WabITWnqkjQx8AaWFbZV66kjMnPoYSU
vkHnvNNlf78ePnH93rT73B+ZsZFZ8r13eOvyRvM5tF3OV2ZxlLR+VHARRg8tyhpNeJIslqeSBYTG
9jKkCYoNC0SQcBUDyoc++9oI5kuOFVn1os3WQptSF1k7u5GU3BjWqqQTM2E9KQNPJLzMU/I3BuWV
wnCNL/+3tF+c2u7rkSAspLygV1v+HBCDGrKSwRf7hqWNtyq6aIhhTFli3uFE/tQ9g323o3CYqCDf
S4xqp/iUquMbenyIMVlt4U39c/MJ9WMBPjZJ11suZz2LwAih3A9znXZbEQzCzewypivJVL+nVMBB
unrmlCdsFonI6YEAkEml04AzwcgYcaeTcIaEHmtRlPQhyveM7eHhvOoF0QlccShFnJg4rNHMyZeX
Kd9G77VKNuY3jAJrqdp80pJQq5KKXExrVBbnuMibbGGTVbnpuiC1Qi2YTeCKSN8l6ia+vZ89Rg/p
IoNeTpEqwkZnRdp1wxCoLVe7f2LEEk3R0OCxNQEGTh7KvOANBZsPLBoRqrvDEoAL2rEoYXWV/rXr
/7pgqhBIHLzWvtn7V3XIkzAmBo/ab1Z9lb3XYyaeTi/gEn6nugJyivttJxZkzwhfTHCcNYXgtsPo
iciJ//lgZ0u/YAn/8Z3Yex9NzjrG9H5j+PAqh0b4fGtbOnBzDn8phYqA+oc8x6tMNsUhn+bwM7NS
/+hD9fkOG9FGp1hwYZVSt4+GlL7OtgnM3+nBeYVNILFiGfqUFv+nHZGe+jsb/TW6fe3hKFED8gPl
tvYz0cAep/7d129o6Wz4dV2CkvaIafM9hSq3H+5jvv2oB9carAF3LQ7Sr9oaxZH/+c5bybKxUI2C
yO3o81X4FmcbjPVsqGNEbDSDweWCHr1Q96MEbYx8T4joQCY/rF4vYUwIFw89I4gvtnzx/R8RBGIo
UjEVU1zLZcm0Oo7iTnE5yFHySple0T3TmkZFX0GA4wZaodeqn9ZKd+VfLm0Nis6KGcPHZZ5lLcBj
GYYV3pkI+/7ydBP/uTJZcvh9h2/HmK58W3j3VHJh4KjdkYhmpdns+OzMYZo79F4sxiOe5VIh4yrC
UK6xd2/kr2+THeV16lLWsXx/5ZBIMM2YW41SzQ87k3Uno3cA3sOcm/w+hCGn7Gr2/BkEzWcdjiPp
EcKMtZO7anljym0B3v/Uu40gzgcwOFKkJ3JgwYDzWBzuT5dSDhu0d8ob5hBGFTtC7rmiN9ucPswF
5jRtqDXLwhOYVDeqmt0+ew1fu5vZ5+wDu/3Yn2fByC1gAhLdwl1StzEb0OFwfPPgrenlKIpy2bly
FjZYZo0M7WRPj9V5AIl//BSofjqDLnx0HJFSsyqOjEIw4MZF9a/HTEyxm3wYByagk3GIOZXTPMFi
uLRLEKktYyI07vmOX8K9ao5pMrSXphI4QNAgvmSCOr0nwh7po8gQlZUZ59lpOj1VxtzvApi9J7zF
/nL8pb9EBodbqHaMLahl++sWFJZYoj/H+UI4nJgtG19r/ahANWcHqTI/COsup0BvotISPey1WEr+
tO/n7FqbRjNYKeAi9qDWj2Sxw32tEDlS3NZJhR4jf1+QvQACKWcjt767IG7aw6tHpC3y370rFh/v
p0Y1hEVGm4WFG2nIF6FX5Re0dFw2MZa08VfjZdAFtKapItG45tk6UhUl2E7xsTJFcOtmwGwD/1OY
g58676JwJuClKy/1cLgkyZWOChumBBJRB40Z82mqr00sFncZZFUKOeB3Qnwu94AXh6zey14V6TxJ
SbwfucBLm/XEtFgSHnqttMu7dJBcGuVZaPmWdv4D5jRpyKx3GTAor6reG50QmKji4mKIlig3eDAM
+BjKlyf+rMG0mz510vcZfZl1J2HYDF5xXneYp9WSeWq7/Ht63fjJPcuWXMrB8TEO4FdcyBZifW/0
UA055jNpvjvw/QAcW43Glfga4PML0ocuhyLyeInywUHUEssDbx3dXph+caHqt8wkaokLaehUz2UX
puAYw1nd2/MyY1hDRYAVxbgY1amEG6hRL7OCo+s8Zz8pLoz4x9kZQja+IjUcZBm8ddgIav01Ow5I
CA7J0jGkU65J/yBCsDMH1AYgVLfntBNtikbO1/BAKCvjImQBc2kmooTbqKIUtvd2IhIIDYawtcXN
iFaAgA5bELcQabk2sAJhkrc3TOfZNU8gY+I4cQmK/Lgjr+mbZETtEcC5EW61fkpoBQ1mEjrSxn9g
oTrn4PLbg3Jb5SiQtYLVxFJZXllwnpCZbMQMy/rX+f4C9+P0mi67c0Tl6bFSGX9+pDibBKnEbvsR
TvBl2QYJWBlXzI9W+K2giLqR1xY5VFslVzuszU5I8dTVv9jY45MDj67GuIjSPCGKzeMz8ryYvkQj
4ixL5362gLvPkab8ovamyFHEj11AEsInhCAECCP+nrsiCNJnBHBzsua+KzdHCyDXbGpFLlkkyWan
4pq437Hmr9vq85dxZTFNzDVYNbr3lmu8Ndl8xTUmVvcuah88UZsuWYyg2VpV5AYwVQcAWEMYrhc4
zoulTHMbhOZNHqvp1SYASRtZBfysliU6uIzN4Coz3YJb/edti+w7ulvHKuY0I7HHNeW5/C4OFzgC
vAx9TrnScdhpiiJjtIyAa1yfYvJGfxY/OewNWUVrI5OeJcGApPei5WtDQ37orc4dlfIg3GZE1Y3e
6xnc+IKYxCPR/407lzmqA3YhcPOUZaMQq0gfRMTvXYzP7FmBz9yXzeFfVjlze8nj3USbdK/PHDhO
HXQUwLPu2X6jx8ja93H6y1Eq2qRAiUxMkdbH/yIrJ//MTvk0g5fpKl7TsV319omiGwBXWi2y6sYf
egl06d9RXnhwgzubl51naDIWwGfJ6a2ahyY5k2hoeg8bC+uqjttHduQ1LsYTzsVgKuJwA5g6DSJu
jr4rq60BibOQ2Gjnp86bChrJRXB4i4DQ+17qZd2cw2zNaaXBcwSLXKMsKn3fDm94hMBiT59w0Ibe
44+F+lJ4gJNw/5DaBHtQe9oWJKrgKLcLIfUilmipcjsPqIkunlOcXT5INnUcm2I+dMcw+BMKojnf
muui5h5iZ5LyPGHk2WDRkP3XONSnpVKfwcqYajTCu8WmXuo3Ble3eQ4UxgMsUKO4tMoDGwZOF55Y
ym84nlBT2dUnaPdZsiZDdgF7LHzbtsM4HjOL9rPuxPMBxtbo8VARs6W6YWdQrCbF0kzvSnsh7OnH
gZlkwdEq54qhTIoWCVPLI2HyCT67EyhnmIcO5u9OEkOb6rssEEMAt/Z9IRl1+KM3gGKWuiJO+C0v
l4qrtnP/0spm/uKrRTQ4ZspK2x84QKc+MhvUpqhI1klbvIr5CER8M2b1SvBUyjZE5h9QuSwy/rdx
ChOpZYB1uocDfJD/8RjRER3rv7TeTmg+pmsQXMrwO43s5QEul6zDuJA3eCjxq7Oou2maLfogvkzH
vYQ7Y6J35CLNQTW2g/bK8gOSi6NPhCXAZC6+DQAo04p95rw1AyWdZvYkhxYJrl5ieIdx24onufLK
toLPmvaVYmyg5dwHfC04ANfpptftKPz3nps662hyIe3gSbmMGvgm7zXs0++Aa4OBhpsMHGL+NvnW
r81qY4eM8tbqSl50C1rb+YQtq8dZZ2/BJ5FPvqYf32a8pPdV81Go6OTLrj5KlUeY0Di6ecr6CYzU
haO82apfefisd/m4TATQzjH+47gWPE49hDPPlss0eg1myqW8bDT2tNVQWa6Wsag8kRuW01rTI81p
e6EeDBKbTjzy9EPBwgNlvuJAe6q+Fa/f45jBfz27MVTkUnjtg+gkg1nS84hrJuQpfM/TBXAVKCwd
OM7hitFOHX9zd5a/mM6HnOCFt1QJWGjPq0x/1i+XSFNY3Y2vtA3EhWec9n6D6TpvQftBgS+XnPLj
+PEuhxP+GkMAygjj0H60aas8/lNGwrYuIX/ReNELF0y979HuV56IpANjexLEDMzb7O9hE/JCVoKp
6Jm0Q8r1rGvftWHJZTFUSQSxcEn8f5IwV4hJ4PeGySN10JtoN2wcMMBnzmP6NVgCCsoefpqkfOMo
MBDtWGaiLQYbACf4QT+BT4cbKs2VZ+fEZ1gAjL3TBEM5fUotHcDB/IANRW19MKmmxZ4PoImoQ2HA
OUAan8nWejsDTeWiPoJIGrWSnkN+eeAHXdfEp80sUkAAjx+6tVjxjPgpjSI2x79aiVNJOZXAGeZO
paT6DY9p/cUFBlo5HSLZ8I8j1lDDKksKZofRga3psGY4/BQBvZKbBNFCK1edcNyjHAAZJnBTixIy
UEP2vr3IQbA9lHAgUr6YS8wo/tTYDcD2lgRFF8mqjybo8OArLybMBvhqGvRczCwQDpJ1I+XzK8NJ
6aJL9k2qZlb34swEIiYmt+4eRylzk+D38FXk7JGR5EleJvQJBj9+nOoy1QIUIs8daY8VFZyHpM1X
U7Sr42jmsQSUY0PU8mOB5E9cGxSttvw5oCasOrdl9iLjMfRObrnEmBhkzj0ANnARoL2qP2DLMAAi
B9qx0e4BGMrhOXJXRwRrlnXeeFEI4nplx/GoHpc/D7rkI1IVwFTE9DHnImCFM3tadMsgMiSleTrs
kFmkQWagmJcUQAHDH+JNPX6RRZVSQEdh6pciml1PTLq5Sb5m7ZFobKIfkXi5FVU5+hzOh9hklwJI
p5mKZZc7Zdo9s4o7AsCw14D6A9GdBV8ZzNrmDNA1/Jy+tbQFT2xA+khbaaBDOeYuxiuY5mPFrw6v
lbnGImlGJU7iBlZiiWEgitKjDjJZmpScI9gEEnfPD0Me9pXESOJe6p/bXxqDj8p1s7ZHR0DFd+d8
mqaCh9qheuXkjXWyLOjdyRmYlAlxFSkiXnu2DCqgkf3clBEehNnhWYVnMhnXqufi9wL6ISNuvxJI
zocJH4cb5CpJGExJQcFcrChvqB99WxQqbi9DWYkPxCxiiYpai6bAPoj+Zy9O+c9JpkmmSRUrJJo2
UTue+19qfVwmMb5oJKpV4d3drPT53O4/iSWs+2todqOWONKqnxEPEyAQTPOrY9JZIsVTzeYM7UhT
OldJRCjXGgxtnLz1jkKkrfZeQOb9FIWd7meAe1vVDIn190sWvSfI4Rq9C6m5ZA31TLkWZw6DvLuu
RYdYVjDKjb6YgYAWCtyuyp3o5N5+fjMEOvPmH4iRxmayl2bFZKl+QNvu70LGMAZkx/GudzsByJCY
iQh65WoRkiK9Jbld8/5XKcQ5Ii5l1snfDxMqgD2xlIM5Kqv09liEwXFxkHGU0EW5ngR4weIaKXtF
+uZ6K1I4c/RpE4iFTs5SwLS0OrR1gFjxlG+oi7KIrq5cl5p1nXA/8MqRqfxfEpGTvmIx24rQxu4x
oPUbpGF7o9uHRA3laY/XGptOqYSajHYQqTmNBHKm84px4VUV1iohe+eN3lpVNMb4AAgqrPOwtAzj
9WnFHQCTllsTPL3a+VYHh88Y5c1BjAjxg9W/K9Aq9R8n1fAA+5HxQ1FzA5B+PWxPBImII5TOevP+
9VF5Vv8JSqitYIMkfBJxvly5tNtlQ/iNJ85uWmxrS8HeNvIjgtbAkPJq4EUY9F0NiqijGgxPbH01
CTNotA2rs3ij09fYuAvR/wBmGNeDg/fNNKfGkDBMF1HKiwBTkyougJoU1dBYJQZVUJ1NoX+bhgMP
c2chZtUYU+JQuLd+AnDXkfPocGTyRJr96/mKRaeE3xYGHGDuX+6L5SX/xq3/oJYh78BIkBm8NpWP
4+J2Hjz//08NCMFdSi0KDE2vnxYDngiQgitYBHNEKlS2DifRlMhw2p6FAyJPOs0Z9479WcqcqTvu
j2tKhST8UkuV/eE7k42r8bLD4hnc6+X+QGI6f5heytKeh4rR0H/GedEWmy2E0oFIYpIb2y87oZI0
hHdEz1Sq4w1tOC/1VnxeLga6ISqoMKYSoqqOf76/mLKK/NmlEy2yl0h6wsDb3A9Csl7jMN6Qy1PA
iSJ8mcqRPJEj5V3fCjVk7KZ3PiUDHGqeT41c2W4hGGysW0YkjK0vw10P9lwugw25kyTprEEQAxcN
ZwylWtBkxAo3ZZv5+fBL8G+m7bunIkEZSQyGdLAgqxTzy+TZJoUJpsX7i6tRFnzQMV4tLhlXTAfu
+VSXR0J4AKIxdHsrrZLg71QcImB38SqPeO3OgvLEfV3vmtqNuunatCeYkxiFGcGTIarojTtKbrh0
ZYTqGkLp7ERU5HceDjWr2IwIE4JJcjcj65+t5xGOCDthiWa5LHH06oeRrkSzfaEJVHJOTXcnqQbW
fb4r+wgYSHz9bLx4OmcadI4SYw4kQOI9yDcplGL0hmczskCYjKGLZkenFR9CMxnYJyR4iELh9Hz1
7RLGNlhv0kHho3U0t79Dqrox9tuXSf8dHmvGOKtgkAp7rxcN3+u9SG1hkbMxF9TD+eJLG+eqxuyW
XjKCmdvUd+MdZSXMh26Zi1mX3LD3M77ZRL+z1VSHDiVBjajC8IKcmI3PR67r4jjHTscr4/j/tl29
y+t9f2RkBB0fqDRMp61dTRV/lYsSk+s6YjbV2zvd4aH27ZcnuMp9e5AyGCFMaOvUmq04EpFKMwWW
7XDO4VhEMN7esdp1rFl/gxoPQGAlozrnjXyePucehOgEUfVxlj2Tze2UDC1tPyHvKHL4U8nKFJzF
GdjtQH26xHM6t/7+oj3krCPQp/7qVr9vl0Ep+S6CAjW5bCNgUPQq85Xhjlo/B/YOp9ASKVYyVD5D
kxeTssACWnNEa3Kid0sHFolazhuCa9QPKIUvEUIqvi3Xrx0jiwUreKzXVsks7Ij2Vv4XEVbitKg4
zTSLYMJI/OEwm6VO8ayfDbXYnazNxriLMB5FPKLp/P8NiWcrKl2XmkRuH1qSpjpDLaQIRi6cCXYw
lY5Fjhctek5ZbYV5rIaAsmdpuq3TK/SpojTEpfnN3ZB2axnlvELtnhYl4o6MgAolk3wZ+dQz2ddi
MPpqEGZVZQQA0qBfPUyfRrfNQ2hY86of4rpGHSo/cgtVM0q4EUGNQaIaXUPQ7XKDXLULE84fUiUU
VTOq+tYtWWqPz1lRhh7zdcCaP5RHEZtCi7amHwC3wcbdY92KbLu3NMtHQx24weIXvxphaAOCdpKA
jCF6yRWyQJ1oKaf0K9y1ndLCyqylS9OmfG1clkhqT1YLl/po/y3gkJEp+vJebSOvvhAhtYbPWFe7
/tQXjDHQF1MdrSHORYmJ9o+TvAAssh993ZC4hRk0Q8YA7IbCUx6voGUQgzIWvB8sXSZRn5v1IPfU
ynFlJksGCgBPDlum31jrSB1UZ15D+qDUITCib7PCfNHka575pNlR/8Dt4Aw7q2HWsXFMC6WHj/KW
boiiEeymtgkEDTOR0KbazMsEAKXfuIaQI6fBs63Pj+WXNiBcg/tskhCDW7KH2tlaIwHpvqAkMaQt
qnWdyi2doV78mJ+sCmFK3oC/ozhXHYy22NuJsOe3K1YHdgmIwpxN8E61yJkVuSywCBXzFShrbh7K
DYjrtuxs5d5BQRq9LXdaEnb9CXcjJrM4H6ziZtu3yDV5Pfni5EDwM8YIvPtaGOHCiS5562aMashq
OT9wL+s7ADMqP5f6I/LmHogEDhA8wi842XN82ADUaKbNzfhj9lYilQDLAOYdDyFUQRDqQ7YJ/t6A
FbLfk8y5MXw9ofxqRKNhKKxjwX9j+VSO+h/ilp27bLro2gidl3xJWoTd/0mLAIpRIHsmv7gZo4RF
E9y4KNyQumcCia2quafNbJ7F9a9PmYf26htVuhQdXREZ0Gi94cV9d1TV8spyzF0QCvti3URdHC4c
tjtL+7x51fxXrsA7E7M17ayCg2mhJ4ZhoX5EnNGXXrfgj4378ylUCdm+V4wzNGRG3MuertmuVwwn
cz5SVVc0spZr3svvRhBv85iy/PpcfV4XzvBUCyQScfQGj3kSiKeip1PzRwZ2e4eWveOGvKo/BXss
THL7Huab2glNAnyQV+qUvj8ozwMs+ZaHX6YUl5PNugXW6DQmM94ZLeGkhw61oBG1CnEFekaHlXIE
QcDzAJPMg+v4VO+jnD4GgGIauCVevBSfRT/Q5/LYjDpk95eqXamomJKQucZETHxLQht2u/ZVE5Ck
OMKkIZCE49xmXjQBVvMUEHw/9YwZiyLWxhtbVTSs4JmqLjc9LVJfWCe+zPLLrVm75NRw54XmNfuO
MWItd/s7qxeyvON5OXGXjzjcGEeehJJSqqQXDxCktpnd818j0du59oQ0ksilbw2vAvNBTa9fOjHW
6blE/7cpXZ87bRWr6S2bZSa2N/qD0EaSa7dabVICoeNQ9TwFAIIzPc0jMcnHldG3zKZZGEc69nUH
mv0uThFAkT3l46XiCK+Zg0kvmG+OHsJj5mQN1wN3zHeyJAk5K6fYgvY8FVgn3WbMHN5dY+DN69nF
d7G3dXlydlo5oDvwiXz2wu2sbOZQ/U08j8D1oLiVyBZf47Fk+k4ZG2iBPSNPTikWjaCQdwQAnNrE
q/V+hWtWx4uqhK9nXO2KMLVUQL+CUCbfUvNXyJPJbTkVcJCNEDIdICIbjCdp4nUckB+WC6rWZLur
u5Wxb9dpq95XLKBC0kc+oVQX8050bIZX+/xu5IROeEqnm5qmPu3r7hSjJ31SIHcrGxFxqhFoEzV4
ZUxqseMaVFYvlxlCFF04uhfPnBqS+02NkuzeZi2BQPjNxdP1qLjy
`protect end_protected
