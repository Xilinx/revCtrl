`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d5VJXu82JfSwswDjhvbEU9He9tQ5/1Rw+4/2nB84LUuT0wfekcnbAADJNd0/JtXdeaCUlOw7Zwks
Bp1VvQeB3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T1a12gH9+o/WCd/uq6lAozrIbwFwnflilDyEA/rZKRAxvRmKOSqBXtjVpxVSoEgX9El2BLPK+36k
Vd8y/iFx5HcwlteYeuYuGTvgQerRA9ycH4Qwt9s5DC83MaSGod9ecMMI8PPrmdJ+hCOX8sXwEsN9
IHAKBa7h08XDRsgW0os=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZE3CBd8eugZohbo93EvXvQkUxCnosHfYT2eG0uuvFgW4E1aUdxFin2hcHpeAodvxBTyPhYz4Lsqw
3nsUxnz9hTb8Lhj5XnlqKx2mVFP8Z35n8lJk21C09QHBGoSukklDPI8dbQUv/KxN+k1qsLBHfCBA
FWz2UAwKlgCaoOPe87s5MUwwDM1/P/D4+XgEQCRDz/7JDN7p8ZFVtltMEx51xjJOCvfGoEeTzG2k
908lkYgt+B4pvwsuFOHwC28xicC9lqwuIR+OiqTI+hvqIl3tijnK9dhEHXmlIo9PqdVp3p9K5niF
C0wKwI1gK4zk+Z+Qv31AV2g5KDXjXxSpUgHlpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1K/c2Exmx3hO4tktdfNX/hsUCqBDw6bH/vDRPja11f/SX2mhefMgy+yYp/XXIVeJlyTPI7AwLQ+m
jPsm9qUsxInkPzY00BDkxz+XjPmDvPZhWK1LaTfp3S2KuDInJ2AYP1AwgClVQtpRFpipBFYqQeNS
QrfV5V8iPYsCh6rtCZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z2R2Fz5uoP9gCKKJ4H8ByaZdL0II83JUVbmmEiqboGhJOssYqqghHZS4Xla1DO6PE/W7lUbFZBMN
taobe7WZ5vLL3z9KT5znQ5u/8vqZfQZBnNTCM9ij+NRl3PRmkUPrtcd6xURukGspBspXFvJDNTq6
HoC8rJF2dAK3E2hXtQ2qzFXYx2JspRBZw2ARE4ENjzYZSYK5AhF3nV89pEvyjDlChnkSNr7Ec2sz
zSK49rQXLtbokqxvvzCHRCEs+NoMqKlklN93OyjJFAIzYffS6GiGtNeycU755Cv+/fAQynybNWn5
4vdHnb+JcudvHzAJFK7/azTzKOJrOSm9uJYTZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5184)
`protect data_block
mvi3i3MBI7n8zvuunOT1BDhfZ9+75ngvsPXxp5+0g3QEMYSUqfdm6zc+CwjSUXFsd6PhvodvCHRd
503JQr+Wyo+muprgXcX+Z32LQiJj8b3Lr41EJJq4AB12Uslyg9WhaIGr7+IRoYiOqWg3qy4hu8DX
oLu/JcdILqKp1p5YY+maL7cOooIxAi5R9XMFwBxlM+haR68vpJmK3w45uw+oDssspOrdG0aHsGvP
yCXjnrMUh3lbLi82LV2uc88OwKOA8m5/09RvtNHDqaV0kQPmdCXfRWHloYI3Kx8PCXVszHeeov7X
tKcsHO1zpHEGJ37Z5F/drI2M+pQcVXMopLiTG8jhO5TNT94Uaw2Wsr0N7dKnum/NeMGz1uER43Hn
5bxfjTOoepMKmGPkyICp8QxnjrGM9WteYQxAbxhSAdcDPk4QUqOXFDsjf6pOltyW9Mstk5NMXWjm
1TZtQY0zxTFV8UYaHNgwcwCZywZvCyL0O+TMc0VxRt4mUgvg7n50CVrwBI24Si9jKQt06rRfUFdF
rlT0anxOSTia08ZWX1EBdH2Vbv7DCY4/V2cYJcvcAyaeS9Q9MkkXqFnxCmYb3HOETFY3r1Yv+dM9
kkrqE+v09KE+lgt/K/D3J0CvvSqyx8P4EIcYTtUG57bSF35tYAO9cLyCtCSJnfjoo+qKIWNCec4K
ShTnRoMvgwYV+NVqj7kHX0PyijJkBoTRmoh24JKQ52jrWfTzxXN3qiI6gpF7UtqPqy0DzJjFartI
/3EPnDOUitpHX7vdoEgVDUPkaFLgBjzZ7A4n1WYU2OitxNmyd2Hc3VEn1eJCiQ56VEEeSRDXHiO+
Xe+/XudBtJ55LpPyvigCXA7FodM6CAOP8uzPJYwfEucZyuTkI+AxB60crHNePZTlrrRMwGAvEJwF
uC5g1/do9lAQK7Qh28ohXUnYA7ISMn2N0DUbMbe5J7af9zax35Kig3/Y3FCIQDta9k0cHEd99fJn
5HwB59Ej96SRexTohbfUQX/2gP/WouSp8fF4HrqIUJdqHn1cj+zikcQ9Pre8IGTAhds5T0VRGuxI
apiRItt1Ijay66NWcG4NXncqmzFrS/fcWJ++yMVyBvLVvuA2Tl3rbcE6lZo+ZRgKL6/O33D3n6aA
czT0/uvLmHFJCt9MgKqAMgOq9aC3JjbGhv0u13ALddurn7ZE1lHLbIIAruWVNVeLsynQ2e6b9UU+
EkydROR+WOK4ZG3dvyjEsNq8AHW3p6NP8cIa9Vct8cI0s4WDj1EJV5RTprANljvtWhX29ISUg5JH
msDQzMR4ACiTLvgx4jV/Xa1Y8j7bT5BozToGlfsvPLS6e2Z6OKCEs8e69fNFZ8bcX2I4fGcG3U+w
NabcQX24TuqX2F9Y38NBJWipBpw/qBp3xDnp2yiE9ZUILO/4ySsFBFThDVcE2+p7CRRDbZzbWPPB
xP214BSI9bEHWM34uOvdiyUkc4lQgZAluw9i9CjrL5nFIzUGIBvEJyHGnzLoeWSZU2lsREEbUyxw
BNX1LmfdfP8BxCozM3Cq4eFQdw3k/N47I2sbgcq/Pmd78+aKkZkRcfbPYhZyl/f0W68lRa4WKRfn
wW7l3KiUNbdd203gydJa023FtGZ4z7bLv/SrSzvXlVn/90QwTxTfzqSgfXhRHCKzjmaHjq7crDEk
QlQaCkQPNO1UeNulbKQHjix8o6DkGwrP5/OEtMZknUnTi53/cuzjtZD6Ma1cia8tabYPbiZ1K8tL
cikLqXYPkLIJ6Q49+dO6r+pl1EjN1g91YhKoHUSdVZVgOwtml+5qHxIbZxsm6lnHKcZdQmFN0UOq
V3o8E0pImJB3lfQaWXxpTUi0yMwnTSBC50l/cHAmnEdTnDrg7dbgvTcRC8xl7QGLf6/DgGhT2JXY
oh43WBtteTayG02lOV7I8Kirt3A/vlgz3QkeSrETNPhM8dpx9LvFnl7T70OAIhySHeT5EtxeJXlT
ntmSAHkHUzmIwSpbbdU1v/fGIvIcSis+auxmWyzqyyTboeUkOT6s88BMSJQniGRrTkJ6GYVrQp9E
w6mkCWptV6C71ZQ7A5tydozuRHmND6sUODie1d2RDZqA6tO/doaz9oCyofdZVbg7fs938YO797k/
lr5vPp5dzOHjAUMUZ0oZDdxAlzO7Owjwap/AtUf0k7rSljLQChmrVgao6aRHopaNsbuj/Dv/2pkY
VxArNWoadKqq2FwiNERe1wyj+FgmcqPlsLOkcy+9GhwjY60Ul7oDJR4PZJGD4P8F/UqoQwom3F/I
OD5X93D6Ua3RXo3KRrMa2KuyRkpQgzeNBTPkx1X5/otrPWXT8DXcTSalsF1HrgTLA9/LQjhH8DSe
7qjDwNVzj9/9nA4441ZNnJlJEJrvVeOounpLSnkeKuUxS2KiTF974Hk7wALUQMUv7fWO4Uw8HyD1
7o/7/eDQpHRXSP1vERVX0cjIl09yWYf0w70HvV9AVwGjhSWmmEGLzswHOh0v229IFmyuNN+i4EBP
RxGhDeDU/lZz4oR3WYkM7NS9u5BCfNejBbOoNBZ21Rgdw1xNaZ9VH9/+9thKuCYYx3uUc8bJ7EM3
BQqOfTv4o3ZYXe7evoE1LiVfbUb959XZin3PGbNV4wmjvIv1AsZig/8uZDu+3OUYNLRUUof5/g8k
pmOnU9ntd9w8FQJaY54MfZPh3XhGYgHAFhyQotJ0QdQZNMcWNjvzqWwdVxciwDAgqU+u7daTho+D
ZMPl/XESCFn3jcXm3ALjr9VPJ7jZoMzQVWalZZRObk5t6oTmtH1/XqJv9bbSOU8LO8WPEq6Nr7Xa
35mvRwkTDtxq67LMdJ5l6glxHvt2ZJvbx7owzyl+gwRzcGRprsp4MC2rdRflOdRG2IodRDqYjWRX
UtWnmc37NTZsZwXlWC2+YtkIOYX63xuzo5YIOz56l9l++fKo5UDO0qrMwNLuo+59ow0l/KZNd53s
nYoN9REKp2G1jp8s4x23o929B5Xit0tu9ptH0BmK1w3W1ymRWC9QbFVmG+H9HyBCgVdh5BGj2yDn
u7QAv90UXy4rbP2jP/55WoESARSUoZEDM/BwSn1VOSVvF2ke9GTim6mKWc5CkzuNyqIYOFoO7yO2
pI2ky3HpSChIXO7asQ46iWaRsUiv86FLVtMHe9uRSfEPqlq/o0ual6qSLxvXlYiXH2Ul0/fOjnx4
3w7qNMEl8TfSpXnjTlHyEROej3pvGvLz+Ytaocb9a7fsuUUJbCLZCMKpOHU9G0q5FO9jznMUWOu/
k/pIVbSOQP4k2xb2Wgq5QbR0anF9dNwmAKZJcPWl3qdxbIOyk6j2KBvlMUsCf8YQDQm3rB1EjLp5
IAs86o9/IZWA8s7PPAqCuGu1CMO4ixzWp7T4H2cTU+0hqvEAO47VmPkbhlTPJJbG75uAQz+rnh9t
tZHzH9sJr8wMlGt/ynfuBDsdtnUFzelLamOm6O7Dfq/uyRvXXxeY24GAoPzvSCBSHFe1TjR/c1rk
KS0L1jcxuHqHiWwi8a9MDk8f4sU1NjtYWKbbcqolnBPBQrwyE0m5aGevhx9ScjkNMrt4eSpvU1gs
4kQL9uSNn7Ji2kXyIlAlKoT50Lhet7zwOZ0R5OmrY01APGrA3yt640EzGzNFtA8LLXQblt3KPfDc
098cwOD5aL0EmM1ZUXfdn3y6bMaDG5AKhuTjBx7C69qKYMI0dmfemxjwWVw5tgVOqJ8wo13tCKmG
Zdh+H0kaM0niTx7nJMgFIlsF/0h7wI+47moHTghNkqeTWncl4g1ogpgj+7sxb/7yV+met3pH+JNX
3OwjB+AUWlz9X2iHwhRpLrVKrdAEZoFEGpnj83MnMoh8chZNWNR4jObtwisDgHx+R886TGE9mG/A
0gCnsfhyGLKufzzHMq7rRyPzmT87oty9jZ2FU+Vcp6sheTukq9Fpaj0DE8+/v12NrHSEXKZ4+tqa
eZQV2wPVgdj63YzEQu2k0ATlidA+Z+wCKi6EiVTGGpiXOxE+/C6vFMz+gjBHyZWysVfqzhfjGUqq
u61mICZ9j1BasI1PaTbca1xFGD+TjswmGP40bBGx0X4IoEHAebGhObXSZqF9Wdf2WLHgfm8ZIiQN
+ExXeTWJJlF8SCRaTUWk+4GpKk/DZ2bN0u9tUyqthXng443IrNiB2NEg6cPggTHAE0BYEH2Va7OE
FUV4aI5HtdIDgdnLkMY2gskSrPXnnp5Gj9Bee2p439Ki82sj9tNhUMXoEUu9X0y/3WECeql+KYHJ
CeDzUECEmdzfGvERhKXhexfntBOxGebAavmMTYfKoVzFCY8lcL0NM3Wu5noLthzO6zYIaGshAv9/
6Tz32LkCOnUWUE3mIx36R2tNpDD+22S0S65PD0xYmx5EdHd53XrPNxj/aWwTkAZ9NS7zQJ9vqgOB
3nyYdy+PdCXNvZzr9JBf4XnkmQRLBKpmCHkdZReC5TuyhCuTGaEjDB4YTwOu9EbKDfRqbbb/ORF+
23uggpgCBHTtT39hzDs1Th+3YTF/T9LLUP4+/sg66lb7knQDjMhLVYnHeqWwW3l6H63wm8/kLcE7
cDrX9TyzP+yJqURTLMYu3brqJCvvH77BmL/S7bOQyriUJYzJX6ZoxcBP0AjoplIl08ImrVQ72QKl
DpspYVtb8zPMZ8OzmKLOMyVmk87FgYcZxt0nAhJs1ICQOfNKFQ9T5772ZjtJ422u9KtP2XB01aAc
jHZlxIW/kAHWgFZuE3Vo0vnLfY+k4GsYsafwEjzKOiLKv+/vHCuIfV4S5XsFsNMm+YmvFu8E1LGL
aPvjg+FCAH6QqjxLv4QrUFi8uipm3c/ds8RY2y9nxB7WbwMv17Ie3sc+XF5MH6zVBrKhmqUQPoFx
kuB9/Csbs3c0qwgQvySX8b3GjBuh1DwGZualoi78pKPuRoHQbWhTtoAOMUigS7t9R654O7Ddjrqw
xqg5Gyj1czJlyDOr7NCLoweB/daIKWQREHHe6yiDGuAxH55QNT6hwDa9f9An9jRFHFKQ1KwWrVfE
B4bFAn0TbvBC7PBvGoKNDCfkwYX8W4hH2cIWjUYpDFfrpZj8pylGMF/3v/4NlNmi++/nit0K9ns9
JhLLdluBFfcFgPb0FJDsdeEafYn3c/r+icCyc6DYMGModLZFEDX9WBSwzD48qg8WkRpXeY1gC2Cm
HhHsOqs2HozzLWPeqQX+gMW7EaKKRgACwjtVfsaC7AeIbzJQMSxQ9bYw3oqh3v6yAlFABRFx2XBt
9jRdx/6GeMcaoI8Bunm+Z1NXrVXIRW5HpOx9VBOGKMnNNo9ocNzZNUhfOLuuVyGvz//rJiua6eRR
aIp+9GdTBe76mvo004KEVoqu1yMLB1tysRK9fjXoR8ZU2MZwYkASbSyyKVSRMHv9lZgh/ijlfUTu
dAt6Rf6W0NnNp8D0Vq0SmhMF0B45N3O284ZvChM2J/w5Ml504GLF5Cj2f5jOnNMiCmc3BAhiDEA+
7oRjiaLFmHwlwhlCQ9JI9MxHwlEGK15/ACKJMKrogUL49wWHNGPYKpSi/O67FhOLk+HMqva6Dk4N
Z3hMKZLvFtO56QXwx9KeT79i8jwN9rp0MPepLNfwEwYTbtPtm9bJgU7JCRfaarx9/QDbuI+SR9vl
ojPYXinng0GdlckyUjGmMzZuwh6zXXjIMY/WS+e+VvgqCdus1DuOZEHZf50SLSRHdIHzWX+TCHXX
V1noyY3bCIx+44g6inDyphOW/PnlEjS8S0BPlqWmNJ4oiFSswVvoYVOinmcbF1QeKvtD1MQBc053
45vdnUdoNbhXSBEOZP69BdbDhIDKkwY+k9MjMtdSGMdlueRcjX6QrgG1UrJPwAvNDaLU0i8g6Fre
59PxE/xgAEB+tnn4MJ4vKZkkK8UOg6eAwNIOehvYJhjCkE8ieDvx39SzaGp2ewbFNwPuqPCK0niL
CroiWa3LRiQgFJtUFSQr9V+5ZuG5bgx3VHm+dfXuKgOhZHSNYF2xz4LeExDc3I+43+ZV28Okq71s
6lEvtjdN85VnKZvNs7sx8s3AVMvmTrbB3pbdOg1XVR1rQa39tkOzOCbx9fxew/jGDdPVom6bDT4f
XhdeYNYWzcNl0qjF7BHgo4jjYjjlv8fp2deorg5xAKxcImFtCNrtsBR75SuHp5hd3mDJ82CQXjdg
ojzHbGTAnnxgOO1MCPNO0DEzJaI6hDCBhpT08y+h/BKA61+3fHpzqOzavKilZc9l4GmPsPqTVAaB
21O2FdO5r5c75EGQ8jWVCSNOYATaRYm5A4eymLvWER3FAerV+0l3uoaxJa8+8spxGVxuEq9ZebDY
YvrceIivV3iaY3ZWH3Tobmm6OxwEVIxUqH0qoFVa3LNfrm8XR2Zj0YpoC2PCixaIVx2mlv2FSERl
1NIiogunh9HdsAsjdi68fCDnnPAzsBRmHAkxT4f4JKDbTNQNw2N/NwLbH9Zc0pLkcGMALOAFTNeX
tVN/5U6G9lkL1WBVfhqieZFd1uc2j89zbPHcsdfidSo4bbaFRSmCQ2ZrdhGXhAXSr3ncGVXDf6s7
in0ldN7nbRzJmAeQNbAY0dBSDBNmGMv0ewKv3jgSV93X9PhnSwFhJdU82Xnfjb3V9tuxT+PJKSeM
tNivG+xGLvd4cf+keHiOfzmRiPbBx71hGqTr0L7oohjzVEsD0rIL5zP1lJZ8XgWPDIHbYQge1kaq
3k359874Cx3tSzx16Y0Rj0e5LfhG00K5HdJ8FMEyFvtBlKpVNZpH2xhmftAZUMIMQJRqj1lJIhUj
m3c8b03ru/ogcP9KSQAuHOQC1SNR8DJXGFh9RBg5Gr59BVw3LXUT1RG/nTfPiVnw81T8mDgCn09/
0rZ9oAo/8fWsl3/Y6lPOHqP9EBMqHV1BlN13OJFTIZl/kfs3Qo8IS5ENoc6rXRrp05qkmqfU
`protect end_protected
