`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 110656)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf+kF
201k+6QR2npVEY+494p8x3Y/iVMzNwQUtTTNrheBLY9h8bbdcsKyZaY7KuUU5K6Dirm5yCA5/cKy
fVLBS9aoQtd0++VTEa8JiZ53ivfBgt7O4dPUrWryf2eOg6vahaqyDuI7QijBHrtM0mffeC4icvET
5KSC073iVZMgw0Z2so1EQzosT66HOudBmWfbcElxS81rk1QZh5OjzgLSlSqxFjzcvu5rHGpQcO1w
qnaGuoQFnWjNoSBKSrzae7L5Ftf920LUqRwwTBzn5W+l+2DkbVEJZz+vOcY+z2jFD7aZSVSIIL1O
wK252YqFpZjDOVCgaCNjmWl+wBEtjhptK5mkqHrYNArkesBAdxwMDfhRCjabFv1GWh70PaPBrtHy
xtLHhcUEyGt7Uj8Fmi1Mn8xu3J5AduHH4kLys8MzyD4ej8sIYC5BhdMOlb3/CzY98m/4CPoSQwyu
sjIOavnwCGYLV7tPkxqjoNPcVUVBnlzeyaty8mR4fTzgT7pn8Wxz+qWAsToBbfvrc6yc3ULGX4ku
9dE8qpMOurf+tzHgL53mUigT6wTpjyH7LRseYHKs/I+f4A64mNXBs+C+wg33fvDl3yxwqkT2ylHS
f+8vkTjh4OjxEX5/khVWDowb9+oeSWkSBf4yBU+yZl1lgHPXI1ZIZFq/JuAqi0csPmmmU0/RT7BQ
su8VulrppPO/YlAIDcVi3KwVtCkmaV09z+FEup4VbeRipyEVpAB9DUNaFCyjAUcVbbvJfBU2hA8w
HKD59tiRvlwDA3gepVbAXFmrkujLlH+Nnk9ev18QubE6mC6zPq5jlIseDA0AissvrVnHro3KFS2v
ILX2Knnz2mrAqF+/AuP+pK4wC5wObPpcPfDhW9v+4Qh/+NZ3GaxrSNtd1aIP5WeTh5n/KNnyzEdq
JvW8IbWoCTAtpP72fQ5ubQmM+3KfXOWRsb5Xu7TDPcqv98ppvoHv65QPJE3xuZo+GzG88l5+rwzY
E2XAaZTXdlPaRovahkaex4mC4sueHo80tLZsZ1tHoxfyfLMWvexPlKcMrUozBrZguFUFFh1H8JmW
z1TQVNjaFSbB2iUtYLi6+jAmgI46p02Td7f9qHQ5mLtxNTVRDsm7xin92m3Zuw7FssYfS3C5CeVJ
7JWLzWONg3oX3DvDQTDMciBVFD/eXOQaLRSWHGlUcAClcE3sRjGND5xHwdAjY2dn9ZfSds6CMCpp
aHMRUs7bR+Y5x3bYi5TKR5XRBJZWQ0oYN6fvPU44XM1m9b/TiTjmDDgMPcpEs5NHbvThp5RTBTFF
fyxRkc3sBJ8sQmnDvexsmuqMF+YOcYItTvRQbUQ7InN8lFxYOBgrqCCcw4pQ/tgilsEvLlp0NUH8
lzyIqDiO11W6qDj+0TG65cgOIp5J6WDm0wh9lRHAez61adh+TsBGO34N+Wa0eULto2Bi9S8cP7iV
KzghSp41zR0YAxhhP39z5N0TEgC3bPkARRPcm9KNf8YhvMZ33qzUb65iGTTNiH429Bdg3+7W44YY
JUsGdF/N0qh76zCkeOItivpfI3qRuK64rYBQhJs5qpWKC1qhfgemW9wpuLZiO2ISTipGXEi1DtsD
BZGzbv+0eG3Hhu+BhVG+ueDD7ssTYjddtmu28zMhuPAPSGdff9v+fwDBAW4jktWT+BWp6+F1MnZi
0zUrt1GZJzUHb6T0BTKaaJS8GoASN63u7d3ceXypFY/BWQfC9G0y3j0AgC6eODj5OdkMlf/HwCDE
QrEGgBOY3qDVkwLNKIkqElL9ECuoTDqOsrCf71a5gYiyVPBVv8w3d415XWHlIg3mSyCbnMrR7ZcM
EIvNSIWsDlbbrLA47zF6C/JwQIJeZjsns+yf9HZQE41iFnhB9XOOTP3iUeP6U1IpO+AYBRhFRTif
ih6P2IqINzPQ4AkVcpJ04F8fgcRJ3j6b00Ts9jVOF1hwDeEWN4EvTDk8Wn3xGOpTDFATHiotto+R
2J4nAQFAJqUY9GF/zah0t8zAecoPynXYV1hDZ540oC0Go/Ohl2fYhLi1ONmJjKbZ+6SIGzwj4+pw
+ULkBGGKQT3NbktDjus7X1kWFzMA89LH6uSwFnqSL2o3r6nAlj4rPKvwzgl2x6uLdZnE/aT2DgLX
yWe9P8AdsgXhOQWdqlf3I40K+2/bnxLT/T41QVADtaeHw2h8sq4FYkOb4l7hqjwLik1eVW4ypnaF
x+iN/m3AcHvoiUoTR3RIfwfx9YukCYBnW15YMKn6/+0BIc5gzoAFryIayPpuNOIueIDTJNrUoerE
NhwjENn2KmulgrzcNP/DU8U2zUq83AkE3Pief3wL0mcIYb2WVKC4wgRAR1E5H0CIFy2q6Cj3tb8F
xx1cV+8hRwH6Tsu3oHaBXs2boydZf2Gp9jisG3qH2i69+p5ffs4aM6JVlu86aICxso4qcTbrxaIH
iG9zSm61JOEU/D0wiZUmIAx3wcBIsyDBoIX06XbsYmgCZnlv0w4MrBG2g4nIOyW3qRSBzryOo9xy
3f3rTjnb43onJ0z4J7TfcPCg+LWv2KA1SOQOa1Lnj2/HkAFpeeW5Xh3B65m0D4o5PCUYZwfKPYLm
x/7uucCYzenRnlPVRoSD+5YVU6VRxOd3pgMLdv0nGgfGxW3/PE3yrMdT/PuZBw5rV5l7zXog4ZCQ
tKlm1okizwuS5r3Ni20wp2MgtTE5Bbql/UErzda3ClTEHn/atSfu8OZbib3IhhLMqgsoNdvXPbXn
tT6lRL4nj3pOry6uqHJWRRquoDzUo9apJgiM7+/CG4yaJieQ9NeyI/0QpcQHzvykvD6Up0J3xPOR
uGXKX7FpVzNgH3P5hHjsW6JjKgKXKviLzLcntIaTb4plmXfXuH18oMrG1QbppJxboG+rbp8KzO6I
+UpmQ1WcvYPI0yB/5PcQ2VWpZrS3kUVRpdCJc/v+csn7fAXzl3ckdieC5ci20tPa7Er5PncqVi7f
2fD8wm0OezWs+veTNzzbqO2SOpgMp4QKZPKVsS05k5YhEY2uXPGe7bN470go0n0leFbQqyjN9vL3
Ba/0Kbi/VwQ3MSLXr9BR66apvnqF1M7+SVzxCs/slP+4ILqzCWV336TqJAU2wt0DyvbiPwZgViy/
ROTa7nUxJUyLyDw3zAVjR5HGPST5eiDZZc9KeQeDGtonnBoRFaFreqDHFd5hyhtE0u7Cdg/ZIDxo
EAqb3Subz7E0d51KhixfA/Xvd4xnuuImH+Xg/tbJHsamdC4K5WJ7iALxx0QEgkNR8TZZ/lDBr6RE
iSsD+s+6kGXCJsRGoJlzwqPszGrHd5tw9DI3ItZbupvzwpMay8gY34RJwBzoP1LbglcPSmDyxWqi
CHyZ4kJmv8p1Ky85cKjdX4pFJH4SEoTTskPU/3JuaLj8n5r1j7ng7vUbVXQsW5ZD8ZSsSV3f0Y6n
XSS5WX9GSRvZTsEIZAUBKQm+lm53fBynV6K6+c/YFaZKBX9YkpY2eYZN9dfV8APHaLW8lx2JQIjI
wmD1pgS1dBLWD35Z8yZrwfSPTHXdeeRmd60fQJK4E1pLd8zGbwAeR5Lrh/bM21mVvxCQ8w5/BVfx
ng7HlvfoiM0ZC3KEyhiMUx8jyhtN+JLj0yonW/Bh2GTS+B00FBqzhDs3EvBI0cCLCR3rWB/KSCBu
LXR72VAKQx2SruIu9sVUvAJnRgHMiWkR1YazA6wqNqa9ru+iu49A6Gd4TPWxeQkZwKO75zn2d7h2
0h/OwkW5s6sfQhkB8iG28/au/rAngTp8H2+VyKKp+rmmL6rB0BXYzuHlhgA9auL6k1faJoWJVlO/
ibc8D3UCptA9e0VXaJdLul+nAy+tD1tcHvBqfON55+R6KSCMyqIIc31QQ2LnOXpWjQlm4wLKZaS1
GRR4PaZOPjxNWsXe+8UlNI6M73/e+GTP97dF6uTKg8jCV3WAl/uhD0IiPqqA4y2eX3gx8mrlh2cu
d99RihhzHFADKx7qDSSX4D3uqZAv9olSQ/jw1tY/3JEMBmwGHU7ngJDnL7XlNep9Z+PhHdl/h8nh
y4Nf+tUrMNTiAfxRwhuaBOzXrxMpmTkm7+B7cSjiNStbJ57+mqdTLTCvcDlCz52wEB7UotTf15uu
BmS7SGBzzTBC+kN1wIF/9q7ayq9hPWg5ev1eEH9d+hBjk859C9WBG6R38qTN5sfQS9rpOVo/8oPQ
r1D6HDjNgKDTE3V69s7mRXO4HLFfK1Fh+pLoiGeQZoXMPyVmkpys4GbPfR7OqvcDIoTZ5+AAPTcE
gO9nzPBp8LpVUi0DET3YiBuTT9MdVQ6Xlib2f/9BGjiU7vI1ahFYA4l/zqNZ/uNh2iy5QU6i015U
FUYVgqHSD1VY8oDk9vyeDl4ntAnSsRkOCiM0zgQhU/dgeMdA2nAb/1kdDz+g6aB+BG5hMiw2XQ7w
T4zcwcxBqUbUVr1C0hkrEFHt2bTh/gX8fhob89J7XlwtvP4jih/PS0fswjZn2BYGiaaJB89pnfFe
IfcgSVegZtOhYCG59nrJS+7aL0SEZZjiDAALHHpkq2fcNLNsfeej7+XPVrDTjhCrw/vH8asoeAeP
Qi7rqViaNsjNSmtmup+PWQgjDPxw87f6yxhzyhlJlPCic4V+9A8y44g4D0194b2wN5AE+kTk0wJb
aKquB9NGM1Au91hJxgyDtFgqGZQHn7oWZ0rPrDTwu6ideNTorhKxkAVDwkNg24aMDmCVhQf8PMtw
b9qoHNU5abnY5bKbqQEdYZOMTXIyyCyoT5NJpAlLeJEXAlITj4hs64SPtrqf2y9jvGjOv3rpYQjn
MnTYMaGEtZzgRPUnrs8Zjbn+ETjjr5u3YhYs4OvFAVyK9adESyJ+EaLT+JOYVOWe+9QXTzPCUVmE
UJpsitToTWaSBmqacdjMMzajPs1fsKKT6aiycPE4Aha/YQL/zrNFjfFhozhW1KPyczhERD4aiKK+
55rIpYDHO51ZuPHiLirdhQieNuf43HjUoEVOzmMYD23b/a70i6AT3gxCt3sB9L0AWxSe5gzzHamG
AMC6bT5EIOFqFp4A2/qVVghXNWWFF6SO9G/mhhsHvfug0V8BwBBNIJXBcLVH/5Lb48rYBezCoCcK
LZ/P0FBtpLD4wYXWOVK1UAc4YP9UTsubjuES95sQWc5SgoW7EwxJ2jtygvqBHYauIHa7J3ZtPwz8
66cFYHVwEBe+cQxNAvWdIb+dWWWwNUSCiU5MyGxX+zqRU4soRlcBNlPMEofop67NUglN/pdWZ9AL
K8tWxcip6SarlUJ9NRqkL35W3PHSRCWgzEk1N+j+jpYhTXt0JhlS1kANSCS5EI2Pqs/zi3+YBoqU
qphKPtgRt0QRGMBu16xglE1ZKbn28mbTHXU1cFRtj3W+3zCRArq13Bamr0at3sA0srsUyObz7AA1
cRfGws4vZeRTuDnS2QLqonH98ShLwaSFON/yaYguqUYk6AxIoQ8MZX2CdHVBc+5rBMssXCwfsBcO
SBN/ReIPt3w+//I0mLf6sRkOzfdUlFi7Ugsr4/bC8GrCCcXdfobPXhocCXAO9TBXC2+XahDs1xQG
H6h0PsnyHoCJkrBs2B8iY/a+LcGMhv4sIhSGdrvoUK2741327xNMlky1Xe9xeGJx94Ef6mBJ9Trt
RJ39n2V+UGwvqwhPj1oGI7DXwYQ/ozhlYkcNPInSbe+fX6ipbEz8mIzNDh9fvLZpiDk20ZYXPmmK
7pvleORB5CrM8wEth9hNiC9aTz5qKLcBz0xf3sbQugkYIQhZiXwmHU1r3A0P1aKo4pGfZkFEAHMp
DiFq8ZvIvPKUUdUib+38J5d84YSmKgltN5FpmiSk10Q/naCFI28RRd8H1syEy/svQ9fgwAHt9v4Z
y1jUZMiOuh5yMxFgxExEr8jjgz0qC4QqYTXlhERwr1JVpNttKmW2fdYX+XlbzJnJjBxA5VOetr5l
JQEtT5F6/tiN0i0W8IFNSgiqayk70MHSajGlDv4ogcwX/Rmygs+3fRaZNqNXBqNu+6t4sMh7Nmok
3xOeOoKP4x3l/S7ZxFFr2tJqjo8XIj4t3Ezcq05m0Ub6buYCnGQsm+5g2AXG5vOpKSaqqEmjCiYU
6Cz4bd5wrWu96QGbm2R/rB7IIZW/v6Qc+NaeNMjVMMpKCmGQOlzzjPdIzaeS7amJLO+hySWcMVz7
aTXYPxWYqDPFsoVENDsinaCXJX5PjZ3+aw2gWGNFPSTGy2MC7zpQa0+vRBXvGk+qYpnGYtpAWK/t
Nig9nraxqOZCWkoIb9jfNZ1tHTeupI1IjVPDU6cKxgYJm0XIM2prbSjjZvvBfemD5hT5H4mpRaMB
lMCppPc7q+oaFSO0zm8w9CUyZU72Vil8gjZkxrFcuvNRrVGoF6gPTf/F5GP6d+MuHE2NJPZkXaqo
v0vE3nGh7tSu2fg55ELAzi3JUeGx4lAl4uehHMD55CkIkyoiRw/hWj3TXBJfQ9IKOGk/HitCHNmI
VgGxF+G6xfE2PW7p3Ev4hnUm/yzEE1Zuy3E14Ed3CHmYzep6Ol3odO3WAsLK8LG051ChdrEbu392
Blz0G9jC84CnuFy2xhHbkctQwq+Y2fc4/32nwy9eJbHjTig96AoO8Vh9bKZuVRt8wynnlUuJ1pxx
SRV+N8Q1FNGA4cAoMOzZj8W4risYjehbZFam+K8tt3THxvEBG95foL4AFOG+Wm30w+sWMHq7hAbx
vJTLAl8f40mEN7SmHhXaz8mUAL9SsVjFyt1On0EF4lxbyIFi0DkD0oeWbuKJhKLDZypmr01cR9dY
vKtYq8N50amrxwUxY6y4KAmldrHvMO5wP7xXOdWqKacN/NXuZSuJXn2hiIgFAbdB5a0EqlNbI5iB
1m7OI1+Nlxc+7DyorEg20NMylc0lpLwBvI7wjhWjm+0yBJtRMvFcq6tkG71Kzc28gEp8M/BlUdGb
p+AK0kj+fxz4oeA1xdY58hsddcC0runt5oH15RzDnHfp951WC0c8UH1ON+yFxU3pMn1pM3Is9UQX
uFBbvRs4ochhD2YpadjoyyM50YWVsCC12vVRVly+EDexHVNe7NtikDAc18oPMh2SWQRdVK92JbLT
OdxCdFX4CZANteJWX5qtGYNoDpvAOH6ahhMAIXemtkXinDZgrAg147oEy2tcuuBdmh90QkHW7cMH
bUhvbPZnZMIIV7V24W8nxkSdLo3qHLzuVTg9VW3sDg8bnmDFXocKyg08RJQnH2fitBlMQjstOzyn
rOmw9bJXbJXdzIJGQcAsflELy6tPPxDe+KbWBNjh6xZa2p2m1tdSGekUxuGBJ3f01+3YkTzIOGoO
Scbw/8DwIlr9HJP9N2BTOWUL30+pwMlXrzPgxLecbEIZNHba7bf+iCwIXzJ4hMLjciuRcDM7j+Sl
Dc7LmCDRwRcWp//7xRn1l3ztqASbMnnOKj765Y9ZsnYuIVR3y48kTSThvZyhBkSMrrXrL6lARbJ5
o/LE3hGyGVhDQA2IpC2jhRbsXpwegG0RSqFGESGj5/5UVMwL2ywwYLscdiLm/3fE3Iagry01peQ7
lawmoTD7oPrwMV8/3qwMNZAr3QBMdv+KD/3JWRmePjkrWbu1a6sbRS7fYunP5zdRvh4vBfRb9oR+
hGluzt485gSMFVp3fJXd6pfOBZvxJnm/jpkSDgm9TF6hzFztcR8cXz6qCf5CdjEkLp9Ed/LcAJF9
Qw5Foyx9gARZ4kBwJ1W2JuufoI3ftQEZdhUlUaFBNE1kRqGqWblsXdzNTpBH7OwoTFM47fq0X7+I
/PlLBVey6w0Jt+byum+vyFDx+qwIw3jNQ5GMU6alSLnB+8m6alTM+RSwDEbwKyAtgIaKdX9rRTZy
XMQKN86dCPDZyU9/k2V2o7IRuZKMxaJFk8XXIBsyU1OBQO3NKwy9KW3dTisDChtoU9wofUssu2xd
kZBI0RrZk9fGd9Uu/ErwJRux1UpFtvkXI1gFzzPzqV1yeFh15K7DsDFPnr/K1LQp8rfJCsBJqELc
4NHH7j6+4ggyc0dX3Uwo0n7eZQ85Pl5g/18fJ+tzBBtl1I36RzT85I9fODKcBtnw6KRkbhx4fwdr
LC0pRSJx9Guph73K2b3w5MrNGuMRlcQlTDSWb7RHADipPIvXQpN0eEHkpc8kvV2fPLWjZa6iKvMu
Fg1aAnfQDueYIxztnjFnIDbqIOhnHFBYcql1yegSoIqy2JTeADlJ3O5+Ky28f3GceQBtAdqW061h
L7wKi4Gd/6jYel92U/tnINpCwp9/UWM5iKG9vlJkI8+sbsIUfPNqFWp9xb1HI3LxhZVOwEdOMMA8
5r/W33ehxJkNaSwkWYAfPSURF2wMCfR5Ng1bK/ljTPvCFSxnfGM+tRADmnwrjx1s7BdXQXlHSlP2
p5jFYD/rEJwOzGGuAQC9Lh9bp250mF8IAjxfogJUCuByOD0GEuU7sCGg22YtNI008AN9eXDzH0Xu
NCBPnoEGgDOxz2hoa/CSfIVM4AyE0crEBeIsCndO3YnpCAGfgMRgfTzVuLnh9oRtkqK9mnNmNkjr
bWiqXOe2WtDOVy7Y5uIjvr/AIU/SHr+vYIn1PyIV3+T8VKKY9dNFmTtAu7ccx/b0yWLm8jZgaXMu
rGSygx5Uqe6Rd4WV0GbDllcoF8cXGTQLHTYDSWfsvYMP5fLHu5NU42z3y9D7cQDp0r978ykXi+rP
ac2VCRxDYzQi0NDXQo4WepamGPm0k5WKGjtAjgEupZ6zxOXOiBIT3CnaCdn3Q5w8NUP4tWKFf8P+
12GtUknKyXw8C8JVupsdKlccTFcPlh8Sme2fljiwFTsVg7MVl+SCDkuo+rFh2qP8TdnYDTUijKwa
4llq4sBq6uxav0e/qrVNLKXo0gudC0nE8T9+PS4Y37770SWjDgR2ZMiiKyvQ0Xy5wLBAByvjTcSH
w0mi3BVkJSmMjXeS/0VnMs9w+O4nXn/yaJ0XhkOvBiKO5vAzyCufcsbU2np9bavlegeMhHyaFQmm
Lduq/s3AjeotQrG3sb0PIYq4E5Yj5ApYleEQ8+8lAIS/zL7GBs3bVn+0bGZpR7qRaudIpVhM6zEy
HVgv2JjuFsx97gKsbheYRR8bR5yG8hDrCr9nKOCI4VqZ4agMKh7LpJTbNLvEYEf2IjpzfaIe2xLA
Tz6DXzovooziwaG0OSuu7ZXGCncTbwE5L9cioPMkur04De2tdPGneVfzp2X8dLzeXuw2GNcuYmI5
PG2x0AsDeyzbtDwzBM7AsH1d7tCNjimGUZUzoxpNpnPewJQAO+TRB2F8l3BBlYVQ1DlTZSP+ssI6
1ksNPRxs6ut8gFkft+lbBi10RDCBmGih1JdHoDZjKXwOE7f9kepdPg57TlqE4qrrYMfjufFZtFSH
Rk1hc4m7d/eVGNFcXpJt8R58Rwd4shd2QP9ATJo/b3IEutyahbfYBtXD5vMNhFjEsPdR822YL/v2
Rgy1Znskemvxi0Wfcd2aB9cw7eJLBlUKi8v5sHEjZLeS+rP5Gl3W7/iMv4qlmFVTK3s0eYEucEfI
2FaTtLNssBcOxDNQGW9I8syyZeZTJGLKDrCn9Sx16PoOgzivFqFzoBRVkXu/uYE3ntAxwH8uS68a
apIfWhiLDEIfEBxVS0FSHDQY3BXsASjI6L3fAlB2fIX5Tjpf7wmLawMq3KrU6wtavoIzf15jIX4e
AJ3n8Kd86/57nK6f6GnzfHDFJBezobJfciUBk80hAqqifF5AicOiYebPxwcnXKKqv01dNYgF3Ob+
+Ps1O5IdNk3S7RFHzEKWsUU96+xBa4zafQe0YG9oTZ+armQZkDlzuOGCTelaDQMM9QWAFzfdyFg6
npgY/XmBOHhMuwhyB5Lk/VA3T6G/PzxLoUU0xbqF5wV3CEskQxDidXTQlZve0cEUa/ZvzPu/0Rvb
V3295mJVqo00mRlB9y2+zZiVIQ1cNQtLAIet1J6vzJjPkeRAc6xXi8Tf2FxOl78MWgHuhqBrYy/s
I7q/bwnQYhVNK13sDeePaJ/+gGaOKXh4H1kmvHEIjiGIYrSVVgr6qL43U5AKG1Iaj7evC/2qC3C3
o883lNeSZgQDREDJfze4p5EOagObW1QCKEv0XyYIIW7lO+Rxeb/e7zMds9A1+3H5waJPXMfP6ITj
FaXVMD49ATvOMnWi4mZPCESOmurOlDJpYNI4tDSpFXjrh32IetJ2ZVOZTr/lq25uDGmLs2i/+q77
xyGnd6+7lnMfOKETWSb//YoqbFsUyE4ysq1TUm4YDzBMRfxiIg9Dycz+Teq6F+uGDFkyP9PDhNdr
nYn+ujTxU0rn7voLZnNVpIbfErtL2Bma/j+xxKWM60kORmdWvcrsIHHY+Zmmsnef9GHl1WST6c0+
M9TizcJx+cvxd10T2r+qJA+PphBoFV+I/3Wcjk0cwgOHvx2D/sCQDfZtzf/XBs/ApCZQST3ec1IH
HrLOXA8wgr2ana0KBHIrSblxs7LZ/dTUEhO9xybg2rKA5QBJcRKvnE6KLc0xCvpu9HhT4CZj1kj3
ixLoEXQB/X0BXDUksz1S23/qbDojhvqrwOXaP3RzT/r2SEMvKS3FYbuEEz5bh4cl5xJS5134FPP+
E/d6YtHu/NxTbUGZ9zTwrIbnny41RDLmnC3owRp0RQpBAdmEwpTfH12y6bt/cEonosYwvxsjv+bL
jHZYtNGNa1HeYIrtRgzT+Xxd30rappnrR0unr1OU8QHH/YtqgRJ21aO+0ljBghkEC5KItCDavBZF
Ll7rphuOh56AdMS/AQgNq1h08ihVmRClj7rErIgeksRVMh5K1xe5xNJXR27pIgyIbmykbS/XHTjp
MdZNJ/nyOgRjNSLyeBFFXDFlyunGDkLqnwO3yaH01y1oG/wD+UnBmqJKVtJSTc51kYlF3aHpJvTs
I4ZVSQwHwWBRZ0tK2lgy8ynRfiDsHSyFmyGecaF7GW59janCQYBs1XYllx/sY03Hgc7YaIKSpeHa
0MJQCEshxO7/YrErG/DeyUsFfhbYgIlVlp0FHbX+ZrlLMFHGbVKdEA/Cmko3BDJr6JkME7bXb0RS
5cxdsxCQICgNbbpxJYs4vCWdUKsDW9rvoC57Mu7fu5xb/ni7Crs85WZCfd+Oa4DBloDDlrPELEBg
YRM19yO5+W0on5ACrje1Xhg/1dYMPyXJHB+vQmUOiiG9KEe3UGe7B0T3PZqdloWzsRixAd234Bmd
/HqKmDs0Qr22qQYbdF0/q3+ZbRSYl3DVKzka+6sYfL8hJ3vUhfII1P4Up5W5gDjtbtgsaqb6UcIE
3LM4INCpQ9wnfCaQDogIlrIbxYX73Sz5qIwr0jprfU3K58dUnYbnqsSaiWg0fpW9wZbq03K/DIW5
jg5Ur655tw+yqUkLX53PvsIVxskeh5gecZ9qA8gvk6VtIhh+3PrLHeIsYI1OiMzl+YsJsTtmmTIT
lMG/MmfL9sEHFc9QU1FUznXwKXF31WAUX+/wMPGIrvogW7N83cvaD/nmsaxj6kZmwBFZT3BXNJAK
vbE2Q8vmADRNElrq8P56IyKvV3UScPMnY0oNMqBDMS1+qiD7CefBuBSz8IazvN/ChKomK4OP1L3V
RAv/RRdlO0Ciki1apso7AHz4hDHRfU6FJMhiYYgV/bimi4Mo+XzWz71pmWI+y7ba35o9EZjjn9Ms
T6S+NApKuMvy4fB00XYjcUjQE2UzWAHM3/LWDbPHUipfUzFWmNMgZJun+1b/j0489EQ1PutE7rWd
IVgjINnLR6b8/v0VCjdoZ3YSlPROm+0DXiWaQO9PRgOCN23skf2rootpCB/JQpKj8aW0OZtvAQ+6
rpP1nb2AYYaAj8TtDmpKdIWH27z3d3+FGVTPB2FmoK0PZ05a3ep9UG/nWCa9EskHQ1wOXJBd+Z6u
OyM4+lrRgNesTbT1WdZR+bC6b8YiGJQL0ItX3LE3UyYHCMQW90w3vCuSY1M49iL7nuyTjiG23aW4
/s3tHDkXPdA7UZ3uJHW3/QPpSk+cD0v66MUvAttsBXJNxjV/nj1j/bl9klQzkDNYZGaa3MuJ2Dc0
4U2JgrEpKVeKmhPQtoA/mdlkQQEDLwFwE/QndFtL9XTSOn5MOC/EzGpyPFBqxPGP+RgiW2l7OBrV
Xk20YTFvzEPgurJpjfZFNdY3ynG+39yz9tG+YKdgz7HMy8Bf2Cvi9JF+4Rl92r/IS4zWJnzLpI92
/PbVv7PRzXCrBnDdvO6nPwEoe5N4Gz2ptmK4HXU/+duuEaD8Bm/4eFFHiALzy76WRc4yLDqjy1e3
lGMS9B4mKaFOFfzU+lacr1LZMYjRvR8SE4SrwaGF+9Hl1hcTPR10ixeS1DQ3LcT1gPy20Q3OkwtN
6nAq5kxTZLQtGfI8DnM0z8GFNU6upzDbP606DfdfTwGqjZCu5L2w5rID7BcA+C/56v4YG+R5jlAA
33KSnQcsbRGtOzx5Dfer0XzpxLV6ULoIJGKTJ2YFAxLzb+jM+RwesGkSi+S8/c92buKTf40ANYJb
Kr7oldrTJZv2aKTFmygrWCBfZ3zk9aam1F/hhwBzT8dDL6LRY2Xgk2a6XMLoCBCHlfZ3NlBBwmS+
DRSomu2PqeKZcpa5F536Rh5Bw9oY7ADTUWeE8FLx2ZyT38bq7vvmcto0p4LzHsF8dc23ppv856SR
eFzPJbuAQbtL11tE9ybd454xFxAkilqRw798kAtjGW44N5q0YlEL1rIVKg9gknV9Udq7GW/zHldX
2sU2JSjgYUZJXLGfEm5uKcRhHQeQn3Qx97+TIDyaFTZRo8ieu8k23dgRxSy51cVmWSQmVcFVgenW
FH9Wf6hOKHytp74Flo/3f1joi26H55GTB/h5ymJBeTmvPT8sCUJIp2URlz/uU0E+oh4Ym7eddd2b
mlkFPyrCe/XN04WGAZ41n5DwHikYhBhOgnW2wsc9StzE2xceOlJNbNOkgfqVi8T1CZSUsUeBsNQ1
7LSavlS/oYsz7L/q2oRNUILetdUNVEGyFK9A+NnIJWsVQrvPrwV1QL8AL5xooU25qYkQKsf9XJXW
hpnU1YZ+unUPw2b0Ld3i+Dksu20EKLqzOoX6s+5QQDzrYm3fak4KriqlNjQdNPonDofj1H0Y0DGf
917r35RE/xc35nApBcPAxuz1pNZFuQjYdv7ZLJz2KOYsS8HAIG4+1L8rU0PQdYJpxqrUnh3OFD89
8WHGNvitb7jmmVG+ZyJYHt+dLPvgI00uBAQdEGVD8hxa5EJGJJWpZfeBmG9h5wcalceHmPT35lFY
S3t2KY/HZWUwvIFJ6/HyBlfg7qrYeSf+Uh2W2rlRQU/GnvXgqLCsdzDuOWu5Je6EeKhAusxEUwCA
QPdC3v5gureo8sN7xXpVOH4kIBqKxUqi5jG6XF2g6YBtcljDQVuFGHKo4W3COgmfGUGVWIsssw0Y
BrKBbZm3zMbK7vTIhcUjbkkAbYoRXaaE+39rDdMVQJvFgMmh6UsIuVdwYrgw4MSM+vGnWU1KsVmb
sHK+q8y0MmaxWtSv4WoiU7geGKCaMqlvRTvUEdQ4gOZL3oKtR04OICIbgleTzyrSvxAzQya53tJ2
VlLGOloYhoxk5xIiRst/cuTJWhqy2MZzYiJdaKd6jl2rUbdT96L2lEe0I7yKFDRfLNDIw2ctC6TR
yl6dU+OEfjV8ndcM2hDIn8xxWo8xw943tfXH5d9USDv0IQzzn2QahR3ZwFgsPPqJWgxYjGs4UwDT
W643yA+lXDQCtUEAdtc6AUu9aY79EQL/zTyARMRMp3s9WIoERioDya5nPp7W75BCrRMAhQO3DP/K
uu8+Mipnaq3o6Gpv8db1ToN7gUkvq60faZf4q3mxTFfgfoPMA2dI3zuFTTqiUMs843Og35eLs2Rt
aB4jW+UKKDQAGKrFBSsuxEjGK01Q0qOuSLPzGmi/347PIeGYeimIkVv4psEYV9XEHGfcxvK4R6/Y
M0fZOwUDO2cOFqeKt6vdAX18uskg9GgLvbnnNxWgLzxODOQTXE91Zvw43mruTNmmrcflY2rDzPcr
mWOJbv2h5loOFqoTFnYnmMYDRhkLEOJoxuO/A7r2ubG/FLj8q0ntsl7o23h+2SCXg0SEnKKQeWKh
8t00u/FWeNizlKA0yJAJZKrm2idpgtu+FWwI4cR8+3AcdL+JQGfSqTgkiLl8uae1cCV9K673CN8u
be4kX98dkvZ481NcpuHPLLRTXMiOvUpFcu2tCygA7GuuW/sY2VmE3RkEu2+VPWuPYRPD7/cHwzsY
1gC7t+WujzCLfzJ7Ai1FkIYE/MxtmvAtqbLzd3fNu+wBZYv/4gcSLLRKf/492mjITp5xrksRqZnD
Y3d4K0bAgu9ZFrxj5SoLfTmrlQIq4i5iNQ3l8YMXbrFH+YN4CeccEOgLlxryhY3GHvTrVZ1PUlfz
Q5v8wRuyHSyLANAxu/qplvXKYuxed87586DHq7JLRfBMpKTQ8z2iQ40aWDWMuoftkBkKMaHWcJEA
kKfax8m+hfEwo69+cCVOr2eWsqL1x+FAyWpvKBqzCIKtU1tFTqieOhZnJ41HOEI8tIiUyT2A6bR0
89t2LoO8dQSQ259a7J/GeWkhOt0SgTZ9Yuw1d1eUZp2ZChjSv1/BrlLWOjHenMtSfSfxs8XTds+i
H7gdx8feB4+dD7uIcVUc681Jn0MtKgLAh9r0sw20hp1k2Gy9XZAhgqZnSXVQ7dUoL560sEPjt6wk
H0F3lK3ZKxjXuqhDmruDF3pfdxpXpKjvFLQ6j9Cp1ipXBxCmeijQNvxs9Y/nUFobB46EPYN2teOF
VBb4WMgBcpnm7DLvc1quTFrkuN+zrWl4UBPQJWs/8RRD8JyjHt5MnN8/6aDtrCSUeo5dBHBqkHaC
LBAyBbJwqf8JWMBEj+BLw15/ytsEmLTLaua7N8+GdAVqEElBnwR5ANFLbZdP81+PEBml8B72BjN/
I+9HaaVJhX9vIUThbu6+nMEz7gbj5h/YbSCrOxlTUtW7uI3Kkfddbs7llurekncZrikNRw4nor4K
k+SRcZKSvGO+UCnoe6obePGRCN6h/xwPH5Pjyn6Mo0YFHB8SdIHOw6a8m+fJKamHQ2TQvnx5BFvq
w/svNbIfAEOg3QJcAPqPeg+dbCP/RUiYr5oWzwDAj/jsly2KnSYHMEzMkabNqaOnqmtB4CYWgpzw
X+coiDHhfaji0/HxNZV2EM1zLr/a1N1MdoB2iXSiw5DP7B4pAwQmxtkR15QROXoTBz1v9k/QcbnE
EBeVDEjQL2v+qtDQHWCjwT3wLI0GGOQeIing7sMPMR+aD1Q95hWhyMSll7dIPzvDyFQEpngV5wbA
VAoP/RngMVp9vto/YEJtxNN3LHC+cMbcxiReLFQnI95fw0YvdDcGXmDheiE5B8AJRY0DEzOORQpq
IF7gt4CzoWxwIT66hbLhTdL18Nn6epahngJk/ukdjxq3rY4eLDdkM4hpbpddCS17FpBn82MC5l1N
jlcBXnNu17yZlylLJneJJnoSBQn7twNM3V6Xhayz+TFtVwvm8U+38kvMcOLzCckZwRz5mpN6yuzD
VdG6syEpbeSRZIwZY/Ob0aj9yIp/O9yE5iu8/4peEN78wZFSayx2hNZI2x0f/YGW6LXvEk9ELb4x
0saWxZYh+gcXnyEfXqKDXMCcBu2TedO+tvuDU1BIKp64RI/G/VPMBJSs24gdkECi2Gu61476zgkV
uuizf343OqjLXPLfSa/EarrIcg7+bNdlsG+vXHzml2MZwKrbLV6QwsJxybS2tTzqgaM49RmiH+Af
RwlpknhXAigctd/zxM+H/MJXKd1qKNQTanh2/BEMQwgtIeS8fiNiy+1diXnd6PrE5J+MrIr4PYee
1AZ9RtUKc0Oexy2I6dAxhVA7kWFcQDsdZs8dMadpid4pdtymCO7ZGIAwwGHh+JEi8KIBLDzJKIVM
WN3DJ+R7oVn7jOa1dYwm7xb0CpWmpj8xiyEXsIV7fDqm7zk8gSldQEPXN1H+c8hAyHUGyC1YJFXW
LsA1B/WdXHMVrbX459FGgtcpZj0Xkq5bPrLqwoDMyRymCeE40YYYwCbRqe5jWQVbvIAyQVufHbM7
n+Z0nt03Rgt5nghoQK32RnMwH7oCzBsFmlkyRjBnkXMlxJ/DTx1o/C7CTd44aRdygY37KNEo99P5
zcIaofqhuQFc39UJcrwtK39BmINMfGsCkGYvPRswxnX61FAT254Y6/xFxixUFq7c+KyqVGS0ohR5
qsK7uLc5Lg1ix74DOnnqxIXM5+29Oro+avoTmRlcgWvsPCIwCGyUAYmPvI8Vrr30O30i2w7Gil8e
DdNBw3StcOzkz+KJZcv6YOfftH8OSWb991JvllnyUxorcC5YyvjuOA0lZmHlliod//jVtc3IEXhv
B6iR+I/rTCwZw2DSVYRH/oxLd25fWu2XqnFGZf8AyXby3G3inpxZ5cg0Lg5Wh5lcw5hVUKDRWcbA
tcXprudS9PfXksW3DNfkIcD8zXbWNw0nwuPpuPkjbPM9ohDdo9cnj0xNVoH043JSiX66nr12VyK+
5BXIl7cG28fuVf/9mq57W86DgpC/fg5599bqLEnzl2iYoyghGYA1W4eOO1j1uIkFAb3Jp+jLkFEp
vO/tXFt8g1/ytm/OlptjvQ+JyS6hZsPEPtzWLxO3i27jCFteAxnyA9g6/0X9fbMkFjUeC/i68PAE
ABCfxOpYvnuFKYdGV/PeuLQQrDdaiPIdWP23KA1zLtVptYqRK9VuV0ZEzUMgXs3Z4ImuaolCficc
UQ3s8bPE72WX2yaJFKcmeM3v62Bw9Wo8NNvTTbWNA9hes0uhPirILllcI+mI2qdZH8dqo4DvyWMT
gLmBqE5qcBavaLo7P7mx20eKYu9ivwYYvdMlFJae5BvYDKiaW4IE381sGTnkQPAdZzXsz9zUKwiL
b7YdX5h19H/msCKTLdoGTPxAJRSJTZjL+QInJANyFllJw8iINQ8tfRzQEu8kNs0mfgf9qEgYTPCV
d2mfD8EybKOmo5uRE4N16yA5MnpRM85Lp0suRWsGnLm8p3HgP4vHAdTHuKESt1o9H4h0wh+YNzAl
xmy545Lk/1JydWBjxt0dJkynAAHLVBhawTps+pOBZwKTRTIJxeLwJ15eMuJx7QqSOMXAlvZ2v9pk
DidnrcarXlPNIhkZ1vkcyUGySrPeDZPM5RkH8HYORnWcB1j5XGGqx3r3sSjYkPiW0Y8loDaijyVH
2H4jpNS7okDgsB2c8zSbapAVrVIKm6WVQ+xmOsIQA5zLIrho6+Lv9f5/gQ1NWXdvMYGry9OQEvM9
EA50mpJN/RRTid7Y0nhYB29U1Bf6pFzZKGIDDhyjbeCamt5Uu+MxLH2ZZa9HrdhU6cvnkj2xQVMo
mRxPccBCfan4YjA172VKZMlUHpExu8n3zrms+rxc1jj74xXqJntd+b+NXBqfSJ9/ZE40Fka4mgps
oHxupG0qHt49SxNIcvLYkulRWAHKnPNyibe64skL7crqni4jrxlg2dtZgq90oOG5ww38ZCBBug4r
fTDMZpfbxZIP36vk+5bvmpt8ISRN3yWmFz+S+derBKiwgIl2XzwpNyusJNH4R2UUXEKFbfZuiDdM
AI9dkFoFdMbiGePapxkPHabayxp66eA0fxdu0+V786/9TUiC5cvQ/rkHout5x+jlyUJrOIp5FT8t
ByvLz/iY2m0VOcLLI1yxQKzwhtFLXWU2aXt0mWARt9UZmgg6b1q/VDG6n+OI/TqUd6wwn/0eLabS
1yDRo8fKPYNVY6NbQEIMtfxOZpzaC5z3SsL85JEXNJi2Cm81C7FI1j3zhY/XtheH2Yqe1SJ+I1wL
w1rcvKxmMtlkYpt1lNwQGpChNJolwRt/avDwj7ShLAFF6yyK8HMmiBsDuDzbkt2FOvnzpachYCEZ
sXni9eI7reub6PXxEr8e8ErijqDmB85RHHXJgOBY9vZoz6TalWcqIsvQlpYgi5NIENQFllB18fjp
1WPgGg5Hx+XyoGchco9Z+rO+LOzw9+wg0PGByH3l5y5slTZiEny9tKALl6V7J+zRltCc7cR5BPfG
dktTi6zJN9qowy3wCIUjknsGndYeNhBjZ/2b97fh+OBCsulxfomKe4C62UZB9wC4UVzxnipI6ihS
j4w8lZ7Prd2SX+BUJfsEnUBdioI6FPja5Z08EplgkgIJ9HD3m/On9EItpHa0NFkQkHi3Fo41UN1c
xzH1602CRanUfTdtlHdjrUy6OCLkQ7QTB/tuZZQthAh4SN9RwEbDg3yWJM1wSiKVRnIVPmpHgDJM
YINvFRKVoC2q46QgCiI3VmfSX5zPZ4ivNMF7isV0EycDIPU7GEiDMB8YYtHkDN28EY3srWAdPaMW
3Gkom4AlhghjYDEYjAXSmAXIHn5r92Awy9ft8Bv1IddlZkhorax/fe4J2xxUyWpMmQ1T/uyIBcSf
cjaOVBeDrx8UpKHx1mBB8qC8mUFm9cM+sx87nJ6Qm0c/C9H7qB8XwpPp6dz0pYtUttVgGBZ3eGG6
kZEwu2g5XZPgb2P3tK999iiHpzeIQy08g+n+RrcDHp7KPgW9GtksfdnUHrNHVObaiTX8ZOOYJLvs
554QmnugvPsZKnvzzfnLp8/gdzHs0JQV40mc6MatFGHgHB4xpofSUaUnB/o9aI3EZUkPy6xVIUoW
TzWsuTv62LjrD/lzHIc/BtGpibX+g8ifHWl/4JLuw5mGwHTlkXkdCf4MOGXSn6GwV7AzLn5StaA6
8oJ8qJWzfeg3cj3QjrNycEbbgjEL+EDJVA7KdnyAo6FPlaCvJEpt3QKi6FfhU9Gghzf/QdJDPthc
/tXJoW5SDyefxlk4B6rZOPflKgPUenPxDR8ClwcwdpGAP6PAq1hWwgLul2O7t3+d4H03SXBHlHjf
UeSi1xn8PhNsS1lRqrNdELZvcFR5D1iF4/h0wlzfAb1oFHh4vCodtH2j/PYlC6goqTA5QkyqLIGb
7fdC7HejR6yO+Nr6N4r4bcsYEUxFi9akAB4eDpfKqwecu+Dol87pEXRDCT3NhiOr5QfOXKIfp44j
yM+eqyqECD+ODRi5yX5ZWRw3GCs5Yv+zRN67C+B0u7LbeD4FRtPTdYxAzujhhoa5UKFdU7HY/x2e
0kR3IzX+2XdCoYyGYalbYfmsj7lahmHwnNisG/fpkvcGE4NRAVtMXyD10iuNupBzqYJ+6Cb/N+sO
NSkzdIREus9ki3Nl0S7BqzMuXdkn9+hsJj6K4k7jjA7uRjH6QA2qmsmbV9RhqEYsnExTIBNQQO1A
jTeUD7ykbACFRjf6X22g9JiKwn573Nl06ltdULcTG5w+Wik43XFoXpaIIVBo9b/Fka+x6uNwLnFp
G7A/RYmD5fTcjGE+l7Lob+hq4j6VCdVZjGD6Hs0ryT2QDTyqu1cnBlcETIUC8Gnlwbwgz6SKm2yf
Vz9BmjHtqi3UhnPufZ4VMeSm+EYxsfouwgInK70cag9viB/9Y24sl6/bxygi+jlkqe2WM/SCczjv
3yqUid8e/B40FNQLjQuYM2qz/N1Zhi3VOU59hZbqGynZVqhqo4XJ+LOXpnuygML/NFwuMq6wID+p
QVcILy0vZI2XkbXM61oKtjS4wzx0MyFoFe3wOZe7KFDzTYNZ79f9QM8fii+VdeVjjQ4cLY3ia5ek
0zIWyScXVgtzBRnVRCstFtSO4TZRWxj5+IBaHjAf7vlPeuVclR2Lhu10wRkv8llRwGM6wsSXJGCY
Kv2nS9G1imOIWJ+JWpJE3suldmx4LV86r3V2pqTQustZyI1vg4krZZlCJnbchOrJMajZDETHHtzh
Rdj+yuyfctzgeJaoal01CeQLECUaGyDV9c3awRsbfHxZCUF7Uabb8tP3UwdqRp1s2bdgXbAR68Fl
N7uhJ0miXIgir3YdRAF+OBLryZRr2GpzBMDI/HFgoj+CPXZw4dbJAT6bWL3A4nvuALLEPG0TA6dv
mo63TE39khlzaP2QhrGtwdaWz5iwUgraL6r9OYkUdbXqzjstxbSpG6V/aJ9jcjOiAsJyTSCmyuSi
9fgDs/wt5fVmr+d7vhzgqo/F7wfSyizoiuJU901U/Jq9bivwDtpwO5ZEXfa3DX3TspxBdOnXnXlF
s5tAnBsLyLCGd/Vd3NIql4V79BoRRRQXxqvCTY5Hbnm7QBdDw0bbUpCgogAp1aYBUlkrtuYW+eq1
JQsjEEOEYM26CBCHy+t357XlCpiQIBO4DX6zz+tynohVNrvMmDEQSN9TvN/nbUnIYaeVv6V3yNF4
gcCwzzjk8iMr7k/ExPkzefSYq/O0LT7D7gPCW263TgpAm1kG3FMe9QTMbuYN1GTodBuoIGuncQiC
xsndY2CqkSa4p2GNpY5Z1spoaeJTvExo2mTIJBxHdC/CsWZiy21Qgttj86yAcgSm9H9ktjC4trUj
06vP/eM6j9qvDCAx+ThILoURR/2UqrSQA0tgrzkc7BsE0Tux0lSLJ9Ap5nsnhB1WXYMcviD6xglz
zhTZWuOTyjOsaIox8nwoUhGTkPLnMwEaWMRe5K4e4N3mYAedgVJtqO8gJy7p76H+b0RXga4FUCmS
uboFqYa4rKaHWZhRSdc1BBse8isgOB0Iq9c8i6318iCVj8qzNCTySvopBng2dOGt1v2JsUwishKM
3jIPZ6mfV5oKhWePjnc46YObNuoMqxvfvh7aqk6+4tRXN6ct7LD8dFJPCc8vm+/vSTjhhmOymRgL
Xrub3q21vfSLnbbH4UyAQ7h2chuExSv7IIyopgHArsjoBTcvqqAzcdzktaH73pNAuI4etcuVPJ2p
4ytAtL3bdm7vheCmET1aDthhFM38AQqf7R/95tI+RbiJWzpg7ZkSKkFLJSHnRnzUc5kyvRXgQ/0q
mv5sSSgFKPSrJRwBdrgRjWO5dpB6xurJ/uTtA/34nuWCknU3LkqYVeWeovQeBRu6DQnXpJx2EFts
Lk2VBMTqxr6xkeLPBnQE25vj2TNpWAazgEM4mzs/BUu2gfiqzTH0bjB4P4Ezp+22rvetBrGLum4n
j1pm2CRqnbUEfeWFRBi/hFsfcYhb0sJnDvEY01tQTE6M4K0V0Us4/wRqT18Z6CudWaeyiq9PNsGZ
zu1llxo83Tlk0QReQXBb63BWc9R571gFe6sFfumdfTwpQGPlTrjCFAtwLLVB6o3kThK2G44yw3Vz
j5yeSpsKmuyi958CMQt+vNt1wBh9LJdz7vRHcE1pS/dd1KKais1+QcWoyC5Xvl87s9u3LG2WyaKk
7k96IexWyhqjRtz0Jeni1K1sLRmce15N/2hL0tpfKOih641gOhQHj17tgIROtQYBhX0nHmBhNtpg
qat2YoW8G6WJ80Ebl0Ld47zOrIXpJrRfhzekBW4aLJ1ffCIx7usi5t3DwEWl21h81RfnEMXmHi9o
QdczaN12wYecp8Ni/laLG/Muo3v3DWBcdHEp3vQM2yteLoNq3zXzSTnP5A5AHV6HLnLp0WWGMn6V
ROwH922jWQgXERbyaeIlnd1/IvoYaPUiwiwZEkV9hTraSW+IZWMIb53btmx97dwOyKGcdcep14g6
sJyzLT9Pm4dZ0qW2XAXcUHB+7JlDLYWSHFlkt6NPGhR/+7x6kA2EnkQnV4W9zvXFaoNZ7XU0WJmg
X7q/B+CsQceCqlYT4rAv6oVK4zoC4m9NQrHFlBFj8pYJx2O5mFQAEglixx18ONTlWumwDm0BvaIw
ohparpCSI0uHg4TY9PH/DqH5HM9KDWpIY8rBIhEZCE8AtW9nl8pfLkYfo0YA2u+4GTxlY8WSc/IG
9XOMyOtIGmFY89ZeZyadVTCrlUY8IbNx1j+97Z5MZ7ttZCBqUQQcsba59muk7dFms01JOVHQrSNI
J7ploJ0Ma2t35rsXmnE07Yf/dKNufLqtiHmOspVUPY6gH7fTVF8r9pbSdBRwyRtSR1pUAvkbTdnU
Aaj1RZ2fRKaKK1QDr5DZ7Srb82x1zWEBrjFs9uGL/3/2mtXeFTNXCXNGPfexulk3pMeSvsaxkoYG
XQ6XfyQiJlGXLRHVyYv2wfdeZFwxP54EvZwLqS2KECVdx7Q+7cs2nkfdEnZMwMZbu34cMDkaV42m
r3I3xam6VZo4h76SeJwo86lOhAfaKgBFjkyskypzLYx39w4G3L5ykxU6zDsPnsimasNG+mClQZT5
8vbjCklo0nLF+NuevqJf2ReWvjIHBPZ4acT5rNCP+XmUpWR7BktuoocSZATSSFUHe2r88JNJEuyY
508FLKcewyUecykkKiCS0cR/PWKiHQeRPNfxFY0hN4prGhM1m/JdzmH45tqxJwe9iWspsgCQObTJ
a/MmwZNhGJRSU95d0Bqf378kRbca//HLev9e0xXnqobDDbvt5T+6lpRJrCSnucIaQP4HygwM3qb6
Vlfnr3J5GfVgCvntCv7H6P+kRAn0oyPrdsvVWZolegGSRjIdNwf4ENrk7T4yitjBryEUUapUJjdx
sP2bKRAIL5YxN7D0zwKO+L990K0Sd0QOkaXx3/4d3VoSNOuG/393ZVXex8Bs1KFxZEUWiSgjxNoZ
ok5I6+sdhB4/FWbVitgcEZXu4OhFRPoTUIa3rOa4JkfCo3QLAyhcee8UyJKDAdFpFx8NUt7uwCPg
CXssqrQSHEVaSY48QymwQ8KTAqiqI0y89FIb3edOCzeQh381/D3mLKJQ7ktZAqDR6KOhTOZQIuaZ
9nCTf8Ywkwcd3kRcopcEhghh5QeeyK0TgCWOCv4/TLh9i/Y22zViC+r9qj7NJ3COSiswLEdaz5VW
6wJqi7XCYrJMVswUHNgUMO7W2lUb+wB+yUlg8JfzKK3+gYZ5O3ZJ+YHOVVDE1nNeASGKh9hDotWM
8wnxAksUV500YojJX0YtUPExlhjptWyCPjVIl31UBhIRZpcPNiE2mOo0FozRan6e4sr2DTAh7NRj
KBXEY00FeISekxMQvnl/PAl4rsF7Ml31tCF0ttbYxj8VyqJBjBzCUDp7ZYTLTXmzmJPqfqXdt0Zs
nG/jGvV98UghswWXQg6m1ZOUuzorsmu8OhF2iHim8cO30vkeQTTvWjjn9a87xkbsQXxWe0lGgHK2
RyFWbh4crb9oaK83lc6Z+8VJXYsFwqSgE5AHz9tO6UZF9pQb87ZRZ8khz1KmFsFj3tOvs3XsZeXS
NABMEckrwmQa4nFbSQWkDZ3mbit18D4HT5uVUN5EQ3evKJeD6SYHkXeLSrej9scfSMUBz1+a9+8h
5eYIl8cirvq+wwy3Sng7MXJPeJxBCR3OqTPSkCadV7akL3EYIoOCLKIuZp+jlzYf22rD6cdAvVqw
cCnEUGj1aHrFlTp3LkyyHuBk/B8uGuyPhhmVPqrU9caE+dXrx38pPGz3IVjCn1nkCrMOfs2Fg8XA
sMqMuB+LQmQbVjIU/Ny42P0mp48kXjxsO6FUDJ+bd3/WSHzpdfShdFuFRii5y1huDPwLTX3Mz0QD
yrdGVKLnP30mnlyMKaN41HtmXSkjZ0TVpM7AN0zVaK+Rjr2sYFd0eBGzWfPdxGhZ1Ad9K1l1H6d2
BRKczT1/okNcnkCbsbKihYrlf6nUfmctQNl1Fxyr4Sg/s18aGcXsscRj/Q76oZG4tbr+Xroew6CF
f9gqIFNZiIvW5W/lmQaVC2y3xU3QwBvct1Hv0lRUn+vWvsF5ZcTQLyiyC5BIncMx8iGzIbtQfzLc
IrloLSilbX+Uk7Svmzf4qgYvTNAvlhqyKh3hbQ/yijf/+qFUS+wCRzZicxnAlJJEZXVt26VAa4l8
+dXOl22p2m+m1+k4/Z8AQP1RHx37i5onc27pyyNlMFqLU/4xQRGgB/ETJ49QH1V01Mhi/ZlL9EsW
5OoT8ekBRSdgS2q7cjoNZwDr6iazcLtrRQoGUfsjrjvAR2pSUX7++oOTu+/4IsLnRgpoAYLHeab2
70OLFsLzphs2n89Z4aOfPTvSIeN9PoJHqkiKszY4uWwPNp2djX6NZCjxGqJpRGcMLUxN0SNEJFTU
zIDMhUTqxOqetH9Rzx0Q93YEqltcU6xlJ3YidWwFEvHdfXes3K/FGeVKR0loU7eUHbbEs01Zrh5q
1T8uWeaFiEgYwo5x3cCpKtGAFSIo5PbLzm6oE6RPUDzOVv5emiQ7KVYTnreYmiGdkf0B7kUn/k2h
bAcmRZKxX9QmAmICrHruAKhq+anygaHtwZjfwlKD3M2hMU0R+LGY8opl/S0/D5uHNVV6E+9lrXRc
MdspEdp2q0pyL84YcFdzE1uigHK8s6mrSdMMg1uWtxiSilx4FU/75I02fW6RLGmk7ngFHORTlsL1
nKAvXpX3Sh5iC/8zlgp0N2xKvFTleAL/rCPVrKVebgrb/wM1I/lhBkwRMc8AIyMR0J4bYa2ngrAD
WzzQNmJ4MngXpcgFN0dwCa/3kA0stdcfFEwMOrEPQlBgHI30WCuRUAus7AxcygRLfB1q9j9C78hw
H/q2VkzPBMsK7cxlbaFNl4iNijR/ngFgpa2LXJX8IxoeMr++3Odin8EhslSINj1ri4vDtj4Erp9O
pKQib4oDIDXisr27tXi+X70biKz0LkqDQVUeRpMWaVAxfq7wvcBGHbPx83X4WdX1N4jCuVZjo2cT
/3ZLcoA8azwJhKws1IhJ9OhA/JTCGmQScyuwi3ir0EiRtgHwU1Y1pIlGU5fpf72jWGqLPH+aE9O7
ciziHjv5x4tsrN31+fDszvEygXR85sEx04Ve1IHNMBuxClVqCQDHv6FtrmWlHnK/qh46Pf0fqRiV
mRqF+Q1nWQTvR7GtnYRqFauIPiDyQu3wle95aGfpR913B9Bva0/qWm9LrqHjZrR6TMm26jbS4wWx
RVtitDkNPol3RkPHE889xYyXwuKSQwXWuAhHCnYX1iwZqwvci+k2nbZnU6lQEl4Esba9hPm+NKtu
Ek1qCOKfr4Hp6oysyTLppVhYA7vliv2E1JAEsRZcbk3fduS93v7VTaP8bxaGIv5L3lRjJrhelclE
ugO8wja7hOaFJmd84QkQtKpoOo8NEGdzmL8IOou0xZnKNH5UFbafX2S3QK/yLqg23UHlM0QArs3m
+Bzl7NYAaSsf2JXtwxU9Dpm6WyF6ePvMN+DRJfFOlbWB5PPZenfCvQBLpcNksvPJnUvJymkr1uIS
dd6wXHGAswSREXiXdbg6oODTDONfKkMIXuzpbo4LoDfLcvvwjwFW5TIMKEvBPaXx/gx7d0kdCHoM
L1pYYhuLyCeb+xmS3XHkp7hdx382InQblc5q13juOu3wLvPH0/T3YQLiqXYcK5Q+8NHDTClIfYJc
UntZ0FWDb2cIrt58NxlB8qcHzZgDtAgHhvcwwhxOGqBW2eP1L2nC68LCVy3PwdLXD4VLlAIDibAv
MuDPdoRaVg0wJ7OLmEvzXlMnQbPH/k8j4SVNikoxaSMgfhLDtfiFlusTBrSgf7wNlX5W6hyJWalJ
bGNXIMRIQ8lsq4X7YtsgNBW2O3gdVQuBN8wiqx9u6ITI/Y1t63p5OhUedTv6V4wIThbeYSe51ITq
ArHVNbiPrUUW3p0E8RiapTx/snd0OeRdbb0lYrxr6rCBBFh2sJjwnUTbRrW/3XzRJH0nJi0Xo+0M
K4TwCoT1XbWPFDrsfMKaXFgsO+rfoDhXv4IJwuhbWZv4zRhs9WpV1Jn9P+a4Hu0KitJiz+RTBptz
ciao9L1KQ8iHMMXP6xKM1LQqqyE56DmMeWZ78aG+WGfRZGH6kHmOkyegIuO6dwnydaxeyCyxRm+N
Jy9QDROT+xbIkV/QXzGl/cE9epHg8LRm/5tnEynpWIH0vzCd5IBVewscGB0tWdd4E69v2BkhnW0o
0EL6RDydIyqiuWYdYiNMSlvpi3cQP33vWNCmcv1TA92ZhHr73a6d/sPyCJ2FUR2FHRKF4lZMY650
CtuRZnvL6uCeU/28/YRD/Cg+fLv1SBaCLVzp4BcBX+mGGRxcANUQf97zSQCpcHMqh+u6Sr6/PAG2
HOcz4vVkJR305ENnePrnEQJa86w1zJwhtZuwlS5eYFLm7/qO8dq80+Hyu1EvNsxRVyyGakDqVFir
T5n/UmcGtlYaRkayXmma53ViwMzh5xiw8F6wrGWWtsnAfFX+80fJY/jv1Wi8qiG/I3CCU9Bc0gYH
PEyxXY/HJLG8ubuXjmihkIZ7MvQEnsvzq8MlZmTGiShgy8HXthF1GyitOpiHWZYSyI7WAdZQk7x6
0nJJudRopAOyVZXLm/Et2c0/iC236RhTq/nX3AZryFADFyxd05zjE4COgcMxrZGBNwlYR65cYwFO
Rctn49a7luke+yFHI0cGwC9tWw95kHJzHsT/5wmJ3iPUqKYD4dglBFS9jgJywxxD1/8wy+5xEd+L
rygQZgk9HYH/TAnUCu+Ol3UwcFx1lPjNTk7/w53CJaSF6S3+IA7rV0CP7I3nSDm54U52KBWZlzBr
lWL0cXOVM/hb4BqNG7t1lTuBC6wTmm8JAVPMXLs8MH2jI5HrlKSTPW9TIaF64CI2NU/CjlIKWnvw
mBc1Ovt7B5VxyAM+5UCU33C/Gm9Q1s8EPN/J1mNR85SZzCtTRhIKIGp8ZbLIzMbst7j7zgYEA4lc
vrwnE0zUwThWYL/HvXb8Ayn/ByqjO/vWgzoP0u1EmXr/i4aCrL0ZXpdGRed8wCIV1fyulXL5cVMj
esJDUPqouBT2zMUXamxk+k7qH1/8Xqw6ffoWWtRQiXvPpbiIVJHKM0J24UKN4PhNsaaGi6vp0xmG
jaDOpQpOtrdwJa92+nEPU45a/b4KCjcr9gHU+b0uwj4ubQ+Ik6nn0+82h9aFqu+zXjAxOX/TqidM
EU9WAArh9VrJOdra7sHI62lBFIIEQeaJJMaBtP/Ju/P3AVft5jGLRjtc2r8eencxG43RmWbbs0IC
yRjBOhuRKydTZdaqlcY/oFdqjtxdQ7nCg0q1MaVfAQ/9swshckPom+h0fNB9qzGecQdU7ZEI19jO
oyWJtIniNjP0Jw6aEmRUNmAP+66EZeAk/Yf4hxi50lV9CmF9z8nNkZVMdW8yCopULUQ19KJ2+Ek1
x9VvUOX5C2lOmkuU7x0eMtzNiZTbV2pC/82VGK0x3cR4+P2DQmuV0koQING+ff8WiAFaeKqtUEJp
HfYjcpPOQ/6seDIyBQJ2IOL5eE8tdXYTWuEZ5H8hwGHZoxXhBUi5g2thMYO1iiYfhuS+biZ9AFSJ
NSf3KB97A+rXiw/NfWXnKq4P78tQyTytfKc9e1M9HfkiNwQ2Trk4Iq8seqSf61PLbcaa+BCiM0GN
V3pVmjligw9IWYSYq2TiAvt72+RDPg82THnAV0dDLI0qwL4tA5mfL9RtQdOSs5DUtAjm7Z62rVUV
H1a8VOUYB3IysBeO6F0zQKA7lqKmPLjgOq6JfU8234IcuGi4wLzO7ZaU4IpA4Tc9pZBQ0eOfm1oI
OruolyIIwpYXQqnTVcv+Swx7YAnnqZxPiM5pjIT4t5h99Ayiab5tqzDnGzbLdqdmHz4NB5CcVCeq
ItyWBTnrS23kE21M0MLDoV2kQHNnfSkfDun27Sz46ePrgV+CWWiPvhnPB7gnMgHuJC1TPtqCwXXl
v11bHX8oFYxtXrBJDTNbL8J20aphxYubvLParmu7z5Tx6TRtlO3ZLt8tO6qTp3scSgdb4lOlM+9W
Zqs9VxilMab71ppR1OAne4EZI+kUOOWKU7b4ODDK215Bpsn+3YTiQHLzPOzFALqGXAD0W43v688i
ovaYnm3idBLFYaD/duJLkpKmO8B8Q8soJWJG12SIP8BtnVtN0VxBQMVT4VCGVWQZ99DQTjPY539L
A5UBjyc9rlpPXuMVvTAkVJzda5erHSn0Wi73IEbks2pk3rqnCckx4U9QD0/oidAdM/z8APRzrGKC
ZpPKdIjPHjlAUOaFsJMhHzfPXS/j983f0QeaMCjDF54dexAO4qzMXze60k1w2VEuutknBdfvE+0L
HVl1XVHFmfS0Nw5ff1cRzeVEshfWyybSiiZikX//eV4Q/Hu4R3X2FoYG8K43XrUUu76rmduemIXs
3xiqokIlZmmh2zTBKzQ0UsMBVWnab+knvk2WtcUbh6irxgpeqTk8jwoKSzN0OpqkG1Oq3HY6uX6b
CWOf42OElQqZxpLtljmAbn7EopE2pNPF7QqTKBpn47KxrW+i01k1KB5Iu/2s8Wj4U0lPA+7/stRF
zmA0yuluoRbwIXn73pVtJ6hqSr6/w/Z5zCjIwIyxTGw5VkbNy+aF0XhF5FHaebWgY+RUc17uoN0x
KVyznKHRSB/TjuhNHQbrygPzdn00EyzjfceW3xGMWRsRjGCIEQpkYV8+2bYEyupD7XDkJNZ7PyJ9
p8qsEIEc2zfTkKwdU9jeGfIjxukCWB59QxRt64EuopeMqgdvSjFxHrkmhw0WciBx+94dy0/OEZzL
hyBbpKfMFLxayh01W8IZ+T3iiOkYyzBeAYg6P09r+2Bjn5mSYOZWEahthz3npOUUp+mFi7FbSHR5
Ioj6pQxSRVlD80xqMt3/kqXthj8pGfxj4t1Qnxz8+KJ4ORHt6LCdLQrcuemEjTRSBTSXNxMPrj1c
ziS9nPjZ6Zgi22lEQWaVY+UK+rfQ7Gwi67H/K9Vcwf0cd8tseSKlQlAVHPs7tFMj5NJX+1bQ/693
gQmQb6NjZjtq+aLIwfIOsEB9ZNui+cC8m3CIGETSh8LXrgA0pMSdYdxs1qJg3gpInsvAxShTVW4Z
2paJ3/le9OixpdSzE1rArfuX/ZKUdF9Whj6BOLpwssb6JF24a0H2MJW5TK7JztXuptojwLX8wKbr
rq23q7w74UYF/djNZRknGD/d0i9mJM5VM7KYcZuoKYg44qO5tMnMp3MsBxYEnGrVUtza27uE16z9
Ko+yTrfoLt5G7xpbSaWLNmfqp9Gaxn2i0c3kXIzW8GgwVk082Uj7pPoJ1ZcPYK881juOG1OZqmZ6
FqNs9PYq37Q/VwYJuo+gHmdlcoD5ACnGtGseb520BQ/j8vAByyY1HMIT4k3whHjzQWxHLbqwSU8l
bX8wDWXm4qMletQ9up24uifNVfCiZnEhd4R4NS28mpaFnMS9C1JUrZXu9GrTmFsi4mYJxFgdhILh
yfKEku92xlS4vNaz3Xjcwob55Yrt2q+gJwGxGMOYCwphFfcimOh20BlvVlTH0HUuZj19ViDn+Gka
+5uJy8DkfyTBn+CDwtowyCtWb8GeIyMk1EEChT8K9mAFy40ict7rT51MiCbECo5uGzmT+u4Tae0M
p5vlQX3QV0AeNVIiaBp7I+7paGa6KU9HR2o593Q9TKFWdUkV1iAiP9xGDmy7Hwhye3e1ITy4iE+n
55Gj77+Q4l4s2PuKP4/RqNFLc3CkISCKMHbzberGlpYEcovfsjlhxbO07OLdBEC3dko86fRZp0jw
sfN9q4IRug09aRYZ5zg2QCHwN1SfXlu13lOtwTCMoSvRwAsvaWYn6Pl6fZels1NwgVaNeSqzcJM+
whf9HrhZURWXES9F3nL+h71HsheeIgyRhYdUYw1ij0w9Mjc13L91TUACph7ECAEn7rj6OSmhQwp3
sI+j05Ft2m2MMlRWr3wXLqz9kSChIcMD+A3JS5qL5l7pbCIEv4cKsJLPbeDIZfflnfxUWesAAmf5
wKBBaxDeLDA4BkXE0HDpBz+qniQLfZ5GBN81u14fVpFKQZ7Xm/eWllwyLELGrijCKY4CUbLArSfI
kZMVyIBBIuiAy95/c4ThtUzFkSB0dai6TbvhqeIZSExRtAYB2et5IK680CuvoeH7//T/q12IUba8
FAvnv+A+7VuHm6NFuuvGCLHdCefO5D3UEyA3fbahQHGi81nJLN1ccJUuaQzxFf0RdUssCwHECGfu
FGqJkM6GlzR+M/H0Np2dsW99x+MGd+4fqXE0HTuTB+IGToNIwUhpRJzPwsNDF57VSqn3nDsO7T3Z
FM8s7tY58uo2PoIA2aqaGUOEOts+yoh1oNUNR7PzkdLU50Lw3dW37aPVYhbENhd+tjPcqctxyBMG
rujtxmvWWoxCi7d3Wx4jq5sY/06e6tb+9xaxwdIeexsR3ejNn9aOqLfM9hQEDnmDL9ac/0tatzKl
sk6ZawzDeLUEX3d/Wm/E0oMN1oDNOXC2mc0oK5/QaFWniHKUNJ7m//vtYjSTl8jwCrcqidJjJhU2
eRumCUZeVgLs2RXqIovd107sLKn8OoBKOeAB1YsvjKoVzqNpiS0x2VH4cdqBQgKCprDkAwygCyFl
hfgoHElPw5DgB6QozmW9zItGtduxo9UJulJujtYvGqCDHeZOsRm6jLYyorlne2qOvEijOsZQaxS+
lH7A7cy/yiIqZKdOqcD6v85Eofr1uP1hxjj9JirTIo3ft2xQs/2ovqO9iqdYzmjGn1OUxuHPE0Uf
1OpzXedw/i/4/L5KbZeAIWFY0myHPNPkZz6Y8n+cpfxLFuMfg2rL/ToH3T4SUEE+YRkAD9rEceHB
tU+80F3UQdUxyUF9Ah2TyNkVl9b1s+zlOi97OOzYG76jE1GQFbODPQGJXyWWKIhqsD15srbXFlYf
3v8hlTOzxvhB2TJKjaVnzF++9yWieuD+IVQM7NVoZ528pSRMfOvM8gOaR1++A8wtGQyftfo4xifr
i7K38PhLuive/FWfpgiBG5Ptkh6LtyHMRGz6GV1Ox3LVlIE1dfckBde9DbB7odNUIAyiO8UgczmC
ZW0TgGNGEknGqzuVuNbXq28kahmL9z2IjpeXzv0Ir5uQJArWX5eW/ssLQZZRPtiQS6hezpgDABYc
j4sGcZ6ADdmmDtdeZf8cZ+Ig4u4rrOSdWP66tlGs9tUPnBg9DVd6ssTUwXpqz260smwFWYghl+hg
bBXoZUUNtx+SdoNKiVxhgf0nK+rWQ4faC2SfQfLNZeTXMktk2IG8+GujOnIN+EwFEjMFnDI65HVO
z0ZLp5YF2D+ZmDCuovmq8e6Y0LLee/wMFmXIxyAeApvrYcdxTxTKU+fc8Sa+5f/uGa2M+ZaQiI8V
jqTumv8C+rIwc0EqBhCt/Vg0pRgZ9HBdvq6wwIXVgHTS47ORpUfCOtAbda5Sq2eW9aVTUOp0W+9m
AkACdKmh1fUuyIDLVYTvxLUptzF5Q7jPywiLQCiBQzNatFwae+WrLW+BLAZFSnV6HA6BVMjG6d2g
BbfGIUwzWxVbN+CIAkn3F6l6zmOfNH6c0hPX3XZZ2srXcu/NkfERH6ojiUbTEphW2EjoBR77p3vx
QvJmHfClWMbEnF5xe2DXxaZIhjt93Hull8Glg3h2DJw+X878IiwpcXVxvOB0zKVTnleI8NIJD+Ik
z/RG61sI13QyVKyuraftrp/08ft5ndjf6CKlNRtByp5g8yQIJ91mhasrcqZ0ktIzcpX2Wv92G7WJ
LMZF605VN75kYwRBnFCVCgDuOFb0a43NXVDOP9D02B5e1PGk/FidGoWNR1QGSio1IBlIZZew6H81
XGh0iwDzI89iCjpM3qoJBZLufJhzEQZl2fqS0V2O03PdYNb7e2BcNSame2NoW1gbNBa58XGCxq+R
7M43aqh4wRNHrGrQFc37lGD50Gbr5o43dTaUS1R9tvnz+VDFDmkPg9zwaSF+OxyXoB3l2iB5pg98
g3kiH+TdHMXNrMjRu0MBf+exfS179qEiLNl2BqZ+ur8274obTwY+4NKfthWCFd1mWOz4keQ07pLz
Gh9r7LniXTE9UVxETLlpHYZR2MfypHyIffAZccCelsTRdikQ3PfYOxdpYoPHBC6iWooqR4XNs3Tp
rX5LNcD08QMx16bi8aZ+0X1wDbj5/t3P60TFWvkkZYMR/wObgxUwK3fpIgOIeYpsWO1+dsIBbWub
uyI/KOw6xzb1fEb6Kw36E/9J6ihE0VFuEPrgf8ArHLpbWCBJ0mmdY9cB05cRaGM/cuH1uj/zekmE
aSEnKDqYYerFK22WmZho6slRY1li2wgHMvWjg3kZoHuWiXgFS4b+HmK7M1cXoMY7A199J0wERKKb
AoJP7MTlNk/BlolX0+ayMnrzTlPob0ngjO6JDx5T6pLz98PIlqKooqjp3AqHXncc3uNw5tPhoJIG
Qd3cueGqGIjD0FJXoZT0TsGapHg0DcsKmetFKRp0Sh8Wjo8aQgBDWub0FU7JpgkiLk6X28d4V1tu
5snEzyKk9vrBGHfOn6kOOGnfVMoJzQqW5bVfk9PM9F6CjcRukBAae/y7PIpcSGLTLlfPWWfpTsk0
zczjTFN3JQbjtMuFwWCdpg0kAnJB9pqJ4f7NV6Kf+TdeIxtCFFZmy4/KAjp47VBHKWypGZGfgFj+
G1/PCtRNgeU4I7SM4OOSb5Ez5/6xBXdBa48tbsHfU1ogZLhopEs5gf4kf9TMvKXDf4FZzvh1P0yE
UEwzSvP9KlSBsRkKYOmshat6/joGmVXqlMLcxtVBhQN+ntcPJ3+iGEf/pfWC/4zzI51Vy+mgF0dV
j2ZUd9ynB0OyoYQwRc2flwDQQT1z6rT2zBgnlgU70xV9zpFqGytrL7+AsiJWWlq9RvgGOMYT1ln6
ZNDJoN81xkWV4zw6MVeRRnEO3oqg4bynvk8MYfMxtYeubEbz5rKgSz8blrrMmuWfBH5zsZ61o4ym
JmbqUDw86E0XDr/kMj9qJ4XSEZdi5WpdH1uZOghugbewjO29a8nrqTXAqgnGnng24j1K/wk5Xw1E
hH1+nGY/13s+liWIgd6sCNsIWVusCcL7I2LGlbY9HohtsxMjNL6UAEPrLi2xrVvpxEqlf+LXyGLU
8gvhnfZr0OXeOOuq37FoRbgMy+I8mwsRv+XNiX0bJnPfNUkHpokmM6Py1D3JvPQWU/h/oeTDJ0wT
ieNnlMMQfsx2twtrtjGACrb4a5S18jfkfH0EJUFGCGNBwUcCNC/ccp7pCIP8q/ojqYn9jjsMHQ0p
+iTF4F7wHkTse0YTfAK0rm80PAsfKOyvZkCr1SDeY4fR6Upp4oqN+VbFc4PXt/RcspizVMDvIMeG
jgmCwmFbxeUyDU94rNOhPRIVT81m+JXPiUjiFcv91WuvFUzwrZ40KIamUeibNVRJ5L+0Pn1OP64U
HGa3j40uaY3l0lpkUQ+jdS+XISAxqvRaj/5E+Bw4r0wK1S4C1KzOHv10VVHEj2RpkmA4iyYmdnLD
FBLqomp7jXg1teWSkTEk2PXzLuDkYA4ECbhWiFo5920/zsKt5W0XFq8iGRy24IwjzDlATv91HTr3
HffDWveeZTIoTN5rqFS58954U9eu5GP1gc6C7aUOgNCZs8zGQnlnpXe4e2Gs8IoEROtIXm5VgVz8
g6x8wfMN1FUTEWqp5kxoqh/NNNPKq5WEWPAUvQS+GmzHV92Z/D2dXAEofNzQ0uf2IAYjT/p4CIfc
Jx4C0wRdG0A4R8ZWUVMVAtep8VFaoyxsX6XHdWBjzc7PQeRmgecxY6umjUCk3c8YK1BWV7dqhx+D
e2kUhZeTBy7jQtLgVGIzD/IG8SqhrKuMtMgDVi7g4UzENyrk5KtzbDWRvmdCCikOwPy8Id9koDv9
SHOhOf6xTPS52ZWvvOWYE90y3P9CxUs5Fq7wIZCVdsvBrzy2MdFDegQ5yxNdbIxydJRKHOgJeqPD
+ClSUMEjClWFU9xMKby70UauOLHoh0+zpw28FEQamQYCnu/yLvty3VVa4agGZpnZM1RdDjYIMV/P
T8Dg1HZuaWdYFgL/zKIlwuyYjHrRNn+gA48KlqxvzgBvbCWkib7z4bqdOl6X77Qx9nSpeaxw7QzY
EuKoEWT0YQiEQT33WbByMz7Owvw+xqAxatvuPzGeDdbzpJnxNEZuduchHQTnN1vYEvR0AfYDi749
PStYNRn4GpNXFvXbIOIjVsLxZ4GK3idB0IVDQabePhOpFeOiifxdMmznlYPOwiWfSFifhugbWJ/e
OUNTLC30dvaodlm3HyLySpW743e/Awgi7WHS0Z70VAQCGPpl7XgwDEC3F98l3/kCePsalY8Pl/B9
DIHoPiPKMsTY4U46kzClaRW1AdIxaSlmzBTkCDzlaxOJJ0OZqzvFFtA1CkQYMIX7zEQcxmgKaHjq
3MkLnyjWj5fACGJzC25dzxYITCvfWWAg4BEaceqntoREnhuC55ZH/IT1bXqtyj0x7rUWtSdD341K
eyOKF+npm4qLIup7rFgSg6SewTdtwXq+L9ciKSB6NIbDwbluSnTBjID8cnENTlV2exXflgM1KgC5
LDN4KRjEoPWD8B5d6MlaGHKz6PqS5Fm5pVtJyaaLfEm+qzn5mPnjxATes5joe6ZASmbCPH1shyNl
xDaJU4/sNh3Z65ipL0EGH8PWLQGgCtGu5F4P7GdwxoEHIba5lvh14zMxjqz++P9/LV+E+/GcKN//
lN1ZVWtg+8vBLooBC2DKW6yYh5BrK0ndbBOd28IuF1nKh0v1BSRJQbaGbbyVYUvsU/kSze53P+Xb
RHuntnxu4LOL25G8qoj4UMkrx9kC8qUi067kbcphl4vDzZF+qxSjEh7rJUbjU2+BssWjjqeSpHZs
hBSz/R9lvr2L9t3D3+FGX2ThcFFHPmlkPYVjDIkL1g1+JDnp5uEnqvPdlmnx2hTyD9bHuuwtWcis
FergUs8RC65Y2AkfOPR0EbJCcpU2Ru5ifnmXMlPjZA2M6pqxNCVEUjeBzyU9rqobEbsb/7N0HJNo
FVDjYG7ZbDms3lDrngCn/NIaoZensIxLoW141YwKgoO+IqTaFN+ZZAmtw/yO7ZZW7vfsSQVfaBXd
jv01TznhvEqzOcovqH/RlI57GljJKswyb1fVon8XPvZCM5QQBKKoj+ezvYXDhtr7tkY7A1NDp5O7
UZlD5vWVA4QlzYs1twVUkGg+Buxl/FZVItIB9ek7clrVfDTPaCGorfYdPG/p1Xd4RK2TJx8qIIkX
rCjN4K/6l10a3ADIJ6TafG7WGvBbL7gMq1rG2FuuuUdYwBjaaxC6KpSRv0sexdci0nakDIneOn6J
xUZhl3ubBuCK4nrHgmbpGbvnsU4hg8PcI9pK8yG+7NrArNNqBvznQoje3X/jZNiPRDqYj3kRJh/j
dlmyrZYcITSTuYTpLSOrIdBCgWEcwGAqiBhwMoeVjGWIXFVk20I1omleDiGxveC/BR0ZkSwy9DUy
fQhEkZElZmhBrK5pf+d5zKbkhw0zUtt0jPktFtqhSVMEEiD/jYcv29amax9L2Hn49xMYQs/CDQMj
47lFT0eOi1P0Yh59pBCckl8EqdUyHRdnEB9B1ISiJuDePft0L+9GyNFh6AFuyBM+KzMvF/btbwEY
4PGWS0R8HuKdvFabweik+IN9uRWv0wDQnFaNdKIOQuX47h/mxdCnrrCt9fxzDy4I/I8bCxDZKzu4
lBbIlMe/jH0BUGxecdYVxhSxN6lxMOdN0pati1Ff2mAgiGuJID2JD5CX/kPTY0hJPkHfISBr+S5Y
jJFm0FR2k4/usvWH4dTFMCeVc2RHjHJ+Q5Lj3j4D2O9NSt5vjw3eYygiMkNVZmIz0Zd+HLS/q4N3
o05Y3W0xGfDyuAHwqe5RVf4MpCNZW1JJU789TgWHLGhEHiHDYi0bDl5zQaWQYDb31MzTiNW0HaUD
Jw2P1fsihLwlXoSlHiWWJXrvV1JY2DOKnvEFDglweM9q0RwcQcY64C6GY9F36GsGGQzAS/PdCuwY
ZEpYUOrS53LNNE7McVvK+yEYKOTo1s3l0TdZrSOC+M7fLUOQcUFxRFMYzPI+Qy9HKrZZTMozK4Eq
bTCIPgusbjAl4tYOsEAE3CkSQfAZpZ6BcQXFJFc+iE4e7cu/0CFkMVteOzmSdQ+57ttx5tsRfUv9
0I5+lT6W8Bqu3QF+gxlLtr5Eth2vF2Ij+DgYU3b1NtwvrrBS0nHedR/Q3ASB4g44FAHyRH4lz8G4
9xKAiUDRjZ+QlIZBw5cctNRuZnID/JgwEj3QFbSz8NYlCVUMXep/rEM1jyMqA2SOkQnHgFfPzwhe
/7Wo/xGKBZs2wVOKSTCc5jFOA61UtWLhKiHtpNYuZKuWO3yDTuQGSnLiFOE5/pWUSmqYXVjwvZnw
KDOTe7iB+GQ8HIJ9e0OUyLD77ko8L/QOhJ4dtZQUzp+aSWebDQbk3ZbVF83NyB7Yr4CexGTlDtKB
qJbiv8fMLLMlqywq2QJOWx+pisAUZjIp9y33LxiWisRR1kLX4WCovljZnpOAEgflZDC0znrvWPzB
P9yVguDw3ADPNAHaA2HnFbQVG5YTL8p74hDlm7WMrbWkW62mKWP86miouGz4JKxwBDrIqg734jfl
c9bLfT9FVHFHuK588Fhe814DVyOhWKBXV5ZNHRwjyH/KNbpfE7rGzKVkoK/wcOVnwLvomzNC7t3S
E7gc1TljxjD9oZCZ5EsNMCxmP/7fNVvHcOxuetYXews6yaMgI+QhcP39yP3jcXoFBssf7aNseQ24
JHr4MVYY9NFAmG3xyI3Ul7VvlvOetv5IDzHSDFGrBIMyIB5m91Qr6/b6zWZ+WhXI7afeB4SJPda6
kOccV35Z0K4QPYUwgICRgk/ue7PwLAK458zXHPza6FhyWAgPje24E/WnKClE1CPMUs14OrUE9Q6/
u0SjwDwFXVNoPV/1rQu5GC8Ht0dbYQUHz5GVTJ5O9wBOpYYWyQ5fAD4xbHDvwH9qwwuOgXFV+R2v
yztB6vaus0FJ5QHfFn9//Qfc5cjkziNU+AHRJI5LWATEJgVz2vIVfpOvM3d0FnE4TcPDeLCujn+I
4LypBtcqFLGpeRvVduFARnDAXgwYZ4AvxCndjN34Xoh/pnf4+ZHxel1aObW8NyJ6F+Hov0vosG+Q
EUfpRQ2/Qcn40P/JnFlOjg4nb4HwQ/tfRboI5zW8cRsQDzOvmuHrqV7ZU9ELOWLE2Mj8J+3rIk73
YsqsMy6RUplHb1W6pYwVYdadNVNSNaMrpGCaxbo15xW9sjtHZRtJsATOBSIcXYrMkLYoBxVDAV9N
QM+MV5vqKK2/ZObDPH6uB8oieqLS1FqLzvIHsCWt8iBV32/LkzwsC53K2xXIss8X8wkkIymb5j+j
bz/RzRhxYaOSVW7rADHko31tehalcoZcpNEjc/BcU7E0Gup2zQp+SVc+NMfrBt0H9xPY77QOY7iS
ye0iWLp/WFChg37yV3Ex5WAsBjuhklurKlPiDi7odcgaTAcO33STDeZsIkQWBiZkRC8stgV1Xjmf
CoWFOzOH2wigA7os027ALpSWyzIxKZQ/SVxvvoIk09/ElLFsq69+7a3sRPhGTwrKH6Mf+XSLAiXU
1AZjZ2LTW996UL2RrzQFCnxVFJoWpNgiCRKnNOW+/ASH50tu2MSeOjlVM1pNqR2RzXEcVKEG7i03
/iuMoNrO4r3TxaM2Stxr3RJO7zSHU/YgC1LKdH9e0/BQcqvJTp6Y8qxDmVx0LL6m/TTnlGaEgV41
jpT4ZPNoMvXC60+pBmztLmxOhMkfUhDLEhVcZGf5sv4kHz+qkhh6shyr5rPWbn9ZIzeI+oDRDWZM
v3x2ZVvfKRjgJYpDCc+lAXibwHj48E7mKUkTcLOKzhw/TIeGrMFZ8PabgJZoMphMqYivfT94Czj2
XyMPRcXJrnEf+CavGn7rKYBau6PA6HTLwodyoSLDjbguZLoq7LbMBbHrXljJ8LgLnyjaSqE7kMnj
Wn3LEI2vB/GAM7obsOoOYjycCf6wWwMcNJ+Rm9FaZvbhd9epCDU0tn3CLTIMdSSN+XUBdsf9aBsS
q1E/sYxDAaWZV6LwBADxdCdtzto/bq2QWLd4hvXrwCZH0ZUKOutTzAgakczoFo1W1qHNGZLCT0QY
iFkSbU+Twedt7kHDQwgjUSLyGJjqSLkb6OR5Mwkk/pdAbvQ7mvL/H3wmF4hsmBXbZ1uyR+SbdZlp
+WxTxMT4h4Qd6+iOgkOLBAicop3UPMsEYIooaBPD3g3dlxNEFc8znPVIZ74ohQ7Y7zF8oY0uk2MM
o9RMnYzpnCDBfY+u7RdA/u8ufRWYmdD6kERzbn9HHMqgk+V4vbfB3TbEI6J4opntdrQWuJGfkcid
rSv8QsaWViZvVNCVe9n9VBQ0TIh4/Odrj0IcM6lCs7ljkLrQ/CKe2aKeQePVpjwjJYm8g36Lcqc1
fdhunqK3J9BJu/FRag1oXvVMtf2VzmRhDuIEWY9YuVDyp3fy/aQNdi7QBGkX+BAP23Aj7uNAzMWh
gjhboiw5wnHj59DBzv9+nf96ea99d+gxK5S4eHolhqLtrdkG9x/z+bTja+Gqo864z3W3GRAr569Z
5Igw6Qf9MwM/kifHKkYvymfASqLtVADDTb+V8GuiuV59MtGMpeISphKYofBmrSDqLLZ8ISaXfVHT
Q2Z3ZcUGTViPwEs2pYO1ct1ISUytjQ1jXPBOpdzwBuS8+ZKipWkIBsXGqmZ0jjJ/5LtbJOOWlV56
7FBwtx5g3ZWWEn6wT7ZGKnoCakdT7QamRcOV8L0Dt7rxgO+N9vxxvVJIB8MLw/oGu98scWneCPn0
7uLZkWRa5CSoz9bCIrEYkqloTM2qVEniU44d05bFKZTvXetT7bEGNJyGH2eudDsmB1sZMSg+/di9
G18CG95O1fLyVQtzoBRRES+GbDfaQRAUDr+NFrqMmzgHjCtimp0OuktKkPYvOa9PruNEcP6ajeQk
GFDWslYYBRn/GTvaPZwPgsJtLk1V5fNUOVJ2Az8F42zWauV/+mZ6E3NVwbZKfaIP5LvVLSmqmR7d
tumRrTVlGlzaMc6hOTzrWwZUhj9cY9bz6Hrtpc6+RHEjKnDvQWO5MT1x53oELYDNUmKKtmOeionG
PGBvZ00V85+sFlbPesV3+OO+BGw13jbRONdQECxqbBD4e8D+XsRuHK28Md2VGywF+QMe/Wk6sHzc
QrYR8Xleb8hDH8KlZbGSqdHdJjfk7+1LE7WuQb6C+yLhaveDgwWDiUr6aeCuDFqWuJnmYVN/05/x
CGCxpfRsd1Wj8+A7Z+N6RYgzYdVmMGQNg3dR019EE3JtZzVuVwftVbTiVF/auGANDE5AtNQqHFJl
D8uInw9d+iIHDE6esMPGhJw5Nemz45UP6Z+xhuQuT8zTEh6ViqrQvLvYRWDXRTwFESp1R/26p7wm
/tnaXKacTa8DT50aQfRsjEW9ft+2ZIJ6n0EHHmN3Le2AbDDZHoml7oLxRHHEnfPIH7eRZJ81DwLN
DKekI9pK27mSO04gdmnPNdq5SExbWfxxVIacxLaD1Qrmy8sl7Sx9WgD3BD7txuYNp+eqDYU1inw1
NfvwHcVJTfH9Ypd694a9XlRHAspbqGZzqTQfwRQdTOu5Y/GRTuIodps53KAcEheHWjxoiEt82X0O
Nazd+0wk+ujyYVHt1EuRZbQDHYgrmxfFMBYRb2BjSRAcTp4rdnKZxEHLhgBfVNhXz7/bbqnEhFTM
+l9btzBsvgUs1fE4415DCFjJ/iuQ0L1mZ64WNLTIUDFtF5Cp73STVOPjaIyJVMZm4uZbXZlcRdA2
bjtaJyXSzxwt+s7cov52Wl5REtj/021e5XvNpgq9Zl8zdFkBb157s08kpJuJBaIXFflMjQ1d2nVj
VWuC0OJ41IDne7RliuxCWlzcM3vlEQM8BNEO+UuMDa7Ss0TCPM0PTKL4kIv5kNEurgRUbpDLT2iA
k2ZcyZRzy/gkwjnWbnyWHVT2y8qIREyFjT1TSyyHqX7IH8BKtE5G/Tw8y5GUKXibzC9g1goj61OB
pkZC6+5wecMMZMZYAM7+RD61lEoKHrCreRN+sB/c29dnfcE5WxC4Q7FN37beQlZ+5ov2T743x6h6
gVYxGl8fT4FHJTClWIhmGt4BeLOR73lIyQwC6PRAxoiT8IovA73kVoFVinZUZeRUs6gfdGD0D2i7
PWOc71SavvlzEJXgR67+13md1amA/PMMmW0kVnfKsUMNgtX92vMjBKW40ACxvXGFlB+hw2EEj9mF
d562upDUbUGng/PqhMql6dTNw50d5gL93GE8IG6j77JjagkvyFiDwfFDqwx/7j0FNqjgDiWuJ7SQ
We24BQWuKyITy1hJbEgLEWoAVBQ5BknW+UKs0AXJH72debqJORdCkv75HQRh35lIvdEgQdREzDbm
OcIrIaOIVDxT8qFxpNo0HzngukAjRu6YYgHKqdTbJwM1Kh6cGcd6m9Xt+DzAzgn80fjjXOoMWpB5
LdtpucVEymFG/S/1WPr6y2jlplBt3LSDulYpnmpYI3kLeFNKtYOmuVSqYrtVBnEU6om/udw5QOvh
pcru4iNgsnJTIlrSiwPbH30rQJjmDdXqU/qmNPl2SVDNQ4OJT0FzJzzz/ODmVUAqDbb64NZ720Qs
flRj7lkcirtMRH35LmgjnDA4ONuqSLQOAE9SXtqnJdzEniL0+8Jn7tfiVPGIc/KB9gASxOtxffLu
XrjMb/5k5Rz5zpXyOS4lcDUFhY29uAB7YtJDZjMFvCCLIJ+O7dXND+IaFTk7Yy88wDHT3oP4OvEA
lt1NaX6s+Apj4Z5rbGe1xocSfr01mXFfMgW1ZZJ7wA5n8MYZIJU4MS6TseGnK5sYE/ltY7Q1iHCD
+b2dmTOZEj1+mTz7Qh75hX1/3CllBduPXFG8nOmdmyaRr/MDAQDsJGQlSNv/+qbg+ejTq2ZFF9F3
PoRljpbbYnRCc5UnhAPbNxYDeWg122nOseArwRmzFZQbG1AZWUZJLTf0NJnztK7r5f5tEtrhuTK0
/cb5giz+uXUl5Gd3ZNhdvdJdFG0QLESG01VajUKK+4Hwm4Ghgw2X03CacfcKc5+b7wCbYnh6S9ab
x/0yjk4M02Pefx5reUJmGCcgSzdV+TugcHuz2Dgg35eafDyMLQrHNnogaeKMFs9usTx+qIMFUg/B
hSlg8IooTX4s5CNA1xED4GuSP2RshMqpBaplWSG1WwZaFYaQuoGepB6R/2BAU1uGfyvHxFVmuy8d
pyvBjy04mEmDzwtR+LI0M8fknU1cvEGcGb9pp23ZhyZvru0V9mp2ZZytzV8dvUuzG3SHRn/l0l+U
8xpGbGmo6xeAXa45FM34xAbV7spzyFJE0j96O8yhSipGmzEOxjX6M1O5LSn+ADnL5HXd5DNvfnZK
EQjzeeLwlQ2MuU62hoxlR0aUDcrIYRIOcIiVwFPfHLIYpl1tA0bnjAi/knAqXmDVCOYtth9Ombs5
gF6TRTiQF34afFFG6BjE2G6AHk9d1VyhZ3S5idPUbvc84N2QsTKTr74rVomRVfmgPiIsnYLkqPMV
ENwJahfLwXMQG0EZK5BRo7zEvmo6QtzENeMEYbxydUo1gi5pnhBwjkshs7/ovw/dzTMlgLOE70Ct
5DMHFEfqvmtFu62+fm+Di3oayCyDQmxx0N3XwOBR0QAlfERYZFVvrhtTmDTD6GuwUZlkIYA2jgjK
+Vg1Zo0ON1k/fB7Mwbx/AQWlA3yjO5V1OH+GQh8YNOkm8+Hz1lyBWn9XoloYY1phZ2OSGDOQTowB
p20yF3u/AMDV5q/4+iBS8KU6aqYrr4b5Iz1aKgI+Ui0TTIFxXh+jXjboEnWJ9nQh8KYmpp4u7MRp
maI8RLetOhmHO8DqV3Np/JDxqqFsyYT/aSHI2pZNdCRQULQ5Yho8XZ7Quxlp0Jd6On2rqQ06BwqZ
jg0VbH/U8hCdooAS2+gK3UUo82PzQDxAw06opMZXfDhJRx6QVX8rcnIW94aMUs+eNmJk3NUqu1Ah
htv74OP84c4Wsci2rFOvlvouP7QtzFYMm0Q9J4FIXDmCwTg4fltnC1aOe0DE5wkG82osXimv7zwL
tamdJamn24sK4/+pog5PaOOsGSUYDPnuDncwSqMgINNccX2+Ilq+vhOOYhRG3S59fmUOZVTTVSGv
aC+jCNfaBYuIZiOJcVLumDB785DSCLps3swEcHsi/8YD/8RMjL06sq7D1deNYfYaYUsQ6IvoSy0P
I4xJrmPRsbpMOYcXZeWHeRrfIGKtvnyfsV8eE64jov3cwaRC6nO+paHNnN3anzmU261P8WC5y68A
NTM82cn2fisMPwgwwl/ywuvtE/v4mo5upjoXhm+5KbKEnU1SaMSoIfuIaGgZoGc6bFrR/DKOnEel
fqiaNaN+U0aMr8PAAIolQc443oGgvfQp8hnGY3KJKBN3BNPnBSIuwWoL3+P8zr6L7ZKBsdiGVnl3
gqqvUbnHmNPctzuwlq/cgXQ8mgt2UA76UDzM2kmtlc9Io1UkfVn8W4Sn3Zo9N2FEdWGW2iBP3hER
EQ/JJVztV4VWxCtJVH+pg+DiasnGMB5Jc89sh9frU08DgpW7T3AoBHTL9WAkE4Q6DNpdN1XtwebC
vdHfTuAna/4aJjOkHE3XJHtvUKkkOJLaxqBXhRhyrNP37742lnV5gJQbmBqUZw3U2AIwcvV6GMGS
ejf/S/VjKYUBx9bq/jwxwtZcv359xWiXgLfa1b2Zg1kqpY8W6j40PlBIQ3mfVxLeROfy7oQMI7vq
9csHepQikabGOD2/lXgOxO2LWvYr7+qwAJRNsdKAhiF5nVqiMj67KRSH7KCvSTZ+rZDgWVEAy72+
Oei57mw5JVRTnEhs9+vbgD8fM0UqAW+vC1Z4QO3ieOg7Jkn5/vI42IUGnid6UvYVxYKHSBAEaaSB
QDU8hCcD+5HqY2T9Rwt/fxirIebjsOZ9rIoP9LKc624oyswzQglNCkeOrkrxH0Ikr1qjdYkXe2fX
GYgOl9rhReBYRjcDZdtd/zg3hlLmQPDUFTUNM/rksm1jlKTRgImUulTFW2PMB9APNPkfdmmeAAqV
O3P1RngmSpmwAZKKbL3LNwlG1dWZvnCDSqCBdgBvkxvIMNSg0/9WLg1qNoSQkRF3mrmtBA6OIO8D
MuvaCFcL21o4eTJl8dR8P9NGabYA+jgbcfAGWebNC0MpM8c5KpfVhB7tQgbNOEFLDGsf2N5XbPdJ
Fc5nKVrjaHr69dtYFw5UT57I7CvBdIaAvBHMh8zpf6Vwf//uWobTRUCv5rU4zrmPmK9Xjf0Mgc/O
0w85839d0orBWLKCE217UAkAkOFWg+bkZ7FpMQJ6VYrz3JlOD2YwK+ZJKKT4W1JMetM9Wz7jjt78
kMtZ3PxBBdPZD7tNU8zE34A0aJRAZClHJK6/x4POyg2CGQGDNjT8iVuUErzJ5DNpOumyYdK+1MlZ
Ca32o1sYW8gXYAO5IvIeSU+wQo8duQVjaiFrm/JaG2UIjiJ3PXp2CnutN2t5Aind+2Udd7bfEhb6
FKHavJSFFPJpkdcRaJeQKvNxbQAtkDZhaYCduNlSPrYSuZ34dWWC3kV8oYiO7qz6b0oxJtmCAVyf
MOu5dNOnXysb7cLtLy5Hq1rPRjTgUAJSubrBwnomgNY0dlTo1uqLLgxDrbmSuBVr4Xr+buzgNoZu
NIIumx8jOz+xvXJMjgnq5Zh3xxY8fS6/0En9/Oot7Vzoc2hR1x4hAJZ304lMic5TT/emernEKIQg
8hdcrf1MNeDKo/EvBcVJOcJwrkXYpZm5cYGfwzTuRfayHI6T/7rNq7SdGaFVD1iF/RGMKBeDNNwi
WXL3zR66tVrbaJdwp1DDPZJTxb4mBs5s40RyjCvp0Yul/MZrvMAt0QJFWFQ8/aNQySAUm0aSo6kp
mGdY4CpdlMZ8rUI3PDeaIBE0aoO2a2fHxCnrdenAv+n/oOTjmSxKswRI5hESdpVA632I+7yyek7z
vMVUIgScWEp4h52qOaYUHu+aAxk9I9YxOMDvJHYiVfFZ8a6+4VtJz2MCNYLQdyDZrqJbJO0XUk09
9bwqTYGBaMX57MbUERkU5gVmi9vxcvPg8jdaJwsg7glrQgbE0YgPBssGb0ChZSe/J74qPgJIEr9P
vg2g+6wnvbp27BPXhsVi645PV7FQW4mB17+pqJqkMtZ+8c/IJdBI2WM0hF2al7hq1LDnxW7mb562
tI1WS3i/RstdE5dmg1+6Sw6EPuPipoAQ3TqFLO3ewCyTfIEkAAsFJoUrKnFEXDRHK4wEhCUR2jjX
CK3apk9lsT/pthTQf4SyFCI8jldicqnJzeNkRYEk/Ck9ltHEJy6E17TSqxa85140IZgBEb6fstpH
dOs08MZ5qBl1101F+qRGVzrLw39NOpZcUmes9K8WsnTK24JM1U7lVUNzumHYg4cf27oYGHCRjkOq
kFyuHuEItmqFUof03ZKFVXM+hZ7kPgyuG1cQU7YYB6aNdZ0I3V4BoOIjnlJfUDow8UESJOtgCu5k
5Wi2p4pSAQA34WYL/4qZkzsUgtHV3O5XGCMlKuwoFYZBCZkG1ZQqdOi5MMRIptUWCqXIqGnxddy3
WDa0W6wg4sg9Hl2MT10aiHas1/Wa4xeuaEyo/zG+VR4eaAnEhrmppAn0CZ/zNI+OGs3ee62NNChM
rNZmCry5QQSTJ1jd+dAEH4EGfHWFvT9oufry5Raryb3kk362vVcUyAyTo/fTjGRhPu/JCWcCOlZm
8VTJ5bGqmYpnsInAJv8jUfmsWFEUXF34qYbrQeql2nyFs/KbDjLYvCG4X2vyMl0irJopFbdDQCPn
8y5ikhseiD2DlnaK9gHMgantIiUI5ZPU0R+5llb+eEWkFbtldmk+5YWHSOOS38si0DXgSVtHmVow
H3eR1k9/lzos4kTkv4AVDXddLQp7q1PZKgAMpb1f9KXgYAIAOMM/IL0m133+oVV3QvzzRvaUiGNP
zokuSkNFX9a6Lqb8rcZaktxXa2s+UCfUJnn9iRmcdl8lbHcXQZ3B8+PG6fZfcWB8Fen+ycLItP1D
XxsMwqsl60DIwKYKHlAWukuonEDUkDKaLuFAbUmKQoElyhHxpSXCSv5evPza2aLq6N3CSr+/z5pe
yQH9DV79r7T6opyWqvi31r/3guLU7whZxhUa+vYEkhY/GcH2ovbXoFPvduTZfkLVcSx6ozv/OIDy
DGZztJqe7eDXJ1TkdXa86sAnJ+o4kP/CK3XJH7KLi2GFudP3q80jqKfGo2B+8d8M4U6sSssz2ILL
YItSBMRJytRzLLwnYA8nremoj9qdGQDSPxPdIMRNTf8mzM+4PJD8VeY1upsbp/PDVaa+lrRZA2Xk
1dZ5yC/t/DJX4Rcs41P5+NbZ8ZD1fggHtt9uhsL/uiWxs58LToGvXbl9peJik4FkWQZAHfk26HYW
K47mJIzMUamd8JZosorcS+d7NRbYfrZT5yDxbccayLoCT6482LGNqPsH1OPu9EjqtMC39es8YUCA
uOyCn+rh5M/a410XEHnMKETjCV8BXJlH8GfgkXZ4By3FcX+py0aDR8ZSw6UMCL3Iq2Qu3PiS+Lwn
ixotxhCwtZaYeafjcIDdKyAZNqZZgOXXb50YzvpoweyLsLmRMT8BZMPRxJbLIZhGMM/IUZgwvqbq
AcRccqAWzPRb9NgfdojkZAsAvD6ARFqEugjQj0rzUrbIqIRvb6VOROwCSh2XylfTpG9BI5YvgMZI
KPdqLkjq8pKQzst+hKUW1FsWlEV1rwSQa9H//4EqUXazQM774G6JY4sO9kZFdu/QGvd2DEeCU1/t
InwiyrVEtZad2L+uGlTjlTAc5ROS9r5tKXvLxn8TRMbfGt0zScjZxvptyzFEg+zbqMfKT0G0BEvI
IdwjT7qi0TOJHeJ5U2jN626RX7NhvvHvwXlGnZEJeql2U7q2nrgHm8w9WkZiTjjC5GvbRp4kYbcT
hDlI+W/tqWAkw6LNzDOkcz5nInol7S7ECsdbvqQTJJ8nZuMbQwG3vE8MyxMQy2OdnUfdsinkMgHC
rHYghsfXxyKdxdP4uQ9QJeU46eu+gQOD4TL+wJvFVLn5Mip2paXXJ5lvPO7NRzK5guRlfw4PTr2r
BHdu55VgobU5MauP01gYjaayvuOvwCeUJsxrkKv/kvJ7vvFsX72vLVmbBYuE5YmEL+o0kTGGeT14
TgbLiGYi15IrNXFtjAKWTgDoP9GLPxLBt+3pXqvexhnGGh7x1DYkTows+KaojV3aEaRWDkx/qN81
KJYUyNCxyWSalG9NoPDf5l/xqkXca4bQPWx030C7utCjOIV/4c0LfxbfZrNv6QCjyBZpCi9wNNq4
AhZVmqAa09+reez6jxoZggGwkpQOqCg26hpUxR3IXJVOj8RicJHS1jKf1UHjEs5m/ndW1G9R+esi
gWFSZ4oD03daV83fqR004VA+V4NH34UHyAdBQCgeXMrFooJuRMYGN0S/srYEl02besgX7bn4aZOZ
Wd1za2LrDY65ggJZwXKAlaKiNmOFOEVwdp2ojQ8w0ggVPNHohDgPzz/bZ7zq335u0cIbWc+lP8fK
PK6Vay/6ilOkqNnhE6QPeL1mL6IM3jEe+6dsFCwUG0teRUTumRd9mBV2eo+nn8r6TybOh7qFQs2t
xGQiHwKXvi30CDtaIal61TifDKvDbzg4/R8sSkq/wBYiAXnXjNmRaTXgeR6/ubJWK33oYL3VT8Hm
Qw1r2tPlHLS6ZPoeKZICPNlmo10A8C9AoXj7DP7Dz+dreUcBWlN64Hoc2ObxhRDvB8E29zAzFYNH
tOMO4Q5MbErpJCb5HHwyu5O2lnyixkJQ2CQdRt/EhmVUGqACC0iPk1tPVNTuhxfTurHZD1OUrqd+
YgfEbR62KPqN3bSqwUT9zOsD3kM2knt2AtMreZIEGVzb7GDpXHUv5rxQAsh3GX7LrbhQiP8Du4nx
QPDf8sWFnBEaAQ4zBrRWTQCk6M+zeR2Ffsp6VZeFOfILJTqrnA8joYcuCBfRl74W0VV61TIRSfwc
oSyK08yTckmHrIf47Bi/6OBrQBMjOD4/Itc3W7nHMw/G/6oMwGHKluukj9PFgl9OUI50KoNxEowv
AfS7UvxEx0deRpZw5Ncx0DE3+qa9PwnM8EPK7/OFe3RcSrQAtNE+2x9RpLZH6H4DP9fexiyihngD
rTQYYzY3NuYXcLcTPKFAuiLq44R0RDXTr2sBQjzJ/fbPpmmTEKOXIZDqUsfFydYh9o2Yh3EOVeJb
8kzgh7R5oA1UeswwGqSMoqVc/ALRb5FNcM8MdroFo2XAemWnZBFHKqdLjKRwJKsnN2gIxhiaYG+u
a9cog0kMhJpZfnYJREOGaViMvusGNuUgPdgQ1L8nimrxcNDE+CBNPgWhcaPuK7quSZMEswk/h/GC
kPEQJ2Tz/AUINXOHmaJjZrTzvEXI5xrznFWotU1yACRoygR44X13r/5+0Qb6drn93ODCFUZBBhCR
T9UkOUcxOuyI7nQH2oULVmKtNAxyd/uRnV6XAamwANyRQ4Oepes3plUFj9SJP2c6RaYDTncWDEfO
j7kQKE109x5eTUdiSXxaLZXxSvqgD2dlfI/df0sMsDjxHJ5wI2SGfdnK9T8z3EE1DokpRIiEF4V6
2/HR7/CzgccW5joL3XXP+2pPlNUoik8I8DTP2GtEpuS39whdNZakpu+3SiU+IIF01+u9Q2S088e5
k9JrlOlmuDJXj94etUjizVQ4WRyyt/rQO+0REEvcqc6gKMf5CqtK5niM6C5LbFNfjS55x8VV+BbV
7g0MoH+vtV0+3kQSuMZHTn6ju3M29UqoN3xHTJddM9ZzEoQQw5MFApUJHli/3bvn3U110weQEvJ0
L7r9yANPxgXQI5vOURr+MwflBmukb13fxhJkf8ZdX0ABlmxJwiqufwkjwfUrHBtHskQGAJ6qcuGi
Ot7wLGoODggEBPxlNNGsUUash5LAm+2F3dkotkdurMkblDebYSaUlyf86OopuyueEbJZEGiaZDCd
/2cLz28+P6THGSLaUqZGpKqNaGVNSLoqwNgL01ei7EnWnIk3i44cJ8KJFAOWjS3oizRVqyhdxB49
SaVk/NLFTLVXrHfbHnlBNv46QgnQU/vHmOsWDTUPNaCnBQbGhYSA8zGsYyonsXLZM1lcmpqHpD3S
CGaAaX9L2S2tYTT9Sn//yOXA0zlcyGPYerlWWkOwi7xs9dh4Wxpu0kjCvqfh6e+xmvy1oisb5I9g
DKgbE2tZPbKGqhglwz52RZaU9ouqKc78x6+5J96L+dlM2i10cfhFzams262U3SXGikzMz22Acm9L
8MBSVoBJtbcPw0s5d9V7tgmGcyg46UGXqqGaAmaUzYAJ5ydaW9ImQRFpgQHX0DzJg6ejBJ1VMCai
06Z1pqiJeznE/w1zzSsDpry2wC1umB4pZjLAFSIzJrgBzjXmEy2O1QAyQIqOTb6EKRtZi1MXHCeb
3oOMM1pvnbutZb8jIHM6Ts7jVI21JAQENj09xYWUzPLyLT+idDmFkkRPgQJivmqT63su6Hlii9Sx
VSykJxfxAsGOSE8leSlTAZKFCB36HV2++jBeArR5o+dy8+Wwy6BiWPsAMyor0t2p06nyOzb/u+Lx
4Hl9iJYCfmpbjWCv9OkaR0AJ7CPTreqYXBVp+Y7q85skwkvlKRRcMa1dHDcWYq7HPU7IJ9D5VpPM
HHmR2VU5lGCq9IG503w39tfiBpBVlzWX+cPo3mHKPv4nh1IbSmjmlp0LFXf72CIt0Vt4V5iIiCZZ
oq7wV9ScrtNudIX4X5hO3PhwW8+DzXu7POu33293nIWxHXnrHABTncEI9NPQiQDpYAG5sU2IamDx
a4bvVdd9QebY1R1fCBiGig1MZ0LGKvXN2DSAvtpEA6M4F67c9Fp/ebyf1VktSVRtkGoyfUKo8Yju
f7ewmTzO1iAcd7scTabByrX/7Hzd9IlAydwv7dhlyOKTIGCn1SKl6yWplOQ+oiXbxBfjnLcTe4Fu
Hzmo8qtI4fWVb4ovu8mUfmmkVkfDAe3aqy38ah4vvttm8Cb9lBk1mTZAF768vr6jc9R+XxM2FnAd
/2OBrzb3/emoRYOcsLNrXYSmE8gmpJXRKXz4b2NbDDXBKprUgbHw5H/5il35SxVjFOfbPmXzFJHx
97dGcjdfQwZjo75EJfpCGWl6TjXBsb+TBwld6qobyRh5rA5WjaIz579LE3Snoj3zsqvBmcnw0nHJ
SWKcwEussu+f4AOT5UXS/3O1goJ0pCkd/CtWNtf7/MSodfO+NIdU7N2pl26Sn3ErBiR33F+d64nD
/+9+gAPECp5AwK+YvyLS2Wy4HALDVBU+Y9M6PEOJsMFQK1vqUdazqRKhB0V+UTSlLgCKMHTSdwag
XMAnRZkitCv4d6magm3BepE4zRT96isW/gVrpU+50e9LzjOiGtM1dX6IJTMlRP8zBHNsJQ777ym4
UyaY0mrow6MLMGG53Zxmfs9rcB8eGblGkTK2LjZiUURE7rtibdRKQ++iSZu89A3ynGpLMTkvrzxu
9XuBJB29BeN7F78aV2ziwrCrkG3g3X1UmeDElzPtkhhXX6VIhF3V8/InJgDWB2ADe7vLzEoZuQj6
0IkiSZVV23RQ3XQHfVWSsPBYrMNTY/2BT+11bgVK3wyNwHZ88H4GA3uBy13J9xWJ4nUoLyCnb342
weNIcWiXiEerL+lW38Rt/0BhL8lB7sHZaKNzRFg5gcSsAJJEZX8LUpcyixuWIOb2VxC0LA5e2yqm
sg643HD1gf2aKGnmDx1l20Cutez7kfP2O/msyNzYZOiOqJfLE/t9G6TLPivbdhaliuRIRY9dITIU
94GP8p9MMdEN6OFVh3WX3j+HOkZJf3k55GyYljTTFJcXcLrvmsdRJoGNUE2XPm6xqPSot9OyW/6q
g+dEDwsbPczmWps4ZvNnulEwQ9g4FiNDVOalbv69cpCmi1VJ9S7DuBiVzaXmCtqvnst+d6WAw/sf
wy8+gdHP3RLGOg5cLuSeA84LpvAv0Zm8hG8GzJesq/CkPQfQhx4LnJcmQYu/n2XiNotqTzF+51CP
aqAX6NpcEK6teB+EGtZYKwNSI7AaJXuak7Zo/M2LiTYh8NhZoyCN2Wn2dRJbLWIzIra1UFPtIOyg
7wWwdPKLKSrNHI85ZdeL/uTq9U4gqPp3GQ9YXsReKV2ZuBFjZT9DFIMUlmozMia5a2fP3d+edO3w
mUbVsMyChCI1FtUsw4AP5qDinuQnDeLasDZUJei41Do3doWy0sNIIb6GsKF3bxRSnkDXbnAc6Dby
bVp1gxUJGaRNvWVs5B00LHXdAjFrvUP8GSbOqecLfVFuq5N3yTeWtkou620QKAUkD2G6CynA54GL
Y4wzww9OCFg1qbcKDewi45Whh9a35NLAKEYRVFFzudQ00JpXa+n0wvuKQSSbdRmKIkPHiBLM14rY
JgOHbMikXKKwYNkm0jyYit6/N/pgBWLT6E7aEPeuBZ3T0sSdOv9P1xZ8BNfeUs1i42SFdrTA0AG4
TVcgYObUKKPsFaW7eQ3OPf0hdsoob64Hj57NEROtk7h0Hq1bygJpQeQoXdKdjUMFK6KaiQo/tck9
zeMYffzFhefsdUdLUuu5yjuHQlVuS7NWu1iHbpTvyh9krOTx0SUW4yx4s79fw+NrH5up0Kc/2snU
jkiiungIqQb52VV93ZJ+Fe/7ydZ1CMCqx4x1GNrLK828jobVkGw9r7S4K+2S+nDuWa3w+o9odVal
FMkQar/9nLHW1JwczLAyk3MXT1xLNl5fP6NVE8LFusj3eK/zKGJql1SUUO7uoAAn8jKN1My64kpH
K3ZdlSQCjrrJfcyYC5IjoWv2PwsB40xnMllAno7A0OqmZGqKeDGb+OZtQfx+YoNtIj0vuTcrunec
hACAwDXbpYQ4m89pn4UcsJKthEOAE/rZ/dYnACfHhQ8vOchmKG1+YAdo7ALxyL33TcxP3d05s15V
E0lgefU8b3/7gtgqQGAaQdnK6iAzbelrDfn18iwt5mpELcxj0DBFLABD6fa1BWMxjlRw5l7gpw5o
he58F/LX/bH4elt3wK6k38S1hzzka2zpacXtvmpeQzTfuApBklYQMWk9YvGZIkoeDPDsqOBJ0DNS
CzoKCmVwAG3EC9I3ZVux6MfDOeNCSJw+9qRziQ2zIP6rbHolS8YDyisvAfZw6r5TahqsYhnNJhsG
jZR7ehQMVoOrIjs7pVa3d1CxAkZ2mmLpE+Q9BNFGad7v2SZ+PTG3M7Zrp56FIDz4dO8ubvcCJEKy
wtXDJGoBiW8A79JotMGCjoI9/I8p8r4zepGQGlEHUr1zH0vQzQTLAu6YGNUVl3fqOOGPRuHDZlin
ZFpvgascPy47zEYE3+jW0WJScW1imxIIYuiOGilAk1aUeM8KrTIuDvcr5E3mgxcISCmcb2UzjK5g
prwizWrYLu3Es6Im/rjzSfoC3ZibxQLPRzU/6F6hlNNB/q5BUH85pSqJxrJcIs+hx9Fgzngna4rz
qsxa/Ecd/zcbiB7LiVQzLg2zNJwvG3UEP2unAgY+E8gD+e2FtayI/I+6WmzbKSa3K7DseaD1lh1V
9ZJXWVOvuSBUul6HUg7Ppt4Y7usptvFsQiWL4qHvE933+TL1PZHelmL8TCqP06r77a/bB+JyhEC0
f4ZzUPVHq7HLOri02Vnz70KPWrOTYCVhACtvMOBPlGh+PEbqDU88ZSBI5GcIEuHaKKDKRZ+5Rxry
gxcyeXpJKScjEP9TfzbZGyeMeM+VHkjYIKqZNd5LeWWow37zZTTXvwxGcqP/SivdT0OxYIZOHXir
8C5zR5/Uf9Qi3mIvOpjRUwEVC0BltaNOAkrnBX/HGPqUzzELCre2uXVhtnjgYGyMunuJ8kRb3YoS
ZhKIBpot5u9ts7y/lPI3zQ1OzLczhT/oqysH9+/CSA5ZGfuV/Pl5piVwzOs9ices/s9cMUxU2zcE
/U1sRCF/TrrNQ9S2MbLRejwm15tz+bNMlOUycbVvDjQ1HR02g/GqSTGLE0QagnLubK8fWaS5mhuH
QWQT5iCpwuaec5bockRmWtmGaOgkB9IIAeiNYBqspfyVNKDKaA8e58lBWy/7COojiixtJXDFMMts
LrfSNCDTDXJdVARnhMvlJKZBA2mvyO5tmCDBkSHfcE3/SNjfaMQSwHyEshSOLQJGAGi4YEXIAjoM
1K1b1tOUPYh+jgVRJ4RuFaw/bKpDOMpNAS7BLJ5pAHQd24dalIIIYfISHlPSfRdznedxNRNjbaSc
oK5EQPzKwmgZ2Sa968X8zfkGN68zHvFl9qtdg0uqEqdps3P5yV+CagRsqP2s/Y5nUq34lcIrO0pA
H+IYpkuMdk5gHssY8VVN3ZgLofMOekqbXD9XpWla82RzUHDYSGh7HYltbXiEVsXx0Zn1jhVutjOC
8Gu/ZmpQUHQLoRXN5roOrOxNpweW24hPj0PCu/w7pH5fmT+rJeyrqIUMOEM5LbmzMk/gDP6+9D6L
OufmaMo8LFQz9+HiDHJR0T/Jpx8c9IxMXnC/UHjHrUuy7tUf54VsjWGY1a/gqzDoJ4ZpsZU3K6xy
uz0LFStbcPRmTWHRoB9nCnxc4kasMYG/4cnR/7W3j/OYYOr9A7bb7vWLE++cZQTPcowoPCTxFmcn
lzg+EyoG6b9PkJQf+X19wX+CTAgR7qa0QdsbYON5t3evWgnGmNdoLzShj+Zqw4FvU30BIcFqWZGw
mFlS7G7BLQPxpQaGjIAUCysSrYlishAnrHDVzbx6nDIptvfmMYGRgYg29bA4nA2aD/Zzijw7BDPQ
Pls3gCC1aZug3oGOTPDwwo7Q7wlYE+APmL0WFo5axVzDlVBkOeOdDQGV8ju9crLUKf9zbQ40V9k5
XyoFUeQxGY49ht1frzJyf3C5gSss+y22P7gbqlRE1gDGprZl9F8lNJKTVbqoIpw7xww9f/WIBnBT
VqhI7Bf+uaHEGUjyMX9lr49y5YS0EvP26h1BGJsRgy5KFmT6QY8kQp89z/gahvDLiy2gh/T4FwXr
Duc9NE8D7A5cB5eQadrBzvCbfrLxpquLoly6o6PITN5ixUF5K4NU1AkW52EPwNpDzYrTj1OkuXUr
xjKhiEarVoxa0T/6IAVT6XChtfnoWiOG8pD+loFhsD/6G6T14nzV+8dipyOWYZLQlxHSpRw0OYe4
9a+ovbJC8sP4WS4b4aE6DQkbpxqtHzv+UIDTQ4jqKHeecNwvVReJZhPD2LBK1Ar0k5ubxkagt/rY
+dNeaPNGJK7qhhNqJkugbmHdzk/1TFnGm90QK2NQFwmDgnuzgolhNpA8XW/4xe7Q+QuiuglGu9ez
RiTQrmCpQdbnsCdBD1adOeNLCT3RaUoU1BW0De3jA0lFrjZBrhKVdNFVK0yfvI+Hy2lomuJKqJT+
7PkFud2f+JQpGlLOkm5xRiCI/erJLV3kMquSxetlBomY+aawqwZLV0/KUcl7hyuZAgQLvu0MdfHP
yMU530pRmRG//i/3DaD6hy8nSXyqcQDwmbHVCSh6AmjhKd1zn6NJ61Yr77lTkJc0AD4g9WcETetu
RsXbgoxpUCz3PBAAP5O54ZPUu/0ugHtiz6eBJJbkFIzExCpPNTuGVDs8OwPo2zaHuyxpITgFmNhJ
9E3cAqe0Z362FfJ+x2ZO2CMi/FS2vxh2X33i/NgOgtGRJrAtSheJ+BvSmxCtsP5bchjUslgFyZGC
yJR62o23lHO95j94AkY7Y4xrGkvRgOecQ5ceDVbnR+OK/CXT7biDV/qfqpMU0sEBnDomhwN1Wmy3
ELkHZxcTOF4OmnSzUNcwzakq8ZXsxItMoJDDNgf6ds45l1qyFVnchDwzNZ12UtyFfJSCQXyeemgE
yKQ2scv0IIZBPPmcLW2fEk4obiR8jF0wlJ3PLaOfw2XD8XZGGSRQxlHeTVSSm9cpB7r0WsUYG921
S7hsE5kN8YTxeoW5Fn+4pMpYAQEYoXdRp/s+yF+C+QVHhubCulpyOTP0dV8RQEXv6aYLshUBhfRB
S8MO1C8chLC6GScz38l5uGg1BeizIeMBLGbyvRRzGsiV8o14eaCLAmr/e/CiwX2YBdb1+40QWiLz
qFpaF30IuFwdUm0q+0BWwo7a/Agd9Gzz6qK7yC6UktS63gI/IaDSCu/b1XJsMvrlnyylawsLTcq0
uQAzTSgimb11efHSkQyWh7BBwmyof/avll0mF3wJMjD8h1DsZMOB+zRTXDQjMOGtTIX4OlKm8zG/
gVXtB0wPVJuodDKljHZ9CE9uxyrs0cmfVHkBBcpPhkm6z5N3l4oMDdFOiwOpImBmszNuDJEfH5o3
pFonOWhKJAf3ytsAbujuW3xk/UEo7ukDTKs4dpPyHavFDNQjJXcNdLtgVqvX0xkf7cwA684oeIFc
V4XbnyzpvHl6poGQduFEDs8/M8CD49vwCyEcfTSZQ6qknMdgxnw4W5XxqVDWUYGTTkKytMelIEzq
Sb8tNeLTcwfMr9m0OGM3yDVXoeZcy3grBtaapyomDsPelp/Ac/dccwYFc6R9bGMGMR31ul/74Ck4
pmc9CBmt/XR/1Ot363hWrAfKXAGOvvuOjr/R5+W2I5EpsuU5LdErVDUCXcRh2ASSNDYwav63hssC
jza51N9YysE8J9/K2TW3/Un31MjLYyVLpDMINfx+hmw0Ba9gp98dSobqg1KwesO1NWfFnP7i1hSM
Mur+3BULJNIkNa6U0gt6484+7dqrzSqggeb88GJncK+X6KbJ7tMAJUrJZQAhpWUz/2BEmz8Bvlz8
dshfEErnzZLKquBnd6Ok70JOHnZF/jtg9QSB6gjeq5TCIikFg2JIhiw/y/GV7XwkrK1DqF2LjbB+
c+lij8aUdUJt+70+oxeIs8ty9JkOJZ7Pr2rfdgk/Omk5A33K01qonFqZUXhGrFV5txwBl2VGCXxr
BGI6Jrc1FIyX+pmPenkbaJVrH9ibMcKZRdyk0KzoRumMvBVatEGaMs7KeV6VowD71PHWem/wNJbP
DL6w9Tg696ZMBuBb3s6u8Gf+iUQSHY5inuAGiepe9gmHw5Udcd5LDJfQTrwTFpFxGbTp4cjlAThz
fjl3AhvFIir4tbrq5o9hEcz1FQkOkKK2ngzRlNozHQ0hRkdgwViQBdZiAeoHL0zXIYOLcff0EZnQ
Rk2NgdMQBdgZmzWf6O8ObTjfi7eXgoiEP+/Yr4J+jbHRrol/tQ868gqvaSWlleAMqnArPF3GiaDh
7bVlZIosuomE1DGz5cb7rHKS8hF2UrS3+9niduKNFYnjUgteYZ10Lv9AQZHC2C1ysnmMyTymZN1o
d9NfxzQPoj/yK+eoQfGVQ4gj/KfnYg4vqgx79FMIBvUgBhp6NQy82g/jH+n6Zk1e7Jw74Ew4j0pN
lprCQnq/B343ABQfFP8u5E4q5pDkVijYTZ8TXWJ20cq6X+jdwsEcqX9KQ2eFsW4nd0dEycx2RAJ/
EQnuZluKue6ER9TUEiT/4QDV/mFtT47blJ5hy86120qQprpZjEjsKYCFAOw+UzlPYUahApYJbByc
5K0RX1iSSY/mAY5z7pGCMJyg3Xj40ynlLdoW2FUSCHzoPMgnSHa0x9lw/aKI/dat9wdjnbkOC4bo
aoAPbngvhNfHIjmYCLbHr01wfcXeG6BlIp2XWoO26bn6zXCxjJBVJCA+h0IasDj9xZB3toSZfYAG
uNe0b1xdeyonb9JXznIiBkybqNX0QfuZhHcXzeLHeQW5wJvT1QScRiMVi++gdYnfrdiFZIUFVmq/
D4YMxcfs4MPNaJJbMLqz/Rya9R2xTBH1j9HtfVsBgdiJjengmhYduGKv7bSYvz9+iH6GeF+vsV4P
nT4ZCgG0KBNdbFCRx5EMo99NPyGiFQ4yZh/DY6+X48cgFlnenXz4fPQLZRJRaQU1m9IEA3PDEp19
b8h+Ei4+g214s0kX4SrLvgRpGydKuCtuvSNNcxgbKjBgB1QKdwJMcVTgw6t9eHEda8f5998vCuue
pwCixV675pujCsxJKpMoeBYC7slYRWMQdg4GctXzOI6A4KOSR2abd2wmthE402o8qrJ1qV4Q/VbU
Ml7hvChIGiHwcZ7U2i71zryQkrT9SCGGc6L6+2V3w5tgPZdkLdWg6o6WUlNePhifjMk3cXYxo512
vvFFYwlpRldY/hGDleWVjVtZn7be9UPHQmOn9JqgyYk3JrGisc5ukDPIXpEyU2wIQfp3NHCxdTNX
a5tuktqQcPx8gKbvjkl9I29QfXM15Cot0tdhQQV/w25u3EM5VglWjZPXeKcJZuSegE+QFjIG9PQP
g8sHFI4FnuHXDtXI5pw4Lo4+gyUxYMloaS8gVabnH2IPYsVK9TjLawr5pAEGvyxNWroAcEdR00RT
7BvZ0/WC2X496uScCIwtWpZ9pG45lmVIotpVC0nThyhRNl2JPyeOe1gRE8iPO8Qahmf8bb+wMzJj
NwI2g7b6xyh5zzkJYsJr9HL/8L5OKUPhKilNMoAEMXHFI5rmd39zv8FSboarbZoQTlgu+51FROmE
aiBDIWI2XfUxOK1GDXFoEOqpfp8r5i3QQlwWB8wuYMfBkz39Q2fLCH8eafpQVQ1O31tsd3FC0TsA
6b4gQ030hafqtC//MypeQsA9h8Y9M+mtbxxmWTam0maHFZRdazbLi903C33PKqL16td6lGinpTWr
ZYd3TTCvXqUxLhblPMViHfzii++sWSsHmfgoIMb8EaptoAVjHPI914jdf8bRAR0poxrVlUrRoK9b
5ddNXaJALDinY1DJ9kEkOPG9qOLptC7bPQ/xDNjvGj5NW37QGDdNU29fBDZmenxDX5n5AUl6qYTF
5Yn1xWs3rYZMtoM1fwhrLxxWj5MJHw9QJFKHX+RSGcYFsShJ2Z6YP/aL3IdjrKauF24t1azJnHbT
y6swuMmXjQFp/J05LG/e4mD5fDBptr+cN2rh9ggX5rINr/DU2zstoS141PkxT4LLmtsH68Gx50Bc
SLt69Hd1dq54cvWnDCepYDEXGkcuLcd8ZhqegFgmx+6d2ZcFjRjEbacRzFGGWEU+71jkJJIxBsSD
m1egwQa6qWgfjuq3DopdeB32sSdQ8sKu9Ee2gvWsVfSSTQVKBSazlrHmkpRGJWAHylLSlwliWj+G
tuJpxDCAKq81hT/tbtrRWoAU8yeGvj48K3AAplPBGFY8V8BaQlIKLRs4OIB8Z6MPnztHxhiDIGfZ
dOoC4qf4t66Nz5GNkf57SpvAXYH/BoS52ujqqes9a/45mK6hLW7kRFwQj5yQViQItnwxDWlrWWJA
oGM1xKrvfQpnffvHdrCOitYbbPuFdhHpxVRnhl4gjzsHRt+EOo0Sspl35D8J4pRFctxMp/09+h/l
uFApFAtB8R/NC+AkhjjNgaGNVvjj4vlx8J3Fpm+TlFTfzoFE5ZgKL4Mj+3u7KA3pExIo4acZcgtd
MMcmCjFC3aHAfsgnI+Rc9cvC3zG5+1RtDyKLi8r0D1OsEGVQW8otR+tElw1hWVy4WhwEBZ3QKTxp
6nOeArItPrKpCZi51P8vuEHUWmgKm/LARwJtCgIfMamkYbbm1sZ/aE9qNPsVF6p29QDsF24f3vFt
z7XKfp1F4ZERuwA3o2Cw9Qy5Rnff59fOZH92zg6GxUl3vfVkcgIcV/4/ArGq5WNfjqd3sN9Vvn3n
aX08x8+Y3lKozu0uVOT3Z6g9y47LSLHg6ScxwqVWKZSFZ2j1GexY3EBU5t64N2ZsTQqFHnsp3P3P
+7HUhd478yT9cE/mfsuv4vuGFI+aFR8uGLTpVHjm/XrpnRth0IEoVb3bmdnW+Im1O49oT5wknNwD
MCiqq9vrVUxllLX1GDDAGFbrcRDmlFKvurWQs5glm2CMhh2hzbhUp3yf2tdvZYWSbTcMpTdZ3rGh
26br2//8E9QQ0VH1GBQCiJZvPOMKmgI24cwhnVr/YX6qEOj6nrJ9M1Qf5s53srdmMFXFnncrZPyX
s6M5qIBQ9WnKISBFLzTbah0Gj1S6dH4bqsVJL9EKYgjyrOo2LRILdg2j6H3l1qAxCk/AuJpMnX3O
fqoES5BNliF4uDfVMGs3YqklKBKMq/R5abQYJE5/tcqorLt7QBNjUABW2KTkxgjvzDDJBxSdKuzw
+ubGqX5H2tiK3J7m52vAsfWajEPo8YJ/EI8/AV7QbVgim/OlTj8tWtsTpFkXTGXs0zUlvI9IXzQV
G1HnAQFljI3gusSxKp7MYolzradg9HhZ4OMvbwZzcCALpFsasoDBJbNnNsQK5CG3N/UBBFQj2Kjk
CqC5weVXsSUIhyUPsA7h+mTX3nOFesRuOgGwNLKgbhdDGZA3pX22Vp2PMxNKK0NIqwtSOjlCHDZF
InUIi+urwtW/I5e98NsE8MgpDe/YTlnSKpd+Kv4D9pj7tUVGlTK9+E6GannKHuwXZsaeVBj1W8o5
hIeetMriG6ITLtDL4dUtaNX6fCIPmWd8D/Kdi3PXcwagbmLSjYADJgggNRPgqr4KMj8INuJP+xaT
Ybjmdn/EI2P4+DpCky0sWv6DzrzvZ3eT9f6Xt8bmJ5Y6lY8N/DfS/WNOuw7/qZTu7Bqt9idXRmFP
TQ7Ygpyh8zErEx2Pp0pmcmtWkFxVRjjhYhMUGvtOHMjSCs36GgX3lylzX14dFb3PqzdR7TwUWdnD
aw6Nss+lnVSuqAbgd18wLwn906OQHHU/+MJmtpXbO7b1/j3dzhVy2LzbfB1w/tafVPPENWUwWNA8
lzZ+u4nS6HgjVAmAAYXaFSvQ4PpipoPWOyxZ4Zv6y+Ewo9YeO/RuT0pZPAYtfClaWLfH1L2qsdw8
cbfUtGdt/57K0pOVnO2ZcYWi2TEyJ2SfKtd/N2kIncmKkgspLr57HPxeqF4HSdW9YpPCVRMisWG+
HWWVwdqF8b2DLRPZmaUsKEfkohMoDMMZPAOm2p8zqqxoVkhfuqNjRAwyJuF0KAeeZtO0kohB0xCM
L+KwVHVmC+BMagCrdyNueHRO8NVS8/r7xNWu22eZLowFlE7IhFu6uhH0iZy5w+XIKZ/KBC/ImC+d
FJ59PorYk0dn0WpTZ8MQ/HEaqHZYxAyni10I2YSAx2JSKOODOtj6IAStQYUx8DjdxqLmmZ6kJPGw
OacmpzQHofp2redkUqfaV6HwOS1GE5SJaUWshYWv1WAmttq9t3wwdiSZHiqbknvcu8xVkuWsy8Lc
q+3HSfC0t0afbNK+JR+9maqYCYwzgIp+gGNbAi9Nt8bwyWUIibXvh+BlvNnUV9CHDRHet7x4EZ2Q
M2dLOvAZ6EvFlXJEgOron10qedTQ4dsyA7Z6ytZA0qQmpCqgtbjnNE3r+tnU5kg3B+G7ZC86RtPn
P5nZ6TutUNiS4oZ9dP7XUJ5p57hB5IW0aCMyo3K2oML79si2A+8O/gcX79iPZyQGaaO4g3y/KB32
XB37tQeT+1DMRUwL4atIjz4O4MlqBpU2Oa8hFLchlNZTPMTGP+7HyUaQMv3t82NyWFJV3YzLh1Sb
rKFBYnDwLwGYxv1dEGFlGZi1YrsH7ouObahXHN34fBhRtpUKRGLb9DkdZJx9vpqfM++61bEdmF83
XOvJ5Tug4BeJDpaaRuyiN8ucGnrXWujKA0H2G2lM8kBQgx7a2oL36iEllQfIxi6V22tIVz04dwar
OjxFuojg1iTguvmWTnhO3czE1GKHvGBlO2Veqd98usSeCXSdZ4Eo6lH1o89oxhsqy7ZMdydy9thS
OBdWGdUp4sU/Eu4f5/30jIJmrBdzAP2XDg+L9NTSr2MTa6mLjWZeyJmmgTm+lyvefORkOnIRgvPC
fxezXzAnKdXSc2XwIVU1jNyJGHlO6nPK0vP7MdLVj2YUiWToNFZzxSG1vtBhcpx0ZQWuQBQZ+dA1
g9NG9NnU0ouhDY6AV4DUf4IyKrFV+jhKMFyuVb8wqm2kiUqfD7KLm2Yyhtt1ysK8J011Gc3RgYT0
U5k18YYiNiL70lKtSnJAL3zTywHUeX6YGtp0chDLHFND5h8/PPQwf2p1oGXaQaHymUrVp7Qo7fNL
SQ01YKJwj5+HEINPmS+GmgTnRzncYCUcaL/M+oRuxr9OH5VntjuSayTvZDXs3Ym0BlPxQ0ihWcEJ
noqkq2VEO3FXP8tREKgkTjGfB+uqtZUoLluxPhmwo9BD/wq+QQD5J1187yrlPkm7h17r82gIxcBd
ywaGbnWbWm9C3Oaif3OcT4bD/XtTcfP4HJZPhwm1OFQPPR3EjA2hw4OtubaTH4d+T8fNOyy8C1fe
ouLxWa2Q5HDHrnl5Ila2ABdVbIJ0QGCv6IaJqJLoyLvcstthGnKDN1kEMFEEM9UuA6Y3+R41SsUk
aQFwPMj1BAwtzYiwqmtk+jr5ZSrZXLrX66G6XaPPiVyF23C033MF4yNStM1T6bVrq+684k62WB7e
gA5a2z2R014MeenKSJlSjNdBgjakMDkfM1H3aEGySAmbA/nR9XGlacRwE9IauyJad06p9xwt8iQV
YfPFtN8GlwtJS2IXSa6xrDF0tpdp/g+BoKRJV9Ld7DbEoE9pAgcirzXAJn+s2XmSKm7JdRNvQuad
k/9tO8kYE0kfTE7sych2QawpG/kJKutJtQYDnMuXcQ8OQRj+z/5Ad4xk6AGjvhLEFwVdcr1R5C/5
OoayFk466BEytQiFc4BFo8GcyZsMSlz3zh+wZNsPv+WBjjs6fd5LT0MrhrNvLlBDixRGvBQDngok
FMqmQQXWyes4UmTCcWC58OoxNUp7dSZJepkrWZX/VuYjva3z1hUNRKou7VFvBvDVMlsQOlQdjEZy
6LS2FKfQ/iyk/3L0gni0ea3EGtOOqQ3wKqQxqKx0NpUnVDmQ1sZt9T4c0wDenDQ5sEObuqo8PK/Y
1w0q9nNyBNe68Lz68jIjKG1kHwD+Jqi3TpiQhN6jGhPuVT1EyXxvtgCOW11Rg4o4UQhN7CKuHil5
5FxDZT6RM8VUq9jhnNi0sZKAdEjx3aqJDNTng+/12L4vbFezjb984jxZt45aVCGToNOwk+CJv8oC
RiQdb7AVRoltE1ESlIzkt9JFA2KAUGvPtifuljRa318okIDYySqRzypZLCJB3rhXKynT7+ZVVVKi
F+VfaxXV3RLoDKLFg0NIciPE83Xgoh5e4pYHZAhlHbNnkkNWdu3CTBsHHGlA/m1/BhQRZfCa1ZJL
mg9aJnBSAMyqOjOd6NGG3LgJ2GlS2UvfLDYgk9hz5hXWstYvHZbBsgBnFgfE5J7eTNSAgkei/JS5
c2wcRdOUOFKeOhf1XTAg4iKv5Oc2uOLvlmgQ3EJpFj7nzXQJezsgBfZYcfOjQvLiE+hrrqaPXcb4
W/DjVckgfHu86lNYfv7GlD/+8LpuZ78mN+UtNKMa8k2hOVSmMPzHVQM8sCFPr/qqpp2GloXEjGIi
EflshfB9jDLZIPCDpWQS995g4pzxHxYOfTrXO1zzOQ0BeYrkauvNDzk2dvIWm4Ih/2Fv8kMuzMic
kLcT7AYyceJFY3yOvls2gPfiWSxAyZ+sjsSfysEyavu8lg+wllOforoMOfNVUXajS+t5i1QUr4LM
5W+3cnNQGNRWUDbgt+84xiziEvuH7NKjAiWLtujLO9CimX7/drtp74PS43pxtk9kvRF6AkztSFoT
uXfUGl5Ph2dT+dGaVtQ84v+2RCCpq7d+TA3w/Mp2STb1lnKHkJLFTY+9ZZJ/FSVqCysVr5WAzICW
46ydBZqPYKpVeG1Nq0XjTiuZtfWu3CZ4/lgeM9RFzeA2kI0uwegTtbWfXJKlXQPLu8j1tKNfQRet
6SMuMtojkoIv3ndN0eSlcuPLUOMmyx2y4Z0KO0p5PJdRrgKKGDbkiox1gV2QK0ToR9YOP7hdDm/X
6v89h5GboAAOm5/Kanq88f/X3NPG2DOxUXTtjUqBUYelmcZFBYLd18Ons/Ljo3550OZSNTlIpYyB
jzd1J7Es1QYanergm7gbK1X/ipSgoxHeVf6rzvTUShnEeCY7NxOri45Lp0wRODMwTW+53NvNu6Kb
7F9zB7IHeD309HlW12PQV9EnzNP3aHrtdCUltFm0vsaeVxDx8AkEko986q/NsvcLg36thziXWFha
PP2LmqXVPVaOROv846gdjckVrHsOyTkcXul18kxW+G527YvoMfKhe/U9/LkeEzPi9axI/AjZUl1I
ovfRn7Nbj2yB9evGbN8Tc49pBLDGOFIR6MYjh2PRC258oQn34lihO2SUZqrThp+42XI70aaeajz7
Dqu0bryJdLR6BWDcoQXMTFmuRAr5uhqY9H83FVnoiJW8GLg1LWNjdzq+dUab7RkssDta95/x4HoQ
YxxJFtU+wReLVvbz0kO2eD51jcAkhjAPaV0Nmm9eRPcEJIfWSmkPUTcfWPZwuFe9ezLNvzhxcdx1
T7LSDGY470vt41l0hQt3Grbupf3OSR7bvFuEk+4YxqwG4CnJQZXgGHOKu5YxJH4JSX+EGcqEECc2
3UnifWqv570IXpSBC1ax8gzCddLjmNg8Zr3FfpxM0D+oxsegbl2+QCIfrUbeZiVdZ+hjbu3xV8fM
7SfQBeTxZSvQYRH/7wZvhLpS5Yn6RUKDX09JqK3Pfv9lqur/K2Jv1mtsrTwWqBlIULxKXmfH5Mu5
Q4HmfjKvW4+NAY270YHV7+feso4QcL2O/8xwt+YL+Qs+gxIwR2MQXlQHFVNOCGlkpss2H4RtUlvs
sKHO9iGfRhYu7N7GC0Qi5NB6Ma6++esjhKKEX9eZFV5T9OKm7zVf6MEvPYDFTHnYavzAMt0PRRWq
oS1G8f+EUVQ/XBXrmGJHcxT3yW5MlDfRvc4pKfVu4w7Eymb6QDXXHwPVUgOjrfCc9ZLyNoPyu/bQ
cl9sjqU1AmewfF9nL+9rMMTCNjvuAVomxBWYCfTw1DVdM/IiLgcIjpXMCSKSmUU9eUq4md68gqWj
gJdIhpGhtoSRPsb6DdijH13k8mAvFqMfxwPQRPlVoAn4D9nD+dGhFPufCYKoGibCr9QM0uzFtCCe
eE9c0UfFt8YM7l1xovtHXmqKXV5ShYbw9miM6dTLOfDp/1Lum54qd/TQQ73pRzI9Obs/AE+WLcnL
zoR+CJk7pwjqqkP82r6FqltmaB5r6Ui15j6CnIPw/RXwK6rOSMx/pQ7VSL4GVWI/1wE2nvPlNieo
5fw0HFiPt9jiL+9N2ne3LBgsUlPrsmuBo3it8RuSawyrL18iuP2bjNFwr4oSeZpZoWbQtPTFhElQ
spfgwSpAaWCTeB353bbiIhD7Pf89IS/Jiv/0kjH74w9Y4EOCsIg7POG113JnOCPJabIm/wkbqnUg
trM/onmg7S5XVakPcPVEMz/GNLvHYf4dvIhzSdzDEz9SceE9Ek9AsjEi8XICT1bjOKoJP232g9zr
qljHGjnR7uYyUwKoDwb1d9hp9k6HTKfM9/RDX8dvQgbuA9cHoUXsK36if+kKoeDhh34DPlfdmKTV
QjSqLVvAGvgMyB1V/AIHcDouYU+q3Rw+P06FSA/AghPFt6UL5Hlu047oxG32WnZ0lu79r2ZKO9wc
1A450vNKzlrD8BP/Wa8R77RlUuLaJpDCKMwv97JgUAu8nyE6m/JYw/tIPnHCGtHd22B+lA7gZ6QP
sZE2SBg4tIRLmspZi81/vA8PXd7D0oFJ4tlaJjAuP0NtQuzJ5p5H/5N+BPBjLrPDsgPzu6gkgxRX
MIhD+x5JMCQ3JEL0MnZdMYytBHMg8cU64B8rbpuXo+EVwRbVF9OpP4Mqrxsm90p7SywaFsZxHADv
m2KhzgnPlvjLI7SWbKKNeueWCcjgdzkr1SzUon3waMWDQhi7bAf6hSnfoMo1R6wIJc2b9WAdmlEN
XYYAssM7Uv1so1h5S0QVlzlM1rqXvO4H/bWN4VSqetyBc4oD90YHJbi6p5yk7+adY2IjRj/lZd+d
K+R0fJKkhgV8w/s31yHj3sGoIt9Z/nf/J1mGRFpaHPzEQkAOY4Zpp7HOidifU1bj6JqB2vtBkE44
jrmpNvjendLMnSQOU3bNq6QuKrbDpStUza9xyp71QDX8GVqzQy64rUPxr1OoXaRVhe/Xh1ltfvGH
IML73c1vxhshungWl+YjBKkOYp4ppoBt8wHKOdQJZL9YwT3ZJ4p3CKRZXU9GHyKli8LuI+cdxonX
XTFwiuOKPbWFQAqP1HabZeilM8MEe9dae0rUbugvMkS8CVLsvO678BmrORtazUXAMqnWG8mbLNkA
UbJu1+HKIwzjPGGgK2mUnMjkhXIxFSLhhQY5O/J9zs/eUIoRdssBDJmG5/SKFllxb+fInJrmJOLB
shYkr91R9QHaBTeFmqtV6cCj5KUNDZpK6x+bRF6aReUIt09VH0IHep9XjBS1FuiRnfjBugzcDvRY
f4wWkY8mkwwAVpShiBSLOWygqo1xeVFDwCnDvkyQE1gAWvJljQSvOo3MQpQKyvcSh5Md/X2fTEL/
FAquF0Bb71rkJGU/pN/Mpt4C3j4kWp2A4YRO3nYNB9J4gkgyjU0Hak460g6JaKLsEu+BewhH2Jfe
RjTChoZ6TLSe1FmiTFOlFWOLRVAFJQ35ubKSWiz+tDv9zuy9fAZTodBsU9LUHqlyEguP0cpY3cCH
qr1RLd8bu3Bl9v6oi0wjEFkCn8cRfJaUa16GO8QLkOoBF3I8NdedurTjZLCS7udOwptXsVlMQguH
s44DRJhh3TAYFG4rBH4u1Qus41Q6EcLmUlcl04BnD8a+KaF1o0ZR/jSuUrpvN4sxJMkYbqCtUktT
i8j0iJVetywyZR/EOZ2HqWUVHJWAzFt3HxXl5kVXKY8q2vLylVGkWcbRksA/qvlKqdAQ/ZCRyahX
be/l03u0t57aj0NdnrT28LIjwpkxodUf+qJubflw/DB0P/9LVlQZv2lik+oSMZj3vHdVheipagop
Jjj+HR1riOmXPdMzqst9UX8P8zypxtD6FY2NlKGo3Dfvoh5GewScsxtdfp99/IITJSrElkoB9rfj
EGFTL6RUWGQH1LbGqCBwdDSYISG5jvfWvQoTi+akNLymzKlUwf6N2tdzLA7qvsFVSGKlcDovL+aR
MpDYmGeNeeIIXAxXjOal8AWnFq0AptzTQ4TUAD77eWPwnmgI9zV2hoI8278RLin9WgyM6tgRwGKd
NKw3N8Eh6yZcoAZ83TciW7tJeLTMIaP35jQPKILfFfwSEESATKmLvupOuVI3bHvFQGA+XzNvdcij
n2ZBYDh79GsDdU6ZYh1laVGlJYhdoErjLbnh11O0xZUiqGYUwiv1YgullBS2Y5bE86GpxZchQBSZ
clH52QbnPkU29ik8RTV6rhcFEggbO74t1LJIskjE1fWeEm8dP5vYHOxi4hT1j1ApTlKHEIHkJr3W
i6Er5CmRUIX3Yp/P+LcyJS0APsay3eL/Tmnqz2K30BqFcidnivsfIDA5PsL0+kksPusDY6p3sn1G
zhaHPsWpqoGmoOitauQaxClFb248hzKJWtCvGjUGAhRgGC8JYHx449/rORwCejza/2Z0IV0fqQKc
brCdtVlqHxr1QdpJKb3SF6/MyfiiTQgnqWg14lv/gLTtTZ81CwYr6yMREL1nuJk+A0q9d3GU0xga
Mzr6Kd2jMLiuV1CODQRRXWaIMwwnsQbpVzUcc0C6K5fk6xUDJv4ZgPwRpLpdhTYsR5TNh9/Pcvwm
d8PVTFt7g3gOIKiflAhIgqWPbRs5J5eCbqgcYSKRHU396npC4ejiFj2/RphhHhxyQPUUruZq1sfo
L+5ve3wbFn7tGWHmVFdrxNviOp/gxlYAfjaO/SEZbkxcyrSlVWp5hyLF3x6yahQjKINd9JjnS4su
zCoSx53iqb1yIe71DwTkCkuSRVeqd3WVvaHixKrhXU5DJTu7I+kmgehIEdZgRW0G8HpSnuMyP7Rm
LV2TjiedR5pQ3rVGiYg7jSfAvQDjQFJC3GltVfFEdZlzL0UAbSWFV2pj+/oPkARl/AySJYWg4fNe
2cOaearGDkzsYXOS71IweTX8tizXSGtdBn4UE510tpRp4VvyrMzJO5g0N8iYshmPWb/zwLw30hix
rpfKN1WbN6IlnT55ngwHH7gPeAPZqSLphVeG28mSOpa6otjDIeHBRZN3hb0x8iNxsUL8QzTvnKOE
r7yvvHDE0vD5UsctdNebchQj9mKrda55veuOtvAI1gFSd9SIZ11B53Vxc/eNOGLV1TXAm2VUp/8p
MVZ7SDQxWLikv2OmwGG5+CCn9kK2dqvWLk1u+fG7mAAmKegPc1wCxtQzACbdRV95q3X4PaesETa3
Fb31/Vdgz3lNv6odDqrO8J/MXFTaNpvan2MqO12JMBonSc5zGsNyd13FAVAWVLbk1JlMgxqfkZGR
w6sFmFyeSJlCooQmNetwqlGIn9xYZ8n1gjokT0b/ADBvxT/zlw6mxlBUsKr91w2ph3HoHHPns9eV
Un3vK8wyxLb5wJQnTobdhsf25U7LqHEA63aLfQFIoeGLHFCCYpIY7J3q37Q7yFbo6KZtrCsit1Fj
rRjaGentkJub3KF6ptoPSo2aMbXvVG0kjvH9ObLrRtk7Js0F0sCuAtNv4oxUsqGoA7BcQEsaDYQD
Qkdwu7x254ql4w32dVQxXhNHkBnUzsukje6Hr6cQ7feqObRu27NKi1N35Da9Mv/QiycyzTLIIq8B
Buw9PStrHMVPdvMIReIm3CqBbARiIDnDBOX+5piNLCvpb+fFQdcXMsM/joZ5djPKR4j/lz/GNwXY
jILO890gJvGvnmpI+KhX8fVtEUwbEh+wx8J270w5aqCx592OwQrqHPUS6VhdcvE6qsYU0GkuL+rd
EN1pC7akVYrSurj5XOZNLMRPPsejgJcwHBciBRM53dnf1tXaFOEyRufHO/Fb4e9Xza7nIbVk5/0A
uPAfHbC0buTcD2S5e0a53EP6d4SHgSj4b6KhbgmLfOpa4LL1ipCFKrh8XSSG11uCUioTyjlEJkWz
piZPQ/f8mcjmQ4lcemKFbIjYSJTx+ViORjRoNpo/VanWVO5j4PjP3+kzA5+jgHkRF7aV8JfiUfFZ
nVt5bPchY9KRm4RzN54LRHfaaYKGvG9SrNkCcB4JPW5IcV/pu91E+BBY1iJ7XxF761sghsLid8QJ
Swty/EG/7rrTglOOtmm/TRM/rNur5YCMPfDG1e67aAjaLdaZlIyySmwfBIJo89Y4eYZUdNtOH0/a
2wNsh1d22r6DbdENk+bYitduaYxZ+j5IxFwRI+0LnEfZv2ITiz6j5NKaK+g8bFvVZ9v35KTOt4vS
uxc6L+1VMbCgD1OlVhb9rAzNBTRVuZNCaE4JvdlhbVf1ArgjHrIOO7TlEQ4x1MsXFJOfr1ekwC8B
2X8pVOU561pFOuEjexak4hXUXWb+w8KOlptcDM71g9IT4jaHvov6Lr3cbSgZ1JGi05QDfOwxcXUc
+ktD1CAIsiUnJkcE0dT57IKZhCpNJUwPZGC8iuttOwfg4I5MRmo2L7uUU/LA2TSSTXMuKcA7lO8c
Kj6LzEvzNl0yn700TWx1SyLLursNSPqZsHLoTqXtebNi5gxlY+n10rrcCUREEOs0ztbDagW+YDxq
IGrmgBH5X0meaPWpUcZ6VRvHOawG4cM13IHwgo2D5zOeJciWX6BsKbSuDlhTu7k5wLbpwThWSWgM
PiBN5zW8/U4MkriNAzOuyVd2nX3K6qP1b3tPWwa4ALnGcywCxCqrbBPMYUFKPP3+J0x2ADGkQLVO
TzyxF7Aq0o1554Nz0cC9Y8SagRqPZ+Rw0fVn4Uvz0aoBD4D8ocn/jNx7n5Omxf4nRteho2HWwFYt
aCifVc5SX+1OD9vEucHYfAmA9IHe2C6Z/91L+NLEtgI2i1Z062qD0bVmPetao+eC6dONpYTzTJLe
PWTNrNrWQRBXsG3lFzchhRSsU9tRjfsSOHCUdt+z4Jm7Jl9Yq1d0n3X0j5VzlLogRC/8wrE3/UJW
77kxN6PElAiY9ozrRkCjN9sOmmbBzD49W934wf7UHBwykLWMDbGT3vZEHHMXulw4xv/QynIjddG0
4iiavzkXLgBVlyiBn6WVuU3QSBKPHsMRXgzusElPHV13PFB+bP0ZGhNYSh7kY2VLRAulAWd2fNO4
1zAV5ehGqEZsm403UNd/qSlHBe3r0vW5JR56m9ZG2uv2nmUuwFmiM3tTr5rUjqslnpIpsqx6mw72
XglJhVSZ/wq0mdRP4Ez9ftBCnpIYTVHR0Q9SyyaphpOwKYQ6FqvRJftMDKiPIYu+F68cK55IrK7S
r3ozr01I5D3f8MfpILzMdsBFEudMtIIFe0nGFDwaR90jsGEvc6C1G2rhn85aMQyOOVJAihy4bbHf
cLWqTrpRrlWdSfKFJC4jekHKlnyCeG34QqxYFqMGar/zODlBn5ukdHAAj+CUMYpd5TbYcqsHkfqS
5/GrD0jjgJMnZpIAzcj4fVbutBwLSoFRYJCC7SK4mJykPTd/WeCksY5hIxBgdj3w+wZYyuH/pYiR
yVdQoX0mbNRbzwhp2Xu1l/v8rnStRPMmhIACWZpKWMnzGQxNGY9uiOc+GNeNf9NqvNDnV2MM6fpn
EjDYyZ1bSt2JBRCUmxbUfZwBbajEAEnNsAkd6BeH37PbAnQiVW0TWM6s/78b5IuhtdAUrVN2xiRH
keX9a7s6AAhvElMzvcjVqu9kPyTDGgMHF5cFU6LlYohCqFiitTS2fuLn6B36kDFT9nMr7veeifmU
rh4KhOEdnBn92qOMPPsIaNs4Uqh8sKz8RGDHVUj9YSb5O9l9/oxLDw8h5Cr4By8ZC0UpWssdZk54
nXjUteNLA3BunsylfBrSJG7UNqh0Q7iHfO9ab+5wv6J8mKGnV+PVACYZ3PAWMTZdqJpp6ZJy/kJ3
GFYd4Jm8IdHc/WFmYvNo9/p0xd6qPa3YS5sgKNzJXVacMrSGTkMu+TjXvepO0wXfVI+U8z3uDjNz
fW3kj+ahHBve9224v1NvJGH4W0S4IomWJS7+/EmzTl6A93abZ2pN6w+Aj9rbJw5bKTaT74XeRcWb
UjRdMtaXIuY0V27G393bBNP7qk7NaTpyQxaJPz+A4Kn2oH7FVLFo237/ZqHoxadDiOhaWi9HzkDI
uLlAW8MZNO0QvSogSSVTLqhHCqVi/tE2WvYBtMH201xdbdnA17CBzVrQk4F6HWFb5F6sWbeDX7rF
w7+6zkYRbk6WsA/88csPWSCL7K97HmrByFNM+uIcpeT8oiJhxQQMSxs7o/UfmGwe9I5P9KnXXqLl
fzCresp32+5cvhR60BVp8aOr9uftQHlrQc9qu8Iwlm0Pvzt0NMJK2UBdrj2eD/BD+C97z+6V/y+O
fLff21yOvSnerBFztog0KF/JnRAKgrL7z8U0M1Aifemf5mk46zV9K+t3cT/CWnXySAEmG6au7bH6
iR/ciG/AQaflRWXchhLnRdKBtxU3irdONBhX39/lH1o3ahFTrg4T5QsMyueEJ1RDjuZ1IoXo2PWf
C51X+sdsNjyfXdSu+eZeyB0DRC6RyoyH4XHbMk0eOTiC8sTdCojU9uUEXvIbZnVkuKttVrLve7P1
KL2ALAX6ENpdm/UjckWgIaKlKjP0SwA/2puJpJ+s0NTUX8AA/P04kzcgQR2gfxHQ+eoCQI4duXcC
dyZX9Ko9sIk5X5xmx9ZwQ0GJ87rNPc5CXCJvoik/tMaFQfTCmMzCbh9RBD+IKEaizsgJbeM9FqxI
3dTG4WBiGBpCvS+vg+7Z1xRB6ZES4dwDIhJB3fD+8hqLOkddBWZt9ri52l2lYK9FvkKBZmCERK9z
TaCufPiy+7t9exYDsjd8SxzlgeA+m8XI7nDcK1vmquhQqmDBpFrOyPsnOrEnNQnVJk0pwyxyHzoq
SSOA9RRfF7mDe6dSsTu9vgfctqNrzplmacKvtvRdpEkoFzczwEaPe0esPgsTKIv1sOlk9bt+im3l
52wU+R1Vc6irsyVJwd69GLSCYGZfsUW86fEpomMNUkgFHHl+N/7oedf4fBD3Fq7Kg3ztLiUD8LIu
obtP9HrUN1pQ+PvyKZwc4BgJl0gRD98KNe6oVAXzhYeM83qk+adDWUWe6DzXCyIleAAanxAUbWi1
lB+V/v8ryLAL4ASa++/DB2ei4yMYt5yRrukSp3fnz0eogQrb/jRwbaRqJVJVwe6p+4qb12h6s27Y
LVlOPIhh4a4l0Y2E1V67IJJ6uBxlJ9nmrYJfWQ+T2OWUpgtMHqDLhWl+2GS5bgE5KvO/v2ZpiOUZ
AIAE+og17J1qpCq6He1+T6NVpz4aXIHU2jprsYxMK/TEz7mU6GXt2mLOcBmZUWXnWhbjAHV/viAj
Wmm2cZ2hWx/1XCbhFtFYY7aXCADbh4XqeGySnwzWuAAxD8rzb/q/zVJLc8sZHGziy3opPsYprrEw
BUyPy/cscXz9ds6VW2icYkwPmYwxmhclT9LLSPwHMUb+21kj1yCxSOsKFWLNHTNy6fwSp8IrJkcO
32WjgxRoG5uPV3ySpPEoxX4x0CZ1YKZkhoa4KAfNryd4g2mRU85xiEeQZJ4TGrqJ3TmUh9ISiTsx
yfiLg8KHDiarVd327ypOQJRms5fUnzvJxvIZMltGDTStKUZONctiLfbM+zEfQuLJmwpNpiZOf16/
BAZ0lDsnAxFGwEfHQ3s88eZw/YGJ6GIVhfaEAOpfWyGLXE6j9rsgm/Le2EPHXvBTFeHK7NhJfJNn
Ava4mR0nkGkF7U7C5D8kxtKyH6NQP71okzNuXHq7bNC2hfIjV04QmxYO2SLIZd+VGxc1lolNYiIT
+knuOw3xfcIwjOeORD1mAchYdBa4AZLCs0inpSSs08tmb2MgNp7/LvwdzbXLSSdQFti23V3WyAvK
/gZcGd87wtC7W8uO6NSyi4cITBxEFlxBdu2KSYizd3CoA2BGBAycIrgH6EuGevQPs6dc61r9DtRh
/fYLirAloRBo/rIYleQQDBAV7n0HOTEvxi4YxaQaQIztRKdjyejbnyrqbHNPI0XyHONcdPSr7jt0
lmdt+4po4NWWOBMhi0zOaV03FDwAMYn5dK1D9YDMv6Sfru7oaSREPi5x4FcgKdi6C1FoXWWKeSEx
CCKuvN+N0vWd3SGdJ6Y0cfqbr5k2SmdCUzreWsQo0eHmdXrGC5C/5oAJSM9jBDFuldPrf2NbRPH2
vclIPYpC+r12ITPrHeKKdkmk1xTAAbBJDugwiRn7bnUofjP9VfV8CkEcxpKC1EbzJsIoN7oMtdCy
hTPeDjz+WbODncG4J2gVGmmZRoLC/jEFVfkjZRmfuJiXeIZUXHJS6cn4+SIYdWYGZJRvuwihpCZ3
4PrznI+eQTMg4G4FG/nI5PwwNFlVr5iyHLR6d17NbmxptQkM9YfsipuWBS7L8VrlBXwXDrKrxPTn
cJVJjdvVrz6nHMmo5L6DuhfsPVn1QE5u2aZ1XSj+/ya3A5jYtNyWKGlqBFfKHvOl2RrlE5QSegV3
Hbn2UpVkUYVB5CoHAdzsOF/blZ6inVAvW7Xi6ndzOBWhNdDXNgSP5rpFn0e/GBXr4gfaiU+X1Qvf
whKNOXR6+KZmc/b/H3VI6lwJf57ZIcSk+cAinYrN+E5BH0eELdJciVeWjyaSwjU6LcasTve6qk1S
KkTMhbbYaeT6BTEbHnWYq0VpKsZNCjRhPrwdmS6FrDuRncTFpj+1ShhumCeTXs64VXnAtfdGlmWc
Zz4HQyboPMC1FhfrU2e3u0etLrDBR0caXCQvyQOgE/BhbzyaW8C4rjK6BhuecJiC3O/nKXri4PjY
QzRZFs4d4FsXV6KQAvecGktLhbax80xAlF+k4Qpq/jmxcvljSH3aBsfAWc5rlfufWJng2TNsmyMO
IsWULl3fYaJ5ju3n/cHV9iQOnwL8cwmJbZl3S8k3BkH1EcQdliCD8NS3i8cNAkQgSdzk9xfmASMh
iG/b5owl5oj/QBzJhYb5Pxy6UL2dvj++lGP0XXyWagvJ+7Gtr9RZTjaENxBeeUqANBatBxtrc3pr
JkeYD7D6MBxhT6kwc8d8AFjWEXmwegQfhop2G4FndJtRhDLO2//8q69H0hwAsm72UQNTuGpwfwle
Z4AtoHfOWbrxkrLtvjtp8gfPa99C8pEVBho3YgQmjPkRXcutjOgE4mROJjG4oxMlN8tvq/TZeQAQ
Zw26vDrc/kGQjziJ0vZxjcv6pIqb25WCmtlC4tWZYk13X1QiIRpXy5JJKyetjPoF1GR33+Z6airv
JGwaNmkJbL4vJjEkKJIlmXM9C38DPuJv0bjI+LdnKcLMSAnCQNzoG2NeJdlz103ioUlWBVnDm14G
KGyed04x4gS4LbgSZkXfWnv/YbgAJK2F4UQKw0Iw0n3iAH+HX1PxtxARa8mF23Mx8xMN1qvXcAJD
EfNz9g0ghqWdPYWs3jzizjifAk13k0WLpNu4+yn3k9/pSzbDRAu++BNUHnkaPSgG12oNcMeL8jUN
+H+MkrAHqwqYGwXBtbauwkW7P8Zf8+e0hHls8QLECkPHtHtc9yRALDM4B4Z6WW2RD6UC5c55RNDi
wuAtzt3zJxxIRKE6NiUS6NmvibCDaEev2WchRmTfxWwAxQzfWeEwY6OXc8VLYLCODCMnmJzvoSeA
OA8gSWD6oZZ2TxYLO3AFXlFFevSFtMTtdKOYokW+M2aXMUNUj9cUsXUMQlSY2qTL0/0mwatBDG5g
Koqrlakgqkb7dYc4o/eA9zY+5A6pqzQ0Gdaoxp1e5HGZQco+GjxycsiwRGbqxqKz7cxF9FBG4Txf
a2EL0G9f9F+XSgQ4fbcGxi2Ei3CcRTBa7Mhp/uFKpvp9JCO2xFrfn02AbrfmAeiCGHsINmsVJ+ZC
QPCquH9vfRqxj/t434Tp761Wk1loZiCaRFvnHZ9EYSkMZdyyqqRLHR2523wltyVKgc7WuQMENO+K
evCfXgC6MYkZwPiHsLNVDO7SKdL17QAvuk3yxxhYDd5KtYifrUkhcFQ0oLKR3EVYzNFsXrvNvFez
MATpXWjb5QrypI26wBwSv3VKbkKCwvF8khwK4KeGVhwGFVN9SbUa5MS+RwpLESfZRlkjCVSzyZ0d
zzGn3tkeD5abShcUTAcgy3AHc8fn4dLIALmFMVwq9pC7CYX/kehFPGQrAkbWDS6Z5IArxCFUIqUz
rfMWROIGO2tg3Bh/amTZWLhTN9Kx9/8rwCcTT2fchAsyIGQjn+zexv/F3VzDyu8ef/+PIz3gbzh+
PFb2DvME+gcJKlYj04fdMMKzH1zIDluoXrT/Mvbhii9hwCp3S/X7Qd5IzZUY/JevhVwZMsegOaj5
r0JZ3ZHIxL4pLIBr4uZkfvv7uouL8QC115LnjckyurK5x8E+CC37cNwrNW8Rfbku6VQethv/GN56
49nDMliXJcCMp52S0vdL6iwavh5109hP69b1/lHOj1NmIcJ21Gt1Q+dz/Rl4dGWi4PE6ff22FsYc
CuuGLVs+fviGzwUA8CfRlWxf+19LO8QNdSCTeIny/YBFS94ULPZztHWMUYZ4mUfRboM0WcGQPC3y
eZHsZAHXvbsdpnolo87AcCN6CbuBVG/vKAjPTD2it9dWrXYNZrup9ND7nIrP2wgE0NI4DHjQfFy4
JEY1bcnhMwkZNk8ufJuaeUvoI51mccyxnWdpfpzO4LOgjjZbaVHLH6Htgyo/t1e/P62mxbEjX/B2
xUcoTJhPT+baalSqPSfjByfQq/GnExKPx7KDwP0EYTKzfqnrvrQ3zWC3HrZd+R4ZpnfuNDXAecQW
5yNfwwvNojtmUoriOUKwfg4Y4n54KW47JQrHCgmWW4zQM3KOV8ibsWrb+y0VLc2z27EvDW8mdxuh
rcFoezWyvM3mZkLdXrviDxcCrX1HcaFRpd6sOY4Tw6Qskmz6AArF4AOoL6QCuzD7FYsF3cOgMajc
1v/WcY7v89SDWfuhc4VluVFJUm6KeCrmLMHlcZ8cDPBJqR9VCCrVY7x6tvP4LFF/GSS+QYAp8neT
UNqUKzlYIMlXtN3qtvIcnF7fcfr4VfQVolQa2K7dC2N4RfC458DtWyIqE4ROpYBQVd8BiUeFVDI7
M+iyHfI8qCIjoIh+FnMx51OJgMlXKtktp2POt5aRm9zkgT/6IqU1kmiGi8TajGQjgnt48p0dK7PM
dxJkmkAY0mtMy5X9V1d2QxDV6Hszxz2n2gCYtUiowDieoGzxW5cYUhiuANQSXk6EQS7mW/6n4s60
BNA+cC4mkjIZso79oKn2iTzXqwcuqxDOkDqUYrKqBTgkxJ5+/P4KFFK9aJakWilNoFxlifg7WoB5
+cjt7BKfiysSM2ZoekS7qnuYFCAYpPMZVpTuwCdpxvsJs9scPGIpYhi8iQvNkViauDBZ/yHG5VSi
zr3wIYO8NXX3B3rv/AAXK3PTQKScBweTYLmyzHq8hjDENMqMFGTlA0MQRre+DthpNUBK9y9XpNfk
vCorXIs+fOIT93GwFDz6mRlHDVCVPyoR5Zyr31eo+MuabVBQbmrdObGixNKETRt3+GXGhJzwPonu
IfEN50OBYV6NPXY5JbDqgRLvwsIAwK+6aksLEbCkLLxzB7iyxCJoLjLmxJUdR7YbTpFl3TGyn+jF
9TWeG+NSC1QYIpibd+1kyAvHCObfrJt0vXkhcVy15oJLU94l0mAZk74+vRw/t0eD/9KNes48GgiR
roRBjbu7hoK9vjrBwz3BdGY8AD1xWMcwHnFfZyd4JIwibPeuwY0CL5to0pEvd7PirQ1aLAM8MyY+
nhcDUlKarpwoUYbbFPCmc0tA4jbvDYa0DXfgUZemmiYKIdXh+fSxWJac4kVSvoW6KH2xMWCLYW91
SgXBMVIcsKs/cG4MpgQkfoo3ikn/PNXj/WKhRn7lC/zJ2aJrMSo1zuVI5e5RJjg2l9aLb2PknRiF
phqzri8wpOzvUMPpSb3RA2f3qrmhiee8g/o8IwQpynGMJNzuRr7q0SZxfKX7Us8I6Gy2GHfFWaxo
Pnbo37tkvjlONsQ5FY9yJ8NqqHBsBeny6plf703VIU4So8PQmzqvdlClSttIjfs7K4D9qhg4hpHo
nDuM+512/T/DNjPr/QesW2oUyPaOBvWEOr4s+2YHW/Cakvj5dn5mTrILcq8YqMf1meG051ZObMK7
XiYVgkdFhRLqa2RA6Xk57frs4LXPfxwWU2OCfZOtFlOPzlT1LUs9zVjE2cnZR3uCN29nIPze7Mcd
YbN+bw8J709hi5qviz0Eb+WejOrwWO4FWXXrgcFMX0F9u/fba0Ve7YBSi5IiAV7u4HkLzBEtteBY
VbsVD1gJGuNOZIK/V4Buhnm8fEFUKSsUvK9pLoQuBvhaVYxCqtAREhG8h6c1qNmCZTkXdAcRZ9SF
+jFdTHlFih6VqaW2d01m8rxFvwdRfYCIzLLdWCbpqF5/gSrFNMsJ2F8PRBNyJ+1ew599sTWCrbFM
nySGML1qkW9Mj8+n+10J8WPrQOy80N2TJ83x5t7xiqHgFB2M8+hY5rAuf4D+d/74ixkjoNYVzDBM
qJty9s7XjGTV2i1BrJOy+Ks4aPIl6bCAp2PdlsTuog5mJezIZ9I3m6aGSDFuaXJWD4uAWCzxPg0f
kvRzr/kPMNN2pF9GxL82MnDQD+zbVqZfnu1KP8mvcuqJV9aO03YtRVHgwPfTN13w6T79vv90Nob4
8PmbCBhVujp6gBYNUpeblWktmF/o7jrrJ/wfKsRZt6hjMiT8sS2enMPwbXrWzcfCoIfeykY3Glwv
jBV2A9YJAkMPk9aC6rNBhdpbq9k64GC5FpVKSl5To6RZPxsFSan1Iliot5XYE2Ad7fZpqU+iEDCm
b+c53d32EWBde4Vaf56R6XMslJOtM4/Wc1RluhEFcmJ6FGg0LtDQLzRhJL9PFenoxfKRUcUWvsXk
aAqC10P4J2+JZAaSdgO+aWpmbknSX1B7/UxmcF0wUDa4PhdPGcVdSFm8UMyZpxhOr35mcObVMapB
tW7UHKWZvsi+nGssPd+EQrINOri9Kc7f5S+qJ7z7L0LSxdy6nKiSARhNvsNMVbWmeTzTQUfn+zxY
til6WB4KB7Mj2M3rlPM6CWwXJ1iKxH4uoq2q24jWbnuw5o1XgoCPm0tFfrq/Ty0rMGdarAKSXHOE
9RZpUjbMGRkbNW7Yj4qGJoTUrPB6wS8Rf2fkvU+ZUqQAVtYho3WdHjVuAVqk9V4RYWI2nECS4FtH
rqLOSfHH6semKrLogpAgZ7lm9vslDMUQawtOcfAIbTs8dIn1IrJhx3AkXTKiMlbhfEufWKAh5+aX
nSeb86WBJ8tCp8uPLpC2dEo5P2jZBEtPN1plTDJXJCZ0G6a/HslDbdjU/QDtxzYYBqAlhtAW5y3U
aCdwTcMAxSv1QVIE8foNdXo3lCBuAk20cpZbfqN2UUhcgLprqSq3mhKSsWKH+uABkKPxNCd3yeT2
Z2/wpKW7ngZNAN/RIoDpw1Nbx0YYZhEbCyMgbuhw/SbhdSg9W/uApo3ltMiXdXAOmKiELSOvjHxm
LHDJ8fKNtarC1FNR0IzzNqpmghuL4My0xuowwXgiNoFb7oRLONe1k0c0vRL81j5z822G8zCrwKnc
raXDyfahVS3LCOnpWS/VP1If6Lda2ayksSjbcmnxNGgvXV7VUksugdSbZFUEy8+Pe/3K0dF0+IYO
R0aDI5dZMtIVrJhRTdrs34GdnLrmSzgAS+Xfk4s+DsXUXddRjrUeTFV3diQ/fhZ4PwBuixobYf/n
MQr31EG4t/f+9vU9D18mW3g4RO9wY8wAZUoyEuywtYQJ+fBudz9XfxoNvjNRKXoUL0tdGwBApouh
sQbZ/ThLIfJOpFYh0fH2l7bp7pJMfdboX2S+mfRJ9kudZvK/LtTjFGbeOHYgR71t7Z8AB03mTcZX
DTqm7CHA6Hzlaf11PMOwKWZ9RtX69hI4yX8z1ypJ4pBEDF63oSCKj3vSJFaa52wjWEmvNk35XZ9t
ZIeI75XQB79GyShnV7TbtJh33Dc71+t+KaEcnflBbKRdVI8MgSpHw0nb3wsR1AC4yVfNUvvV1qim
BLEgV9fzGcjj0XPF1wjuZhQbj3xXqEyR+AeVXCURZZQhIFykGefnNaRq555n6Iz2Rbl3PDzuXip6
hxBuOrtrpyeLSeHHuSDL+WlHADnreA5gBC0DtJOVuDMoNnpUJJULdlQ1e9mWgygBVVtPe+58Oki/
tzIa6hHZOC0C90xcVZMSjUxkIUWAC7hQnCSabMebfKhNDiwczS6lGe/dEplCjHmKvnqmPFsMuj8e
vIXD9DA86FftiFR6D1Gj64Em/BZiDyISaLyn5tHyfZvr7k5RfvE0F+SEbT+gzgLmytoEOOSIopgT
mSLWBUyzqmridEtJo4vM4/ee8STrG0LrVwnA5Ojc2kZKfvXIygW2w7lfC+Ryy1siX7pkP5HDQGQw
Cfznvv8MUgfykQ5cuTMGBZYK613Nc7SQyZiudT87PWbeWzTfdnl1UqjOAeHUHUhEea2H5ALPLtl1
nWjV/T27yuihKaWS87GFe3+5L1I0oNu5B7fOY7HVBi79pD86ht35R10oYrzt7MyZX0IH0C8z868W
jXa1DYt2fxseYgmZTsx+ui2P5RA45pXj78FWMINkhJjiU9Fh1tVQZB1v6PIiUBtBW4kQXIO2uNWR
tQ/poVYWnHgDti0hPQ0ju+dlOTgIngb/nTo6YxLfgni8pploGRzuAc/CvaXeM2OyxWYX7iFtnTFS
dCVGVHXbLGkx/6aKZrIeM95h7bZ5STKwlZwg4bAoM2JCv9RmuwB25HigXdzQOsBzoUIaCzTLN8nJ
7az0By8bVdeyMBNZ/sCNeH6xsFZ2p+0qapHVTNCqfhAeMvhJutkL+BscWoEgxX3LsEj2JD4nu5u/
wxW5ovs+A0EiQFJTkOrk9qEcfFGAw1Re7FdkNWhH5DtBBoEcbXUpm6EGfI4iu8RLJCc9IVmJVV6S
gpTQcgnZVs/5Ntb9y5rgbpLjLZbJTF6nrPfHZU9iloQt/PtmD5gmClefwXKvAKxk4gEY9LiqCpHm
qu4CQjhniDXm1um7OuV6jl0LOHNvfU5JHMhdJ7hP0HbmcyyitJhQVClvmzZBIHKeBSKIX0x1hLrc
dULpbPrLKFE/L5VLcR31VslTzHmzA4c+OGxm/SJUyRQOZRsQ0zRU6CX2NNb6DC3fkUGfMRlv8GHQ
5oNYs3zevpXwqH8wyTQdheofI2a7lTTEYHeMjWwiTka6zDoGYEG+yHjB963oBVBeaP1llDHXupP/
VDk7XtMrt4lt1MjZnRVCnHX0Hb5sVC7K0CqXQ1fe87I2stKKfD7khBFJBDL42X9AYO1qWWUxTOjv
xyZApkXooQ3/gdGnjr4LcNFtMx7UVeUzHpmiYV19W0QyndG0oQRvTvL4EaCrpMvE/DYGRCRa2GjK
C+K8ix6qmGKYpLytDQtVgAsT32OoDKeD0LBQLzabzxrRc3vfGB1THsqfP1NJ6PBA2CtdoJsc7zBG
Eb3Oyx1JkE6hGyWCfd9W9W4/mAsyObnvn9EljvMgt6Vb/t2DPUl4OtEMwTrpjH4PTf4w9d5Zin3S
ceOvia2tSId8MhBX6rcE1Z9lA3nSgFeCCbyROFjLX4wzk8FdoKFVSEOE2Ia4+BfYviDs7E7J8DQu
sFJ44pEmjeXKrLQuO3aW6X93isuKSFYNV6HuOyIV5URvfWB8+htM736KTA7BFMpHAsimjirGSMte
26oDcWlsVdvMlcUCVcpZ2wsBVpXEPVRUWdjEJ2hSd1OIj45vsG/nn9dbWtwcxoewdPSZI9Lxl/nO
cXEmA3GyRx9hm+8XGflatdtaj18kvINoPB3hNpA8dVzLk/5JMi1CDM5stqfjDZrBnSiie/Pdsdrd
PrmuF6a6DR3l9LsErLz/NdMiKKLCLRYVOKSA24HE/hRPrDjCXwjU1rSPSUde61cxZjcoZ24jHH2H
T2IK+L7B1ItsZB2BWddi8yvhBn00s8qh+DHqHUxKN6pKQFy9Jmv3EsT6bsCnPbPHtDYPsCcAqBlT
3p7sSIbymBU6Xy9zA3xmBsmUE1DfgYf3L9dSeWRd3RSPKRwwaV1aduK9LRr5GUFmeMBUaGNcvr6H
RaZLlmOaavo/SMk+GqEGV2RKOkUaKiuc1lH+K8s2R05zICZi4SUlIrmUHFe1DrN3SRZlwmLGkP3s
E+RLoQVvghCEZ7Ih89IJYn6K25TAP7hq8Itl8MfA2qdMjonpX90n/boiZ4CtRNTJ0cSbHZkkiet/
i7gAejt2XSEwfX7D/30F6oAyhCJ1jXJaQ1zPe1CBlJoiprZpY/t4TZQ16UM4uK58OSnnTJV9VA7v
1lFL/6/XZtFNVOAMKYWu410vj3j3n4sFOaa6rRkKyFg/euOvYSo1Lq5VskTrSeWzNvyjR4Zk1I4k
ATiDadc1+leqCW+LHsetn/yANbS57N4nlA3EFmJRFjFzXZou5elGyM26UHFE+jqe8aLxC0sZsoMu
mGmrgES+7WD55KyILaZMy8tQt1Tw2AYqFS0kUAWTQpBg25FDFsTWy5sn8vQ5N0IkS2J3HxO9trG4
Wl2nCr7enaMDowWPhL2kuEUIb8OdLlb9Am44aDbrdpulj7Xg2i331frkED5QjXWS3ZKgWv/4bDqm
tJNHgTKNMbmiu6qOYSxCiLbUip3AaG5vQDSU78U4zrd8ofyhy5GV4iU637P/p5WbCN4EZJV2apMw
PsGVMwi5w7Z8Q/OfEWf7h4oJAfU+JFDKm79YeuLwkWn2UKrXCzmtE7NdaCZwYzrg1/0ITTSUTf2U
tFdGs+cqeec1Yz0+Nw6ZMH5u0lhK8qFrjuSaSmumTrwtBu7ns4F1frU8lpLYMIGyApDS54Kr81zR
qg43iIQ1dQ3Ob15TfhkFAJPECW8uA70GlMVlqKT8R8dNStifpDwb7r2qF6hJft2uRDsQuU1+lklm
gUL64Tr6q0kaiH8L7HgRmtCQku8w//lMf0t9EIZD+/InglZ8/Eed9yQhlsVy3toesBSCHyQnNyhx
IPHvKnF1tuRkMmBGnYHQ9/eyCffvki6PxE8h8T29VByRLyorX6rUiJ8Qli1ud4DqQCrSTN4B/0ol
w+9F0ezdG7hAzR1FvsrEpaE5LAUPlXERLqWZy/LpWZlXrekqEoZoMXvqM0PF9vyvhAPysGyLCxjz
miu334dCsoJfjT6IkbeF4ZBvD3zbFdpdtjUNP9XZJqppcWOefVv3He3R9AuxTAlfgjBGA0cSLMrF
P4OVGtu1wbw5hEiXYBuwW0QsppcbG7QxrIDGangPY+nhmNfLPyETUZEKiav42+hGHOVt4X4C4kOK
y+Xz1NW3KMmrANO1Gip7SPBjUUeVeeYaub8DjHfLY+kB7iQ9IaMb5ZOjMgaoM5GIOHh7LkjkYs6Y
t9TU5RC2x6Q4G5Z/0pzwI+mlZ6n6wH2o6gGakio7LgGs3pVzFXUQMAfAUUgY/e6EQoFZPemPNRlm
Q+a1WyngqdbrNPTlfq1EXWiFcK1AAAWDe1jy6+jEAr4HIlHYFE0Uelb/9FxAlurY5coxXWslGmod
J51NRgzAYGsNr6hyM4CQ1HPYSgW2KgruXTQ0Ol05X1RvhxC4p/KBvcYv17ICcU0FXv/l+buLPULu
rKGhKtgkJqUvCqtGeQB2UaFomFEQRPURw+Tl3LIVUtETqt8qsqPTJ+Y2sp8GCvveTidU7fRJ8TrF
E8qz4CWWZTTuY61BcydfCup6Xhc7T2EzrrcqMKgUuCUKliCcwAAWHxTcihY9ez6QHdb0qOU1Kz2x
yZRw2XGOsjIUSvP/WPFrSS9YedXTPJkh0JV0MdO5jwTBb4SMXhlbp0rnelaAqjbnpbuk7UU5zSW/
SbJ3c33rbNfm02pca2KEtp4/i8+FR+KPxk+URH6fKNz5x0x+k979LGVAwgXDeUl9dN3e2D/RUg2Z
J3I5KlYx7H8GxlbbBPGy9ov11+ij7oGgAHtM5Zc3VdD5SSnxgg0Ew3RrdLLU5FiWRuNruNUcFAmT
2SrGxYQEGTglsagaHFq/OyR637rGhLXG6PyyBW2K1itY7IZYtxbuTrUA9j5PjQ3I+RRfpT0GVTH8
0K0NlFuWNoCLsYP9HuQXZg7jQnn7AStC0I94meY0SobHbEJP5vCkIt8RfhGiydAw9NwaAnwz3D7O
Ew6skqzUq8k1wFiouj7J2RvEjaPfpbbc6YkE0GQAYCCwtAfMDJZMDqPAH2s1Kor0upya/8Luas0d
M2B7+OeC9DGXQb8d8vuC0pxfxV37sMUrVJF3NbR9IpgQYpbcoeybRiv3NykTSHckVzs7pl3xsZ1t
/Y94AlPgRuZqU8rrSzWdHSAHaXlZsHqojoEB3TB8TqF6tv3F8toMEC8a55ds+D4Hoz3VO6CnTH9A
EMQJtssMQEeDa59teKqnLA8IQCNNOHknVwXq1JyR3d494X15Ec4rbMtTIEFmOmqIBhBo5x5eKawX
dM5Lh+mFpoP75Th9j8XsGZqEawzXVhyOocI0re6lYKI4WQUxybqDP59/vflqZ2DHa9Ul+qExXaoB
EbjrOCRRp2Oui9rEGmqw1MrtN+GsNwnomjMEpXmpnF6sc/wMfeO+9MUQaiGggBnrwVdwgNNGXcT1
DHzsbemmxzQRTbKOpyjt+9Dhv9dpNySIi1S0bKjRrksIi1g1E59mClnqPpdzqBdLFjRNUcIlVvfM
Wj4ZTT6VwP3fqEX2V4+w3mLO5J6BSctI5MvCrZ3YgUlBk6KBTfNin58M2YvPq3NUsP+cUZNWi6FX
NBnANumRiQq0J9uIyQg3WQ4u3c7eI0A1cJEzicH1Ff9Tg0yq6D9+eXaMSmFCVYM0cfVOuZ0BO0gO
T2E2/BVmZmpm1/rZhm5a+D0mrzRFfABZP6i3hRYu/DND+0UwSwGU60DJVaFt7H1T4fPc1b6k37na
UJ49piCiW3vzV5Be45L8F6ga8URxix1ZBaYHEFg6F7SVHqo1rlj+aqhDTTSdvbz2CX0936oaGGka
WhiXMD7LROiiGJBG40MF9H+2XjlPssbyJP0+662mN/kfMd++almqk//oE47zhS64kNH/WJjKbEQ1
GSvzy1laAfoKEYDwV9gQXg2pZK4VjEr8WhwA6V0cARJHp614FfxkurBbBGvpvmfw4V39+Aviptxa
XPf+warI96UagWHCOAUlCUTui9Gb2eANp8cVps/QPb9oOeg5xlhUavPJ/my9Whe3E+BOyulz7FKi
SM8W8U0OIeYCW87q5S6OTid8sZxJ8gArgbbIXnyH2TI/8qQVD1CBcljF1DVv+Fei3OPLaFWd1a5H
bDRP84qcO052dhzi2MHWzCN6aGdlNG0I0s/KizL1YomLFzHUPdNhp+dDJol7MyvDTUjofQv1piw7
7jDL0oOxS524gipdObNm6s9a+ZfKzGYdow448xpb08dDaKXfhCn+Vo3vyLLoGg/2TIQPBMaJk7uy
8EOXeNnjdtf9mS3SY/7iWcVCA2N4SYgf6H08VYqE94qtDMMSa0nvwPSROYDOHpt4iQXhNoiJ/hgb
DiPyy2Necwq78pVyFcMdlLNX+V8X/rL1UcK7ZpsViJ8m7FQQ8SJw3fKN+3/AKyRUYQbsh2wiotdY
+1TYYXkUEH2UiFcvTbD62f8dWRxZQ9RsbFoTzbjAEdIee4sgZhxeNZpvaUJecEeH9eZvilYPyQgI
EIuGzexzzYbqSA9I3uneLKr7c6k4hh2Cx+ThEYVkgoAo+o8vE1hxFosQtjw1Um+E9K6cibMLSaDJ
25YwMOXtbKMPbKCXAZ8tyb6iX6msr9FvJy8wlSQG/jC0m8HwWf9pzX6hyhQdlvtMvfziAmkz3oEQ
ziS77g4c1hXEs0QaPuuqxvE6tj3eRpfQf6320eBZwx/fyKXR8pTNso6CoKy4a3r+wuu5cKIpd6pC
JfxA8mscNalDcwENLb1q3dYVNTbFxL9XkawIhNMRE4w+Q6dHXVOsVqDyeWc6kyPzdA2wEeV7O23S
ojQRLfbrXZFelc825QnX1NpnKBLW6MPZcdPzVq1XkY2A8XCFnGHT19gNVzg1UJr2Oz612aMOMFJq
QGL7OtBnzCFXHQaLlxYoVxg+gOoofa9oQ3FevH53ECnnBYQkd+YfyQAnT5VIcZOLouAED2kI3wSM
+G/f2HxTnTAETKsLYkVwqli8wsoxn4ICKF5HRBOgwTH6/zk2kECsLxFjSPqD9INEUoK2rStNALo5
URoVRZHoRwAU689H0woub8Q29uOITlSOVaf9FfzDYPljZriApicg+RypY7ZnaIgru8jw7m1wLh9V
Iei8ipPuOnt4M9kwuheOqTmxnoSOkFHKgX7YDPNId8hBsKgHulXm19x4PqLnDk6OchXUYxuiCOor
v69SgDEE5dLK4yRoZ5ILRWEzWFtmyjkrnvwQjfGFvUtOYs1fbTbAODcqO/TvlRBUoSD5TB6j5Oj9
Of9ayjf2vqfVz06P5IAurVxVxOpPkaFvU9JNlJe52dLCfUykObj9pQOUVmVCOvWIBAIcR3U2WnaS
LBqZbjCxybycBVo+SsshhVBlIKZpKhS8Fv6CU/r2AncLBlhGewUU8D6GZDvZt0aQ5/89TU7k/jOR
rNR0+tMVpOt0qM6V63L3/5xYGZv8ZRlCThVrboOS7Wd0ax/UTxxxhQ32Lo+6B45kXlbJCJcdErjx
/7mtMg10h2TJXlx3Zqp9vk/+/gfhwpNe31pEEuetZTBWZSix3xMxXNeEbssBdH5oRYSam4geUku7
VgOihTheWfp1b6QwcXcj80OM+joAoBu5E0JD1aR+8jbS2zV2tuNEOSMR1FH/s1qQH8PoiXuXwQg5
jjRycxdGB5bOON7jiK3mEbr9NwxphQcXnftn0UdFmdG/H8v9nDmWuSymAnqZZhuQe/0KtPNcEf7c
4RwRgmHYewMxJWPFmgs+9ixy3PQgvLUe6Q8pvI6ldu/zACsJksPPgWVbFywXvoNL8QdVSghLE+i3
RNmWq2oxzduPHBssur6VyB4ztN0y3AHXIUOCBAvDaugNy/d1WNLlGV/vtyvMhj7Qyl4guAPilEU4
0fMJOrN2vQADF/M6UaVuPRzRlKKIM/M/9XVxXoLCO65++aGCWYwqZTwti/jnkgIwZK8U3LnB+P9f
ZLgB+3ogenlbl2A5iXeMqiOyBKdv8kS4tHYgOunsbxKz71qZdkG9UBTgmeGVm9Rw9qucJGlGz5l7
/rXaPsTUwzF23aln2cAJIpTblxR0q5qXjyLfCZAKu5LlWJOxBPb+WD3LHaqjutDA93YkNwxjBDti
a7PP8SzS0bJqDhaP4DI9xgcjZiV55UTVXyoxsfKh5cryELTSj4bDNyG6dB6hU62o/rljPon7xisk
vVryW3NBl50k/dTspslmsiKqcQJl7b1kwd4C5s7xbHRWHboZG7hEAClSfQHG7fklW0m/QfxNuSvT
slhHHSDkBgMp3unu015U3rHuGIaBNvyXAzoh+DnG6dDXXN9s0ARW2Y1DYjYZ/1k7i7O5d0mmEf2a
mtrSEORlRwEecx6CaDB0XSbl9VdyDPCVEUt0GIvWy+8XPLSTaWg5wAByTpU76jm2DoEwbaoJmk7F
hGrnWzc+N7IF8uRVe4ZQkS7VA8SzDRjXL3aAsWFTBWIzbFbY+0sdKYtE8GO93+UAOakldIiapbvj
lgOPJVtp5KkgZReNfiQo+HJr5ThxN2oxWMFs+DUPiQx4pMnPsYrWCwKwDQtseUAXQMA21xMiu9Fk
A9uUke7rkzvyeFMQ5f/oVJW344rzlc7SP6Efl5eciXUlXtdwR4OjFeNYR/gL7lJJc3kWjbVQ3Lyz
Ht3fcNSmdS7Gr7HhM54JL/ZUXIw3I25RZGMOoVoS70Y2X+cn9xT7upEW3KWMTzlkvGZyJ4GI7OEF
Wb9beNLJL9pue7ZU22bQZL0bMg4u9IoGMtmzmYPx/AzPKHNiWezlW8kX6ZVtSKoKJiudbSJL76uh
FALvwk4xUnWsl9si00RyHSz0OYRcRoy9c0s4iYDCno8Ne5UqiQ05DIM788x09z8KefeYQ8tSBaui
Iq021bz81qWwWhir9PFyJZ0NDWN57L+ClwEhXSyHwKolP7nY5wHj6gV1qMhZZq4r6lba5VN5WjOv
Gskz13+ebez0e1w0om/IwMhFRw6aOGr3lqHwJD5jzfcjesnD3jKfe14ZA1Ksbq7r6Cwmf/tsNF8h
41cVHhE6mGbsHgWr4BUw6P9OUWdiovCakTcu0DO6bliu+A1SoBCztvRsmStQn4+KA62kZ3ddkfj0
kESykSHi6g7JT06iYC6Gi3WcZscds/5B8bIW+VRfSCIy6ZII7VDWA2UPB0PWHZU66zkCH/cbc4ED
+5RLcxNnjV3B+UXxpR4VWKqPnynJ/CSW5GTZtlwMoJnzgqouRdyjkhWsJEkqs8EvYvhEYrT4KM/z
t9iHTgDzn/39VhPA0rOrKpQ9s28x3aLUCWlWvJS//6ViPk3JyaX+Jz+fOjsxJcRxjaLpPq9dhQc3
kAqW7xwxVrZIlASEu56GAEZKvnjYCCbO18l9VRIIDfyfsZDZYYtXqJFBefRPDMS1cpag1XC1KlVs
rPeoxVMUyyORUorO6sYMtee45TsiOjNQMN21K4YBNB8azNBTUnVm3AkbEMxSJKKUzX28xIrdtx0j
Q3UxjUJPG4kbzrC1f6uhzSFuv3wdMjNDIC+Lcojdy1A5mfamMvQXDRgMkfnbX4TOaP+EI1kjCtTT
Vu0PSdtWF0nGEVrxuKMzZs08myIWCofZCEM8+RDgA5mF0vGLG/iyfrsqRtECICcV2tmYNQDlugKe
KyuGjVZUzIj3Xs01/2MzazoxnGPRhZwiLVxTiqqYaXDAaVPnJudNNleosy5bt8kjvj+b1JuNDdgF
kWB6kJFg6ubH8jMf6/SdNFuGa4f7jMhrfPhE5y4mxkipKYVFkms3fcjBNTPY5Ij2JMi3JT6PgQXo
0nmXtKiVLnQkjKYTSfIH2Ftx5+X/hYZRG54Wr9NfhYBOhfHx8S+J9w6Rlxft/9GOSIu+W6cx/nxV
BzbMKFxX8vxcjfwBAtoiYzgqMa6TFpS9PzYstCcBar4qAy/LJrzbZgqIwNbo8ZHpBqhXrnKAcabg
lBMf5nfIsgKAVZ/S8IU3SPXqS3OvKmWVVgNfv86fB8+70ZD9XgUKcM0d2eOaRbbe4UUkQIcZXaxG
nn1AmBpkzV3AakY5hbdUNU34TVgB7NQc/2721zp+zrVRRcVykCmtH4JsLGKGX5DUq5CRy+oSMpXe
riIjaGzQ7N7wEG1ibP6WezG7uLMYc+IvttWynyN4iVdXFATUarb0UlXJVOymgvAbJ5eOyxoFF8pn
hpYWeVw03+C1RmoTY1VNhFUTi4hmLXYeaSC7ENP9DcstZQafr1gZ2YLkgFfy0st1JFKVbXdowQNB
Ui7/smpM1oogSy+BHf2prncwFli4FgovmBxQE6kNf9JFsznqU4GRRPFfSqiceO1fIyw6duYXjZX+
Lc0WLled8L75ZAHa1RvtDX+EjDJ2uMjJna17ttL55zdQ/60RFicHe3v6MstWVHuLPLpkzPfxOUl1
jIeqQcBmVrpHJhUNSKSBHR83kF7Z/0werxue42g3ISqDInRMybK2QSSGf0DhdUqn5Bjh2CmdfWaZ
lyGtC0NiE4sIpgUYtAIcNWTE1Kymql+vEl92D4JOYsToOy187xProAPfvCfJSveceEowHzAyS2ov
YVOd1QPEWKapho12U9o+IwVQEZq3m7MopDtURsGYfPRsT1s8CcYclOcI2EutxP2w+kidVxkJuIVF
VjaQTXZpC/5kB4fSYSGdpzi9URolLxCO6G6wEKkMftkD7b/0iuRKjsx+3AJ9vDd3flMGE2X/y66y
OMFs8PXIT8LCJM5yzEnjXCo96tD86iSBWE9dOH3NxNOd/zoxoFfpFld30L6Qi0uwtG4Djn3YqtkI
nmHbb8kAvCWE5HCN/QVN3eGp3jAnEbbuFqE4dE6BLvDHFTtHieefMksCTSrVyeZ+Cj3rlChHMFTd
iT3Zbl7Gm/6YHkezYtv6zbP0j2By+eA+c6JC6wtBRzbLFI1AnUaMibEWGcBAbgQw/4Z7ZxSpVnMl
di4Dh+7PG6RcmcIWxvAHQVA7qUmSU3Wtlt9r6pOicHQdJgk6OH70xOV915EAXedotE73SFHBOhh+
94OGcBZ/LQ3+EWmNB9+UjvV3Nu3k+mSlbOBrHB/5rtz45U3IBiIV8mPotBDubmtASKqeEHM3bxlG
LpYAiPel+HuyKE/hSD8n+5UGIwrM8TxHAfAVK7eBpSksrU6VLZn/e7Sc/nXkBqG83nH653A4+0Rl
U41IvNvH2DkznpItnTTTbyoJs4jRBGdQLf0J0NPw6zdMwQtt8iUCXsmajvrEgrVybTQ8F9tTEslh
LfOJiNy2Sacf9ulKWhWuwijP4j7D8Iwb6VriyU7a+FWe4x7AgZwXB0Q3iMVcHJFPq//edzaXTojj
Ro+nftvHeMA6Vtt3m9iiIxka8TozPpDa80EBIbob1XvP3QfMRfPEC5q8+Hkg7Y22W1La7MieKIb7
AqHDktz4VoQ10+ikqD46fCYPSTX2Wpd3Kbiia8EXBcrchv4+lGsFXFRjCWtDtCWlsujZWchFb/9F
bQvVu6rTTDhlORBRkE6yNqCpGg2RHSpFcJaG5U26N9TuayP+E1Oe06sY7zD3FK4MjbRmQFc2JRsK
9mQUMKbu60GifLAvspmvpl2QKQCLNlcRM/PhiUy4P3PrenSkENMWhjccz03Qq4ptLL0xqn9eOpKX
PIv2bbh6otD1J1+KZgjlSx55NEdpax5OINBthFu9URrtaS6sOvv3k7DoxHFNMXMG0Eo/gUnjaRH4
KR11Coc6v6zlOIE5jhBcCWdqfUfRjGTA9WqMGuYYKMSrvANswtxOqiOzReUrI79zjm0icYgO4D4b
F4JnOhv3v9ClmA4pXOsHqu3IIb4xsQdT3EN8GdUaoB5nqrWwnE9MaGKh/S17/H3w6mfNSCirX3bE
eC6imeQ31vxYV8cRdL/hib8Y+gAJXS00PG0qBqowi8Vin9a0IEv7jJKLLTgBPp89+zf7HR6buCGU
TOgPkCfqvrn0Oumu/wRaclsoKFVXPivTiVWvzUHcmWNvH2zXpyzFoRXb9pftQ8ZMzYJjDhnUBumi
2qkZEzW7Mdat37oVyiJVje3e6FO98KwYo+TbU1bRnCoym+u9W63tPbN9kYf5hbOgNo4v0j5HI5PL
FjdsrKaxaJFJCDeqx85HVzMtLPojARicxaj/caMwqkuXa0M5zOHqFMBwaqNywmQ7fZvIdQtg1Qo2
n33NqNbXx2AcYsthOMye5FRc4Mn0YP2QAgsUTCDekvPGWFMd4Bfk8GCANBtEeaRV0WjZTzAo6fVb
Gc65jz/t/Kt2QTQK6I0Wr5cUWsIUTakt1V3ClVwF4rm25U8gyzeWmU9rQN+CDvZfE3le5vkdh/64
IdnAxt0tT2eFnvoahh53xfeBPx3oHKz4/dN86clWq8OYflX8d7pT2sacNTv5718rKNUKhCmupliV
SrIeE2mXtBRvHsq5niFgSAkIn25dQ1TFMLv953F686wgLoQkyWPK4rNqFaI0beDOqJKcXJSay/kn
/giVpyIVb2DzEbjC4pmjb3lYmengnj+XJa5s3Evbn63Oei8A9jAxwjFKTxAwvBdWY23K1vy82xVC
9TFnJaD4CbdH6oeQ6GlorlUO2/RSjBg46VlkPmhqGhls5pMj9cyXauklKoTdYCVGZjjw+26o0cpE
7XDiwcvauZJxQOl+/NDhsbw07x0qvLWkmqpfZcRUokjQzLwRcf0vDxy3tGy1AqN4HD8IHiZnv16m
SfcfeRfjhbxIDyh9it86A3KgYqhZgPCIXA9TW2Y43D4eWjsGipz3OLr+GIlBE5U/nVapV41kf1Kw
YTYOOqWEnTuCHj1IxjyYbh4TzEnGRwOh+/e2hW997yJc7SIJqERMZcACX2grpTxEdY/VXIgzra5b
iJmSVmxaXogDWaFc3beiDXz4FO59qOHaXh835uKRnW1tQKUWXccWrX16NtFQxYDPrs8n2ItXaw5V
NB/vszQbaFoBaxz+B1ubWX/3Sux36CdTRUhZowVyPkSt5EggVxvvOhFEUvIS8PMAvYOLqdVz4hRj
FPSbYri9gdLfScWScgPz8yYdDz2AN+WutRu8BKa0O0oGYjN3Nr4jwG8dIAPvQxazynemuNePoJ/5
UF/rjLU1p7Fyf+W1kPty86mJNUfQ8I1wnbKTgSzOj9A8dg8z7OEAQTUBE6a9i5LC/dY0dcjP6nTL
AbYeuSZU4FsvG3ZATkyRkwmIsKSZQYrrn7kXlKH6euXJpqxAAtcBsdD/XakdLUfHjPgwYZgNujWN
L2M0DeanctK4anozARcl6I15V+DlFl8UrF2tBScPY/XTj+9wO5sBgheCYmJtjurs1b50JE3uBdLD
+3KHvnfceXU4CFT1RMf4S8hW5ce2s0LKsnzVYOYkCf9PNRguSpO2CK7rfKYdI8/F3xhf5PANXzHL
Wwp+Jox2bGMhwBPKzi5PuUBqltUDKeY7S7FFy0r0Iqtqq6WeZUplL++DUUECvSzxagRxDtdC4vX4
Etf0PgP8EiHMq5byJVVa7Uwk2wMhOoa7XU7wv9O+jNHjFLPZotsQ3xAitNJOnLC5jytGonr7zNyP
XMxj3WG2LDUV0idtdRWiZ97s/OmbrvWENxFrboa87qwPXZnEYuPVdZK+0TUqsEfiZiGmd75rMP+1
LPCxNcyaB+xYahp1nma14MEqEQByPqq4dnUuf/nNDHeZyOlE/hIfO8XNcAeSVhbTByt5eJseGeKl
kwAwxYBBwQZ+pKOiNHLSlkNnuRz7hXErjXG30FXe0kJLtFiuy2S7/dtfKdQ7I9OVvfuRPuAgijU4
p5SSVWpNzDx1C4Xqloe5LL1XeW48c+EzToj6TUZ9qA8TC5m7nXqnPGpPlk51l2HgEusVxmzooiIC
mCmUjx9lIpcmTrQPhhrDpKl0ZLqsC0jG609E4zRXV2WMxoR9TFPoOPmeFjXiibKnoTZ27jKg/jwU
lbbQfjMCHIv+ZX/oWAhDvNWq5aKVLlyQgQycDXw/xR9yc+rX7PBUsjH/jkaSqWjih1pE4MTbEyoY
sbBU6TR4mwfyhiH1eyAgLbc4nMqlLFilbsFsClMS35Xz1Zd0ec9ra9p+tC/gKs7CcBlGj6dcYHuq
FIDY/B5+onLoXGy4EbfRID9jnQrc9w6582Ua0UE0IxJt7j0qvjoW+LMhYKz6n+JbWXTUM3f42H8C
NpYnhKKScTAmdzW3WhnXVwPIXlfSDjMukLAZYvjVsTxVTaIEXwRuygQegnAAgNUS5XIw1BdN4NZM
qSq/luIHOj798/J1rX0N45Ud6DRBciTU6H72dzRvwxCwV81yC69a5gubr95ubBue95+xBVm0kBby
fanCQfAV52q7fVUm2f8gmPup/ze+vx284tJdqN9rPObJ7eJDxo56G6C/0OEIkrvdfWfoGnxOkcdr
dDAtjNmDTz97Z0TzuYxmmQmMvhtjx7yPqND5P5iB2jzYhmvdvAYTXL28AOgPc5fDqeSEC2Y6cG6Z
hU6l9D6O7G1A4lyjLbR9D+6czzvtBNDpSlECZi8upXV+qh3e4ZZ90+rS5IKLbcPb4699DdutlplD
o/JMWsh/QNpHjQf1s3xn8Agp+vRGllh7i9TpSGbbEMuRMYjRo2kyXL7MfxmzrOJYZGatvblbY6C9
wKjNJw94hXa70qimaa9dbm+3AliTVpJD3g8hQ+otlbwpCcGWbToNMJU+qECbGwP31M0R8gNkT0X/
8k4Rg6eESwei/MttTzXLq1x4ixyRTc35lGnO1PtWYE6A+jIc1eDSajkgZxk/p/TOYaUioC9yi5ZX
KDmH+XVv8wSO87IrrAms7HcPZ+KmFzY3XD9E5NLCUbDSWeILeZBtCTAMYDeoIss77VDFAWLzFrVI
+4e1RzxJ1V7Xs82UOap1vcV6GTWXMADmsXMKXGU3p3ShscOrEbPpchmZF6riCqoWEyxWAgMsgZzj
0yKqX5b56Bv6u6oonksToOrvO7E+KPoFnIXT/vnK52fhv9p7BanVTUzezTcEzP59TpCdB7EBt3aN
/hDr2OzMhTiK2xQ7wJpAay+qKNnBYowW5+6pJZyX9K4b6euDqh+2+eO6iAKNRYltoagdWE6EfZDw
BVRHZ2EI8sxKrRQ7e7FOaTc2ntIzva786OOuG72CZzmATkMD3OZJjKgkaz/NLlcsOzhLP/wBc1WU
KokCUMoMJ9U2PZI5xVULzHKya2y7leKb50ONVhQricTks1ru30I7X6dimYoDdLvk/iJ8ULscQZDX
5kvTHc/lnqJcAgh7FQ5dDJey7LkESeT+6CPcYpcxCh83XsoPOpSz9AqHrsvhvC99QdmqRkN+a84R
J9VP3bOyhjqMA92XQKzb2b+x4r2pzgBtsKDvg8EbNilmI8JkYy1qBaSSiXQHXhajlzp/P6NqKCw9
cww74pf9rB5dZ1FSzTkUEOHNEW1dCrPWYKQxxzDGGdZU6bf+FslQDcSPczI4fXd+m1oH+kAhV45+
AaQC94enHL/zO1aR/+mhhhGIEHkh1KhEobFyksX/exR5qd8388SKFQ6d/x7NH3LAtab+IfMpOGw/
EZEX26TGzKw2sbSgHwYN8CAP8zU04YyExD+iG25mL357efIsfyPwlce8IdGv291MR0iLs2y8IOb3
2VD/IOTQ3kVho2O8b0cjJAb/UfCosLP92yVPOxpd5o83auk4KpDyVAfTHxTVTdxe2bNwFs8yLQg6
4+zdg1uRPxTBk1GdG+tx3qcDOEF4GXeqyACvt2uzqndyAhvhbFbtfphAI/EIKCMPEv4H7PSS89k3
IB3NiLV+SDkOptsD1at1VyZ47D4DogidkfyPkXVAmYP6EEGablvGXdZZQcRfdVsaIWkTnl6NKlTt
NvTQwWBKXbTH0sgQvjJBQPJ70HC9l7+1nbE188vWd/EEOIe1h5TAp0mob81KFukM/2dkD1JjNKdq
YRxLejLKn0XBfyC7xybXv858ZGuNOAQXdF4Vq2eI0n++TLEixtd2JkTgiKMYcb0vn/ai3Pa6DHuf
rPafrhNUmbsp0xMCp9uSeLgN+eKU0C34MBtgo5aJ48y0J+X3eAOPZTLWUjxzEfHJSmOloCQcLFO8
DBv2fnJWaMvUmt1LoCIQca4Ivz0QZ2DVMeeTlEySboPxBp8oHmIrpMm0ASiIOl2FPcVYDp3EO7Iv
qVgroJh20UisSygzMtYa5+Q4WzHCdK2Po9h9bUMq+AnhXDnrOLx/FHhvibE8ILhBRUh00A6i2H5U
iWVYFFKCZlaYp0Gg1sSqGnL5GD/Pd/4XskJcA4WQCZtEmNerj6+JnZyM52baxc+EtROu6CleJUWW
wZ9sdZR4HTmp2mnkGTdfOl3sS4Us4KnxOiyu6/Emg9d4rFJxC3OE7g04gXOJB4LMfs3HscZc4064
K4K9WNOopEOZJLBuXUrFrmDsp6LWZxeteMSECJ1nSNtjwhYk41zH002YVbR0gIAcR+GZ27qTS36u
zZnU4ycZyhtW/on72vi5DWt3FvDRtI4LTAUBWyEwXfnQ4K1RQfARDtPTiOZVF149M2XhDGqR0Opa
L7oXOxiRDITw/r06OG+kcBavEjBlApp/DsNjifwBaKR/LI1HT6mJ5TiTT43YPL/5cyP7MOnsaWcH
Wyp1KPnvndoG337ETVY9s/x7IZ+o7A8rr2MKyQusNJc7Vi1Z0ddygy/5yNL89Nplp+XF/uBliF4u
vxuY/xmKMWxwRQ5cEAOb0JoC0ATgLBtdNqQV4NAYg3HxEOo5n8GdpdBhX4fsunowZEC0ZrfxDjW8
0sFtYZYxi38qVTZtvnQfFgXTjdzNerkCtUubkWeUcnQWogpaT6WwidI7SUWcbdDqqm7lji5QpEo6
NUhtoQ48Q/fds4mk7t84Y/A6jfy8eRNItat42zCf3R1yUwFS7lXEsGJPstuL0e0OPJpKWjVevE34
JwZ8Elbe6HH3q/nUaB4ecsqphCp5JR2DNIP3G7FybPw9gOI3N250abpyyb4YJ1cVL9NxANO+qStP
9O9/AFxWOoTdK1s2sCA9eyvzGG5jVY9/OGFaKqw3KoGWirLKKxCclD7ramt2O8ChfrXfPbtTrG/J
xQEhQAv498eokfdaYdIEA/waCVybekm+V+1rG43+w9ZIYYKcQpGoct6KcwHsKKefqp+UAK4xdJWE
zNLcsTZ60X/h+2u+JvPoWtExvLurC7tmD2pWDKLjRZY6YaiT2LVMaVt2kkJRAE9uTzvcqHQ6XYur
qd426yaK0I4hOdz3JrWiupQ/z/6c7uXDZnrPimJKyddSh3bvB4kjTsTcjCkJ/nMsisYWLobtj1lQ
Xgx8kOh3cyBvs2Xsl2qD2coNhER/CPhbRzpOtrH+mJWqsWCDPZWXAu01tYmN+CJJ5mCKas4x+IzP
eiGM5oBFVU211fuevF3ZcDwYPLNtrqBhq1m7OtN81aFa3KBbici+UChrF+2HzWLPQcyZIxuGKO6B
OuoB9Zw72okn5TbSMnYt60Dt7GCVAoANyuix8zp+ELeMu5vJa7Lr4+dlG8y0Q7bFWaHqBZxSDBpq
OyMOG0pQdxb47DyF19N5rdOIYuw8xThCfBapsppfEt1l7HHQJ44Hiv9ycIpeTECBWAaxK230U6Mb
2OplzbaRH7G+PtAjYhHt2r0HJPA2lp0hqhYGXqL7am/RTisUc6UwN36hgPSw97rosnNYzn78JXWy
iP0+xcuDLGMSPZuBdZLBAZ2tMfz1NH2ImxZ5m+v7diWiNAyHg3ivOXxVQRNVBAwJZaaAl9iB8zHG
nwXtKmhDrJkbngVSxcllWZr5fH2tF6SP1oyFiECLHxA+njJZo+WaJ5rTb5+RwzQHjsMH/zBK1Exi
/ndfpXuzotcpX9vi4Iy8F2Lrv/CzzZesagz/IFcKaEVBCFSm9Meq2JetXk4yPI78JvULnGh9F3SF
JJBJSE4YvIpEkRwmbN8NvGj3aT6PltTAbj2OCjKk68Qqwu0tS4j+BktM8OB9Xu2n+Q1d+fFYiii5
Zy0HWUud/tJgYOnKwaDG3n3H/K5sbOZ4/Tc7r9Y2FklcZ33vl9D6GVnQj6KIiuBR/OQ5ytACn7ig
DDl6HIe/vjEnG0SVb67g4RyYnIDh5A5MwRcLGSw+2dHM5yj6nZW0APpzkWpJycqWiTKnSKYswrTo
ytB1G+BGRVR79qwfebJdUgG4eVRBuVGfYXaKeKztC8K5yR3ks66J3jUrpFaqA2hb/S6d2AUdMLtR
iZlNlKV1xL5PQ3KmnrgxbL/XL7riGQUxwLbwho864+RynCmv113Je7Gp/bpS1QKEAkyUTd5HQCeB
tmCLxXoUMIWWxy1NGaiyiv4sEOAmZj3qv721v6o5M+p3Mn5QXOSGe56oEyC6u1gUiHBeTPV5tSam
Dp8E4BTIv/Kn7+BX1c7JbYk2a4NLjV9grryiKC7vnDJ+3TTQep73eKYFHPRSToCw54Rxkr8syAnG
8xH3wcQBZuA89BLQGU2ZVSSc72aHLeqHpVNioDrteU3X6iKBC7Uxq+PVhezrQAD2Q3qCulJcN7vc
erYUI0Uqjy5aouh9L+MDhofHp4SUPxG5vs41jmiAip4yueznu/giYI57gJyiYqYECTUNiNr/0v+t
EUKV/wsgwqWZhKG3ArXzehLMofMXxqcMf9U56TYCkeh45Posxe+KmqaI99ZOjk344ZGOOz0usCLm
N5V7vuUa43tDH6pSVuYNMW9vmyApbr5RDz5z1sCXOfgO9Jt8mhvJppwyGlkAKlQBOsZPXehZA/7V
/VLgh/u/485ff0HmlhJfNsieZBoxqE7+wjFEkwyO5eORsw7qxUW5eAtt2XSemOwvJVhcwemlYmAL
zCKXVWYwNYY/wmJOCfPYSUNSGjRtbA1R61TKQokxJPQdp0gkUgDjo+XrEF8iD1keKzwLTrtPf+7X
fmSERpYIpyS07stE/uGFIpZORu6mehYkyX7Lv61LNZJqhitb5HEeOIzi3EZBm7KvGbjl82kO0Gmq
FUoRnEncetMc34T/U7wF6Pc5XNIhi9pbXJeMoLTFDAhEj8qyX0oox45tMuLIzPcnZMnO62KlkUJL
2D7l0agS1vNbB6a97O0LhyDk6J2Px5A9DdBDvN09C77RiHh6aK72TtVPf9xmFGKxIOHdfE0on1w0
GLDJOjL7qKJIBfrFjMDajajNkxJaoxRSnvhoRrBSXQp4xZehwH/PQq50wKj8937YHN6BLSVtREhX
3xQfcwu9X6z092+Ce6514kGKOfc5lQ4vg6gKx/xnCD1LOVqJkXgwrbEPg0OvXpuOceojBlH5qy4W
8nfAFsunk08f5NxFbGP8S+vQtO4FEUfaJ2IYNCfP+QX5w6q2btl/E0CFERZeMNdBTv0v7/QtreMS
hb/56uD39xy02J3UKjOMwIJeTugbTVlhbwYxT/t3FS7spaFu+OV8GqJknBCqMxDAeKPrj5uljV1D
P6Q5jCb/ZOoD51R9/d/kqo54y0ec5JuXMDltMOMX+lodffz4to4PTX4M/YTg2HEZKsmSuc87J8th
OBtAWK6OHdEQPi1rqSMH59O42npi+D9lhCnUl+EentCfXMgu9sDpv6mzJDUbX94WZxh7kbpGf4Qi
aISdCca0rvVF9w9xI9jN11ZXLVIKOCQmnKVOQ2033PYfDRXG6GV5LTVlAsrb05AXbLtuHk7SKj2N
/EfxhxKZs2LYmYGncyfeJEw+1JfhLC2+Aq2ZXZjcgZcu4FzJF6t7cdg6of+ZXJ8Tlrxh/e9D/9hT
Du4tz42SbTZdnvIVoK3Hx4QCwzbAJkuATtKriSd/VJc4VaFDo5OoOq/MgM5ipoXBrK4EZ3Jd0Q3M
lrC66YIcNxGERSnLu60Jjcs4wmfgirBhfrWbOijKwum7VnGoBEYl5lrKz/bVgRCR1m3xPm2vsBZn
RAR0xqRdMrKvPRPAlcmQoh+RmmUzOxfSKfvn3yfhKmOpJO9ceUW3XTUHyO1pcfoG4NRkVgcu8DSA
xoG1f3xPNSyEA88n7wDfANqJ8ElcR3gX9HNBZQqWZFowz2JnGFQg1jd4MjTs9HHBm3hnf1ViXvZc
3n1UD9gogOyEPG1CF6ohMRhqGNASez8NeC6t5q9T5NOXcCC9pTT2yaKOD0udhxOOjJA/CKr35v9d
0o6PvYBZTX6ieclD8QoBcFIQ5PjQlyTX6W6trqwqxmWCxky8KNsZzLGkZ6NQ2pbk7wRCw5Yuts3Q
RO4+kjl9G1XO0EsRJBsKC0V8SmL+vtP7JBrm9X9xwsPqCn0UANlqnv7CYKFWrwkFMz/AJ0+Uf1/C
cnDHfgzpuSphX2/z/iorYS/B66zStu4NMq8ou09sAi0eBdYhdbLhEyOiAbfw8fw927R9xV0wjRLK
JCX3NLnQYtPQFuvo0D6o9ImM6MG+fatZBRtpiP1ntwIt24PcTJHS+/GJLx6by9wzYZr0H3rdrjQj
cw/ZsNUdMSh75oHTohDwDh9obMeEtoTcYzFD3/+REZCYQO24Z97JgQc/+DBXVgQRS69JIUF1o/7N
9cfAamOcAqTjJK9B/VLQWA8JrxStzaUbiYOJUk9hLWqV/1qzv8SGxmqR1SBq+0PkfM4Kpkyq5l44
t5EeM3TzjKuKR7lxb0ma+cRtzTNgvE3vHwJCbDaQjdt6YcpI8ovdNHKy6yuq351KAkGG3nW8ta2D
vT864hVpdoiCiJsEubxmPmcQpIC3iCzrZG1EuSbUVhtWmE4g0D2/2V0SGODSVoZa1N0cslZ7mXgZ
tdZ4YkAehVT9ZsmiXiKGfvX/niHdRIjHbEEi/SIDRe0b9DVQF5zQFMIVj7S63dscm60G3qygF7sX
6VEMVyrtjJ+cZZsimeCz8e6roOJs6tZACdDWVaWVaXH0DWLu77hbuR4u+I4nc5RZo7jEiQShSQS0
2+lTg+Jtx5baRv2Fqek1D8oQd1GLX+ZmOemLZ9rH2GQ9ILbV5DXR+bfrBLIM988JCOiU4mTH+TFc
/+VZxt4vyAaa0jOWgbBQpfrkHwk6zUvEx8ict3i8g0NdMEOsvA7sing60CXh5pR8TC/W3Uk16rGY
NIx8BjaJVsPgmUey8TQb1iXPGgb9CHoVmbIIM3jseDAJd80nfPUkJQkN9fZIjxKQnXk6whJfPP6I
j5YyImV340jApgv02iA/yr9DmYgK2lBSZRHXBqRQB6BHQRnij5LRWRCMXOm1mMeAeEOFEtdEGnlG
RclNV/ylI9m342H4+9JUO0T2MQ4pK20/OfR12UU2qRVYVl2z9Jyl+uYSCqFjtLDNQEID4ZEvBm94
duO3BAiYwduPvFupMqrrKqr/XgVdefQQf8PkRIgFiK/VkrtkmQ+lQxBkRxtjFKq2xDm7Za/39GZk
fkynFRG2uJ+mFk5q/CcNToyphCTB0vXCjoF3PpKq92yLcvzsL6C1i1st2FXBZzmsAOAb8lUZNFWT
HpRcV4IfkwQwxHwlgRmKmfoRv30FGzhYg7ZuoqiNBbmve67BHFZ8mmnb0zMSWkyDZD6PnVfiJsaT
QGs7ODP8MRHZdSS4ZQUA6K0CoGBbp/YW9aAmUBqcvDNyxIzw2nkybLUUvKKTlNhyw1gjss2wmV+x
Syq394h0wcY4g80OEfUXqpn7r1I5P5e51iLAVJOX9+rU3yNcDpAkztmVe6ABccbxxEPFQKGdTS5v
klkJFxi+4YC4znwtH3/w6zY4aejRjCmbtoLPFcFNRaRK0UC74GMejtknFsF+IaiAaIdE+THsQZWV
WLiP4hl9ZumM1OAcqZaPUEY3aUqcGKyFTrMbehUaEMVjCkaO/SYuZAFOdnjz4xU69bQfZnszug9B
bjsZfo0i9we6U4XUrVmC3leUZK6ap/yyfUNd1H6B3dLrvP2IaL6H4OCBNNKG4+Qz5ElNpCE8Wezp
dCiYxFY9U7WjoPQfxvLUh75pe92RGBm0qrcP32kVIoHq2HJ3n9/dgbOnw0suTCIAc9wg3iqO6nvL
HCisJ3MA86uexbfoL8D5NFjxbPYxldw5/1R2YvvlB6BiGaZbIFMUE0ikx+FxYcpC3D2bbwXlF1v9
lHMH90yX9U0QDuxwbl//YCajG05n1Gx+ELFtWn+Jnul0Ld+gqlFvzdUzq7aJkSXf51O7KSHcIn8G
HRcAkxUDQE8gRSUWdc39wJBO+uO8c5ymcI/kZTWmHy2CiX1e02n836sT5X2Ag+gwCK+F1ZeTSOon
YHwsZJ9vIYMLGXAKfAFIXs0Zs6WJ0yqd1hxC+brL8nmZTDQ4zu5Ss87VVH9mdVJH3wXECYm5vmJ3
WXxX6tLy7dL/4PQX/wybZrJWw8bBc5waLW3TrF3mqrumRxiNG1cL8iuG4GeS+n376cWEWMntP+Lp
ueIXoNcr7ROfmMBo21K2z/6iN9JCvdgV68T+IVwL3ixQc2umwXdnhnV28QiLqadwVpuS1ylWHq/8
Qo5BbvrcFIud/xI42s64BECumDeWR6tM+61YvzyF53zGrfglhvlAPharITF9W/Dr8e9ITmjVa6uS
oTLsSjLlmuBQ02BgDvV9DBy0cDu2mwTBxtJnim0chxn4cU77PjzzkpdGMM5idivEYoumzEwhGllX
1F5IGs1psw3Hnblw9lB8LZcC040uu6JbUi1y+AJ9EdV33SsWjUOK9I4YiHkbtdb/QMv+zvqelSvZ
hq+7vvad2cw7DSOJOASQV4SaB7dt/me+eT6fJmb+LQjrjkfJiK0VTuINolOh+Eh2u/tV+WRd/T/G
KhJNcJsSMTUXLHrd9QZiiihkgwOcVOlX/a3jPgUm7DcOtDq86C49i8IX8VZA7U++QfRul5ZFWvVl
8YH4fh9Nx8ne4fjEpRCTSEfFmemSiID7DX3h+bBUHOtrrdxFJRfV8s1JS8nxmQwHky5SQA4z3BQR
rOcUXNHJKraMJVyQ0EymEo5H7oC9S8D7eoqCrqil3R93DUuAd9SPQQiJvjIodWQL55UzQLtUFyEy
q8DgoWsZgGlhOeVl2pf12zzkCwGnfrod4yxS8dijaef2qM3BoQhyHRRQA5u4ZKc/mZKTgLg1uCCV
B7vfZXDgEAQURAok7EeVTiii0qPzFtPdfwv9gxIX8/UTcv4z58RvgAHXdyOyZfJiDTmw3Ek62Crp
ADRiYFZ//vk/wQ7J6uY47CHB3AI4VVkkK6WtdOxRfdaDBTaWUDwC3ngF85gBAvArs8CWYEJZ1wq2
XP43wJ5YQSZgUHJEkZ/hDs1i1n6UG6mVJEuSqoTViL+GRZVbP0qjAq2/uBirWJA69hHXsBo4b9SW
xHn5bzvavQc0a1aEVbgNSxgxDrymALW2dJ5nLWnGYdZbOC3SMz+ii7mMG+ImoHsdpmiaeEaY546I
fLr5jqPGKf2qqN3af0Sl5lZExeQSjFSbBsf32ruWUNYighhgVhLD1v436c0YNduuExHUGI2GzLlX
pJl+UiNnr4bpNmDvPmk14ltm7PW+EnW7yj6VVHsSxJGNhan1pKPbR1oq7/xyauYizeeTdEqru7Di
B9G34uT7vS4bBvIP/EC6OLCPnHPLkJ7IqsRVlKuzVzTNIc9LBtGsotCff9GsM+rZXgHIlGUNeGiS
fFrfbEO1A2Z0gn5KbaanJP0+CHXroQccJFQAH5l9dNWERktsDJl7RVG0yvYqG0vC2LTHiqq8hdix
lIEN0oMLV+xkQ16pBr2AUwsJPpRoJCGgnIEiPC2XrkM2JGutsXSgqQnN/4/rGfXz/kYyHkXQy5F6
4W2XWARrwiHohWqmm0kvDU8YLG80RvC99DWpDPfcFbpC2ffnG5/n0GK4B9ueFjAIr1BTCQA22tgX
dFQXAWxvbqQU8logWES/Q2HCfotLKBQAjib3rtovEbzTuGnw5H6hkSm9UYgY3VtGlmsSV9JQqtHS
HmZ1Jn+2pgBTgMGC6IWsoD1Izr1OEfzUf/OIoUibBnyGkcG+4j2UOZYBtjPk7ZUKatE4sZ9CFcuY
+v/VOAHdWDHjdPyL5UX4uXPLFm/M9xPEQjlJQzMlJaTwt0u4AQ92D6x0lyZsMIUx62XZy6yaS97R
WBm8kq+gP+JK9XrGBxct6AydGZer0LxMysTVKP4K6aABJb5lbj0AyB0wWdZj6PeawpLonILlbqBv
5dXH/s1I4rXLwbpAuigkO+zEaphnye5bICGy3ok5qmzvlZC6sQzr1HhTfw0HYp/++cPfxqcXlnBf
P9/V1I/uHzU4Ct4BxK0BBbWnBWDtFT4b55SL7IEbbNOfE/X2djGOzKfUEwegNRIumHpKqcZhANtl
Ay2xMRS8c0TYg73dwK6tWUNpkD78GIi9NB03K0gD+N3yS08/wYVCtHrgwrLI1V80o0wajOEQyCjK
L4W48YGWN5fmRDgDqwlfOafHHuono8LO8+MQs1lPf60mzfHAtbW2+LdYXegpXzSHp0P7rh26aaox
Wn8TNp80K6lHhJ/gMMzygk1mzQsTzKYI4hPsCXU66Mu1VHjBLCKlOzl6WZkH5t32c8fMSegfDiOh
osx+KuZ/JXTc2kmbzmNukdKwkTz4kVG1QBRhQsPFLpEIfKd5lUhdSCUICjoHW6k6+D98FkOHtx2f
aTCBxtn6g4sadTaEtrWG+2eJx2eHrbYRkjRQjD/oVgK6kG3RHnF7m4MUTtazGZdIxeI56WNq6C3P
ee4+FxR5EJlAxujxnmtkyebx7OJpZ9bl9Cu/nfRtbKpoQtQSUT55N5XPDixjqtk+L5gkd7dPdjPs
iA2fMUKsh+tVDN9wauXmrGuECg8ycguE0WFNecGeXBzw3Uio7r00xOWraG0rEFUZiMWVsZLNYwEP
0LTJsWNAyS0P2ijbODbPe8pGlPvuSUFHh6Bcgao+tehu8OIBrLYeZTeKh7kYKkIxrPh+eocAMmpR
BwUht/XnYzeItFq6zJ7wHk6rHpg+1WDUHe0RERFwCOPFv/6xgKcXs8iJr55OBPSuiTKKWMCqhlgQ
9yfhkr/QaEtlVm5Zp5e6u6UzHf4WtMvp2oPW4qYGIdwkMD31fsxCQF8PwDBBU5ipOBeaC5Neqeh4
HHDWk0Jbr3cV9F+R1hIrsK7u3bQGaKHPPY+S+0TqKHxHyR5quKg2hNwvr/vgJth4XXZwLoj2tljn
dLibluI884BS6YnC7URr/P/fF6SOfbMMWLi69QJatt0ZK0QmfOGoL8lUVvqv97BjfPYSdjdnb0aH
gL4xwE48znzo/LZWwfa8c9ERaMwQTp+H5tgE03/xI+4qQfs0B2Urpnce/Xl+z41FS/jA88c7IG5P
XfK+sgFKZzy1om9e9R5g6PItqnsH63eX7XDZ8fauSWbF9FDnOe4vFwIZAZ5gudxNNuSC5bDuh6kC
U471q7w+FwMhQfKz64jStysJPVkXlTRgn/gHryZZt8W5R4otLSrdIHnrWjruLi5Poh3jwXjWoYGP
PWy3+WAgV5D/1y5OuyWszdRMZKZVMesA6awxKC8u835QyWTbvMwqCi4nDW2zTuS0mxu91TaEYRDJ
2FS7aEIpuok7IIgszOONj/Tk3mswTs1UGscvaDsFVW+bdsQuRk2hNF5pvOyfXD1GNVBXiM2lhLOB
ZBXvUvMFzz7ymKeU6TS/gvRQSWRJP+9pT1gg+5Y24+i6e97Koe8KsR1Ds7D6/4U6JGGP2KifrbxM
ehYs26w3AvN8mjAkUzRCvxYIYIjBLj/WkfvaLUlydu4M8VaqHarP01xutD7DbHUgW0UW1Ir7Uz4K
joS2CsrG9E0IIqanoOYkRmOMCEgmZ98gqwzeRr3Cf2MKvhY+fyz3CDXogVEbOiKZyZovxJnZEob8
4IWgZ8+AkcJ/RIlUk46TYt0e4ClyBkMFvT60F9g2NZhcwMWKbu82otOwfyhCH+0AjUy+vjtHTixa
5/hNJdoizhfQ7s1noYtdCRgzte9hvsHYPc/Dr1VGpN0dqX1hDCd9TdpRZl2aa1Ei7LBoWayF+/7l
5nptiJ/yiOxiqG+g6RomBQe4LQRTH4DXIoyShqTC8MQ61YqviXJca5WOhXZicrhexsz0un4xai4t
UfmRw+rHp+n/ioZvstLrTJoZjoz2QzI8Jl31pKn1DtHEigdzeqJa4AY50nMVGqySoFTddn3jvxOO
zwRMhIimwyo9WAHs7gznWEEOjK/+MQqhZ4xVpcEdG3Mpx/9VFbulLBpmcCiUgSKhJPENY1En9k+a
6LA214LWG4ZwFOcJxYEOkvjCjFDLEEiYPUzIZAnpu9Mpi3raoT82fJ01NciBAF8ZB3eh+PM2dWWf
yL6i2fqrt/14h+pr1mtHGdGklZ9qPpgKXSFQondQWmc7btx88WOgBng8L+cZDhiFLq4gWKUXuHvM
810CUUrIpdUK1OBTDsQ0i28bWXUIm5x1vmTD7cPPKK4+ezaLBac7y2bjw7ok70ttCRBw4zcgAqdG
2q8TFydXHf66qmNmjSqx3VW95zFOjbm6EjVUSKzO+Rd+umF+rbM3asCzlJCf66OptO0ZZKbIDAVE
xw1E2PY7l9MVBk+j2S9uVKXAe1Yq2PRzEzxvtnV8AAhAJVAmTA21SYnuoIf85pT96kfRtuTFavQT
YtD2wVAU79GRG5CDcsDiZloSOv/bpksnnhmbN0S/u2GwdRrRzQuwyvvMFZ2t7lCJZhOzMFE6AXKF
fimLgUd2hhgfKEsRVKueRqR3c5GrjfK1ve1jRDnpRDToYG91YodoH9wgjU1WMnmlwejN9VE1dT7I
bsgdi/TtC8ufDUj/GeKth3AyU1fxqrgRjM/6t1X1P/lBKK3SZCtmZw1FWZov+qzsW7xhe5Rhnkl+
YJSNvTUyWpCzv/Majky/1dwURcP9X2wWd3HgL7EZXQFfrzSEcoWLbYVk0x5YWgirlHU+tm5C6nCn
IYE+tyGVq+QuoorOxCNTpNsDZ0UVlTp88W9lcWpQKs5dIJpJfOsLnXVfYzLkP6JwIOB3439JSwde
+vTeqA4MhtcG0VkYCwREKdGOv7fuuTt79n1OfwX3mb3A8TV3heLDy0LHcCYXSEwiU3/6l3whO6eE
77IDgpBNJGXjv6ivqQBOdUZ9Ujo4biEOhTyOH4hpbcjejNxBd2nETQTyX8UkuZy8BNLCS8mhXXwb
9B1eifSErLDwXnYazjGokwSmZ5kat8hrUf2hsLEtgE5MAZT/1hX4G+YnwtpZ4GE8hBfKrR8mGigp
dnpyDclyMySnPhee7iEDWmoHzOZaaFmntoQJfAVHUdy9Cvz8KsZNoE9Rg8oI2Ksq+VNgaIRV6qFA
t4we5qxyjlK5Ig61j65il6mZ2hp/KM7BZA5ltIW8GY9qROMW8Kzz13Rwm9IlsXpWCJLrmeiowVrP
sf5XRO//5THynIKRk78cEWoGA74eA2yANFndFbEdVueef/3IOqY7ULc1OM+ef5q+8IuRmIMQviXY
suVhIBsvZox/Wk7gO7viuUc+buI0vbHxgzERg8JGXjsOvj8J4R1SQNot7lwEcvshvqs3r383S/ZE
QzN4HTWk7TaBi54v3hDmYoSuxibR13BEacLtk4Pf0+vi3in6fYSVkEUs8UTBCyJezkEgzwg8HFaR
lkUPL5AhKcv+SMIVHzZOgYm6+DLu2wq0Bf9h4L5kFjEoNRvjJMThVMlu5BEJOKQR9BkcyzYkPyv+
lWGYpjW1SsUWZoINcLS06s5kvAwfpUaBmA6xvy9wpq0VI1Joo8FJlJipcrJl5qd+/rHk8GGB/VO0
5VR5g9AJm2nu87nE5aWHccaZq4DapFaIB+B6vr4N4OPgH1V26RbnhWg1tnRbMlzhYQsn/aroGken
eqPEHTG0ZUjeBu+QwvmtXpwaL4PVFuggiYOMfDw0dF7K4H2J2JBmKYpCnyniJJ1YE38k5TPwj744
g7Il9l2vqZQp71eDE/Y0z4OUcwn01p1GZdrnAuCU766TZRygR5+g275XVYDZYKg0SJJfECpQJMVm
kZlva3NCAMewgssdrWOeDQFL3SdQEo0u6ob2jmS4bknX13QgXyEjPJUSs7tnP4XO34S7v0YrMnzW
bN5zqLT2D1qMiGMZbyrV056eRdYrs+P1cDNKYbAL2X8e5f3NBU3VVmIc2mWhTI2X3Q1EW/0Adl13
7/5IqE8UHHQk3VYzzgb60J5CS7r+j4SWlJvqNwClwRlkt0TlR/gF9FkeKKsarWmTCZIFYx7eKErz
U8UuONXCrfTb8Ve3JBeMjcYjcJNqIHDlRU6fJHr3MY5TBt4bgr8teff//DJMg9wpzNzFPazHeDd+
sg4tY4ve1zNnNxcxzI2LQTcwdtaX6WlO94toP8VC7oQqq6fyHQyjIwS+95qdgmOY4A54ICvw0+ak
uiQgMLEWUIC6hAdHdy/NTYWVYncukyjxPFRp3Ku9EbANvliAYVvbwMXK7U/Kq+Iz75V8NoXmjXnW
C8v5ToiqNHjXdPz7wE0hWWbucRrWYNM6kISApkmMW7CFz4QxFsbvku4ehoC3k1NHGDje9SoGZicb
W6hPH3PghP9guk96reMFmOsBo1V1P7/l+W3KPK2kUP0zuciTrpliEF9QS8M+WHhAz0QsvhE0PCQ0
K6sl5jqjk1lVS219Qv5rudqlwWfUjK+u8c9bDAWG3Ev2RS1lrgRxTDsfR0o6Jo0wAe3KzUI+D35a
8ScNGRwr/ZZPIwmtSvePoN2aHm1EBNXWhZD3PBBRfwUjk1hAhFhYRfrHAEX5w+6Wan3qNoWG46Km
mSCulvG+ihHlJWTcUuAEne0e4dTYC5geQHtbJldDMUuSmnzuYdpW/9pl0WMwt975Xgj2H9UjGNSC
5nbNgIwkPzhOFHk2S/aSu7HyjmetXRwED2U9yIZsHanvTTN4q6z2/zZgHeA/k/ajTpi4ekfEYXdH
o4zvqUpjD9sgLy1kfgR5OW17sB2NzATNCo+VdWLnbcaGNn11iDvWdeSqWu8yFRcXcLo/fYsEfl3y
X8pqu4e8NN90CdWP9pdadzwxNiUcLphDyIV+ez3QbzgW5pA+yXy9v3oKeGLObjkgfYPl31FdsXMF
7rfssUD3aYaXJ+w5EgNNPpivcLTJKw3JZCbytBIkLnxTHGxpXiFC8K6ec5Ilz9Htn1h3GS7+NJW6
ZwltH2DtyrNdWACA6Cfn6tMd5MwB0bBDLXyQ/iBlya+x+ridIVzlHSeaxm14lsnt0bgIYA3cZpC1
By9uDoJi40CuQycqJGWQu5XRdnsRmCHlRZf5y/wASoC5VsX31DQg0Ogihb0CBhOhCuGHDz4zXpME
WVAiCHswR786OK7AhPmpREa5xfZ3tNlPTTeMKO6TLDOxkv+qY/qwgQMUXM5czpzcYxXjUSf3/xih
XUc8zs7c05W7ztfM6qCvghGhL453ERvP4kDkeHgb3ztITtV+Hi4fwAf2uAy3yOGVgbvxB4f3P8Kv
ADDLhkBfGlRZ83n93G0vjJ5qSMeK1lZLkTlTWdqF18hD32EJgvdxX+jyAWUfcdFn3QzcjlOCBZ07
zggnNtc82V3pc1fDN/fwn8hglNCxP2eokt6m87XfjeEMrGLsoGGKVMqspQbsiHPgA1A8ctgKirgn
watQ1nQriJ+a1FSIivwiGDG84PMD6OrFZ1dxmRCi1oeefMyFsJ0sIbJFo7+zXaZYvAzCS+MVGLD1
1XicTDH+MgNz25km5/F2uCMEwLgepTznqM33VtUk5hA7pPue1r0reFK5kXkcWiNCKSB0rKvvDpiD
gIB8vOw7VTRBcGEIaNUTEe7LeGSImLpCLHAMmkJHEGprD8jXFCcpvpRtEboYrHWT0crl7FJ41xVy
9bHZqxtGve5V7Zhfw8XACyo67g40TaqXdNLSgho1uHEV+UcJPBDJbaJAP3j/g/TaXbK0b7dyI6bR
d6cnJIWXgUfVmVzq/roMlNvB0tUNHM+PjgrojvoEo/jlJSPEDER94ksZ69l6N79lD4QI/EfP8QjC
EBZJkseUPo7u028zLuozcirCIRHyK8BnFl+8O9I112DqLaxLwX/hazS2f8Pvw6Dr4wQrq3qCtZdb
dLi1ThVADKp/EM1tSKqrZSdFVGLBkBXmUXYn9xhpvvKfsRNBbTRTyuUJrcKbhZ3oznLg1GT5S5o1
1zDIOQpndtRuOHkjBnUtbmhdcnDHRGDtE0W4wf+tTxfUv+A52YIXdDB+dfiTGVZxXQLDZPe4n0HJ
J85Ltf9X45PYdOeSyAJu1lFZPFmRzOdA/r+4uzcrYVrJ87HPW7ofJ6bnmIaa0xwODxkVHfRq15lt
KF3YTRXqbpjmdzGmJGtzj7rcLcwkesxB9Ye5PKIigVj9wlaAUc2de9MqybE4RxSYpSnWutvS5wGK
TwBZl6Dhu75W8PMM/325Dw6NvqgZymljkEjfTNhOCi98xQyWp5Nyz6TAEdugs5lPXnnphTUX69vF
B4G3KregCh5djtu06KG0O3fQ125AoRwfeQB28Zap+7tsW0sXlyfDgD4nqiGB9vozju7Fi8OXBjXM
FALWAZTdpARl3gXWLqB+SQytNYjXTmC2mCoLsm557vYG7jj/s0X2G9ZVXwnKkud9gIyL16MQT2Hg
8dg1eA44XVD4uvzAQj4hqF76vbedhDpjiNb5U9VlYSBY15n28GA9Vc3KBJZBndmJWvctJjLZe51L
jkPAC5pRM1jwMSBtcIXty1kG+c2QCjCptijyuMOim8SUTGmUE3RFNx6FqwchbHNp1qCA93C+exMO
84h2nrvx7mIaSTJnUy94qyMV1Ojy3VjIMz4agEpnwcVp8/Mx/4NvXtDbAaZtiYTOwChM7Z8zn7XV
U+dkcNSGN21IvcA+GKrtz5NomMuwHz/HmnMOcLpkUWnwC8PyMkS3uwgp4kJKOZF/dVRw2cFEH02q
wikOfChvT7YqSGfkB7g51CN7fuXjke+quBM2tepqGWvwq4DxlTOTmUDcsdZfwjUISsy4zsqiSe0d
I8E6/XSX1zEfnG1v1uKMGi45uuxFwiWRGmxKR4cBMGMqOpynEtWwNi+L7D57w5QJ6X1ZpktTEsAw
3duKvlbfhqN5+GiRMxp3fUcPzgktp7U67QTD7LjxqN462IjZocWbWA1FBmF9hIlD6QrWyO9rxjJ7
MX8bI2U7Kea/Tn8rXG0Gc1hB+ye9cJbEMs6wFcYKpR3izb0SJwwtCto3QPqGmrfq4pLziLfSQja3
lOMKTxG7ZqxY7TwhN/gTUrdx3NjJ4g+8KzzoKHgP+HcPmsxtvilUHEff1QvBxHk9B33dxr8rf+Bq
1MOCuGsQZK0FTyyZwS3wzq408Uqi92u2WAg060dJ7okDoPobAuWsbnaGH1rTKUk6FU8kHdiLbf5j
EUQtA2/yIUVJu9Tm+NG7AUfIedsfgbfKjQlIuPn+ay9dVJwj0np+kjs2Du9EjKE1+XVkBrfYsE3j
IL+YRmalumKRUq2Cc/7Ldze4XSxWYTzbT0/zGy2iF5AMC1Yw5HWaqXj4xHWotrwI0XtftmnzZs6H
G7Jz+1++yBPefPk6sXY/Dn3LwlRv6M/wSDraTk9HUTyN/HiBQQt7IKJ+Rd2GVwpTRIC5e5gpUdDj
XV859ZgYKU82h2kldqlVwYqC5bL/Oq2PUQKsqTFhhgMHE8qYmlVca0OYLZsbm8u7CanXBcBr3b5d
189ERuV4SJf1i/NxM6uMrAThAHuOnDb8jUU+tzyA+LeGMnR7kRy1CJKfYpAOTZcY73+z8YKR/uiy
HV6MAML8kLH6Le5TW2S92fykks306nYvd1Kzvoh/G5w3Ply/qO8yymv7npxUpV+bSgBwTTZ2Nqn1
WWstnQR81wTjknIN8VdLdOWdw4ISHUEuBgGoTshQRb9ZuV86TLQiwAw+KEf6/GycoLqV4784Y1wK
71x8DF+TUZePNvT6oUtqMHdC5xMRZdTHQSfGC8pxK/q6QAuSVbgJhocWf1tJKLDvlyEHqBVSaapE
/HIpoP8IUuvQ2GL4vCQDmJuk6VoAG3Gd8ZaaxITZqFtSYfZd0ARTYCbH5XLK6qm5CeMzFa6o77tO
Au8Z8fSZR+7aXlcjajvDp46haE6bwuDxcRsfVWNbfD1oyRN+tFWEwXinIvqOfWJvzeZb/wECOMC9
0zJjrmxRg3JRwVZnQQKCDKWZPjp9jHOhsSl2sx2yI5oNfTxCl+NcHGoT0nZWYxKt3dtrPNWfTcMU
nvBjREqrO/go+d8InhKDgABDrSImZaDzSnpLJziEvQ4omHVME4up/3gKMCJDB7Z4nDLWUyaYsyM9
nyR4bnJ6++58o87Qd1kdZhdzC2qPYnJJJfnUBWUma8BPV575k8kCb8gCkOis5SVWM25q4p29cd3M
FUuqu9yjEv1fFIE2b9JgrVa4NCRTRcPHZ5FcKd/qIO+7geQkdZv9HNDx4Jantu3BMQSDuaKYPK4S
r3UBriOEZnO5Aytkd46u4835FpmMQ+8uK7Cimcou6xP47BZVKaacVaEs9pd7UAP9zgjvvzhGxpgn
9NunreiW7HNPaMe578FmhAjbvDOH4m/z5Hkt2tPvUZ0rGLfp73wPmSC2jegtZVPsQCGl9gWtmCJ2
n246L+Tzr5uzEhRxCSzTSkDV4k1iSCsgMGRzIQ4p8Gmo6I5zVmGo1G2EpooTeCs0AjTkRJKAw7S7
5zwbaMbwRx2BWy8NIdxlnZn8jJIFkgFh6k7EtSf3GHpCqz0ZRc9RLy38Mon4/JUzToyOZN6BSGjb
FDPkknfb7mMa9KvgXE6wQxpS4Tn+5bKcAqEDRD+foCW4jJDimQshrOxnvRTGGlfrO13oE+m9zWku
OaGPMPTP3qFME9X6D11tTbxCwQSIInPWtGSGzf29ZRElorADMaKBljR/miWjWyo6oQjTbKDD3m8A
ieVmuJyUw7KD51X6WJOeCYJfU1I6BRSl1zwPn41J7rl00qrUFnx7i4f5MhSowWpYLyfJgkD2RN81
3VnY22luxyokTOnD35kr6ChscxP2QMh5JZ75WAVmVIQmKrASZ/BtQYXkY8VeL6uXdQlaKZmJYkex
Jm+SDjpVAdtaSIeEsgUvjH8kzZHJZPP9v8vsH2iFDvuYy/7ziXdEN2Ho/DGoaYitbLZonGmCCv9P
BhiUJDC92bthMk9CyHp7gzpvgAn+aGOFYWWrRcq4UR10dLNWHXBYgskhkA+flc9x3/c2nwtqS7m5
+nrNk8KZB1J/Rr2us8d+IiW7cc3nabd1/1jzZT+2KsQlS+qAu24nNlSFvUKCu+tVi4+PrKfb9yWh
LFPc4h1pAkGpNPj///p9+qhWmKgRYt+AqsXWrDzDgnmGNM5L6p8MZVMIjBDuZiFAn7BWEAN8N3I3
OEdCj+3aOgCUGezv7SlMVoo2WXFWpPkFZxBmVexnkIqLcPFAg5OzxGtn7BbVunpknq6rnf/ua9sA
BFyLrlDKEJBYbF8RFhTfAr9F8UEUDWp1D09Gc0Hbq6IxMdG4IY1mog2IF8TduPWyMcrq9B4yso3X
ua0xce5icd8kC6KhMS2qBfUAIIMiu2vmERW7L+qeGFHBxI5pbhKJOQxix9AdCPnE29U7fcY7UcSa
JTCDl1O9ynLZ5ZY8A2hDjdKNLFI6R5INLE3xB6Sa9OVvBLceBvBKb/tarLpEU7JVkVW49wcJ1Jnh
O1bJ4/SS2ZPcBNBUQEZAhDop8D3XnFGXHUb8WFw6y6aC88QlSwA/XwRkWafm2czlSyJZpqR6mt4l
n9fOKIh3ZVu6qGaoz1Ue3N84No9QFSFFmFTNGUCyRqo4pniAP9DriLjdsb3Mj652XOk/7vutQqLW
CUlyfEppvDmieIos02Epj6gBEnbl0J10STm5Yc+sHvcmLiK0HgT6AlqA4qF4jbHQ0hxbfAOIFm4Y
IB3YHVul+rYnBhSyFZHPGU0tpO+r35sBd8upKSwxuFejrxoS52WUhHW2NmwrAyly864/LeLMi7p0
u8jCn4KcXMKqLhwO9+HWA0gVtV2vC21Q8jkFfyOBUf3L3FXT50GkLzWnPI9NV8jrQKU8vWLmrjl0
OuoFr7yz9SxnuyxIgPBhXgpzv/zAGTXbJqMXUxPsEX3x0o1BLzr/OmGwzCAVGD/6ibKEQe8K3p7d
rhjW49h5scFFrfc4Nd2TZcnLjIJtQIKwo7UmIXEc4UuoMczOzeji3HpgKYM/JpjPox0wyOL4PsWG
utOfBtq7gsETUg2qgUIM0tJos/sRGX0+wUDGFQBSVh8FqKu7rZjQi374uTzwbK9+nngyRsqHqcam
wau1tUPhP1DAElrkVPoKQoSyz2P59wzUCH29+7FFIUCiBQh+T1Wf8IUtx6wsY3FfnQeVe961IIqQ
jqDBzj49HRyzAnDOmZvItHBJOIRquZY0a0OEiLiffoPP9zG5M2m48UoSbWuHxm7q8pB8i1lX2qiJ
QIeloGDYvWn5FkfWNCfl0X8WOoL+fbq4s+rPff9+ObcOQ3qIYgMvwNNqH1EWr+XvoibNeYK5BtqY
/UQFMvTlxMfu5rAs93isbenhZ+RhXqOuaglW5Fj/F/thwaWQRqnsaoDPn1xKEeqvJNbkqT+mlvvR
tCWiO4KgbM1QoemwBPrpvWiit3+RHUhEZhK56UO2ln9YQ8DJl1NPhgKJjnBIhBFUxdJDPdKZsbPH
pxL82kwQfhHiarxpaJNuXVr7izM+k+n4ktkHZvczjoiAFE9IJPKw9OKl+mWi+Bnv4qBpvVqsoF6J
zxaZ9iaspYo0BfKKhqsIkC/b1NnYnBc4LBcH9j5Fna0k58H/dX8MKt7zhMvQI+4NNq+anj9HBZA1
OXqaSC3C2e/7kPIUqOxMaIEGeytmXixsALAoCFe8Oat58fpb5Q6hTqBPEcSrG2jJtxNMp1ZKBGlD
kpV0LKr68Ae2UOJ/qj6CVkFoaRTdtEe8qQgHuY0YRJuoAK8yacD/lCuJUHssU0f8EX4SVOzUBkcS
+IsZk31KvjTJT1zsoSkl5Fz3jgYTXmp1Wq/FMacx3spvPP0EAOcqhDO3Dw0y06+2GKayF6Q1RcB/
3viKj/ooJkmw2T4bwzs9OZvA8LlClNQRDDo54EwFvVFScb0yS6VdJbSvN2/HfQ/sgkYk2uymoM2I
Tr8IEyvbgfr00z53Q1yslwf/oMpD1dAC7hIS/DnhELjllnQ+NBgaJxa5kQV0FDLbPbJKofs3hInf
5jy4P5gQ9W9r82NJHosRXN9Is3dMADAM8Uk83aBIgC0JnfoHYa6nOty47QY+fbDGqSgOFCA/NjQt
XuqXIXLGtEF6h/HsIqgZJrqW3yLX7jUJ/q0PzelHxoZKyw1yoUEKPFR1cNuflvbxNXxGA+c77IQE
em1rOT03QpyoFxbBglLrEd3Wa72kfOgveKZmk6u3A41NU4o7I8tj6TpQiqsY6JZ142fbnGpynX1n
2C6N3I2kPGIsprVUGm7M1JrHA3Pmy/vpAD8OMqfvR1fve2pTKlfDyYFXbMj7bLUNGl3+kArb24NL
i4eReLF4wqg1aYO3uL8Un5bu91wAWR9NYN3BfK27o7EmDClOIDbrlKVdHVEa1Y3GXngaw0g9oi7n
XeCbje+q9xlY7FjBgzhRovXCTXJiMK+HvveNCncNqqlNgEX12FZiS+hLSsSKOfA04f4r3JTTd0cn
P71Q52OM5WpJaStIetbsyzqLiyx44cltj8/7bvcOLpwzufNnTTbiuolLE4GK2TSI40h3gBrnr+5B
K1TWkJMsd12GTG7rSa05fqH8w61j4Cgy+tXgI44qDqT+jF/+JUrAj7DyVkT0p0+NPJpfm+kiH4bJ
CAxzRs5a/zvqwSw+GkiYifw0h/HuMzBAO2YJGovO6G81aAwUBN/oIUE7CST2bJ/zYSR4cFVLa+nV
8cgtFZ3WTtY/axl1ukasyHV5w0cfID3PRzEvAVdHv0Cja9h9kqOsZawrOabDbqvEQCYQ8TD3ndi6
UPQkz0RwtLM7Ppyo0je5QEd5uHD91wRSLot+1ps3/FA1cM6pDSH7sRCkTxPDBXzYEBjy4CPxcw6k
mn6HjbkjaKmgZtfzzBvI8QubCyzqTEje8bc6SU0F4d9RapwPYgu9lftV9jqLNdlAypBggYcYgFdC
AdAHLEyQgXV7Sl6O3E3EZe6NG24mgzl+aybe7nhGKzQJX65QXixeI6ExDtGKFX8GT9koAAjOiGdr
ODoS5V5uYpWHYv7BrOnEcvIRGNUJyFhXDjV40zimWDA/BJv3CrlvmS44MUY5g1yzhZ6RM8UU3t4d
5foN883+0mSp/vfMSz0j0YC9nVFii+R9dlCZRiFUDPDlTxeuAHDmIRnN5gjxmxqiJIc1YSlPUCLl
F8PpEeLz1h7pteSjO4yxtucHOgxbYxIblVidQH1CLWvvR0uT1srF2qWMuAcBaZBOMgHL4CSTu+ks
D6kdcubRIMCoINIv9K/+O9M75HcEoSQcW7Lg61pjTk3x4oVlIHCK05jJco5JvS9/jBP8iP497FYe
f2HUG0WOuyp14rGEnQL8V48GeBdaBRpTLbJYqLL1/pQ+GUKnYGyp1wVXKOMknX4ICV8XqeE/jwie
KNRKxX9CKkTEOsaj4545mJdP5gPKIKjlJd0lxy6+Ung9wO5ZeLV/e7f35jC83v/UlXtBkdiF+aVL
8094bLV9CkQqrmX2/SfCj4EHk6v6IPXqRWXEmz2/dsjud4OZvI0Q5vzhq+x/RQcXxMmVxmu/Swuk
/Wg4I8p3hzBL8uQDuHu498WiSLDsNDCKLW9lMHwFtZTVtzgiExr0zXzu4f89U6EK5IvybnxeO6bb
JjIr/ysLVdncFspPnr2k1mMbhOmlMkC1pFW3Cu8K2GIkcq9rdVqv8d3CeVSa43cYnZILCrdRUde2
0+Gs3sLuUeyhx1KipmgPCiPe7yajNWtGBQwkYJd/fZUso8j0Tzx26tU6DY24+o+mZemrc5gqoVJ3
WCSDv2+It/4+InmeMHLUU81re+0orY95McoiXfmFzIvoyP5IBFjb42b2uJoEZT54exuKcDajTPTr
Z36hU9Do0cL+I5bWaHds0PKdoYHgP4Ceg/8J6x8fguZqFZAs7j/D8b7wIftUeF7t5Lr8JPLy3X+Y
B4oSpFxWMNoKjrs7ew2Ae4EKDqV3fIzz3p6je/WakSMmW5zQ8cQoAN4PdePQcmrfF8+ET+7xcwvZ
bI5tvY5jDbHl4XgtKFPW0w1LJwWRytcZvuDw3uV+z4rlQu+oLOQjwB19+VGv/HIl6V03IseVM4s8
dyFLOpFkpRaDt4hP/fge1j2L9RukkcCbQtA6PylO9/X8ab9r2oaN14wli8T6XjKh/n5Xx5Bt0ieK
GmKuOFdov/QRCeiXEivA2rqMnKzLNcu+bOiPg01Qwr0lmwYUqGbeR9z0mGTJ0ylTGXRqlddSYz3V
I/k6iGGNhrgt7foUnwpcankCnvya2YHINhXetuG6H5t3EXpTiTkxPZ//LPTMxJmkbDtuaIM0gE9T
IVU22lERaAN4YMY0hFQhtyGHBP15sKaoUcjkAySfOc+D111HhxHuMThCm+mcnLW6kbeXh3+0W8pi
vG1XK8Oyu6jiPO+MB4rcUudOu2A0IuiMBvJN7SxagmilXWr17cpFZx5kNL9BLMfTvY26qRjkiJTV
afZ1qeUF2oPpIiWaDPoY02JdY9FplKYn68X+ZcsIUaRwBLHmb0Qd49JthDZ0WpfvKTzMobwwxjc5
HebauIr/YmjLmeGafcflNjeCE2An2t3ltZFpsIxU/HXdwp3gZzfSU99Fxbtn/pjkaWjHYDTuXkG8
77PUs2nVgoOZ90dODbJU5q3/WSHiBo7x5mILI9al4mL8n5Fr2+Fyvz7U6mS0W8vfyDHCPvH1u2FE
AnLpslPU6b7ZC16038C5yuRr2vycR0mOwcP2Da/iCInf0p9Jy7fnI9BCA+ySEG4F2S401fra/12y
t0LIs6ui/u2N7p/YX3G3ULqlIIU5IknbZvl/XxVwh5P8sO0wHILtigi7NJYCDrqxCi3vSN+PfNf9
Dn7pTgpcx3kBf0r/+ce4E192BCF2JtgVmexmB4x9WLPa/SyaO+uahxprvBv6FuZgNfYJuHsEFbi1
NkuLWWCkDVXFEEmvCt0TcAqqBGbKK/OQjeNZRYMNc4m/IFKfihd+xuS0SRC1bQpwwZjlX7k3NNNJ
eSQdMA/EM3SQ4jAKO4jIWP99eSLRVelOg73YP5T/ri7JUGNigVuZJ/obURPJfbsJqh/jv3JesdrE
142NILuY42ZU5Dr6l4E0aE6vmRSAdLBqg+BJl7hYVbQ/P7GI/1qYs9YR5OFIXzSiKcinv8mAvzYE
vtdJVHPjov+cgWI/xWyP0h63lx0glNGbUYKWrVIDL2NE5qtDzigIciBGjuPW5gaetbnhZKPs8Z1+
6srzcN6L5nedynY81chGYIbjN20wjpNXxAWeWjucd/qBVZjFihDoall/Hv36JNjwl/pVphz3wpHY
+5abAxvKUfDtTjmpXlZk6lQjey6siluO52OcrHv8YirWVV6Tnn14XW9Mh4PucFlixmltfPIoWhFJ
3dh5syTTRMuPskhcMPwtL2RU1qmFeckReITXcoMWNdngUfB/yElj5lJoScCDrK5SLXxYMyTSa/YW
7WiX1Zc3xBEKAWFm2r1+Sc0/HjcCdyePdiJQv7VvK/Fybv1QzAJaaUvRyPcZQ3wQXHaXk7VeykEZ
cBSFLPLgfXpe9Qqmm5hACWMHXbDDT85vyTPiXqpbsJvZFd/LrgdeZnYKd8Md2QtNEv6M6DoYGvEh
JbNjRCjLwlIn1cLtHv9WDJhX70rCEpAQ8ZhXgNXcbTIMT4zEvkIdyKJDdMnP2+8xXEOFMHI1zlfs
AjHy9/+GLtwdBfeFjnThitLv89G93TUIFpK6CKt1RSpyzrU/edQRp5FMsBeQwHGBYulu3SU1YLpr
sph6iC9VGpHv99RH2i/vRASdrtGQv0ruOZcv2idBc5aSJG4FPDj66RdAVp0qG8YRFLnKx5uSz6SA
hck1/mXOsGtFxShLdjUTr9fqPkM9YjTM76xVCxmGxy/g9QbE85eDuEGM9XiCCTRV3c0lYHmvyWW9
weq/L+plj2VvicFzxMpStXJNxPv6FtpqCbPRYn7ib8nF0mbejFTAhfGn3KIGKKVy8/3Qs0Morn38
gIGIAsdsmYH9Zty739pLfVN1wCy0YTDAjKgppM/ua7yNUnF3oBHIyR8GamZfsecPoZpNJMOWjQKG
eE3S468CdqOaIZ41gMN6V+wKzGbsjC7BcOPmQQY+8fiTJsmZyjMjEUWO1w6kay8Ne5hIC3nOustA
1tVcS4N4K1Z0TEeH8usnGIn++J8QDV6MaULzRD5nGzc3wfjWIVSfGF8N3CFkiBJah9hl2KA1BhpZ
2MTP6zyO5Xa+wPLkiZyTFhDa8auLr95ik2cqgk7lSx6/OuuZCvWy9M9lmvB5vqv5iUt4ZGRJvVaP
G4qbvEXknh+s/Tx8Lt/OUcKU6Aqh0GJhYEX5mGXLTcDAoZEzluxLHB0qyozidr4qS4t3cDhPZ1ZI
g8QOgIXZd8TmgdNfYMYwNeRGdzbjx1s0E0U/trr39jO/kfrwSXvrJE8jrEVlXMx3DerKhcZign2x
lF99xJ4uZ3v8n8cEkeOjBtHyWEiUsW9lRedQTQqpzCqWVBF1nJCyh/D2RGCHL4OJjuzyV3Q7w3XJ
hjSaYqMm7xR5vHMbE7UjqF5cjZ6l4bmrSek/AKSX+l1/kjqBr1oGai1nLSMapV8q2b6CRqYCkJo/
0XGSKnu/dfZcm3G58TAkmkANsFQJTkJzHcj7bBDU5tNASfUrxAb6dLAqohWW7mwlbjGEsOuPqoqI
sq70PcpBQuxy3y5KL2ue0ktGpEbHS7ILHfdu8ooQftXMpCvMR/wSipUpm43vpTy7AglKx3gNResQ
JhY+9y6BE7veqWBgKwJ7zTbDUwPLAIngxioOBHznfAHjQbQCfuYP0pmtz8i4uNoBd6qjJ7omFA4e
hwMRkkpGr8TqtdYzTwB2GuP2hZCAW+60WBEOKBtxKaRvf2Y7v8cjQA+nRSVVvRnvgNLXMPBCyTs8
DGx2DQPPO/nx+hx4cpj1vMRBVJnYBRFPYfqhAqbVXc3YRMwQAAL1eJX08pMVi0gZq64YrGUk3dyB
WsgwW2kDCU7eIvBZ2DKh2vPzlv/+L19Q0msze6N2WLbiwztdaQwnUkUVTbPRBlxfR5RaNBqMpyOq
gb3qGLMNL300fYjPn0Kx4Fu6hMxv5AYi3PeSq1zIifYR/VKss5I1qfCkoPTT4ZFyoeY0GjFNuqM1
wFHoGfkFcB4ep/b0ioqnPw2Gr9fxBZX0ZScxOYpy/dhD5Xs1ygTO1IsODiCyR/TPsqkAKVNqMBa9
aeSM1BsQloAyzsYhMVZ91/vG3I1BHrRjBdgGV0I1v9E0B9g0JoiPzyAf6F7yyS14V8LsdE7OA7N+
/L1H68BNpg+DP0mbOJzY0IkFFeDOyLPN4pBCkIPBQexevu7o2G/4H+4iKSk9dVPxJHphgzXwhP6k
4+fVh7+6br4DEBmTG0Vj0PhDr2TS/ZohA5uC6ZM73u37u1wuYpm5/1ybFLkxQczryOM1wGFABR26
NLCpMayUclegxM005pyhk2MSoiBgGqSB02/0kTmixOisqLpDHCsK6eH2UyksZq7GTbavBEue+2dn
jDOvBoYeipb4L1xfcFaNMcwa24f+9+zAf/8TdjjIDRUleH+fAYC/T01AXboDxiqcTd7VZV8o61Lx
7+GMFZ52R0yt7I+s/ac5QTp6sAwcJ477ftzMdBNGRNLH1NjsciVS3NUFOwwhkTXT5fovQYhEXHin
9ItfKRqMKr9F22OgxfkpzDKt7DzBO1rSWQbwNPaS2aLUEwm4e0dLNxxHIzy4O2ebzhRgbtKUVUzN
UNJ05OJ/A84bqLErIgVMkucmP/AHeCy8N+ar32evwwoabplRDQqDOkZyvADcS/eGkcumwCu+UNNI
+gBUbvdza9vbwk1NtwuvL1n/NeYfF1sxd+cAn/CtuQlF4F2IH3P6T+fUqxhOdrRb7WOJ0fWOG7Yu
gG5GHCA8grlqFtvoHlZT7dLR9gCP1A6FCzThKBqY6UQdEJAlgYy3UrD8xlhzjhjlYB0RBSHNhE90
YYWgh3uySaCbkSCwnflzJlePprpvOkTC9FN6HjI8KS4vSOYrSiLNPbRlX1EtRbQUC0ott4z3Md2l
rji5V2vyXglJ4nU76bcVI+Td1vD32ycKqUVbHzKKrzJ/Npa8YlMKzuPuKOZSIIKQo5S+uwk9KTSa
tkcGXlO6DDAeEljfj7BIHLGI900nIjt6TPEEsNzZiKWTki2QqzpPoNfBh/U+uMkZwKAOFcXJ1tuq
rht86nUsEY2HVFB84BkCNnxQV6K19ooFZpBrBCz861yQtWgDqxxCXrpOb2DiFpO28oXaLm2Km8ok
XsekaHklpF5ny6W5FCwIxEwwrGOsMNcWaX5rv2/zsPidyrkTPKsOGVJdMUpwKE2FcY5DT8GGDAJR
9dyh0zgwQsjRZSmnQacwPtMSZURUcBpyPWiAitV5+hfFJdq6QL3YALD4ChxQKtN9/Nk+7QVFGaos
/iPzk7qjCm85z2hPobzsLciw3hneQW+I4RCXtkKg6t7h2B9xSc6e1CG63uMMTWo4Z/J4QNZaYiD1
xOSal6cFqUPDeY1Mvq5TAZ+VbxMWLqKhyjEaX8lh/Lz3Y2iRxzO81XtrDL21Clv4ACcVSHWCVYSR
0eVD8smF8NwdtDs+wc5vBxUwJdDVJQlyFz7shi6nZWzYJM5dW9M546tRqCmBOk1Jrnrw6f6khMOM
omS6VvqVxoJPkKdIeFyJWcOS2tJSILGVIpgD6n4f6V3p2iABG9jjJuCg+rU54CiGU/RpTVYURuTh
aa2BJLUvu5q64WRPT7balY2OXH6btwDwrqEJkWNcTIk6pKH930mC4c1IZif0GJfWkWNepWeNdSDs
es2nDhOgCz907IYR4CZSAsn99vAZPkFodo8MPp905/b1WkhyVCXVEm+H5rb2O2fdIQsUGO3AK3mq
sAAytbpqFJWrS2GOyoDqFtToUs7pUAgsqn+5UbzGZOGQZF8WVFaDcL7ws/1p6JhLvRPT8gQcbQZZ
72HJ62sWKBcYnZ7cXsnsxKS1F1DDORj413nAnsLgnACwus4K6+BdX4RM4Y3/08nUsS8zrlCftqRZ
Lsmw1BYaJ9g35Jet2FX6I33OetyK49rhQFr3Sj4MbDdEwjm271P8ob9N7/cVGzklYAkNP7Xt4OA3
6WxypqsEH6pC1XLLo5meucsimG2gU8EqMbVC4YlEJxEiENnHOzuJAFLaDVRgtwFZ2WRb3U38SV3l
VHIUiJ/X+59HrNDsk0g5rftceE3U/fY6cLIwm+7csvD/ej/73a7rCLVqfK8ra3iVUKQ6OZIqAJNe
E99aSVOkvo4gQVkbXqoGZErLMjFCKbAk6y+Q6djfWQqjIDSWJ/39HUBxiwXd1fTReqJiT91+bcYV
ve1a9tba611vdtHn3lHZikfLaXeXQlHSheSHbxNE3YpLwkBJwVjYozWScQ+qn8R43VA0NSTI/xc0
Fg37A9SZCH2BK2VT3I6SgyU9lOvgNAarL0U2czwqWsgGRkMF0pvNVk9U4g0Xlf0ootzoR56qfSa+
n9tqV5k1HyA0ZOcoMbUgZypOu4/yF82AmsbZnkWzKbwk+xY7DONAvfLrOw28K4BNrheGNo7SA5IR
b1NesdqyTXd6B0SkgtJ99WGxFLjQZLuaXeYLaAKdswuwIEtESBKpfNr1/0cx4Tkw04gke00lhPLt
9QQbZ5ofZj0zM0u6fZ302sUOaGII1FL0h5ynxxpI78hP/jmeshuBQOh9ggoFy/UXoBL3Fj4Y920M
TmChwbjeieo1N43qkP5S6FxsjrCj859fr/W+rx358GTdaNLRYPf50dEGYUcWaJwrBJF7ifSuVfv7
hmxm99Bym0g1j86YwoRPxCEwpwYsiavSEn8UxiZJkiQxpiwvPxqygCJPNFbBdIoUVaYoKrQBVqjv
OD/La9l2BFrH7ESNdtG0qLAE1vxxYV4Gao+8PsENznhpZ/8uBFM8WwfOywcQ0cwpoa2qXJhCZEs+
m25fLY+T/fAPvUanP7niBZkSQQ80q8eOC3kW+WFgutnR8tnGEe2jhZ7cUro2kOC9/rGFBl0b/0he
TQ19MhYot3x3X+pAHIST1Q9EENmz26JXJY7qyCSqJYV5Wv6aVeIl9VU9pIf63boClmLv1rdPcI/v
UtEnTe57OMQCLMt2KBVJwYp7T6+awAnSZPHmBIFfhZgon9jOZoS8h15l1FtCPrWQZsHqBVVZQxXQ
6XjId0h2xZlqoUDcRDDxuI/r9cNwlP3aYrb8WPVS8EhQ8xeJmiibYJUCXDoP0gyXFkZlmPLh3WrE
C89bS+VlHmw5t3/14HUOJl25UAjKj1SOVqNX9GIGwDA7lDOzlG05/Zjh95pwF1+BGVOETFsQaMNG
pBBqXAFbg3ZbeTwQeGvy5XZGx/wtPhdOXLosrVdE9kvk0gBB/vqnZRuWX+1DVKDRFsb3PhffaFSw
1OtkU6ctHx+ZJTtxkwwNtQ/nkkzXb6iNqhaavJAGCCKqP5D4JyuyPLbO0in6M4R2bwsydjZarMEg
espogfPu68aEws43HI1O16OVJJnt57RICGMbelI+v+TVkOjcps6Qd91vVfhHMmG7Ea/KhGnaaLXA
82FrsdBWWHeva7o82iN/f3sNoJcYDxLLqXxxlVfXEdW5isQhn/agu4waxktEp1UlsqfXzAdW7SqB
uQq/sGzf/yZLtYXXqom7o7ca3PcDvfUaasMwmNoXOs2kWxmE4t+thDMVSTjTSv4D4n6U9GeQEOnZ
XJJSp5npKjycYz1bzNpUkPgWKD9IZiarlFyaY0l2hXdc21nOEvDYQ7/hGwgx0sh358VFL6aPQPgk
qpyh1TO6DJPL04rAXEx9QI/pQrVsMih+986BHbwiXZFiorRirULZZY6YvVJdrCwyywrjY7UjTkSS
7sVtKN7yMkFfFjx4by6MqMAq4fXJYXr5A6Shm1FDkVAMpN4SuC0JdkD0D/RFb5+59L0HTzPlplmD
eFPJ5mdKomnUQ+vZCTQnla69SGIMGPDVNSNCIZUl6B9RCkQG3s10xkmlGF70DpmOpK6ALeQnghvM
lfTD1XAL0tWIvNkVNTeef6dtNzpR51GEM5mDh2r5XWrfmZL23Qi1lKuC9xE1yu0im+Qm2jPvLEK1
Yhoi3BbkR2JaIFYeueCT1E50sO8p4jPjJzqCzCLGiF0e+d8hsucWHu+Ob2/3AvP6ojmFW83kXZ4C
XTVErmBrSOo3pv5T+su6xnpQeaHG8zTleInnT4nM1MhDlpAazuK3qsTE2RJqgThu1/ZGSnzYk3FV
Dv4U9YdjYAFQ6rY0x+ySQP4OcS66v2cY6xC/8IqArM8LzT/u+ayyOSWQL0h462Ko+sBV2TTukBUf
+IsK0E7UWdNv2ZDzoB7zx1fvZnAgn4yknGi3zGiVWwTQqgZ6re52pyR1KrdHF2s3rXComzMXTIL3
MBjj7O/UnRSergkcmY6MF2eKLjh6dPaiAmBnToTvd6XiUsTwqAQn/DR2tUNhKTC2WRztKfu83f0F
zm19q9vEdA6fOVqGW8rPFDrugwkfd43l5mKI6X/oue92NGlwW7Ud5+uDKS8o3HmqGm2knv8tGqse
8bOCtG0CJfmjRA1J1Mi1/nTOeGX3Yjp4jYzkwXtnt8DxNK2UQ+wug9BHG8IQPaehapG6sxCmwAeM
0zrIDHaMJc4py1Ogbil/PxXP4TfTwmsT23um0ZPY11RPZWEA5h+V7GpmbQlc1FTh+4YRg2iPIqCB
ioWzFfQMGtdb9UFJboIFn2fZJqMYg2BUlWIeQKd7dOObFgT2vqHkbBfGHssxuNfhaltMof8447lg
UQp8OJXV3qzjFF/RDkwLHjsMD6NMc6ZLzFf46Lx7MUbOxWc8anqWBe2OJ62JSVXHMCGn9HtSShmM
yaFRfe1ZMbp0v30Sli54bx1kusxPYfc0RAYGFS20yvggdFZlo5PLD2QhQJTCJR7eEywgwrgqNzK9
KANsfhjt8Wi2P4Oc5hPEhHaoSnbYviLTzsG+NY+y7xDBT4w2XqAkah3aCUx74IlwEoWY65JuDUeo
TKb3c0GxFdPEew7dXmKUWE7IpzvOFt54Hvrm7t2j0NhwlVv7/AHD7Ir33b4Ikgv9Ep0igJGhTYGT
B5+57KZAKdcDzJAo7AVzNF/nLidgcebQlOiyRvkq5B+GTD86enBvOEdkrnlrT/8jsV34k/GtEO3t
8Kq+x+gG3O92jguo4Gtq+J/OAQlOCAATU2MI6o7oCKiobJjixjIZEoVsYFB2oQGMpTdbntTTwQeX
LwdiESqTWMJx9qWZQ9xTJz0sldj0l6sPq89qttIdVSBfU9TVnIfsZxYnb4PiGm+CYRX12Q93VHmR
UkfxC/r2P+LXaGVtUTJbio7WoJ8OeGCqwG81h36mP9oaYtNEH+2WM7dqIccUewHq6s3fWLGxGm3M
L+x56KUb6vS4YIseGZQeNx3z+DYmtlAFdiaSLwiqk5mi7VNN+C43n5ycSPzbX/hChVFD1MgBHAr7
E99OArp+st54j8oSJORxurpReZrKiNgnyyvfLdKuJ4hir4a/n6CT0kjD2gG+0M+VvASCE5P4lsHn
Pr5QX6dCsnkxfcCBq/uFBmfEesfmNqZHdQhkdV4cozwZ4Sv9QgA8rJ/laR66OMSgEfbfjbAsY7vO
MGcmMxGkRzOiiLfhKdQnCPed/1go2/HI4+flpq7h9GCwktnsCEIcivyGsLp2guY3jqJJzitJZyow
zjSJ6sfB8guvzv6uZD6dlvhtRmbu7jRL38t0Q/4yUkid+erSGktVVtA/jc0Me0Mgmr24/Es7Du/7
ICLDpALJAHfhhBTFqx26k6tetz/0lZ/PV3Sv1BEJ64zVHzz/C4xe9h9iIzOEEZEQz/y1dUORqWTp
O0O8Kn/7scyzDQEgelHItAaeAQu+Io+6aKNSW43SMRv+fcIhpT2X4YMdrgSRoyiiMgxNDq3J/RNL
dBJjYplylwV6+gocaXYW/VyT97096gMPdppylR4Sn0BZty7YS83Evz0KvXKo7khkmTmkR4Ut6wgo
i7tKGdt4GOZZVKcxDV43ArKG9o+K20wOLUn6CM1FOFJuvsFggdT7XNZYMIli4eo3Thz1aFUvIGtN
ii4CwOrMAr7YpljLNgmkZF2UsUf9Nm0YLEbY9uHo+nwe2wFB+/3VO6B8IjbyQgGtnc7V21mlOGhu
7mR2d11Ypr4a8X5iDTuVL+V0bCY9eBJ3nhpt6zNcqD9Wmju8FvJuALjFxkorsy+Mb3IPRqTy865M
4QGSfSZGf8Fpu+ijrHpQWC0p41Ol7IE6h9YDf5jVXNl3uS756XOzDuBMpGQ9UMieaU48nRJjVEqc
CL7glQhLFciXBk/5H4e6LJDfoPVPHez5AeB9wNeenbUiRhW0czh1PwH+itDqjoMzn6oWoT7pm9nF
1kwfj83/9FOR8cuEBCVQ9c+GN1ok6b+0o0SYdZAMOzeWbIBOyORhd1EjIiRLfGPIE+Vwrjb6X7rD
HimYOwKRgUluRvhIMeX/VqGGbYmWtzD6BJcnt0Bb8EalS/FUdWcGTV1vvpqW9zmvI2djt0TiRVeP
H4C3MigpH/9Hq8BUIPDGgQTZmO0+MPmMyK5UnR9pzzWUPQCT9f+xoh5HRCmrLw+rYzeQ/Oa2wv53
jStkfDZXHgJ7mFNNALjqDaDJQic4owlP2/o6vbbCjywtSFJoVQswDE/++lMN5vDsx0QwcCz3nvny
jMiHoIvBQKtS53S8VjpJT0qtjmXjA5534MDMzKcwkVPcH6ISENs5u/03+K6/Y4skZGDJngmsuIdn
m6Lz5y9Rh3eH6fXWbHLmrY/1ECxhxbfaJlrIPkCJTvJNGnPLOxz7Eh1Rk10AkDx4NgPPwKUCnd3r
4wAXHOBtmqq9glZ6Lbjb1e3dLYzBvd2UmnddIkPu7lBi4Udx7pMUc/trCjZ3jEtBf4k5DjSgKKl+
WlDGLMVRfFok/26Fwzv9ZfRejdp62Wr37gktocQ6cREQhn2jQG1yGyZQYimLznLKQhgbghFtDhkd
GSaBJVvMD7XWRJ/HwkgDR+b5xNJpLR5GxBVnc8yY3wPW1ts7/hlzBv8/K9oIWRGgMVFJdE7up/Ne
r2HqYNlnQgMCL1XOWyMKxhc3sMX+uB1FUIlmEUHia1EAYfs+iQ4l+dzr2RKPIQxhmOQsSc7P1BCi
LVxtU67Ujkto9mVoQKF9T3ztNwfUxeSZX034PJdczNNbuethbdKoLUc13DgloEPESS3cmUlVAWgr
qsHefr5nv+QTb92eNxYVvgcQig9kueYmoET8I4LwYgQjsOE4cT8w6Ko/eDUT6yNbQmKiXRuC8T1T
AHHiWoZ6Yd6GRZll7KJX/yVd5lqn7oNXkLr4YbYlL6TSza1M1tjP4RneHUqJ7WS37bruIvCjGJh3
DFnwGXGgnwupFtx6QSrLC5cTJcB0cLjOnluHBSO3wrWOYL8kyfJv7SUWlIeHJEYTthsTMVI920Hk
dp9/iooAy5gbHVK4KGriR2rGygePpse9FQrj8I5VmeHCs0cyO1PrhhF41GotAlj6O2AMQb7MZVdy
kNBHGnGPqehLcKfCnduXYRybZZgtfOACzs/l4Cir4aZgM0EtPNqOh4wQAFjzxI52IL1mvdtwbNw2
5WV85/WJ4zQdxWogr7SUR/ZxVbzKdyPTrEpgOCST+98orHx6PHteqQ3paf1g+zdWttQXE5v7g596
UT26Z5jfnaG5kHzroww4GMYW5g9TmXWZE5n9jImaNddk3c6tQnddLRREtaEqtIyW6oslOQpRG6v0
UQ6xDttSCIf/2xsds6EyX8bJT0s0+KicgKhktOFaCmWb9zaP3r7JY72beX9yYBY+cZBqax9kPpEa
XkceEHIWtbBMWIhMckswiKdoQEp9idP6vo+rPAarAM5WDCPXY4JmhmjJFKV+hTO5Ihy9y4XdiMfj
Bj/0+kr/YD6Xq/rDGxOH2R90QWgrTY48lHMwpmBHrtSqF3HJQhuOC+qCMvrjUZhT7Q0MyK6FvL29
rDSqt0XpHl/n8BT7slTBP15sU3lRvwWM8QBAySPJpIB6a03EcN6MZqy4rJVdiv4/yAWXkU+fLX/D
6L9wcUFi0WTMRt1KXF11MIIdIxoq2ZjgoEOdqqp0jlQihJIdeip9FvSEHA5aTK4S4uacoIZArpQc
v92LdIbdkfntqmkPxxs6kLSFXSs6Opm1ozEQ14pBgTmaAGlhnsLYV6L0C7ny5IdHuf4PxMyOO2y7
AHfHRNznYQK6ejA4++3n5CRZEdeDcFMAKhYQCW+3bu9JhpON2VJ+2W9mj+dACBq1qrujys5SARCf
4ByQnZKXW/60ciP1b8pTfOgzKJmTHtZ+jw6VUX28dJd2EBPJLOXw4pFo+oI+mAmXRrQku8ovYmvR
8sIxUiCoi3a7T7bHW4VS60JYm1jUHbtnZOue1/pCvwejWAgoq44Nhs4UMKnVP08KbQXc4ZZODVQs
FlYa9qfe1BRaUAuGzQ+1kbeNjHt2vQofE9YgXuUc5HK/Ag0o68vwBPGq8ojT4eFPx1Jpd4/rWCv0
YU53fpTW1P+13SeA7Xg2pzB/XXz9IBVtuiMyhmR3Al+t3HUdPPLwsnLqlwse6cOxw/uH8ZtMW6ZC
W2xLYv+HyHzhb828en+Iolz6pENBFI83OuDwzW4XAQSOZRLooPEUqCQUSt7zrkobIrEBXSLHelpl
RIMc0sdZA5QD7dWc04MUjfIZ7iHleh6Fzm/pSV2SU9O0jpD6qswgPkhYOI3Z4OBtgxYtRW73uEmx
/gNZSh1g3gm8gngHAjnGpBrqKZvNgzaCIQH+K16Jr2CuHwguE1fNXSI9OwBunn6/curNKEQcWOt0
RhU8jLMmshzNvM6g6XNl3pQoApKFRTv6i5kVFC24Af2t9AhQmYtjYu6vy1OBIFH7NsOXytVitlSC
66UCg6Yi1IYfM1epsBz1OThnEgTglsrBp9A79sbK0/t3jTDIJsbkWDVcuV+Ad87SiUCDVjeA9a5y
0pOJ1iX6vc309NkGWzYz7G79nXm/xO/Xf7ygLEiyC0fEVfz3MDfnyRGhgN63HGu/DwYGEpDiN2dD
wW5OeEaQ6hu6neX5t61k0Kr2tSPc2eMm0f1LWmJKUynmXGRk2FNMKbfWfd62cWjRe5Hcr12m12B0
FwrVaoFXvbXRfUcm3HwFnm0kYeeSazZtvW7/e5jxh4nSIcH/yqwycj2X6poa25K+0hVl4KnwN2mV
ZxGAUQqAGC3gC3Py2TgNU05igC1Y03kwR6NA3tRgOGpPacnNIjn3ro1m9G9lG1Q6bhTSiTdeZHsH
ITsU9NhwmgZKiVPG7LXl7nvIY/XAujmLcr1Ju4jIeNzggryVjNzIneL1CmRsVHHKs3hthQqwWKyp
6bNeUGMi/mOSaD3rfI7St/V/yFdtZZEpD0eqJFwSnDkxcAMNtzKlr2Wh5Fi2eaR2J2d0gIsccmMG
mquehTN4AuW9NG17Oy3KwmHrgrWm/A593Au2eWXkTofw8ombjf8I1YAVCT5x5KxGwWYCX4h89/31
jEmGQ7vwDh5CqeRntICVDr8AUr2HBdiZPzjykwcLoCTl0qbvPyzaQHuEs4Rs2uQIZg1zuRfy14mm
efo440PDWQ9CAZzPMyTXo0UBnuvvjJdhfRlfbuE9T40uWdt7EFahd4g+PsX9SyJfnlen27V66Wmu
3PVbuFOsj218rZn1jiKmqMFbr++vui08WL1GepK1pbb7amU0xpNpugeNLk1TXAt/fV6jdleMZ8qW
haDc2C1cCqcpq9hSHzVkSIWMtDKZL+QDRcKZSVsKnjcV3W3pYcMPq+MKJMUQdeoLlCX+dTRX01JY
xgjJ3+f0Hos4Bp52tYC70Ured6nWW24CMvjrWfTHc/xSntdkYd1aMR4E8bAi19feBNfXY7TY2A+5
jzy4JBS7m5Ej2MGx5X51LGVYW5Q1+TYzTDc/j6gahT9aeTAsdbO4v15ZA56H/TNRj9RgJV17Db0X
V8+rk4c/ABrrWE/Pda7pYjlLG0s+iv9G5HxEaxOuqAcVGN2HvyopYDt1pENaolRUBNad5gNkIIMM
SQEZAUBfh5r2r3MLgc/U791gKXhZz+W1FvHeWGx8UzECbbao78CsW26P1GhI7pdDhEOEvfkIqeW0
B9GD0Jc8cEe79kh7dPGn0m+1NFKjjuyMm8JldGoMhSHvzO1t5wq7+aTtRmK1Zd/+vDF9Leteu+Pa
/nJpgeM2ZjJYaa44WSd9fG83vBy5uDtMEBOTi9SwKY3Tv/XrUslD5N7Hn958eH3OD76RSdZxzPiU
qDoMuZe7IMMYGFI0Z+S5bxTCkhYNNRA7AfyXHh0VbXyFLyaRgHQM8payeFBszLUZXDGnpUws9g6m
MAC5AxdyKXptWlwT9DxZtZxT7BuYggY15VGOngRf5ur1YUZmXNjUVoNJtQys6EjMRMdu7q2VcBLe
Pshn+hFD8W/QM5mQgD6bghPxi3P2KS7Ga+kXL0nhATlra6xXcxAsk25aMdZYDOBDk0qAMX4ZBPcy
fgE8sSwR6uxX6ZjegoFolrxTo0BVtV/Gho1D5sVesukG1TH7Y5oLkbSOLNr30FA8Qu9zxS5vGBB6
a36wHQu/BwMYYDwTQkKFWe69v5LqN6BbsPfmkElJ47MnDdA+gd1zp/tMkQwYlZb6qMBf6nv/6nII
STif3fs0jXSAtBKfodqEnldz2aCHNYjgwvjvFnmBZ+QzjU95NBaBGbW21Vl7mynev+UdzEkj1OlE
oVXxNRKtKl5Cp3RWeIuvqfMwSRGDL4AAmKpXO3cLVI1cztzpbOSxCw3xCwTiU7GZVLhiuN7JpE9v
qOcVaDRl/eXSzakoSfpRMoqoRfzZ3G8780WjBDw7xQ6uGPu7VhBR/696vTCuHpRpBXCY+g6yojru
H6ZyltNGcOI6UYmscUdmsPNsuBXCzH8zZFMzVV1NoqokLJZmbgDJe37kPDcmf6ohtRRGGRcfyaH1
H0imvdXzXEeUt/cj2g9p7iePhPZmsjWIFyKpn1olxMPwMs3PAoltCIBFj84RQF0naWrm5VgSNBeZ
qSd4+vyIXTAu1wWonG6hOqR/ytuToTCHeBs4vjpM70WYfua7QcJ65V+Y+0e4H0UdSUBwIuYTmHY7
jj1olH1j9RQm+Bfh7ZglguOHxbwoU/whCnDP8v3z5rIfJwW+vIj1lbaTVjTfKysKSp8toq3ETZyq
EQoJu1wpr/SqrDUYYsrhRknsCYTyw88gR7ND0wrJcBH0Nm+ORWU6rBxZnuXBfwHTYRCfc8nF+H5N
bIK+3QfOTwp4XJSNDS1IpReDNAwr8DMJmiarDthWdoOSRS28GZzEyHDx2alpU4DrIBRflXUetqJ7
0hLwypaVxJi4LtPtnvFl/gwsH+NPxCxX2j5rqOWYw02Q0+nAXXriG7nygF53JqanLFOQkR6Il5b5
4fhB10k2Cwb49/WfCLkc7HQoNtSpaOFX8HC+a7cd5FAyvmylSQ9XzowEu4V/cbjz2uDm9GJ4ueqN
5MHjTds99k8f0oyK0X+mBHhhB4BlWpaUrVBA5trxtobxYqZUR6tIB+NnQcwlTXDA7P80yNnKl0AM
WJRk0vlj5/Zslg5Vu3gHQl60dtoP8l4XGBPFLxseQRgd2Mto2bqw3WdzLmfQ00DONFrp94iyxdqv
Cd4mNEfHiTo0zsF4q0VISiWdK5ZuJKrWHVVBReS0fmHG4tDszFhmV0H3OyHDwUtCg27R2j3JBDMz
K2A1PJRv9GPf0+zjI3/ngNwn0FSsRbqwrPxDnp5QdHATlt0vFqgxL62bekmXGpxaAyTpYHena5/7
OXi/GA36zV0IKbfpozBqrezw75GewxoWRr9Z7mEGkRB00wXyH19v7RHioJNPgxybV9BSka6W9hDc
i0Vs0aeZAm0VoviGYJhLeaL5J9kDSkX26G8rjIuS505ceqdjZ9uz5tPCfG6vqMdRtvwNgZcqgpK8
1IL3SVtXo/5udo4djbclmtVgnkNprIRF2fTSI1u9BuOv4Uw6zj4GdqN8wQJFhlNkKDLbm+A0Fpz6
h8jomM+iH5msX0wbikMSHM/oDx8L9dQUhS2qIUgNzyXJe66H5Dlip1jX07gFnNbh6N8Tr6QPPijx
dxA2uruPxvCDdIAKhZZmew/k+E6g6LQNTlpPBt/q3oYmhqUReBRMmKtq+jqO8fO0ASXUDR4Q+ah+
+Vzq9xMSe6tTtOytugB2iAeDd6Rj7Kui/m99UmJrNo6u2kaI5WGS10geWCdaI7gUR9IeBKIFlWvq
+KGr8fFuYgzuM2Oy6FjXrrNTsbZo7I9mUuzepL40I5xuhbY1sGx7ga4Iewj+6d/7cRYinrK31+Z0
jPE1+oI/G4+nVYM12ySnGKbS2cWk9XaKPhB72/C5awIzrRsnjKTOdPqvwRCIYSwaUE3diHbk/Rk6
buMawkPJnFVh9QLQAloSUHV+ghfkon/sN8PK8pNn1uqIZ4NhErXx5YFjjdSLNa2nKiCKfw10NDzr
fT2Pg04wwJXfpXthbruNDphJy6I8E8aU3Ps3aHxGNJb1xXWEQELnvEEjq1duZNX7hLBIWAALof1H
nDDvyrqAGV5zxQtPVpWK2XLdl6y0rRxls8JnGONsHCpIGL0Liz6heCJB+lP5kYxRKG7ekPp3LdJ+
uo1oApZ4ZceZUkiuzrlfvTFW833hRRlvrUohVuU/KAvBs2XFDf/cMDP3A/4d8wedRuqXsjE/z9Ye
M+U8ygXYZ1QZAwFt8aP2yfTCXIBz1F2QGfQyHGcYlcLzn6bJGpAwZxvt6vfRZA6Ij/i5o7tZnAY8
ToMshZFR67zKoUgs7AS2pVp/6MrAshLwUQMyn/IA8iI4AsRYSq0LRX3b5qMkY2kql9PXuFeqffG4
ila9X1fRxUCdix0R7UmOjIvoyN162VtYTwZn0mVhVMsc4iRHx6Ya6/B46jpQudmHHZcnh0eaGyI8
zP1zTuj2Ltpe3OAbB0X9qFD5Oq1WLwV+LbVfTgeqeV2dWtp83fwoDD/KOzqKYLv94sRTfmeuHLlb
O/qknMki/N0ujasPfBsEYZXiRfREM3qE/Xlbp0b7pidTexTPVTwLxbVbpQ1vDwSw9h5rEI0Jc8w3
QO77x0Yaa7VFhc7AiFr0igOX91wsvMt1+MXBBLFhHxbiALdqGOk0OIgM/LLaM0LzMvYbQheoauNz
P+lYB2uSDNPawcncsTChH/KogPx2DE6daTIPUA0YMSED0IgYY0iVg3wZhyAjZorrDIexVEaB3RKV
EAKZ0YavIxERTKL8wrYp8xrt3+v1MOt149NZcQ1CSZDaeAWEwT054QROcbo4u4UiHRf4aXUYrQuo
0BQkGvA36PjJUA6BXmlL9KnDqB6Ybfre/j3vAOStJAoBGppxh9ko1NmIjEuCxNqhbckkCtjzmyQN
oD7CvJyxNLhueof5meQ0mRVx0NeihUbm2pY9jTxkGPWDlRz0gTSiJg5mYLCPvWYO5VwOYfj7rBSw
GmlB+G2BJ2LpkYIQfBUoof1FGlo/OZN3Z261ELM4ZLjyEXKnE2bYJCjO9PT124ZMPGhA9gn26vjv
e86N5voupflJViZY1OIDuXRgR+4dbb/Du2oJ6sRadL5DBUggMslEMwi8OceSTry9GtUf9kJu4Jrl
Y0fNgMHHlfF6H/9CDDk14Y2WP/FGhgJR6qimMdAeuAk7ZFj1qL1M+sjvcuv3PhdYvx99/C0BsLWf
eJASJGN0zpys1lNJjVTMB+fBkSeU3tW/NVWnhRrzk8RZAJLEluEXP9sCtT6tkMyEiC5qVemlWYL8
d4S7zFd+Znv8OXnzgkQG5OgfaV7uravctWSo/X2ICbonm+z7IgmVhHj0vG6UHx0DbHlI06GLt9K/
7EjtE55TuJJNtHkw+L0eQMtoyXzOC+yks16G4ll5qJDrKmRH+m2CwHQirVhTjc+vZzZwQc7O2z4+
2aCfqIFK98BLsJHxS1x9/U1q2xRZh14DKWzwxvDSjL/rF7SawCpT2tb++CpAkF80NETpMkKxCVl7
vTgBB+m9XlwzgJF/V15PyEullTTBe7k1Yi+Y3e9U953d1G6XovXYYpfkq3hSi9tlVOV1fBkdPUrX
c/ueGVIFz5biV0pybr97KDtWYfNsaGiqp1YN36HzsPrAQPhSZsLmMG+ZUPPIoZnWZVlGSyQn2hnD
TklUQDgieS+lSu6MVmlhBDgJkzXuPBNqigA/Y5El024fRR7YWqi+H13xNostWsT3pQAUnKbm19DL
9+wq/jL/fYt6JAubzhr/ofxq9OwUEfRPDnBSpGLkypJ3daBzwyPvGQISYEI6w1dx+2lkYinJCjYx
iz7RHb2lHHwuxmtV9s4ObxF33ilVhqtqZMUQIMOrKBLJ3G4m5TJvnNDAEtOHuDIEw1KYqodx/oL+
kO5qE4KrJiFxuRwY8gnjmQQpRZfTLn7qQ362208DX8EjXwWdcylf/gsKeCLtzn5zqz82RKAeTqum
ifugyK2Ubz1ol2k6O83C/ubG2xhKfoXeCv8AgR4sZ8A41NJLC4ZFM+Zr1rOMuaqlQ2SkTwl0kvXW
WRrPEbFf2iKapxiylhLXWdFn6CFpOwhSN7ZNso9rRLW8yt1m1wUpRVCw1aQdHX6y5qywmzVe2b9V
uL3BxSSaaUzUQRgVTn3lGvLl7P1zkXu16I5Ql0ALRp4ZSC37/wn/EMv7gcFEm2e++k0xSTAAIuYR
/FScK17F63/OUng8HxfESow/LxrH3IzYuEgN00LuiOzC3ACF8dQcxv9Nec1PtaLDGKOrsE+Rsx+S
qAIz0Cm1+iMU47Eyzg+O97DHjGUUDcpyvPomzb6CWSMJFAB5RFZc1Y3JzVPCFZf0aUTVQgni8w0d
kxfa6ri2fXR16rbDhP45IqEnIEorWUBxJcHow75OglKEHdPCxaqR7Kd/Db3ca71quCIi+vGXCiT4
U8eTjAeVHKPH0b7PTipxMbnGbgt69IjZzmh29Aw6SaOr361W4Pk6KZ9aJnqr35kUVSi05q1oi2np
Yf60AuNpnop6r1qepzLZh1um/fDp8vibtThapTusY0Ix9I5dkK7R8EJfdzP937jgB6i0nkF5Jf0k
HuuxE3Q5SjcpWB/KHFYg8cSTCCv4Gw2W68ViQuUKzRXTcPwEZO2L+WioaSzn6D5cfm9rNvqgm/rA
sP4pzIG4pHa4UA2JIsZY/G7K2YpdI+wOU7+gvesaFbwawsWsptjXJ3/aiwLs9YIp5Lk4rpCFsmHc
WpEEz9zIvCZasRNM2dIMBHXHyZc2QWH5lcAII+kJo3CNFcFUYNiQcR2gg+InF1tZbUqw6fPQmCwm
z0iKD7qsC28vTKAdrJozxVI4fc7Hae07UKTnKkBEG2HMgYXE9sT0qdZyYKPaDl/Tmx+vmdOcfGet
RKWa/hNoU21HbznkN8m4CFZTC8kQWFNQ8L18yKtCPK6oMOd3dzMFkoFptO1Gny/CEn970Egieyep
thLt9m3fD0E6H+Vavu0N8BOH/RNT07MXJwCgzIdCjlIXKVdYlqkBbcPoSRvGV9P+xanxzbwG/wLV
qJzg6XXAHHAHFJ2aGcpAnG7s8+7Bc8jTXvdDxlI+8zU6JH/KLHDXXrwVRa7pqt5UcOftQLW0JRiH
4KE4S5+HlRzsnmBDslSq/zzfbProxm0+Prnsjfb5OYTnLuuog4ztonDOgc8jhEtwM/uq+ST4Al46
uRPuKUQqQuMyc87hVTWxR/ySjXM5lTVpNKPmOem28W3lbyfxqIk2WOc052y4dnvFJvjRCSCqUY6m
5rrbEULe65HY00ZEiYpE5KMx43S9eakWoOzw8ZpcJ1fF/WTIz9wW3EVA0yp+x3Kii01BmrZnPXuV
Auh26iq+NvbutJBylV7wwGNAz9PJET/9K7wHUGCblVIjdkQkk4zyaDsy3tiXIlqKLNCiZ9DI3fzm
hI3SV5iMyl/XHWvggwosd1TEW0c7gpcptkSS/cQKOX4zvIGgIIjuH3ZjE/CCyhrmWVAcXpNh68s7
K1dGc1/oV2ALVUp5Ip32yKhgZxXVNd7ow9QbUmbA1uN4sqmmFlABIfwJVFbn7nNVAzIoxff4XTRR
11BXl1/jN4WI2Ahv361rS0NI4zIZYKVgs0DREXgxB2LHl/pJhEkB9bMwr01lX2IDbJgoEyHyMaSJ
KjZINQeOe28uNKgjMpkKGueAUhp71AbhyKdHSwUMFHQwxwJF0kk7ky18fG9bSY0CeUqMKg6oN41Y
YqA87P05txnXS83RihYwD8ic5Sl0dB1+v9WjgR9VygMuEXYIgir42O58FOjRrRwJdOZjol/2PMeg
jtpPDU+Ndp+8eVOu8LXLjT3eUDWZUcy74J2/xtYBQ0u2sTBxIVQp3RezMI94Co1ju2p9V09Vei7h
sR2Tg9n3F32j/xby6zgyTTb/+8ybHYuiX6zx0T8lWr6nfQYUEpZ5APwDPaqMvfrLLFi9pB+2VUdu
MmYvaNRc4VhaWHfVVRExgQYBTvdZESYELDh4Jr4hdBSPao/GaNxH+rRdWrgiDcqRLYQyLrMQvMjV
9d9b/z/mFlG3FSqxwbWFsz4jb2z3U9e7tLAOoGqlSE51004/Hu0FSa+edijj8QjLi5obDtO9NWH/
hBwHY4EYT0x97WbICrBtQUGuIHz+eR78jo3NmEZaQAgqnYrP6SpkuE/3NdD2JxRNzNm9mdqz0GIs
Zzx9t8f6Ml1fj9y7AeV2FgalQFFCiOFEbLrBYqj4xjqKGlEVDr/w+AuR36jJtaLmTf09yUKfpZIg
uxQd0RlVH4PciWrfq9PW2JKqIAlhh6li465cOBHbxnGsJ5TK3uCXz0peXiYxEOg2iZx+3oV44ZaI
ZInaI/0Q4Yh7dii7GgigoStRDQ1fOpAbuVOHY2UfQ8RD9Y1KB2ncfTUGxGZ6M1Z9+0yfbmRUARqR
NDHcLF2SGZdBMlRbbACAPDl9oE7I+vU4Iq9JWidkulCoXJtk7l61QFg4XkgH4eMK9USWZdi1a18G
KvsOuGx73/PYww5COWMkBFzDttpC9Q6EVa4/Cqw+3ZNTfTNXIY9ciy2AQl0+cjWLuB2sh+f7WKkN
shCZQeT1Je47gP0i6SK3fngboyqyyOs3k0pw1GAPBfsVmnTR+9os5rWppaKMjiCPhngn7pFbBAot
N25UXye+VxolCceHBIuqP0drP8w/1Ta3CnOq+wBMA/UkawbtWoPYuaVLnq+vOvGylLPc74+vSQoZ
XQBzhU1VXdJq2QAOwh1GVvANIjd+3vPnGeOHQu8doQSN6xh6GBWRZ1UA/+IXinge9bgUw1B736Tk
9qLWCNbktu9aiDskeezJu2i4Ygbn+mCslguYGFCzUaGm6g3AiZeasZqyIcSKF0KoUdGsO3iv3t5w
2KRJGxbxQqpJknVen+evd+D7FCVAi/zhOruT/8hZcLu59a/szrK/Ql7prZgOah3IMcPmYB3Msqre
s1g0xaQTIR++Cnhqswc31lyFOob+R914UyxFlQNIrdSJ83AESC09W+ggPCv4J1XPJMN10rxZ0fqi
TeMK1tAUbZuxj+ALez4GEM6sxMnjco2OkB0DI22QhJ561y9LytEz7rlaj2E/DRMIFQUTyqn5nura
FPXadLYfwJ4ZVugiQDTasdJPAoLyk3Q/XjQIhq+lekyH/pW/3TU+fkqX34uuOu4NneA6WFrqE4FM
pMocTUaFI7ej5CcYt7B2gN0hk4Nysvf/a78ns6+Hzy4ghUGBzYK7Y1LilpvtHgF2org3S8Jx6sUW
bJD+3ZDVt74PoMBwhiIX5FYa4+KtTRDND/ymUqYRfxNSJddRZUvRdhKq18ReGH4oOeI1ioM1q2/V
lVXFHwxpxHERj3fBkyKInNdzLCF88Um+FupiTuCDUERVb7m/1obcGjcFAGwVmXuV4sCd7C11JO4X
twe9e8eB1qIMVcTMz167SpeQubXAy4Kx6XAkjcMbotH1rqtBIwD9QvvfE8IQBTXXHU/b2AzlPnrH
p3VWFrHaTyQayp5BFEG8RUU5luJF3MeOSgTXXxNr2+C0PBsHU4SbeGU5OGNqwlo/8IHncILnxgDv
pMRWcWsMfE05r5CKJLYDDAODafNOtSZexLeZrhJntsW5E3DnMnEUbhZe9+y0bXPXvKHeANceBjfh
7B26WJ+eATaJzX4A1U7JsgH36h2MlYqOeaaxfBd0MXY5zP39yGY32KIZ49qyNb9DH7twL7hCNx+4
fb73GTf5EjxBfwQH4xHT4VEOFJ1FaF6+tH3/NOlsT5DnuPqdxNvdqsZTDia1V/+DCai0Bzb+255s
0VGW5GDW12+23zRn02tpHqX4i99sfjU1vkCpaYCoIGA6CPBamaLMrJAbyr6RPMR+EftEYcnusZlD
0Fh8ExtQgFJU6XVaQnGEbamm+FYCUEnsvkqXxdc0TYhcvcc1CntLhVyypJ2P81c7YFPtR8ehF0b9
di+dUJmvRZjboBJO9jUePxlIUERW+mzS0vVJmZ1iagCJ1jweVXf7C+ZxIgLZP8YKwnayHICoDw+A
WFQopgi3ul7HJaeRbdIrokYwlSJshNpeEg+6G3Flw48mqB4ar2PHy+TBiK6qAew+Vo3JJPD/+ekC
iuydDnPko2Wob+0vNNKpJ20tojYFeJVaAwNBgL6ZzBmFCoSyH9+0nQo0k9eoc2vBfcan1YS96vUq
KnlrCi9t+J+2VzBY1MP66fgKqQYFOEXAazS5AeOT8LuN86jpKY2QcojXnNF1nTnc623XK7/uuPZt
71gcXgg6VEV1Da34Jn+SaW31foeHYMwS8RnHMCWh4eXBP+FXup8wdaKjFmuLIoBblCRx4cYzbmpF
nrxbBDx/I/t8FYdaelrYg/SC/YEB8cMmFmBToWwtBhwvYlH6Ad4QuAdggXdFZE7wB6peGodZ/Jsm
o7DQ5q07zEYwBj1f0r56d9vklm/BYC37G+szL6//2M+wAf7/70Z9JtDbhehk+fXGyfyBq6ee2+mB
hMabjq8oFilr2rTc7JMOdm8qf3JfAF6OjQhargKU4dzk9fSsKq4+eRttshPGAVkcB+7LRDvl860v
tJlOsbAmK7WtdqI2q4FGZo/rl4PPkWTSzRznfjtPRLs8uhFz7obU5w3TL5VaNVPvd17Ypo0I04OG
H+E3T+Oja7kvyr4nmVHhTX2MFehRoDu+iXLwxFP94Rmh5vR9FfM/FI3zwzE1fPkeyi/8wBXU771b
mgccQJTXYKJP+JB42horamR5/ksOtTSIr/W81+GlLxFdFpjrUkgBQYMaal1Azq+5pyPPL5HSJctj
tW0FfOYD3sc/DXy1fhE8mAnPqOFCUp0KxIToRpYcjO171DLSA33Ymo9ZxIb5/jMW8mFVpNH3xAYR
/qa4HzoPj9S9l/So0EcpdRrQ6hSScQTXGDutOzWem5t+Xk+7+vVnmR5n5iuRjdn1+1d29+3t3ChP
V+dthc5FLU2ri5rqJkLuK83BH5zH+SR5jNJt+rCpQXp8KjA3nkYWfZoLFVn3N2jEG80+IGIL06LI
5uUsKMujyxZtMrlCemMvYaY/9l9rqFvOmpFaolmx7fSMVFgi/mIqLRgGBbSEukgG8j8IifWgyaO3
mXzzBvPejF9OCedgepiC5A4CJ1Ysvj6nzdo5nd/cYVHk5mQwkkcr1Q31gSyDKSOitLyem5FUHhMd
0mvswOhHwdyG85WazikXs3WU8WCqrmO8S/Efquh4Stl9hm89TVAFewefkfzNA3n4F3jFzdDyEUdy
1DHVtlKjvCCD5n669DO7wrsXuK6i1YIMb3Y7vfpS6LVyDXUWsYw8tjFx6Z+qnr8dwMNlTyxHG0Nh
VYSSpC87Vb+738nxSehB44+x8BqIoB3soASyeXkH5p3/I7ie15s5RjEbXcdzBk0wWgJjGTeXOvkj
3eFuZ8QTE4EfC5hy7S3Qu3JrEHCIljhqmOGJH8e+EwY44zPmDBjbGVvUMBCpHUBw8XwYx/AgSA0L
S9YRfs95MDGa0G+DUYx1FdwL1IoY3iz8ZisREkmYIeJzi3wdpV4qcfgsFenBuTtqBFIHGAobMnt8
Ela2Swyk1+PD55H4mfCEEejg7+DVC+qCBx7MchVcYUCEMAoc/FaPVHVFPHbEeZ9NchyFeuz2DWkB
dJVW4KJBkLtToLmcvoRV5pNfaNeKW95HcS617/Q/nRfQk+D++kvNfKVbyG7bmLUBGteaOqYNe9oP
+EdH9revvGNwbLGquT0wZjFofkpbF1Xx7zIxOzQ2V06we8Zl4aJlme0xAnLCGTQQo0fc1ZO7bVm9
zCH9mjcqmcBDZ2p//ENczFo2AGpnmKJzZRyqJqB7WkaUJ2TSyxwBo1qEipyg5SA7w4TNLSECkGIp
j6A7oyzF4GEuaJNT+qJ4tYXculZEs+NijrOuMBD+EQgGj/l7OgcXOVdsFRGZUk1yht8yVQ1KmX3k
0fXNoNyPferq7fRLC3PLJMk3iZVeVLS4yU5nxkgAm9uwAjE/F77CT/Dyg6hFLEDIUwgBRDTAdenU
w65lQUmbQJbco+fXEtDZZN7KEtyQnykC4WKFEXv86OZ/8ScRTpmrnEW4GYS6zB5nzljMF3B4sahQ
NvdALIkR99/dlYrWVthCXjmitbkRcDq4hiDwSQ4l7qkd2Ey50ItyL+Ox3/DQZ3gZYOO23xC0P+BF
9ENj3g9Ig94XXHrpWuN5MChjUUPv1OGLj4ZpB/ft3X1jdUpssc5wGfdSnBOwFoSfnXDBdcREkUQt
yxAWXwn71sJcgz/pnfmA6FRxGGojrNlWx1SdPn8uVIOgJeLncds5HB65i6nPsyD5+FWhOoZHQ6ti
CzBn1WRT2dpKh1QlJuzCICfzULH9jGfs/jHr9UmcGZlxeXGtLIFC331+G1eh9skZZhXVXLCDE05v
CHzA2zFgac06APK86G8i6TDA+hUNPdfAOj+NVzvQ4M+eBBNqGdAplbgVBjNczQfeJ6VTYbGoF2mK
DHTdeOM+7LHvu3JM/uBEZprZAFAA+HYohjIAEA+vS/rJojSGOwVnOhSKyTN/jlgmpoOistSpzWK1
Nt2dBzFRCe5V0iSRgWdhcv8MYfcFPzpQbpgDCoFalSJmtglaUCZ1is4OfEE1c/KcS52ERRh6JLXR
V8VR3LFkJbXxBZQJJTdm7QGwPUPmOiEwG5XFviRIRmJ1utn/ci7s3Wv9Ck/Y4f23KRusZEI25s+B
MMDAOlP2PmVsAD/NN6Ts7tQcLPatS6kGB5TXbaimhQNHNIXllhX7UlGut7zr0Sq82n66IL/r4/7l
GGBZ/63lXiVqtYy7JkhqQG4xgnZ22Z0lwsLZYEhlGgpUQImBMtcALwZhxaoIW7QfZidyJQs8+cdo
tOxz1qQPNwMzrRLZWgCmOFRXlesIo+36m64LFuAC9Lzq3m8O7uULFo3C/mhEccNPpWgV+yzmzM2n
GLaQofVT/nCCz9WCETcOtjXSxd/WysAymCQyo2dTH3nBVAFCO40OlYgopiwBUoZKinzL5aGj+8pP
tft1IdcXGdL9XNFFC6b8TZIwdVW/Bfr9JfcDfDqiUb/vzr+PpAMlwU957aCNimr0FaOX84QDP8tX
OZFPQwB3kZcJEFLQ7rrx2pqU+wbCfpddCUhXwLc9WzdZuIkiecoz+JaYbOoZkEBoC4eAj7NUIGwa
hG8tPwL859ktLh224wtKLJEi3jTwgyOpibzxWeylY1vm0aAA51mm7VcpkxCMzwWwdiMYT0EBxSwT
ptpkPQDxlPGelHsaC6P5n+XKs/gSCX/lc0fKUAB+8VVFSUxS58slLLGpqPytyMTfAlStaks9lzWV
c0KtGmwljH0jKDpBrRJYGVKdHtsKKG9UldknBS8KI/mMXhBKi0rGk0PEZ0GqS/wynu9BaJ8IJtF5
juykjUUCN/hC/cFdYVYTf8tQerP7L4A68MBFK4LD37j2Fet2qWCfIL1WVv1UgnHmPSIhuoh8MLg/
S3sY3HFwq7Lg48wKybjneJ3PgcpjLn+YEOktLFyuRYCMgcWlv3Y2JDzic+cJpj3DJ/q/m5UJLv1G
tWQTwkARqgQ1hfwyTn/vp9Ay3wUxX2XjAQFpxOIbTweLv55HkPYpwPT5g5kr3F7k4/v5qT7c1BHH
KlLfTCLMGgktc6p8Cv8B9xFgqabpWWhA7HypmPegYyYdHKeuZ0JKpdoExBYLyQe+VFMV+G/8oaGq
DWJ77J37HOG18jrTsXqEid6cDShBDTuIJkws5JK4QmKr2P1vtKSN3N7gmdI5mobyq6RoPsXAzz9M
5Nzo7Kpi8wt87qR9E8TIeVHfOhaOHagOh2KnzB5zsHATbMd9pEU+1aKdyCHTQPR/nc92nQY2D6MH
cXb9YuIc77IkF13oIdbVHMaOBwTnKkq4piAk/LzbYReCRvJv04v6uuGXlzTxb6U1y/wzi7aiTCah
etXwf4NFdSVFEiiTX4jReBRw2Owugqi65gO0DAI06+kg9iJb0f5s5KxZgvGjQulDtuhl8X/ajAJK
GRBgrBWtL4LD61pv76C8O1mZZoE8tjoBtypxSf9sfdXBGwYXqRjrHGHrLZrBD0xtaDokWuNrr2hA
st6li71PL8T/BEqcEGqtSHYEjOx20G2HP7yocFpl9SgNasoFykFDh/HeolS8Erv0wgcRsa1ciawG
6NDGEDfR1rwWPCTx0RZHfWCDnpu5XoI6eIVyCxS2hoIBzqIQt4EgiqhypR+153G7auo2ppEtZ5FN
2gbCb/17Z0D9rr00NfImr710I2lfXru5exAqF0e2ZqQ1kqqLL5w4Siyfuor0tnRbgyTokxBrvutu
8sxKAxOp4GJB4Yr9iF0eUVwPzO81pwydu1JMpqPyrQ6fuUuM2TaRO0jupHd+ezoC2y7tajfcx5Ik
SR/rARly9zewztatbRcAlPLiHQy81/DpxJwPb+3PuIF0JUTvJspWW9ba6vtNW0GfWY2duUnphyZK
FgsIJk0sKCh+LUk+b6Yutx3PzBtjzz0kqMysLMcxMJ3sQVREqQKUuNn9Wbo8pL0MjG4DDftcEiI8
1uOhv0WB8p74mRUzPYztCgwGtZVxU5aUFwC7f9DiRDRpwNLfqqu0GNWfMEiuxaWA092g0RhUOjGA
IFY85/3Z8gCO1QlaZB+BXCo2xZtpkGFDcjEg2anSCK1Xf5PuirnwnhG2ABc6l2YbDxcSDxFS12FV
zPjXSQZYjUi4c1qQJlA+8mrMZ0cFhZqhSsrvj95YSdqWLWt1O7OYHsxhB+CsmpWYufJXuCEZ47ep
YHEOFAD4VQkkF5PUUHVX9ojMce7tvXwtnw4fyj/kkFBtlQ8bSX2LKJlJjKbipAWP/lm5OlePgtbh
8oEkKTqfZgKrEraecPh00uathVhJWJvbd9ctG8GSCxqKzv2tYkonrsunPnfvL7Bo6NFkM34zV5CZ
NqPxHpTZLfZIxPNR054Lp1FEyvLI24cBL4ipq306CzqF3iCs3EXTxFBsrVNA4M+B+fGY7VuaFsA2
hExmWTiBRk5A+4e53anc1I63llnvzGOBovaL76UUzUe4QqFwHBpWr3+ya76q0+2LeXbyfmtEDIlK
cDPO1Z2b+6p4iDtzqR5dnJ85rDAYzuxeVvBdMyBouywjXjmyshfJ0WJrYGWoykovQo0yyOLH+lyu
1qvSX05gU+SbUOe8frrEQBJoevtBNTTjRmKHli5v5fDgfJCJiQhE9rabowqki1sy9C8hnOcOz4i1
9JIl/Lmp/6WJzoTt1DEWTCHV/NEb3HMMcGorwJ1g2wwK1UOMPKY3y3YVllAkLwK3t9D9D8f4Ep4f
mkZ2098H6KYTBpqaUx2qQCc9Qz4/AQSut64nrTu9XPFjISLVtv43LJRbtEh6L/T7xjQFRC6ydt4p
+8HIWZQvl2iJaj1BmK26u/xvkOdmym1nd7R+heSQQeapZYdz50i8Hq6baIaVD2JwuR8A4/9RG8h0
jqNPZ0Jak6rZUoYJcH6dBukhiCgsWU2TCDWErH/iCPF67peIhEj76F5v9VqTG7QGfazT0OHEXluS
jFttP5QdtI1JQHtqKwJpuIhJptbHNq1Aqy59KFsvdCX4nW9Suq/nMfu9FE8GU3daYZiQrszN3Uc+
MQmH+qxgEY886Gx9PGcoT1dzPCimvhZYystSqkf1xlP8P1yjAMuPPpYGx4io0a3DFaguD/38V+rf
2U4WlDP4u6DO9CdySuXK9E1EdFo0aMX/iKULq1JW8p127qTzrRfQgTMbPZ3DPv2NIkPwZzmXDH+d
bde6fIQWSfCk05UleoMiHR2uacdFqk/JZodYGBPVcVSkYgUBraD2VYC0g5QIBO0LwiNhcYyI8q+S
tw1vHAsT0k+jczkAoWtGCtGha9ooKjn28QTBhIeaG8KLpE6JabmF6VBLWRJdkB7Q0QjydzOL+dJr
c7gABOqeAYICpLBTH94oDOQ7mKlazPAxoORYjtunuitronQBQ8mLIrqu8TLhSgSJQVRzb25CbHZA
8l6HDtgxAvsgT8rCF3CQjE2PSTWAsRs3rkcf308JjOP+neISNboKFFZr4Rm1OavRqK6DEaeL/cq+
fW2s7JsHmKpkx3ojl1m3p7i94yQhh++WtaLzn4P9v0h/YTB1ZyReiIa6BFEWr9TUYgtpmfCtrSCw
YGcL1HfRv/Lp3w0CWt8kooezGGzQ0FfGxv2CaGpfe4dFiMcsdqTZM40xxqczLJCYx0cgrR2noRbO
fsxgFFpGEBxsWyCrn9VRN06XH1iGzf+k9AXr+yGD8dO1OBQtGVh+uyP5EFJJuQ4I8RuyQrtjSn/m
ycrm74zY4WSgMOjBjc5KQxbYfwdlPBtroolcMC5+h0vSJtyF/jDUtMO5N9K2BupjGzKolUj393jz
Z3p1TRfDuwbpwZ5ynaYAsq8F3RfUKV2xaqRj98kQNBHYd8d8eS9wnTPca/lWyT6HRWbx6L647Do8
/x9TFH61VS4/2lWriSn38nc3BnlyCxQfVrjlxmBaKJKAb2o6mRORM6lYGR+jXZKmKC3VgpBz8r7T
Utv8cSFuU51EgoEQ8LNJPa02qo6voi6+Ochi5vF+8opMs8Vzhzk9bo4cu+0yFmNWiUW6Ubu0UEb7
mEqPi15soCns5L+YzQ/UtjLIyI5IV15Kv5Qgoe/VK5MemWHUWy+RqV9BdckFZo6KyTR0x8RfiDG2
P4XC0g9xg8p1drqwjhKjCjtoDR2Gc0qc3HgXUwxSZD9CTRM2aYzbf4U0p6CD0rzwdUTJ2LOAg2z+
LYZTiNK/e4DHP+mCkzWw80bPepK2wvUe7fLLOeAJJWVv92p+OiL0hpn11hlXpQMFTcG0kqMdV2ET
oEmA+cRHd7boRqrc8mDVZ9kbW+Gzkls+NErZow+5ZzjBfWr1yLc0r6UbYyXG+d/a0uDTrc6+DgxX
dspy3Qw7Bv2kAhDQRjDMcGhRsdXhF4ltEy3U76wRGyhS21NHWYrPIpQT6XYxvya3MZ9Vm1qCqse2
OQ2sOgl9MQPyNi55dqnWswjLUnDxNR5H6l9zXcZxfcstyVxXKTqKQPSF3c/ts5GQX/L7h4M4fldG
eqnRHMZZUO+gkaJrwdmv8aA7OsD0KtyscVB6ZYzJkT6k/dAk96AMrsujHT9Vwxu4oZGnKI6a3lmQ
+sesVzY+djLFP5Ma2cpnNzlGbs8giSXCHfQ7SmMmcfgJXd7yXW0gWQFU7HyF3lr2DJBs9aswFRQY
CbzV+XJA6EHxxKBBcxR3JkyoKIL08ZL1CZXXoON1nXg9G+bBXMdQdCnSnQEx+KKwT0ycZ7l1v25l
t8sWJc4tsNEAX8qBnNiHjC+Ue0Tkr8nskuH0z+7s1XiUOrD2JbtpEnpsMUKZlUvaCfb+8mTZaR8j
G0gaQbcVvaZf8Z56ZBPaWXDGkenhYKkRzswD7BJOn7oCIVEXtYHNh8lWypNSbiucUoJeLf32xhWF
iUH603yw7zr+A7d9m3bxUwr6zXdrMiUIS7uqVhrbv6wd1lEEq9v29bSb8pdAeldYcIj7IAlSz7cT
arUaOt/w1gMHnifuVA4mfkK/M2eTRMzRjjotVbRESO3swkllX/GIE/x4/N7yVjtnNplcrLX9SarU
z5F0Md3/wP1qJPq+/K9KCTdi/SsoGx7yPrJSWbG7Mbp7UwWZzGtPXzRgCqkqKt7YExYPkBlsjQZ2
VoEHKfWCl+S6rLRQaEPCqpsmctIfBqg5JlnoKbhxF0wbEV3UtDCEaUUOFm3c0SmBQA47nkp8XqfU
F/AG5JtMoXqWIipRsPUx8AuCQFm3qOivZV88MwokgTm0uNSIELdAQPmc0eC7M7x2foNExMj9dXJg
8q2oj3FqhjEsQTVQuDiPBsbynf/djgzBQbxUi0jeWEReEU2sxDouSzdiZC2HCQq0ZwLtNQ8EMKS/
ap4mj25GrnMGJOJmxuyOTMocftiIPZKBwtl5QC8PnQ3CB+vjLBF3imTtR7D1vM8h3SX7T6EdV4YY
V8qsWg0iAOtDGQw1Xq6zCIkeh8PFu1F0oNTPTlaUQ7PInM7KUJ3C4IPAEa5XvBPvzBF+9iw1aX+l
0r5sxdBm1iBIlHPiP8HSgfnFWKaUHKphP4slSY45igEutCSt9ts2LKOLSfkzKJmDUdjjS5q9Wes6
b80CVf4JWbXEUdChbcK1WLv1ul4GIF7xzDxpemaG3olCpMw3jACQp/3X3TvjCieJDIo3rQ0uKHrF
cwvN/Aef6E9b8iXKBYDVYANgl19WplTO+pw0rlzPZsRPBw9pUgbgwAtEeaEoHCceD/Gp7S6m0c/0
8iGdUvM9b7mEgivkjFXYp5WGgX9upEwNSC1QYRBuoxwpruZ2O0TUZCBgWsjuLS0Jtu3iOeCY0/Nd
WCHGZFo7cWNYW4VhgWUGNGR4w1+gpqqpEQ+45jkfJoJeYv6gRw7y+l2zHhBCXwtez/OgLkPD7f1y
MAmxxHjHLUOkWL0gRA88nf0KOHzDZ5IHilB7HTwXKV6xPEJMSTvqTSHx1TTi3K4Q/1kM+ZumIEyv
jf0JyVQXb4oXPo/0r8QLPl0zdY03n3Znc8F6YLUsdQ5qbaL2X2DxfhzyVjDiP3ZV8yy4nI2lbs1y
SeOkj/S0JbYKN01Bl9YEmZz5A/MzzUHuwhmllgDdeeHnluO6PwHbc0PS3q+nrsFCTNo2pBMWXxlI
4v1FVR2x8gi6isTUEidQKWudAs6KCIurXjr2GW5hV/bmWOT27UdOfogpN1IgYpr8o57jXda051V8
F/YZBy9tCmkyES+BNTGkPNtdnGpHMeteU3DRYbuvd2Ys2vz6qjrtzVjWARdi3UCP0jblSumh9vo1
nTKJG0mg8kuds4ilYJxzN2KWg/DkT6xGgEvJhp0F4xKOocQlq0QcUtzf2MghcO00XVyD29qsrbug
vAq3TdF86rok2BwygfGSGiRmOQe9LpldOG8pHRh3ce+9FegIDCdjpstS49siPvopXQZIeImnb7+P
vdbEXYXuX+TkIiSqaaSmv7CTIkkS9mQvq8Ajp/5Zkxm+sPAR/8CXvsvmHoAISKV+HTAOk+VZcJc2
AYEP/Q9EBzoAto0HnTc+BQz89IwGcKHK6zfU8ZsL5hUprBTz0S2uUcDt5S6NX69Xm4sR5UDJQGG7
s6PxtZ3Ws0evvn9qeInmwr37234bbN4k+DNcSkJ9CqbwB3y30zTEBLPByzGhOd8uNpjjpnNtdMl3
mAyxk9f3fTE0UhxghSrojjZT/uVv223F28CbtqqOlhFjBfoR/Wp+mLDdYnCK4LcREU9nChWwb6g2
/qWNDNbQEpZOLCTMSh8dbPlWG7P/je2j16tu7juOeEg3fQJFQhmnsyo6D63cxfNBHjKi0dKc70Gi
adt2jnSO0wLfEO3aQlAD/2c+9mZehUPW2BZFa0MbS2CGrS/BCYKrzegAha0Oqsh9KpFEyJ60CoQi
xyTraImYvm1UlTD4hsPnv+pjh+vYpfh69F+SZY9RP4cwHCoVNa595d+l8w/1+abcLrMnq6thzMIQ
6RjYjZmE3rztGfprLtDWP9rX7w2Y25UZo+d8vyLyiioe9KZLx0IJL6C4dF014Btf6pbcwI/AYo05
VCPLhFw/Qr/wZUeeBO6su3LDlksz9xIsGakT3igwuqXmauNYaBt5AUfkB8c+WzQZQLc78FT3//Fp
+55f4luGq467n38WK1wBaGj6x7SCPoieNoiCYRb0jGiv0qGTOi0/tyFBcAFziJ88a7AikFZw4+BD
4G3VPNJnWDnWpNX3K5smYDDrFqa0HjHVdg57PsfnNFe1LwMNM+7tlpfLuCiv0Nnd8OsqyBk9wzzf
k0TKHWdVbcx9Pq0XHoqY6hrIF4uJFfbTd1QEFGCRyp8S86mK5Sqc/tqHyDmzZ7jCfbQQT27XQ10h
PWxdptzwmZ7Brx8rX6mgsn8WcFB9WhghZ643jn8r/zne5sdco8BCgIKwRj4Ktp9RT2MF3119gTwp
UHY8NPaDEwbXJ+NU9gv9Ss6NCoqxU2qEy8A9JymGLW1syGZ3QhMoiy8u7lNX8IkLFTtPC0KTH/OD
7VTgpnlLOCNzPUG/Gcn6QJpXZiCg6AVJ+wx8lgx3EhKrkXEAivTVp7E2ELhFZJr5EAjiBqIESdI0
IM+NnlYXgNGEcEeoEVeGp5dEKjFdAhK0xVZYNLnslfCSsOpdsh1iKlndYhh7k77nNXvh8/t8K9Fk
jxFiOyTiTzXtX4FKsK8US8LpX/Rl4RNKhOAfi2GNXOy+SJrxvOCp42fReyNDr/iVUmQtR53W+Rup
eV6lSCr1Zc1pceFWCGbzwOP+MWSSNw1q2alM9qNTvMzmIpytbUSmDJUa0rdhs45XyD8Rvz/jbsK9
E7PJ2ocHW0u8FnRo4Mlgekl8qOoQz0UAySpqvQHPXTWPmbGt1pjlKdnzoj68qFKCYCsLMPOOiCHS
EkvMry0DKZr87iicfn1gBzSNDOK3xN1uQNTa2FlUXl+H5KDt/nQoVSRy7OykG2UvP4sjXwsUvJob
O6Qwa7xlQnjgKNnBA4CivwjWf8H9dLGe6n7H1D9MtBYC3ejwt/jCHNrZW26E2KPWqkrZkr2hgkx5
t3EgXpqe4uXYoQsYnGpGcE5FJGtafcfaOJcRXKMWfyX3fpW3uIIJjrNYW2TKSOF1QAyjdkUfsu3/
NoplQS+3eeaQIj/YeOfZQPt8hw4VbnVze0+/IMKRkO7PScy/ktaNUUQz5i2M8Gae8qG/CENoJqnJ
uIPTNYWfZkAVjXm8iwxbZcAxkaJaX2hsM3glHnkqlUZcvolLku4x1Fm7P/smWJUWWiGAeo+gydBE
Q1iabbI26SYkU6aqSqPpRr1/cIK2sWT3GVPJ1TeqbX0Zsekd80aiYT1tp51oxDF9qXz/Lv1/C+lK
IAIOrZ4OcoD/bzCAub1G7TiaJrV5Hm8w/6k55dS8JVp2X0RqhdrUrKpoDJ7Rw2uy+RI+6gcGStk9
gGVBCorqnv6aPDx1oj/JbjDLe4oHqy7eR2IMDjSeH0HDoB/xjo6zaK5NROOxkb7qPZ6L/bGg+9gI
D94MPgCDakMFC2ZWgIyIrzYKzw9S7CSxMhI6OoK6Bj5fIDq4kX2hk4ZN+AvIv9kxKFjdGQyPtojp
YgDrJdpcgKm6fl4ISTHZbmZehGTqQdWgxh1BrnWx0cP0BKTIsPIqgK5wbHYMza4MYh5tddTdsMwZ
dtF4B7kzaVsrfN14jtEAhpf/9Utxew8PUJlVrlc6vU27l/uMyUOI8IDRO6Q7jO0VUNzto43QevzP
nRbM98QGd+5+1wkr0pQtjiW3HCcCQKfeWSfxJkg44cBZLbUb9lvxhlbrs46BKIRJAdlfw1a/NIeY
PxxrPyWvmvuFWwjY+5eEp8IptdCkX1W9SouVqq3M1PtYBF/X20Y3BbKJS8YMrRAlnfn+wRYg06FN
XZnlqabcTvomTgO2x9bKmmF8F28EJgsXTzsnpdnIolOjFNF0lalu7YR5AJdo1j6pLCD9tN51Q6l6
H4Pg10x/g8Atv1kywE7U2J0FU2+ODI2C+diZceq0Wda0cczGP8a3w1fV3iag6w6PEZN/YxlCrVU0
yHTBXXWN5sq4HUJRJLQg2XgPrXfKhFjW0vTNzxYTX1ZCw/WAuzgZ7iIgi5Pv0feSLZGAW3l7zsIm
jxUZ4ZQMJMClJwOvUANbUziws33Ir/g2vRPz7Cx9gbu+Tea3uu4EKoubwlmuCz6jDZZDerHf7COn
ALj91vvXWGaFfZZH1hwbVZDGB805BiSdIng3OxqRgjpwzjikjkRAuQkFHk/oaWPldOr1K+SXwV01
gMDFunfiMUid9rB+Rd9sx6r4PQi0XyJUqTAbns0Cm+VqxK/M7Fb1/R6+Q59dRB60HM6DG65QRidy
xaYKc36BpSjrKn7TEF06nhkfu+i+RSRjn03eKYXjW9U/NYaVrqzI7FOovj1enPv8y9xBtlaP7sNm
/DxeAtyydw5OV13fKwpPSls5oMfoRXHlUhyIRCM4YoZPKtPgwMQmg30C5lIUcijSGOFXN3IPqIsY
JApBJHrzWQl45qIIUDTXPuz7s4qM8RkLfsUi6wBHfhOJNJZvoA+P8z989BSI3GtVDDqm1XYyJma3
k5p/gY0DjX9UcemqI/LwJ9CSzLMfu5iHNkm6iANHMjoEX8rdWAiR7rpbPkrynaBjwN/SpYuqOBQk
J31uH17wLF7w1kIQR3Lppe95SrtENc1xio1dChdnYjUlwaLTSxIP92oEgXxyywG39m0wi8h31T4j
cmaf3Rtp2HpqkTPEGYBrkaWqlt9yZRksgHmOvuiyutEGKz3LXxUBi7gobw2Bni1HUq0TNWdS7I6j
CJumCKeQ7Ly+8/cx2RhbjoK4kxX+Ybf8LdcIxEjKDK8byY5ei1ksIuQgs2Dj8f7clGG0EDBiq4pq
BYaC4V7sBW1BwcKSwWoy5Km3aVQnz0yZJEEb2O2JlJVjZbj4loOgIgxBbZhvS4Gh8HXNCRD6Htph
jzbwcqx651nxVUo62ieLiI2fclySCQtR6AXtbURT4Av4RnzjlPTo+tFsDdHO3BrR1fPSInoo6vDF
eVE2osTVoq353Ec3gR4T/lUmpAzKbfCZB576edCcDvPQh+5Owkkga66Yr4wzKZDBFrMFMNd3egJ8
y4huVHHcJQzn3SFs6Yv+rIszDMpNmsLPLAMkICz39uUymlpdazPoH/BxDtAFDMC2hc/TTaP0L/6N
yuv/k+9ce1XLFq35Snkbq3yG/LosEuOyyQJm/qlV6jBzfXyHlF7d66Kpzy/0oZNICJq/x9bluyAZ
ckLvKNKKoa6qzi29GxLJYlHCaC6e/Ys5yw9BnN3hPse7ptu9kK5zedvErNbF0clhDibDx6ej172n
gzB6zAI6O4qROiFjj08owGnlRX4ATPM0jIHrIjiUzB1hcfdVhp58leFmSSxlQu5d2LaPlU4hOwxt
DeSiYLG/2mYlplNLN0muOMMdkNcQyVp9G12s5nP8x6WKvmbZVN0WaiFjWPHvFv/UlVfegwZyLlNT
CtmKVMONGqNmmIb/3ideCnHCqoDMES4pgZDC93le2WtLyfcAUx/qdZbcbnK8LmGQ27kuOEkn3y47
Tdj+DbbzeaxfKULFGYZF+mWB5WWFF1eQEM3ktJiTDeJw2UBsCFxeIhHDTjWNGZGe1YOkeywLoKni
sDzkzda8BBCbuM3mDMc0tqm/Bf2ttXV61mOkbdOtpLLRFvWA0W8mCiy1yBJ2/zxJ+Ejx7yThj3KD
pSBUwxJVh55d2fJMhEOo+fia3FkJQScQvc1SpDhGVKqVyFlag/8pPGzdXiLZs7Pdvs7kZy6vlErd
4Fsao63rbtPqUyQ2Ft2YkKeS+2hYWOc4Cq/u3Dh05scHooRU7pOt3/n9UmSfb1qa3i17I7gzebCl
zPzfXUMnH43uxAw9dE8YNXgfSOXebfxOZXVB+IhNQ3+m1ig8SBmQNJnaN03Ipdl0DClQBs4oTeqI
lt8xEF2Tv8qoDsqTbbo65HXRYw==
`protect end_protected
