`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10976)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9TaBM/i2ZgCPEH+TSdpehCfUxIR
eMubJuopP3JP1tAf5+7viyfGMYZ7LtwtVTMklksfAftE7xt+CbDpGa38bzxsPvMerwg9BtDObudS
sQnZUjvZwjP0zoPcd7m7AaIrlvAzElpdyFpWVlp5mYD84Jgy41aubt1hyOHbs7uNIXYuAnge8gxT
ufoV2xOI0qYIXBlJ58MpPDEBKZS6cdEci1K2Jl+GLP40Wm2xaXEJhxviN38lyVF5XhH2Kcru9jsx
3WBOfENY44+UU4Mg83IIoewMNA5KmHuJUQcGkMl0JYzKnaoa3BRhDZZdW4P1hOo2ZA0fUY85dG50
5Jvzuuyr6wEpGbdUuJ77lmVcLuRjB8GwndILh7yzVYe3uql5lKFL5VZ7dCJ81hCTo/XBOs3ThIvP
b7s1U/K3lhyaVQRmM/Xd9BRB9ACrTpmmGetIkX3OuuqpwO6bY4B4Lzh4z9hGXaREaKDvv1BkGr5R
IV7N3ia7E3aKiZ2wUvYGDX21TeQKr1pIYsp0QyvOh5/fv9x/fGnrI0qa2LkX5waajeVIbIY9oIgd
K4aESwjkA7KOGaImvazLzykpi3ch/XRozJ62U/GFLyLXu7F5mSabcDNQ5aeGB6TuTg3+K5wby8h2
/GN1QEFxsMeO7SY24OOdegU8cSD8og5aa2adt23VSNq1TSonckmLNvhvXygJcDI3TPCs0UX9WJHT
lwKgmjdxTwULLrvPbTTH5GpvjalfG1Dalgim64CCS3MgTTrUoaERM0VAje8xcJC4oMwSIr/C4Nnk
U4kjD1RiTx/gVptzUn3MNN5Ca9NX556ZCI5F83NWoc4z86Gvrs/g2Vw6rTOo2sL8OA/wCJzGJliQ
Ko60OEuVi07mMtlaKTVNjzD0snSQ3VTBJS9HZ4AKXiht0lCoOu3nbqxUpfBhBKEQ1J0JDe63nVHZ
wE5XjunGjAK6qj6raXLdlz0MAokwnn+zUcQgHETqJe0BMj92NvsFTbN403DDVI3HQmN1iSnm1Cra
awS+uUBSviqtrqE+KhtTLrh42S1+Dro/91jPO71lRwCLZx9Cs/qF7rnWK0DVw1muYy/Mq7y0cU6s
kb4YQLPaADbpnjBHMeBLr2eVTq8riqWjyLdRUkMhfaISBDO1SzyJDkLApAg8MSAxCAyCgXDOg5BA
VHaN5b29GFSpZ+8Hmzt9foJ8ZzLXSI4t9epg+5XaZLFfUPC8UZXLsoy4ARAQ3j5a0ddyE5OfAxM9
qnZxoKYHnjc5OO1mjsTmxFGlBt5tInlETHtlbJCtRa8852vjCejgnsa2wQGQsUdHJbn6XWAu4VlH
IS/wUgNWWUbWEplTPlbcUQzRZ4Zi/tZ0/lH2MpZqFV4SavqQouXYC3iXnVFD6h+0JNz1J3prhAbb
WTUf7exc8SAJV3PxhAtpuhOhL8/oebiGfC7fmGjOGoLGAWhLLWoNnQ11P9QvstTFDOwt2TWn0916
72yaMqEvf2sQJbncsXew8/GfsePv5zx63RCDrBEIcYvCzkulbS78XsIJ1+kqdq672OZ3QgZaH1cS
HJDhrgZYuVnDjzuc1plll0BZu1ZMyHCFazLhe6zUnU62hKcbbzjJU3Iil+FaBm60DbeX0Hzjfo5/
lKiAXPG26fkKFwHz8aTw0xL00ROSe/1BqA3AdgxEPDzc4kDEKi8jyE2N8MN2kwvXQ5Qx9buyAz7l
OBUUutg1swA7aFaO2Ko1Hoh7vxdYTwDg1zpo2d5HwUaUqK6eOz2VivvWQRW1i2FcAqkGa1z2yYen
1F0ywa1eQMpqPKCXuhmrp87d2d1PDAgYVMjyFfruQTo9bI7yTXhE8e2Ac/mWZeqlx0AZRT6YTn7m
1/ZqOt9sYicuDgc78EjjI5BjYzs2BoDU13HPOWI69mqjyz+f7b2q+ZvD08PlduTGsdYB5ltuQZCB
+H5CcspixuK4H8uvs3aRNJQJeQLYbQ9tsRmV9e/bdtsaaRzf7Pli3RB5q7ZSA7JQszJ8hycnoasg
QHIZjSI975la0BhuQHT1ExOgTYsZ7ouKBwp2WZ+CvYdsEDto0w8TxVgAhGyzkR0pJBcK0+syAcLp
9S+QfN15fq9ZPIzh6o7DctNtr8x41ra+mas29xb3qiQoyowd+uHq42hZ2MXk56fHk2zaX5TMghY5
EqlgML4zBY/K5M/sDaXmW1fgG9girJQdbDPmRQ8lsotelCp4fzJf/NuK8sh/BvHV1XUwHALk8Qku
50PpquYxvO6slsyp2uapGfdq1WRh5YROG/wTgF//n+0KeIYVDlg9iJ07JMINzVVZgiy4tfStRcXt
Zs9Lyp2KYkjo0f01E6+jXn337xhl4gB8LSQ0mrcHQd9Fj5XhH9AAd7R9XSYE0Ovuw6SvjcfOUlNM
AQo+aJh5liezz5Oz2yt54FFm9Csi2zCAyHN1fucB14o8pC2zMLHFrvUJ2jPjtqxQ3RpnrgVcMvAb
R4oYEv0fD03ydtYhBQAWR7qAC2+/eRVvBE0NF1btJBopq3yfQhHIgkFf1Y2ANMew8Gi4KbN5PYcp
GvZB6GH/zUpH0oS5hmRgWZaVh8xBIKV7RabxLOdNDjk88Wk3jN+XcckTnwG+Qg6wPg0axfynOjfW
3TDYENb+NbvtWTtI1t5wXohGjv5M3ApOzeR86V1K8Erm8G11z1Fzeevtt2Xiv2HKgKpPv2wLq/eS
oV/gj5HMnLZyzXMGiSL+GK9UUw/DGcEFBnoFvFJjgUnVW7PSUy1aCK4TcRr51Wt3nYleyPfmwJO8
mIVKzV/DivWLnXBtz+eFnYhGohUEo9YjRDzCrktpIL9bULfKLNUeHWXqshMNMgvcEMsRqmb8LLyq
L64SrScjLQMGjJ+Q/MO/79g1NWdsgqmaD5KVkEfSIDWZ3t3ytwh4oMz91ocWgTx+g0K8fMv28geq
pXAVowlWToJrFa8cZBO6WK4Jh1VkTBbyzXMwGlGwvvL5OfuyBEv+U7t2Hn7UzMJlsZ92vYkVDjvy
UqdprpXcHm1QP2SEClx5b4C5v61IYp8pIyrCiQRGhl/BofWo7b4YdhrJzi6DfTJJq134F5PeGz15
5mYO4UyfSBoeEk3HVAG+6iq/0eF8lryLfJKm+v8Jf3vZ1bOzmAnutWUM7WTWIVMg97qJL72nqAJL
4edFB0Noi6F6mxiyaU2KMjcYCh7VGIjYLiaB4rm3d13KNDRrHWj6li7Inew2PhCWHoYYoJ+eTg1T
/oFBb5pKJptKom94I5E2r1cB3iL+2iMYVHz236Y4ugW83qRnZbMZE8qD463//YJFFhWktcxGx2AL
m8Wg/guQEtmR3vLvhs/3zL2/z/uwguTT0AiNv4KBUt1mKjVzDVBXcyr+ZaboJfE17be4jXv3ruKF
g9qZu/uQfIZhGX0SxB/00EprenPZycRrQrQDFVj5wCOakHOKr4x8554p6zJ3UfM/arImrYLBHdlU
72RMWwBNyJzzi99FATp9Mzx7e7d49Y2EBgd4/KckBtCyobYm/gj6RUy11As8k1K4gtSPhcFFuSz0
f0n3B3H5Oi67c/rrLJGnCbU3a7NUXqAKEuz2O1IBkGC5oFWZ3QWHfExeyiEPxS24v3Z8Z8zCvzFN
Cd47YBoWZzDYYmN8Wgu+PvT7vnD0DeWyx110HMwAm97Z66cV+ktagFQn7ih35S+Xaue3605s6qVB
q9kALDjD3V/rtUM/C9IRzeS7Yjisa6wVPOnlHrsLr8iug3YCi/fTHBdZE70elk877opBaJ7kpRFg
wLStggaOkcn1vI1KOTCNLjPiMUftAdomLgBM84lOwTMJo93N7XOcJVbe3OK47oXVQ533R8vjf7Yl
ZysA2O3UCRFXc9Mp6v463sXYeyyVA5a5Ww/zc4nv7eOg8opVxx89z0JqLkbcIrbGMUxxVOBDM/Gg
/+Um78beVHDuA4z5uK7CyWdf0Lt8SPsDD6WtOp3Q3+qYfV6Tw0A9Fi7u2cxxBiOfPju1KG6sjqKs
4Wj6wy8NPBhDFcW0ACGb4jC3h8J9NQ1UzXMsWLx8CpbNn3CWcU/WIGWyim2iJolYfSB9ZLmE+ZaV
nPsGr8qYLOiTomVhWQ48YkKCGkmUnAAZtEMenk3USCkXbX0cr2mjde2T1D/2mTtMnYgtJVFRrq0O
jbGaAaemc/ZG1ZL4NONPog1io2gLpoxzVMP270d6wLeqVX4UgI4wSbzkJEdIewk5gYeQ2B/ETe+K
KDkpJDTn/+lqzkYVZagmYaq/QYMbHi+qQh0iCE4fF0q4llrRe7+qNSOBQ1CCiTVtIAljB2tzNnBF
z0xhZgUSC11XKutT9Fez2Ovhbdloh1AN91aWM6FoTRPgOE4s4BKcKNmy/mdJFTHdNhQuHHXsyTiH
CcO8ZW+I3WxCNBsskFBUrSrUc5/iS9hBHr3FljiKNOAq87xl2SbnI/jcBSzGSX1fUj3Vo7rrLmPP
uR8cCeMjNPwyHLWdOKRESBA9/GwdAxoKOieXNiwNHidroDM1TPXs+9dMN5qUBJAD0rX2Ptf3q3Z8
jTuETkj5VqMX+9n8mIveJ5voTcxPI5+rN8Tbh180K8w3Fk4CX905RnbSMgLnWHd9ZE4UkrUmtise
qzA1QUVn9lmixFGL82FMjeGmgrJMDsIie9dz7WZvC46XI/uXtktvhLAeGqF3Fm1A0E3zXHRkM52k
Ouma/jH3Ynrf3SYcF2ECesJg+hU7jUxsu8e8DxE7kQ07Nn/mJ4Gq5X4+2TI08w9nMEsC3zzp/+Hz
4j/JhwVX7mEttcM+pSzGF4A0fCC7KATcHqB/QXhkBUAm1YdSzvg/qA2veIRP6/FdgjnHercrCCCD
Lk9uSjlytn0YOeb/rS63sBLY+1lhGiHuIgnzBmUPtXO1iohnAn9WrGDuK96t3mPFeedHKnm0j7iy
K/YsAkTY+YB34QPg+cAZe+xPtUKiMHlo/T8Nj65XU6WUcdaf5+J1RROudQ1TtJtoJ4bczaJadPAU
U2iDDJT5lja5m/ukTUAmGJS/w9cZXNuMV8WP7kpcteoTJFO/Mrj2ZsLV9WWsMr/zNujQfzfAlh67
mFsMY/a51tGEERjRSRZjY2EX6AH6ZPAPqvLhHPD8w4fcGOx2NR3p3EbfJFL9115yE5x+imH7//q4
BMRaC9k81PSLEaM4Jc2o2c6o82vePwys8qvlvHCVWF1n33GKWNy20U7HioT0zyluRKFSfk7FZcLH
dYExiD2X2U3TeFni+wzyYbO7OgkvnPJb2g0PanX82jUJMVBNmTFnkmr9uS2qK/K07hT8BxhNXAdg
/dN0DYqRQUfbO80ZGzniPmw17Sw+G0P3sqxaV5vvBWG1A6jzE6Gh5CTKFkN0GxEOAYuZ1sxcja7l
d9zYv07MtvEoxqh3uawH00GFHoOiDU7ZtzoZ2xXMz5uSP97FE3EQ1m+i3AnHSbuDYb11p55ZbhC0
9fb7ltB/PQgfMR1WKFPbPHVXlwY3i70gXRHdDPyF9JqDyKhNVSIK86r7PoATwotUwp4Ijl1VdC0G
z2lRbsslPet1NS0m3dCquwoVMzV40XPLXCgQMkXk6Mkl9nYr9FcPa5j3E+AWP3D9Os+BWWOFRlC4
7wqvOIeNvma9UkCZzljtFu/vZVeFWBWBi6EMhB1AgSD+Cf1/Mw8WHyH3QgZ2aoUrgxyE0x6zMYnM
/LY4GfDQ8aRiGbUOPZu0yrrMyZOghF7Qo5WzDBpAVOGAxPDiAk9LHtWvEcNjajWvC0c0tsKyDZS0
bRtLhrlgombdS/SFRM/zFkrPHMLQUqsJpXuJWRkGeDzQ1dqM1/HCZW9YifMlm1c40/ozehvERnKT
DLcXFc6CEUsPh8C38nrVEzm25wC2bVCpsNLlivvLldJcrz+3AfvfBleqpXng4AWVh+tw52N7ZUW0
WPuv/qUE/iOxIheNQ3xApB0IW+bSgy6qeiL9BN1ghSHI5SnndLzDYrr0K5I+o9W6UoLw9j3znxyn
fcaHpXSY5YDUV20TF+S41Vc8snMoYALxyGj1MZ+qMTekX6vfK99rbhhnJMDUBXI3vV5kRCKghKZC
/2ug5QRCVDms9/yVhc5CFEpuY8FlCYA/BNpZFCcxJTaPUFYj8aU7oaC7Paa3jzDWaYFzz6Hl9pPh
a+j7jkxxWMkpk4lsR5rms6PVgCAKgiE2Qqfmljl8zre96wCSzxT3gjg0wh3GQMZLkgRYZuaxEgB/
9gQUOMhBu52RqoU2oUXoqxhTgaI+ltd2thxXYUdRMSzWobHyADJXNaxN1/A1EGJeze0JnLAIGpKO
/8IZxBhyiHap7q8ii2KUPWNp/Lrce9spFG5ARRNYpTYtW0BzxU7YSz0Esh5vbLxBNy7heJpe3y8P
5mmkvmG6RhsVmKtlqX2yZi+PGn9LxoRBbdVBMzw5UfjczapcJXCtwexnTe72gYjpytt7QGnaD9Wn
OVt4uEamugtexbiiTIdQfB+Y6aXMVf7PFuOOHEvBHS4OtM4dk7/Huw8B/7VL8yUFFewA3MD6nKEr
QU9yZoQ7Jj3CECFnt3pPGEk/kjlRhm2LSTrd80keiE9pHE1WGew7ITSdDVuOxaNFBTHv4vkBw4f/
rtxW244K5NOXlpIho9WJ1o3Kp2SxDh8cufaB0tgrlcF3btzCUjZ69bUYS+9Kzs8qNpV7rlsAtPXP
uNE30cRcd0Kz+5cVIzpKC83l6BQjwtcQf6loDAo4TfpQo/S3JDx8146UKB2qoOvz8pYizmiCARQm
HjiMeIrbHOEDiRP7/6SeMLHPC5j1u/kxT27zp34XuiHLxc4xr/q14kvmTzjgPIiDlXWKNP63pO2y
6I0upjdxgRz8Umt5r+ZzI4cMzlHaDkY8+VnY5Qd7PxQdoX2Kw52lW+Sfno6OxH9qoesCAfp4G6sJ
23Nc0tmmTLTPeC1EnqOA+xK2Gy9ZtDchygffKYVtXBW07j94TP+ZqnKRuiXaTOqJQLkxi/yCOiv6
8huwAkaIQst+X6+o5RPnmPh8ARUK0S3PyB9YI9mRhAcxnfGB2AI2kMLPBYWfsAtBRQ33ed3FFiXy
xXFfkxrhCwPS3n4QUTj32RmCD4/fSNjNxNp+DOxrId4R3ZBSqekl2OenGtYqAgk+jrEKLLNEaZUv
uJE0m/5zjcjxSKvPdDM9wA340csCeKExT3MHKf198sQX58ebM6YFbnJ2PnASx7rKhk0dFnk/rNNv
OlYhE4ENQkK5GxLjxYCLNN/JmhUiFTT/RvWyFryJM5rTjNJ1wzsj1TWjB23O6+K0wqqHHDVFLE3a
oP/cR1fjJq2XrhEnD/lsd485+pp7SnPvsi6Bg9cMv3mbNBEShrF4fBRoiNp+lB0HS4P+aV8nD7fz
tn5mbNLZE5hEADZwN1BU7+apA70dJ5xacpHm1unlYQABSaYmVw2IpB5h4lsYf+J98LaY2ZnnhDSV
C41yiul6rbhS0aDtwkaGddJUHsIvcPXp1M57TRE+c9vFTL4Vp9nrZ//SMrf/wh8HUlSkg9qiRI1V
tUQkVubArU6Vb3GQHSUhLB+JDFYm1EuqgQER4aiuZmdf+3wS5DjEZQ6/7X1UQBd4cXhNOrwUTDSl
1iiLGX4rl8d++udsi4OjyeO/cpoKWioSNdreDSuRkY4rt3e8lfxIZXWmCkYx1GG7IO39mZsNAnKW
3UebFNFMObS+EZAaRK/u8M1rcimvN35ffDfoXLhx04rBluMkdqa6LQ9OKwa96KI3O4dZan9Dw6gM
JgFCGafLBeSekLDCEP9ESIXbuisVw51Sp0ivF8Ly1m9S0nFjPd3+ZvTBVFF+IwlcPHbaJgGJhoDo
NmITpnED2D8C/EJP4D/68aPZJPtChtGmHlGdubtBQVyd1q6VCKPtKDdT13Y/brL+iML9pU8Bt30X
Rp/4P4+HQvS/X+p8ygZ2mxW5iElAQ+cRg8TNEt9VJVNQdbOVcs7MLPaajG1tqNlYh5YHTpw6kl5N
8klA9uUzOL3PsG+t8cLvF3ES7w1j5lgIu99YM7fPI9q8ksALsVtMGdJfMf7lVsU7a27f7xci7IRt
Nf8WqiWSfZPAkXEbCIMpsvLRwWsMDzFMjLNHr5JmfBFI0KvJmroCTrlXEs3Bylt6e7PGgPFJj9cp
11u9Xa1uP5riIm+DTFtC/nb3+YYCwmeSS9gLr1KCzrULRFw5ZeOrrk+k4q0qXpYTe/y3/gxMzeO0
/NS0l1swJpibcW+b+c4dFxUnk5DM0UngcKnUVivYNwY/zV1VuP/l39b/9v+s1Gk0QwSEswnJTvTi
h0P5UOYEZierbqVWR/FJvppIwzLAqujLpElexPC4rZcYLjn8GHahjBYhpW0T5cpRr12N8wWXuP+E
4HOU4y9ZIaualk81tPdcOBAj0Z4x2u2A/fBT1vbrbEfudAEq0LIhgnOHPWfgDBVv9ppndceeJK80
hoAm1eN2+TEmaErQ0VTxcta6/z5iWwBB1tFC8E1S+Z9p1TbrQCHKx0ZzP+V4oHC0gTqjGTvxmpqR
QlAw1/00kEoz5DY9vLQcOjEg2dTdtmvermIqP18kOD5qxDljmaKhvA8F3/XyMicvwV22xHzub7uv
PMKWKPrWbz5EhZ447AaWoLXeLLWn3k7CRqtLniVgf6cee1PSk7hTU3FZFwSmZbcTvNwbVx5hCdKd
SUagxOgGZAp60dzaLseYJKLDqiaG1F0/RI39m/grinOYvbc/3EDTvWNAz5Gi3Sz1UelrNObrx8TP
SVV18f3BREpXJIGU2t3uuOsEJb83BzoF5PAag4hI96tC5nGwQC79uSf9mp+qCskpT8ifDJWTEkhf
IkbwCgZ3GthI9stXzdiWykHsbgYI25aWceQBp4p8AUmq+Dr7epQJVUK3QVc0VhjiDPvLlj99s1h2
lbdZuRU01T4LlYku3Y1u8JScsL/wXvIGkQxNW2ZyjYpBT1a88kedDPUG8iwTPpCOrkwXvJ+9PeC9
A0WbjZZYOpfzyX8N/5cbpsrGi/WsZFmewYuVYRCWc/WfefXAfYNaVETDAP0FgOixzFkc4GLt9fLe
o+z35ciD0OM55PE2OUaUeUsZbAmC2YwLvJRm9rl3Y4m0h/EP1ir/kfc4ssECPZHSBEE+ldI20btm
AhENjdwCSEeFc8dWqm5CnaC0kXjIDIZwBG92j2/fBpx82Zt7C7heU5QVNBZxrfKwa6NbOvecHMqB
V48wsLA5muzDjXDJaoBGn/agiU+7ArSvwKwV2njWtl5rdBhx6o00UoMC4ktRnVY3JT77pT6LXq1f
3FABCkHFQys05lluTNEfIHliw3PwrMkhDGl7zL0uQ3OtHXKTHCtSyWzZZuuvuMBhpWy1vcJpy1yu
SY+cNX/aQnelwL8JRcHKjCl+XYWLPRmsNBOuMp3KlCP67w5NDASeV31c7cELJ3FYC81B2WtBU/o8
4SkhaQVJ76zYY/1Q0qbWOixcE2NbMLTYaWLSPjTU6BUPOwnkq6H7zyEK32o0iTRcTFoGcH9cwcMm
6pJb9xeXg1Hu7UdvEt7Z7X3y8CVuvQZosxeSOMih1Q0y46AyELRGx1D67jUCon9F8u/XsJx/k+TX
EHzPPNwV0vOxAwj2E8o98mX/AjO7MFokxXE4ntrUwuAq3/EvoBYosB29ye5NUVUsw+d5XyjzC+uL
kIbqZrRmoNmSmsuMrHSYLedv+n/OAIVvkeHB4ZLjKm2PBgICxV4+sGrRKFRz0lU4+AB2YCsjn0a8
Cyf4kaWmiTuML1vnTd/Aj57CvP9G4bP8XY6v8b6U2+JvXNG4ODEIxvRgS4FrG6kEiJlOYTzp2jVu
jSvt0t57bQT/J5prsfDlUA1h5mRkGW72lAqBM5G/5OWKUv7N9BS+9p7O8GGkE6DwVvTSFE5O/Nvl
+ohQX/x3FpTDRMYlcNRmHh/uOafTJYZeA1/29RBF+lauhUV46Oo3cwa6IEEFAqcvy794s83kBfi8
S9DP6Z9xAIlLlp7Cq3xRI7Uf5bWh4RJt2xX3Wcrkw24PBlXfM9QFlDWh0TEpz8D7qGta9Lao3c1z
yFLzqabT3cNDHRzAPqIcbIafEVADOX9sM8Qt5BLCVxfc8XS2joO4SjEgMTVPKLcRx+FIU9louJYW
+GrZhViFrrujtP4Mdb0bjp+a57/WmbzQ2Q3LGBpVV6G2Do/E14TLxqt5yWXxdgCdIRvkn2nuWEui
CTaRhPRNdZW3mDzF3X21lg1cl/e4vLqU3I8COW4ucRg6oZaABf4YbJ9FQptyqQBkuRnxjGDk+7C6
E4tPIUaWOakcCsdGk7++KY1wGKkqM4w/ZG4ou9prpdeLrzsc0gSL7H8+d3FgM28CY4Kegf8gZQty
kko+kx7in9aGP3vMF121GleUEjjuy40XxQ8NZYA+xXhA+fJ1hDh/s6y/7iuiSnvtoV1VU6X/O7hK
ywub4TogwmuKyXoInZEAtg9AFQK9WWVA9nMDiJ1vbIKumQsY0EL2DpNBnYXKCWkMzaObAgT4wfsn
2hXQDqv8gQg8beqfZAjNGtNLcxVRqpjA9lZE/FrdCiGPJW4E1wfOzCcNo/9GWsGC+cIxjscISuhP
819fvWftwDQT2nUyvoJhJ1btgaUppr6ZtvNg/4x8tOrnVqkO706Z/uZ1HKc/nYz8kj4+PMYP8bXg
xeDY77x9xOtmwH39mK7ushlLiLbsXNG9D5bzDiLmLVM4hXJ6pQMxf9Oi79Lim3ndXpUqRIe39wRW
AD1u4d5LX8phUry5UBAUplIgIFJXk0ID+71ZTIjIkHv/nfKpT5PimKQqFiEtkGsOMQD2dBlSbAdl
2txnFpVK5d4nYqFY/nDvb6avDXsLHEh37HSJP3KU8DujG+fiTYaoDkerAtv/CvE+mnzLZWTR9ibD
6mvMRFTcNIzhrOO5kr1P+njwVXRjY0FSGqmNBvrjbE74gEfMM+0A0cxgshuGWteZ9vVFAUknpg2F
NMC9dxXypCXf3gHMzYfJflVoFNjwTuoYMoRxGANFPCV72d4Ez06gAy0PJGz/aDhYA9KQv+9gWnkX
mJrye9kfN/F8VctBcY6nxSeeMPKuylCD3d7+uB5+W8Ur4CMKhbyGJoFTbVBAQns19pJS2jg/9ZM4
2xNA4RSfU6tXX0407LxXevxx/Bg1CM5EanOo7ULRe76foimNSAFtf90ZS2TrOctLb9vOkuK8jkf5
R1MC2X4gY4tzqxYIfs1K4gPytmuA0l3AQs2Lnhm2mHbb9SC6O3xn1Zc2edm4qSnz/W0M/oxeHqVQ
UkMKE0SQ9BAW9kSLbWCuA36+UEraJ+25qDlN6GmO0888OGn8qG7f9nN+mnNkBvYefcse1qcwx1sa
svqVeOBYIAnAzfYknkMVMP4v+6gKLXVTyqEIhwMeaUBX0yobLDxyjKG4hFmROZcH/ZgHqFvH41dT
2DXpTlGSUlXBUpm3DcP4aeBtJNCI842xwzeTGBcVpcs=
`protect end_protected
