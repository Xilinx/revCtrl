`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24864)
`protect data_block
td5QFuuLITbKOtkE3oI0mKF0qX1YlG0qJOuKpYVLALLrLeda9QgwJltUXCInERXFD/JgQu18K8aR
RHHxyOJDAke19pKVSlnenItG+oZBs87zizaOCc28M8Beqo5TMOSipKyJw43F6cT7hbB4mdd+sdI8
7EPtWsbfpBeGlXkY5HKvX9nXI0YbaWkgZazFWr0jMxnJ+uFxTS9aqhmEhbBPGqB5glGqvXLJaMtj
2nRP6Bz1ULHWxcQaoQcCwZqtcKZCzU4TNEki0qxIKssv+KuVsaRQ7V8qHTeJNXm1/GRgoo9v0gzg
0ppkjRMSSms0SwY+BcUKrLrmHZIr8vvrxam0T26TF/bg407C65S1acb8/EGQ+xNfUFGpKqiN8Bi2
HiqwKQPeGxikRuhNFazdZtq9zwbKo86g37/SfQIWCdvYqjkaGoU265plt6M0ZBxd9O4YMLXI7VPW
Mc3sZvHWLq4uY0RYWpRElW4mxN6K278TwhvXQ36haphX/EQuVK7j+ynCbvMjxhZA2tZ/qAK4dNEK
Qfg1XPZ3yi7HJleFNjMEVHLr1sujWoak1NCk4A7Mzmje6/6I3+AsIo59KjYQ2iKlEOVswzr7QxnC
JUza8CyxWv76ksoEDMo4bdddxFRHArj10M709ABQGFn9N939HLBVPz2WnKpko2eEcjmJskY3f9yh
xm3RsyWGWphFLgf9A4JLBCisAco0e0H0tMK9gI7M96pSJ40PsJ2F+aSlGG7vu11HumWRhdvjtRlT
VSr4SBWYZ+1BksnAOtkPUcvmgzZtrNQqbpzPyqhohzChRzEbgKTyv00nts1lVGs0bZH5IiJ6TbLr
Jnm5NSJCE+HZq6Enfb5VFfBtfWC8PsNu5meytqJUCXqPa6OknJS+ljfktYoBND+O0JvOyTdTe8E1
tlsBC3wUgtJWit73sFiWYS7mEjvtREi4aGRPCZanYW64ea9p/oBBngcnu46hhZQSNU7ivJI/m0FF
9y8Sw4q7kJf85/ErdIqwgVKec9cRjba7rZ00+iGBlA6B0l8XRI/6bI/2eovmCHyueWCSJpXQgv4f
Uoz/WkVWhI53mEFa+waW4hqRk1oqozKLAQWcEFt6yXpNBx7ltniyEdVBjGRHlxYTO9oiZjb+O1fl
tnU3qmwRhg/V26mDYbmJNXbUHP1uoWOk0marWaBTG6oJcD0eR8oZVmxZJFiub6vYZnN9964luf/L
Pnw+J+TJv/uSjLNV60GcOABdwstynDkIpBGvTOtG+Q42uJNvPxN2nnAU23XJpvDHDIdFbYMzpdiZ
YNrNI+glAhGBw0yBoAzACqU4ToAXZ4CQPZY5a1AbEhQC5Pb+N6llmbcdciyhxAreeEAI4rJQYIID
qOtr0cD9O1Z+Ki8zbLYr3HETYqjN3d7yXqPl4CGrvDKJV7ja9B/5RNj+p54np6XAUUKJhG6/qhiG
wpy+3DEt1t4WbYshiNcfv4IUY4Gbh/LwXtk/LItbKmEq3/YcOIRX2QRCzkoP7eCt3ks5JWO7vuxH
8hTNzawhBZe5pcZXDPSbM/fNFuj6jVjM69LaqKcQwnrQ+H2OA8pJ4sKah7kJEDHfUj6pOvXWXiHV
kFJfwqLwXamNzHRVqHj1H4Gt/xNVStwyGKEPuGUtNlRAScwN/lOA52hULqQkPZA+HBaVLTWeuPgM
DyAnmu7WrNv9HErEgeRFXw26Z3j4gyngRnmlNCVa74CR81upga1t95sxvrx4FMsYE1Y6z02L6UWO
bjez8B7Uy5jBTMDshbPO/NdmFfZO9GBtNzG+NdOxDmC8PvUj2Td9DXR9f0V6eSZPgOcQxnaDkGax
teK6+iYf6cY09T3GW+HJ+Ah4GVMz3S6ntZvLjkd6Eyjec30qXnou4V1K76TtKfmX/o62QWCwQV9X
77WD4r4RG0wP63K8tyuLf41ZcYd+XcgfYmG9XqvgiS0IvMLQrMY6oreL1paNXOT5vJJAL3WmEpOW
+Crp3DcDSqajouZJCAGuSYNnrgr7anvmggeMsbWLFFi8wsgURe4FDqYYX1BI0zEFh1dhY7mDrx9s
lnZHcoafZD4f13bBBGWECpyz4rtl96xoxneS1FMiOdEDOASr2jnA6tA4czQIq2SdHh2F3zmocMhD
LH0S4vH1fn69JxO7c62OUWtpHpGO583WDPe5AemNB16aOvcMoPV8fH2IfCZdQFIdeeEO0/wwm0ZX
DjRxCjFSN3qAe3L0chSEjfUNfPPlokUHLUy6DdR8mI0luCuFgYOmU0KjUi/+MOV6wPQmO7HDaH+4
mD1S/QZiwOJCNjLO7irXb3xvCcebUwTTkcW2HIIiNHDymDeaf0A+WuUTPWQZJskT1ImA78jy3BTq
uV8gmxBumQlX0FgIcYLp6NojFImce6NYavEht8DUiLkuL7xNr6xJfhkDTiEp1mNyxvOwSOP+GcMs
2AFCWaPpYMqHiMFGpnfvsKDvsoV+hkY2GS4d2NKSigNFewlaQYcHKT7SPCc/+l+4nmtnK+EJBncP
n0unqxZDKyZQX5ZjZ8DtRT/yXexndLOwc3FU6aD2CHbtF0g9tk0OvcnefE9WPWlcO9OyyoiuNlil
TImu59LpZX0MON/gSgZR7Qr+w/Z+rBitg5skH2+5ABlexfexu1nc4WMIOFJAdr4l5DMhYrLxscVH
2umJGNhxu9+JTPMpO1mC4iksCWIZk8O8LkDJH9KSeOyBn5CX3VP6VzQHKtPZqtYxtqh4zbZB2mpD
n1qFnf+x15PD+UhzTXOyTsxGNEjgaNwGTDE0WlAVzIxIyyhBWsMxWF0Tu4NVTA4K5wHh3et1CkWp
LNfooU0GHUmk+41+E24nbRSRwr3SRmzKuw2ndyn5DwuTxI13+33fBjwV92QO+aaZYoVPbL9ueRZV
cgxxJCKWOR0dXVHHEveSFNbpN39uea7Zn1qiKa9ZqPjAdf8C/iG4mBFt/8OeyfeKB2DCwxhHezRZ
v9cW0oRKyTnittftPtQSvCErww6EcVrNSQABONhyIdlOhqz4+/w1Y8ivtYStp2iOXHMVZbgpEFQS
m0RPEbGehpSsQKFKoiAUyV1K6fiBNTCPagkaCErRAa/fMAabvISdFgS0pAJHbJaIiMSOZdTwCxf/
kjSsjYbVxhzDjtVqtIRQCbqewpxuhaUEE7+dnsk6OegZUel7sMQSpVyADUPMDyDULhkVzdWq0BwP
kxLbpwA7jUvShqEfJydvDUgmDwNsTYVGP61/gNqwMuwh6iGB//HTDClWLBWyPO7poAJsIlheYWOg
HzpC6a9qKWbJMbeI62FuOyQZwopDk+8lSq+PIQDxmhA18yXiM456dVlbaAoXKdLTOE04NpFWvqq4
O41TenqKeyDjswi21Td+/Va5J2UXdOmkLcIgrhBtO2PMPWh2ZQqvIzKO4fCVqABkdLXDyjXQ54y2
hghsgJQcch8hu8hfSHLVaJo+i/enm95r4tFTiHTUNSeQbSCb0dcGbTf8grokpc2YQ/vbl6yKYZR2
Nxgqbw3lzwX1r+Go2LS60sUippRvhR+hMPW/M62naIg0pRBdC5fPiHY+uPU3DKobPxKjBeIh1PY2
FNfd3IsiDm2zTx56JnqshdnRa0EwhAl1P/v+gbKPC24I9uszcKbkCjpnyggFxnPmvZ18y2mN7ttL
Nwk2eWsxXB5HfWiuqYY4LIM8lDJw3fsjIDPgZ70pDavQK71uUFD2HtslRudXF5EP8cqGbO9BTkBJ
FnPlJnvN/zgbqR/0BfM0AU2Lnd3OC7/CADQ+kfKTvXz3EIx1DlTGsAN19UiHO60qt4QtiWdczWE0
PZFiXVJYnMVmIDbj32dvRJBCguRZPXOm0nlhsGpwH1CDAZ1cH/gUFdGdvFcpWzxjLfaYcDXpo7iW
R06aDpjnPfq4+zClnhw8qRSspYmCYIq1AUjExH4MlKNr3VLykUO14vqx5jQie+HgaFPl7VQ9eJxT
S/m0S0tjUNutsGI8I4cv0xx1lf5bb70s5ipGL/qG4feV3l4N0G57VV+tG3Co14s63cQ9QGlWEH2F
dKR5/NhS1GcmR2Mf4BFZrH3e5ZvEvMF4vzKQBDkMra8UjBhmFNjA/PTI17tuBkv5KyD640ZPJnQu
WWbacukC/Zw05OTcSapWLx+u9CLvOz1jpy4qnPFCIeBoK3n/gG2bmmc8dz0Bh4As55WZB1+pviTn
/+JnaHnoyKLftI3E7S23B5PXirQ/oLoY0ZGdbETEHATTSk0bSMx/qc+jUBbicSFeWR2p7jQBfKle
h99dHLb4iBGnHeaMijaERgVADBQ1gKCrveoTTFTBunbaKOUl1HHUsJMY/HrFGjfrDX/e06ttKNNV
cfTi07juOuynRpSYkCJU0kBkBTRJP3e1zVG0s32cG3Rn9O9KQIYNsywBLfabTiinYr93xkKBPUNb
wyTf2TEXUu2h2h2ttSwojlPSzc4pv6Fa9pk8HTs1z2wiphSFkjjUkul/cjR3hEIPsBsUhY3rrgyp
C6I8lTeU++g9wh/w4CEpY7RZjMrq1yHPLqEQXtu4cLzIMskH6F0Jo9ZuiRHY5XoCedHML/a5zC/K
mcvXZXHdf1wK+I3pyi0BaxJuHfminaRZxQXDL85R41yOAHfR7Ok2Oe4qa5wliXPQCWZOugmft6Ln
zTVZMGKswmToAFgUQ6DsGwAi5Z8tJPB/Ui7h5bS8Z6qGn+11dxyAUmasVx0u2X8Au/3qnjF2tJMu
1IolQZNrLo+dMneVHDm1PHceD9z+rNIf23T4DMeuHHZ7EtyU/w7I5pSADBskLQHt/uqWSyWOQfHk
C7ree4gLZ0DcKbwQ2uxCtMzfNeIVR7C1nY0y5fuwQddkcY6ihZBAGwSDQYZJ6heeNSymrOUbJUKq
jBMXLRGiBmHh+RiDUkxW5YKNj7lYP23XE0hHbHUIvj+o1drPirX0Ps6xh0SYaQaU3rFUoPCYWD9E
snQSwo0QacS+fhqV8JVyV32Nyl2+bqe++aDDRKsHZrg+QUuBau7Tmm/GZcmY/YNJAF1Lf6HEqike
baQmn84be59mahJEBEuu6RsX7iqTP0ypE8LuN8maAEwbQ7K7i50XAV5//iWz4ab/TOVp9/tI0BbE
YiK+VarnNpGQ9Cv+65JZ9udnFOCzKpb7i4zlZiYaXEbNt9ROHvwX/SpdhbYE2/lK3iVEiz8yHQy1
+OKcNzr75cAZ6ZenmgGilwfISTmxEZAXKVmfWxCWAYnYvCJ1suT4rRXC1VmBO16yiRKG4WdSQiHn
vQGsrWIimDMoOnQZgV18VbJTCU9AajZHpcsRAIiFBCgP97S5OwvuefMyhIc3Ax0oi2a3VllF4qpe
ZurhPE0RCnMc8MkWYFNR2qZXu4kkeAs3+1081SbXoxV0de0YpaJSkndYusdlIz0qCB4st35LqM1J
Lsc5DEuo9jie6z4G3KLfh4rorZxuq0LmtHFLFD0CixXA21eN0ui8+J93EwNcZ2Lc11wriFRvIjyQ
4S42IDqvgx2SJRqTAiFwYye/xHdTIYz4hXuWs/2V393zDA6koJNplav+L8RCX7ske4ZWuf/7AbBd
0+1NpDn1yRw1sK/djZtZpAbP2UCnNbQqgJFWSr47xhaGHsT4vz5FYnGjsnJ1zNZWkqFlWNwq6mU8
VPghGl6VhPFwbDIVDTbOBt3Xrmm0iHRjMazXxI+JFoBOhfEtI65Joj/5/IsRf7WDbZW3g9sClpwS
YUNOQmq6OLs2VPg5W0DMBOD7Gk11tma2yBL98GBuJ8DOotejrVdRzUyVWmRg9d7GsGacIVr+Z14s
9yeBbNXk9wn7Ev7gggOvHkKTXB2HyyfME95dmJSquzWmBXliKZcHjvPxUgvGlb8T5HbkhfE9SseU
Tq/43NUUh90R+T5JPrsDY+SyKlKqT/7zK5hXn2721rTFI7zBF8L6eIwgPd3nwR75FFRk5tZRjU0E
N1dZukUtovhKj+jzg8nkWz0V0vpwoDxlI/H6CSV9wlEuHp0FPTyf2rE+pRqVxmfk/sihD4vouT+g
hxi5wKcE3sqyKzzOCuB5sE7iQhXKLau9xmnmSCvztSW0s9cs4BMYrOPW1oc/VUlXx+0HjKT6E1Xa
uph7HnZMhN7kg3VjxY1iajKUu7oRukCERep/mfpVUbMFMEBNuqNlFvKGEuilgwHItADofnmkOD0V
eQa31US5Inm9azxrkCq8hmBV3QzQtPOiYQQeQTBSTX+G6SK36ZB0UMrWPwsMLfZCIdZpbGVflchi
U9yJ+yDjXav9bAVYIwxbPE65gzrNSaJX3o7eAzG8xGGRhqpf54TgDs6Bfp82DNoN6PVvtTuabpxT
KHNHdCnCqpTtYkQnaliuWBxxsIbO9n1yEKt/c6tqBu+03FjqLpjiZWWBtdKsJs+1RP20NC9tLxzW
9ibcGceQrNRnhtridPPQ1aFQ+6/L0sEtyNhDTzBbqoHFMBUnSbfOzAWWfiUIcczCxMerstx4befm
2CyMeFYJqbIPsIyxFB5FLB4VGqGTaZmGWPo/OHagrfa8yaEl3rDKo7zWyNuC9Ph7hLZZMa9NZDN4
AZSKuDbaA6ztdykWIrmvUqJu/OUJ+lo66rkCqv+zkUKJqKOujwUfBRzWOpYZTvYN8f5hzfZx0A0r
jJp729NdXO0i/jjbV90+fUCzgaw6iFfBLR/HYtgEhIQ3nF15zTwfIDTJmWQtsgYu7uUQ/3i/8Up4
kXUu1ByaEINAcdUHvLyfNZ3fOmcGpkxZDjcPZpoStMWhSrBQHclFI+zAu2Itmq8jvEBkMPp5C4ji
cF153BDyACBUs7Hp6FL+g3IwCxP6Kl8I1QBCTmJy7S3VIy2eiTLApYW42osSMTBmMwgM3pkknfkN
2WYVSjnA1MVLiNKYMjzPumvqVQ0/2XdYl+4IYwcyrEK4DlBnc0KbIXAOSfl/QiY/1mfahWMfhS2g
oDSlUbOcB9me2EMqc+0j1du+G+CriZHiEAwBdrEiy5/d5Y036d1HbUkEOOvDoonTPbZbqbIi7fYZ
aHV7lCApUEgK6QOYbaJtnD2djlnozQLzMdEPBawyYLt873ZfAssVkDTnHah+1Dsbv2DmwXgaXIsQ
9cDHY0yi+qCWtqC5f/snJaE4LZCE3RCb3rADqwWhsbXvyK+hVYdGjyE3fcfTk2bafhfdzmuPdY0B
k1TEM8aoCfh65p0Vuc4v9ZMKx6uAbFq8G3kpnyrYXN0oWP/w9I4P+TvUAnylN5u+YpervVLYJypu
mIb4meSv6nUF9ZLS5fElTRuTVyj+HSx9Aw6Ekvk1S0RZoNxQKjRcSSe6JkzI9ldAscDjPz7bBxh+
fsYOOoylvY6gHuif8aywsTzNicxASVJXc2huF+KL7YJQjXYlra0l7SjI1ZEw49CbmLqyM9Hs6Nqo
MBX1NzzN5kDS5yJTYAqpTpEUmQzrV8iWVvqwC7tSay/EiOKeO08tlfHrrC+dogqxqtc9oAThQ8A2
1klXd+74ZBFYDzTSz0KleBKjhCvkJJOYRG4suWH1puSdLF2KN4C1IKFxoxI3LEJqdnHwSTize4qS
VydkdPh3pPDNKVd0IJgGG8HNy2Lb6+ln83K+1M8TcDt6aZ/1EYG2MVoyoH85xBbiMfCpff25PmmM
ImjmIRiBlGbES8+n2nQOvs3sgaqXpYPag/vRsKrYlUHCGHuZHNQjy+UdCoa4q338l7NbzHKvJtyw
HiFTdcZNrd8X7y0KpwCaEgy4rtYGRgZOKGcyAc81r6w+6FMtd8YkMCC3JdLe6CZAEShSS+gPVu06
O2r54A+/SdGzODZGDrdsY5roJ5IbhJs9qPh0vgngKy5eQG6g/VYzAEEjK8HwXD83+BW/hHzownBN
L+kpIuQPBCN7uFtU+r3EtveKBI1NYqHtH/dlK4RE0c9m6ExpNBWRFWmIClr5pfaB8XL6CsxmVe6+
VLu2CITZtymg5Fa2M0Kkf+LMLIzsI7YktQ9BPYAlL3DVBmoIla5HqbmnnTzGnGoetJxvfOI8bmOx
ANS/j4o3JJ/rhMGGzMO9xWR6XBiOB7moVYUOpNyHwZB3Kdqhbb1jKHHk379UukSmnYfLFXKpUNno
eBKKBuNO3uWO/0j9e0Dg8oXS+8ROTufej3iwOn1eHeZ//RIPONGxt5fmiDcd97jvS+5cMdurURJn
VHIcjZgYk5GAzfdUgvRTUxnJWF7DemY0KqgSlktPehR+haCRbLzk+QsybLMWK4UQ6WivoiW8fnw9
AT9RKUYUFqnq+B75eKd8QhNVFaYTL2LZOqy68Qm46mDQjMeKwMr63Hv4tQq+uT3u/DvSU1oAQ3Em
YI70qlJ/J4Ycz7ap5IyzNORrh15ok+tddW2f6+TgWwo5oMgLZJ5onWL0Nh3n5EaI58gLi31rYnnH
j20n4Djh1Rlc73td7lGhHcdH2akwSrDTQdpS9XKGI7mMisJFFHfAUOw3Hl1Bo7SagZIPKt6G4cg0
EFzA45A7sV7waef9GnON5TqoXFyfmeMSuIcJ35mVMt2eyaXgZhv0u0SU6CFo9uvp5CRYjUj9Sz8J
497qeK16k0DPzderpMm7Ep2XUdJx66l3VFTdy+mYO0CntXnYjhwFcjyJ8nDFbTU5lMqyuMo/7MF2
OfocilWXGiBFK7dw7eIXwRsI3Ie7RzGORDXDX/pQl6uEQe1NK27KfXb1YS7nATmyxH+g76gMk3uK
2aek04s0UWHgPw4Ad4j0NcagmILAmbSughV3SRrqYGp9WdCABEtFivKj264130NJW78cftywnshu
I5P4+p1LUkm9tmu3JtBsXrYVYYzkoM6oH6vHi3VWwLDD/IirzMhkxlY3UJWX0V2Z8s6jDxw5JpVB
H8EM9/nekhbes9+bD9R+suVowVApSf9244YTsapXXpMSjTIeT5q8J5FuzvPUEKpfj7aqyaZSc4Vh
F8SwIK48fov7MWAFzmU5eVDEHtJabkPS8Ww/wlDgB7zcY3G7sVnye0Ilc/0G1yrh8kzrrg+9BkYJ
PEZPqsaeIfAzzKY7MahAgxFFYK5KczZpBGi5tuTNdLRXnZqUXN+RDh30UOXihcf/6ZV/u2OPuzqe
d3RkUARqMHwalsjioq5tUF5Flb8PCgA9hS+qkY0tCnmD/tl8dwFnK/fDehTcGtO6RXMCx1/BBNPm
fiN+2VWvULA+CRZoJ5aDZgqsnaoXBtnuW0p4kswoqucrRhl/aRymDEME2TqWFdja+tfqtz/wd20b
yRl+s6rAFjW0/kuk11bPQta9kx/NsZw5EnpIV9yzpS5KQ7mgD0kc1X1ZI2Q9Lq+wTXWw8J5vBICw
hTK0ER5KcSDIHQfgZPrII7AxQcIButX9GmRj+mlXk1dUV/UY/DLHuZKjdmrsma4huYgHF2BvxXkn
BC1FoZSYmcNVTgMYySRL+XJfD4dBJc+WIaijFfV2XW0/ag/hW66u4/bHHTLuiDpBhGdjsJuxFUqQ
i8hbnQM8TYfufMlF6KjhYuJ17lP1GROD9vchs9Y6pwhpeTyPWxw0NDWF61LpIxnBimtB9npiPKZ9
H8+opf3e1gw7Z7NWZOwDJqumIx7jxvqhCB0xsXA/d5QUO3Z2DKJQGZczT7W6jkwcVlljNrBbG0KL
OYnCKzTAdHQ0AgUiCSi1V/utWC78wL5ykS7TmgVAstUTgZ0jFrsiNvP3WfcfRB+T0vmjjZ+Zo50e
dVITP4sFWuOyJqJqUeSWju98qBj1Xh5vxA+YMUeUnX/WArMFqGC39Fwdq4cjfxk8FEQ23DjM7O5K
Nh/12tYYx/KG8xCMOQLl9V73Me/q0KMdiinDtxVcS1ooJVEf07sLwnh5SDgTz1w3sGEAT2bWzTxi
0cOREwaVuUf7u5MSyoh3bzRt8G5jHwxRvBJNQkwU8T1b+b++bn/GEizBhjRv98Pk6tBlI7EVMH0n
p3ekeRK0iKJ+AraTpE6KK6J0v4xbsUWma6Q7sHB4aSLsE55lggo92M7eHjDiEcV/uQ1EMcQvmpps
0EQQoDHThXbFt8rwGyJfB+asi8QbUHnzKmiXprdw8yM4TergubDhqc4m10LcdaMgZ3yPaPl1dg1Q
1Y5n1OVTTpn4edJh36m0W5KFbopzdBRBw87V5H9NBZUP0iemcLtkH0Inb7LjGAPrWjKAaNfHbEKC
DFEFOju5eJVFD/HruvxrZ8mI92QIPVlsyqaORViTfAQgTcwxNNtpOufPaHLEunvkcnXmasD3sH+L
vvYLVDUWAKokXk84hUFXWTTfKE0pQmphMiDGmDVjUnsotEX5dpdqj+cVlF+azSmu29tdmb8ET1SZ
om7VkrDvTJ0Fs7TKnR2flT9tgOrkpOJvNak39t4G50lvKu97mUOwWOlwYlX/p9xxkrMMx4jvTju5
ZtVYQimDGXGd9We0w0me6ZM+6jQRGs6xsMzAL/bqflTCIEr6s4jNro2vfXMw5PQ7lF2tV+F0DCT+
qYDzXkiLy216Pn5pU8rL+UWk0fmE5FNlZqsn4UKbRyhUpnazcBlU+zBv9p1mnPcOGp/pOY6cbgKT
vXnIgp15W24+eoLhyFYykzcFPllUpihog5qGpomr7d+sFJCIIH/UpPWeZ6ic7OJzVxTspze0uXU7
dxleNxkmOQgfffi2iiYIWEpC3c5E7Dmief/eJVpp2pWYRdQTwMN4Z1XOeZitzbekW6j4Zv4h5ZMm
0s1q1pUqCvt4y8xZHVJ4/r8me75tRJTxIe1q++hph8RyEG7eOBSB0H2qsXdGwajbs50frcQxxp5/
Uzkp5QkAtjfxuuihcQycPmycdEvLpKrvDw+fh7Wm1ZFUw0Foxg7U0C1oxHUwX8BZ/4ruXzECMF3W
SQBPUmjmkj1CNIFklUh2gRj9Y81T/uHxqnZSR2FcmczEsz65SO1OjFsP96Eg/AfrahM1mPRsGG1Q
RyxcnGpvqvsMJOnEnPAzXTMfvBaOv9d5cDs+OHvKdakoYS/96rL6UrRhSh40ipkg+wML3cSATRJW
BIF6HEx4mrXbwxya/Cdei0lTAQId8wI+HEYhYxBl77jX4Gpt62HxiQjmkKk/Cm8wBM9pG3lYrLl7
0EJSV2EyuHOesqbW/LPD1QGBmS4IFBS8DKaw728xdGG15NevEQp/f5FJykVkxYjlNlUjyqHT3kBL
g+s49iYjsy9dMnS7pKIYMKhffDe1nLT1J20CLPJO7Pj3a8k7Z0YvyiaSUyJE3LhvLCibAPouwa7Y
WqSP/aFdeBB0kQF9KzvBJmW1ziTxX2cB7B8SPx3FQpOqr7A+xVp300wsjQcARB8HPR+4SRWKtQ8M
w40pnGEDM+Wv/NDR15d42Str9vZ/IeH6YEyUW2C7Y05xmlb+a3URSnqtu7ppsqe25ZtuHB+K5mwT
q9UkRLpGKUmH5mWEV713rLPgAz07YduLcTlBHdiR/4RJUo6RI6NR/YPWzPMp10TJvprk6XSzu7ts
ePzGjRxwu5iSXcgMpqP7tzR2+wkT0CIdZrixrpgSbcFsz3biGXypU06ilwbeHvidzMMgTAmsjGb2
4x9snlPSlfUozfo3x5+lC3aTL1h0/co4SsPvyUL29WkJLcKgB+SQuhe5/K9nrzuCG5vbX3h1sQGw
VAuyAr0l3JpQSYfqubyZ2n0aVN4Bff5Ux5INs+nWIrL+OZt3nwHhMIaBNeywMuvtyNn9MOn+cyco
lS2ZTn6a+TngWROtEKzDodCPPWTOPr3HRVc4G0TooKM9eDK2mHpQCyF40k/AuwwidwwjywdWubxu
lXYxGQd4EgITeakeo9npQIF6u8QmbeB2u/wwCX2p7mMnoPUUyMsEBmswtZFaWNMJ+cG5Zo942pEk
feNcFTPpFrodqckGXTYM3+427DTPWm49p8DfmziyYykmQgaHJRwp1tBt2yqci5CWrCqemfMDt1OI
JL8nE84rTmxLtO2+VxKJtePiuUp3ZEV3WtXxsq4wFi0mmHS+3PC+bTYbyRTcDx8kM42pwfGKpI3u
RPm5EbYcOj2j2ZA5XtFhf3hA3PB5xHjrHMYddS21sV5gJTwUqM2zAq4u01uVg0oKtBF84gvJZIYI
we73vrFTWtxZEngR1XHXvYDkpsAEqCrEYDAbMUD+ht+Q2se03IW7RF+AbG2Rw4PvGRJIrkG9aNk+
BpDfN60vFlAUdqUxXOxsxafBNH1If+7PAeiNM33XGaQsHlgb8QiyrrYbFyFXn1AyEBq9s08Z77w0
d6bShenz16BB5S5gFg49Av2VeD19IQpdOA5NLUCps4oM+GCkJRXD4hB6D3N6ICqAZ2cXA2cHFKgi
TM5oASTARiqshZx2n3kQfwpIfLmVsN0GM2q/a4LIQsoe4oNi6wd9ZmRWTEMst2nbRvrHSiKypI1H
jmkDcArojl2WHgXVZdzkjO3H/UV7OUF0a1a7cRjs1L09OlXjRsWyJUjBycHWWcmVnQQ3ogR4TgSd
uzlClYt1KQLyKZC7z+t1T2EDRw5MHrR6o4ahIB1j+UNvHL+r520VR1nxuauavzh3X4hvHISPT70Q
mqbJ745GQAlOcxMqpMmHHmJmAjWMVDjVjmUk13L2QhudtSvRWQbtebtZNG2K5wbcJEu1OHXyyRlT
tR6J/m7+Ipv8wvSZgbJKpDKtZjbg77Uy2aI74XMr57+S75w3Leno3PWEmU7Hmkoyjbc3Gf4Owkm0
hYqCeXcsRgkv1kxhzLEfXDde2SRSFk5nlavVNXAApRD6W11FfGOYlcK9Z2Zy3mlUgauIinunC8uh
oSp/ez2PWtsL6dssvaDB4xxUxu3RoyfjQg2e9avI/+WlyrFQrMDELdZ8wCrZI0OkyO1S6x3RnHL/
J3GPR2xT5ZDsT8PXJAZkWAJAVB+X1616u4BwvwIuiMHWNupUwIm142VJiErYNnQZCgeVZldBvQje
kwVvuQbezZatT91FStQRowA3oP94fjp607yqL/FN8VN7CGDy1TMQGqkqDA+c/xB97XrCJoX6aep8
Mx2AEo3y3ZJs6dLWCmpoYaSS0RlTgZgQvKRW85sI+0djAAYU6aloLri3tz+M2kMRIBo6LBrk1n5D
0ip0smPT2sOj1M9oi02Kjb7SWb5kG9WxzPxA5e40LxWsdYk9LUkLBBLdbOgmBmtXbRapuCtgzylM
xmBQyQjSBm465ElGqY/pzpJQ+XKkoNPaC/zf5kt9PlI80WAHxQZu4x3i88omKgg6f3mtU86aggsn
GjcaaPLXmDI3PKbfxC6csNTGH+3PCMB+u9FX80vssleS9rnQZZ5YQb4vW1MDNrv0/QHmHqnhlwPX
KA4Z+7QHOJVxjYS3r/JRLnfzoAjvmI03tt9zuCLxg7AWN71shc5cf+w4r0kcICDqLdNPEOad5Q8M
lzhjJhqzS2FWcMWWmjmTbwulQXD4Xq8V7kpEyi3X05VLLNNnFnw6oeKLcHRbXDqHrBv78tOtdaqi
zcBDrKDv6YzchB/clP5U8VeuJCtNCrm9Xpz1u1AIsvOJdXJRCV/HeJZR436OvcVtLTfF+PSgltvD
bys0UwMkVIkRmPDzn2zDk2H0u64cJUXWX/40HF2NVzzLC8WOK9IXYXf9CqOkxmkqeY6oqlahmGIr
y3TyfoPZdjsl39AtGNkE+0ueX+rWKEM6BE0IFL0tOkF06A2VA4zEv7m4yzpi+g0l4ziCSpjh3eq0
LqF1q2qIJMwyDYDlitbxvH9Zf/aI0pqbTiIHXqPyK3TnfewyIBzX685TXGXIG4BSaVwLeUCG7x3s
gKRsvizgExplj023tlV2TkSB+8IdtdWoz46lC/XkVZRlw2H9MEyeKIQD8+FeFIEStNpcUf5PqT6c
uXTqcEWFw06vyx5vvAxbhP6whGNADSnUc2eAJgDCXBdrSsar2xjbmou4yPWEcVgkmDGInkxuHLKP
IVAO6hWaSVSmhtf29BkBPUwK98FqmuRSOo7PTKgbgj9Sj5W5GT7Si6UR48IcSFRltXUxNCTUgLNF
cx6ABtk6+U8nGgvCwEd/SIPcriYfrmIxIQS9gQscbR1+aXuqhqVq0cgq5TBG0kLzc55otTspByQv
ZVColhUMa7e455p8PqvX6kwGD6F/PB8r4lrRlsDbh4JnGBjUK7+xFLlqmYuEkr7vdkMOl9JfgmsZ
heq+4HVPZqRc4XqDBzV1AEI3HQQv0r8hjFYlLKeIFDhVg+FUmsYoaH1cn48RAs687GgbrFGHV3wJ
nbzmrGxnCslHeuldDgIF6CWKFYO7sI82etprjYpOwnBiweE4BQhsYmGSpw3PrAxt7xHGhEr7EFn9
z5j7YlzRowrCVYvMXBZSosYD+jh3VbiPUySdjzmsynru5adb/KUtY51pzi2pmlB8xd1DIZ1rHv/2
WQ7oO51PSu6xADzw5JLmwjIKdjaOSg3jrMaOqBZGWq4frANBmT+kC3f7IZ2yAzRbrsZ86dlcOICV
FxJMkNQsGwmdnmPv5s1nMIsxXm6VgE2Xqi4fH3a0bjSAZCT+ADIMGT0BYrlKv9i8+meO4keiTQCR
CdVd3XtLBqOAya6ir548yzhbSysMMoj8PZILuwlC0worI1QcDrUAhLF5p7b5KFjwC2Gxjr2Revec
DLhyszczHoDswvFZsbDmF56K+toO6QzWiMLm1Jpjy3Mx8Jl8Z/Mj0hzM45Si+Ts/oJkTa349jSEV
ZQvuXTeALSLFtrmEYz+ugq5M/Pvjfvw6dD0jevGJEowrIFhkAt5fmVa1qIU/rJ+WaQoTAmoTQwDX
lBQkBerVQMC6j3YE47LgbaMdbuYP4NWcgj6yfV3HH93xzJaTmgqk8sYHYLKf98R+67JzMFUBfp6U
nHcQ43Ejmgr2De4GM6q/2YnrqxZLMpP2uqO+P3zV5WMUF1pJIqftSc0qDw41+7+DtpffVZYedxqD
MxY/cLgjyA8bmGqfS8BkVPm7Q4Y6T+7uTnyYnpZVyc8XQePa9ZdiYDDQtRnqJor7hoWqe5IyIr/i
q+y04M1bq/NIfAEt7Zx5WIOhdZyHbzUWh55knm/gQwbi2rYlyz3HjT7YLosrkR98YUHysmB17Ao+
l/49HsvIZVrOcZv/pJG9/QdrAoad4x5wWFH8+E2Mdxnl6WFK0I15c9CPxhuA7/Sy/3km6Liz2N+9
wxTtMhUH/tezLBGc7I3ywVylR46nRBdhnfEXp+UEH0bjXbrUQC+1Xfgg9AjdaA6HnvEoBA7NWuXF
1YTVStRRqjM9iIc2DGDI2aAAxukAVGYZrwUzWQihURr2nslz82MblEOkzgHhtUc9O+Xi+NFF3uMZ
KTQigj/awOb5z5P5QY8zTr2A4XVQYmUW0EZsdze7CXV5Qc/zA6UHJIJYlSkmy1yapSqVQvNBihHG
pD/msl513hc029BQZsgl60VUtNV2S5ptNeTFz37EQJ+YYw/ySc/EaMDatg2Idwjrx4U5EUEN+wms
aDqSUQscbSBK4QWiNqbyUhwzsIUwojMd4A1HvuiQAqhd4vZHpov4OKRA1kT8g6BUzRC4oejTRml5
MiDEAmfxY4gsYUf+rTDVDi9vtq48a/6gr2BLPl5gV46t7TwHIdQJ6UawPK+Ah5HLaFNaMbkZQ65a
EriHy6BGe69nNrZlGMU/UkIj8R+8P6iQJeYTU0WarJaPzg7KxwYZZ2azzEzVQIvCY+OCnXICytsM
U0HzwTUpINDGzQHGH0vWeo4srAwjupddLbR1l01CspVLrLvZ0hYEO385+HhsDmaYOEMlEgHy7H62
WQ5xwUPS3WSROGaAcJ7OrHquUjpnfm+7cMmGnkQqazo+GVjDB4CAX9b7g1X4oYluwv3AXQgBY5fB
KZeXVym/sfk9OymEmTlYT5/gUWtQUtGJYatKZzgfMUMLz1faVYYhTCO8s+TzyVLt3SNlgYssMc2k
ZOaBMRmYcdYufmEnzry1Qg/iLtmh4jSJMIFlz1AXA8H2Z4AB54bMSlGK8IEQYuEhnL1WhZbV6oyv
Qd7QrO2d7Zu1Iilb5SDYxj6pzVtAi0X/oCx8gd/Hw6ABphMDG4cwQZci3kQtDOGSSiqHkPnSJFwB
Z6leHXWILGSmQQMNJpD3z9gS53G6xKlDQLPfkSwl8RdSzDt5CwQxQVPVlFDtbhtUq618qxvqEGZC
l2ETkg2ofMpN48O6gqK0UBAQ2mi5oeCKkKmqWsdsIYJEqKhqhbLrzKMQP7ebzQ/avKlkEuyLbNgF
a1VIM+xD+S4jzx9vFvdMs9fmvHNlimmNAHKwKonQQYT6mAhHWo1mrS4av+T7Ykh0nVYNmDPMy0PX
NG+9MaUrEvb8qEBqqgvGijIPsmYR/+OwSky4FLWWjGusl9yivu0hav9wMOd0Xfl9p+5tewR/rwcI
WOzPmWwUFhGdwbJt4YvpilcLItkF6xoiD/1cAxIUJ004o328tmFN8rNDBty11NpP4MOY50g4VPky
M0ZzO0FmbAzODeIgxZemIfTgRsFLZc/RoJecV9/v6srzx5mCMsU1nVCyOKeSctHZ1oH3XvdS/31c
8wr80PgnkJ3b4B5TlqfOBQDPrEQ9oXeW/q40lxat5D+ar4aXgAEXueYwEpMluya5f/2jURG2T3QD
xvULD3FO3U/KZIxRJiqjaM9SsCeC9dKX6yYNk76wHoXgszuM5F2wEOE6iuFjCje/Xz4rVye8AeMf
YgOcQ6T/crilZqv0j7Me/y1y1EyiDKFF03IWAGhSAKgm+5d8NGXACWIgEjOzeOC06GIs2czH/sHY
BA1GTF/vLqDO1zUvG8fC7wqEq6sfMf+QOcwI2fGbYgszxcX5r1IlRTEPFmvzl66H+pxBDpuYP4Xt
SiBr1JJyh1iW1MTH4FPxYNWECJOxcV+elTZa9ZebYw/a2S9opEvA6vOqT2oMWRJQhfpMb22ULKlx
xDUeXoVAroogoV9yQyScC1/RCfWldj0YGlN8pDeX0ISfsLTfHQOR4g+Nfh3sd/rrxQpXB/l4WMsq
MkCC2ncz/ipNVCrRKye3lT5z7DOyOGr5PP3qbtAQmdVLu+67XVFajvxjzXPHcujy4BC3IrTIiHFD
aoNb4cBi6YEABpBlLTL+mXFLIBiZ28h/jKfJzMzqiAeaGtv5GS7lk/Ab5SmmmtZN4/IW5G9kKfSv
oy6SLnx56jKZtu4vLR3JAVi0k5T+EKeYYKUpZhcHXRi5JLOadiM+MMzNTbCa+/BrJPZl2plvUtWs
eEAYDOO133Qx6r/8FiXpoL3xJQ6Vh7FK8CLG30uaWoc3LIlQHPHWj/Nht1qajD5LeRbZmrZgtAGx
LE3dKQqACyZiZzLDkQUBiR2mAbImlGQ4yaASIfCTducnx3km3Z5B05cGHxc5/kfgWPYdK2MR8cAz
RKhuU/CQsOZjfaqeJBd94Oyhn9FIVu2jFAmkkGmaTRAF5WABIVcJ7Soqef23Vom8NOHDpoz9zqEJ
ZwBdmTpxIVz0tdqApfCLs4eXBR1RZxKsneAs/vGIgeYfxIh9O+SvDfUleYH7ltwyDO6WGViwGUml
TVkIEwAylhuXREEZxBGWjBakZ5xnEZJfiD+ShrA4wuOguhzw7vcdVUnl9bPKp5WiO/qFU2gjK9KB
exZlnQR+Cjzjc9Htvr5NUw1DkN8/Z0Muq37otzqVjDKjprsu8yJHbZCQ3dDwsjtv4tNW0JcjKrEr
Qe+L9gdl3qAqrRb0hz8VooyHsU5dx8KxHMRMWhWl0YfYbkx+XUDTtK4vKesGtHSeiwIvDBqqUpbf
Ok22dXhFTqjMxfXCRjL3ZisjgyzYOr6j9VXUWRgKQdIod0mxPTSULSC7mfGANP7nnNamPwQeAXpp
OuV/1qIqEikkSHyRPTguSAjvh6H1RavZ0WZ7mLMAdP+hdbhHWzonk52BMnukaegXl0pSL3s6rNIm
QU2Z3uMgt527QhOUrCNDQDr3Xbu3HcDK+Z2/SykzfQXnAAJ8jHmnWn2pdvADa3G/4G4ieAw5ZtZ7
MJqIjkwIMnz6zOcIpxAZkq8j3Dwl+M/L9sCK4eTWrYpOnEH/gVn/GrlLa21g9Y/2qfHng6m057h6
QrA+AEa5pea81G3dJpl7Eh+eeeGfQFbL14Ah75YcH+l4zZtJD/50yD+MMr7mS14NjFtegFxvcSXS
SL4/+paFqcZWegElJAjH/21M6bNx+L/XcvZ7ztN2o51wpFzn/iiMthAMnP49im4pCMH6Cfa7RqA/
Gnf6HaSgvdRVIms6SkB9RF5iObQsP+QweodoTLXwZwUcDBJ85TvLHk9Q6+nj+cvPqlHP/eEYo7GE
n16sXD+wQAi32K/Jm23cCaf1XRAUUHwkCtJkRFTB41jShfGXyAg1CmNbeBGKlqY8Q1oOm3zRMc9a
z3Cd/8EmVUWh8G5cL2YmUYeIwf3c5Dv/GbN0RmMGu7VfKSpwv2iiCSBHDbyDNSfAm6QpD0/cAf8b
MPfYcIIbmLBKzNhhl/mR6Y22wHjP8V0z0GFFJ29gdIPKoSy9JiJ1SOmI/Cmi7ONhMqi1K503JUjQ
3JDmDviTw310xoCcrdgIyelFqmxQ0rpMuhYp+3HKuR/BAehOxCWyLrcecA8GuAZszFYXpoqc32Oi
ineMWX5QxgteNk5UOqS561B5lRV5DmX1XVLXbYG64LF5Y8GnoalMnD9KsEnYZVQjVdb6Rdo7evyD
dbB5eBuiiqYSV9ftyN24kOycQ8otbSjdI1Xb2D+g8PnwzJh4A3BeN7JjUjPww5v0Hcen9y1c8a1d
TDL5LtbQkee2mWquR3yfPud3iwhCs6OmN5ueqamkWRbQDbvsEsbPvAfP3mB0MLtgQ7Ou43Cp3vgw
01O2I7qZgUp8H1ziCHqqBfcfLG7XGJn9qB6voJvWVrfNcaA+5BDBRAzZ2NCcFJI2H9vIN3LC4mSi
wLfsyIE2K2JCSfkWZXneLLZ/Z83eYAbJtMtdoVlEfWv+CtFYobD11V5IHJ9fKNOMIRlbWChE5wjp
a3mNuaXt7pm3ggJb38k/3a+XKCBvWdNNZVsjsbLfgG9tsMoa8SvD6pDwTyKDYAeRDLIj81izI7Uz
GXuGR10Ub40I5+j4INPX0WOYLbLi0/xF8zY2WN6dd/zuRp7gdb8S8RLRYJxk4OHP1b6rxNpYQG+E
YCxcqyXB1RBHe2XQQf1qRJYlYkjpzXEKQaYTziyvknCWQCJSakSm98Pkk8ISnBPetJQuVh3EWYIF
5nLWHQpUf47/mid8YRTTUqa94OAbOnMQvh//vYsrGWDluZMcucFmhvu1c9kVfSmc7RKeHQz+aOmv
/uvsOh0bPhtHODeYMctl5GD6QDBdgjg/KYMtlYKCLGtlLBds1uv9wrsrU8hR/tRgp7gaPreKPSUG
z92YJw/ADpUUhp6o/SfpV5odbePyDZemdzgxC6mdW0Gvz43KncLsDxTTlHG00zdMD5wxZjkdUzzG
Ysq0aVuUYpDo/NUlkdXvz4QLeES4QuUQ3RgSNkR/sy4v6boNHOJR6weh6NLLgWysa3asmgcnUkQ3
VllUBAZEp878tHK4fjVtHCIHjpw/5Cs64MSozKsZu5EBWhgnFsqXxc2NgC7hv5zH09yDb8uPCexQ
SOWU7fhwaRlpq2XV9EVCxvJBBd7H8TxpAcWot9FFEqbqbOG96sPaIXddVDenwVtii5RlAf7N1/8H
5PZbcTa0gK5D+GsV6do0pFOFQgxj1fSzvf3mjREErkzNxDA3+9Q6tXgvsDirvV9IGueZsclhQpmw
wcibs06gdDw+HBWkeE5F2tUn24wR+QKpkREWY5ZMv4PEBHJa3vWGM3kq5EBvvmVJoI6jBSJztY+e
VgfKIbZYwUOjCLh0QM2OmNgemIf7Ms2nMr8ghfao+OaURiwhzCf6EL8J5Fc0DcHkNZnFXWSpbMjz
/PPjyBw9YZ24nbS6BQWRuJxT9VSuVhhOw/lsZ/3++5w5kG9lNG2FpanZeZKLm1i9dIvS0zGZ7eYt
+S8dx7S3v+JYJqwx+AHNJU6j/7qPmJh9qctXdShqEWR5r/1+Z7zXbnlhFC3+Kjg4pWk5z1HVIzIn
doZ4garHm9hA6tJ67YGQ0984f4cY8WImLhLtXN/D4b6ugUQpcgIgBUe6ZXasMMZ0OjesfsUbYCiG
FLn2NwrExQqtYWfVw42vCmf6VZ6sOm9j4X5CQ2qJUcLU13KJlD8YFfrbtldSxN7wmkQvuvU8HS6o
ZLkZTyhhWEvC2uaNt6FLVffa0uUut6zWaN5Bf+Uq3+zVNW1z/OFmXs+fALTyuoXPyvXFXUew7M5h
WnYCqufvGXUf89VIsZ9++ZKN+N5g1SbHs5HP89jb0mmoyhA9A0F7dmjN1qTKw3NyhRAQ6MI/O2M1
WUBazVzKRYg6ygVG0xerKVRenUBBYyLnbkWurFotxESXfqo6tgZzAPJWaMSvXoXR6uOYFjfsYNxq
SPw/h7A34j8w6WQOMiztiuws4T326VQL7VLwiVDVS0xhwIHN3JQeiczEfQXIn+ejrqamjaXGKosv
qj4JBgJJrM/RzR7tx1sLZH+uioC/XW+7MXATtQNUt3xJK0qbkGY8hRcAkZU7mg2qotBJNlf4sG9m
8K4MrqhfMPloJCSbrjUmp9c7wtYalJF6f0/jnw48oQhX12xEVMDJGZuU4xUYlxSSsIsQ3oxIchAd
/pkic6w50TlRICi+HLI+cZ41c35MRDnVgYbUYf5juyDGcT6cQE6FYad+nKUzNG+lA9VIcNTg5Zff
HHShDAvjgqBcBS/83c5msj0I1AZLkevBDfYHsJKeQrrdL6J2+KwWTYS0rdQFUJpE2FtxSef45tsT
kJVn4l5whYEkWm49FJtEM2VI7laafol1j/MHFIRVojamkwYMPDJZy+XZCbR0gd2XZN93EMvBUHTC
9jcTRfTVr+tiA8+0cZYJPdAL35B400plK752Ec/QdZhCt0Dp1eey9+fE2VyUFrzmQJDbZJqheuEX
pxobVGTLh+OKXjb8fJAwMo3P3lCqGOxAkVFSW3hUToWrgZpXxwZzddjI8v6OFcBt3odZe5ky9zr2
nI3dJIZAADVpI5b0Tb2FQ5CZTcOIjxWJHmesDYlxmvkb9XBLCGVOmYg3xwiCT2vr4w02E8dRF6T/
qr7XSAIsJuE5/QGQK8dF01xvbsf7V0JiylhJI749tr5yG2PrVbJhzLNW6F8sskmaVNebS4wk3pTm
kN6176t4l8PH3mN1oJmMhlbrX65ZUu5yivAzkelGbXb26Lnz0QwMEYBX7igrS6fhg0nicZrjXpyA
by5tiSTjyzQBt50lIhZ5Gqx1iuN0aGVeIpeZ7b3IpM3ot126TjJvM46rp5tVFzPU2Sg7x5SQxvUx
Us8E3W84nO/aHfXZfMB33UnaCqvOUee09MLkGS/GQ6ZM+qCX3ffsaUzSojndYoGSu6nE7sevFlV3
D1s7BlZHO+fCc0jQHfgrtle58LS2PMoiej54+dsRoIacpAagUUrwl/cln/EukfIcxhlyADYUiQsH
glXoknp7l3q56Qx91Xxy3rhKfMUHv8cJRO3SfuErT+LDT9K934MWm2z9d0vKuwph20TmxZbDcwEQ
GRC896LJENLenST6HHvduR9edpaBuMHH66Pr/7f9Upt8QGRr5gYsoDcCSxMOxmMnLRUIh1pllYz0
B2IfcxyxOuORGcs9qyTTX8ChPgDN/BXpxooSanr5OAm/1xDYXphxMu+fvF7yV4XwBCbxk3f6mQ6p
D1fkyD/hiVwKiibTnajw7dBXx1APQ6wXa5Z7CqtFHL1t1pK16wt+iEoUWO9mbEnXzr7abpcCNXmM
+/1a8XkO6hPQt/FGP1MobUQ7OJ00HC622FWUEnWr1N7kcy+N7ja4IHUx0LSkwCucPMgelMbM/06v
F5kBPD3lQB6G4o71AS6BF0QDDEkjyUWykDHmZ+ANn2qVAU468stWN5yNYNQi4tcZmBxr+HGzxyAE
uRN5APQc4TGBBZaPrvNNed1N4kld1tTHBvKk34baW6cO5uCS3exTdeXZRPn9CqQME1b5GJQhwHqF
Ocg5kbxTp9zBc3vqmZs7swb813E1b23s2TFOxitFC4ElS8yVIrhSaJPCt/h1lRdXczqbOqx50tv2
0fTEHSnqtsYszuMdz7k2VGtTtnLUkLVdF0xsEp1/qGZqg6qDl/z45YP8QWFOmDwV6rCWPe1DiinF
B1fWBiQUVwAMKzflzV4CPvo/zlQ/thYqWvNroC5ium6fhHubWRkzqpSibbXEMwioEZnXSFIROwJs
gFWabT4EJShbswJQZVw0oznyn+H9JbPwLxXSRlZVmAQ9FxUs8F7TDt3uew9+YerE3Ma8HWn2h17x
kUn4P41CJHf0f/qaBT6zniI3oSHQKnwGXc/Kdu63VB4lh5VuHqNkuNQhvb/erTn/DOOCOgpbbXWt
tIycl2jZzwrgZPjrenHyLVfJvYyqM9wCdUsOzl/n8acHOloPNTtENyImcIlBjQX7+0Fw7tBl3NRI
27v3A/IOIwrFLYjfunTLkf5/18lidg3n+irs5CaJE1cpf2q73nKH2PN2Krnd7gXpvJvntycD+VGQ
mvvo2SddbjorJtGF7gtpNBpyWrqRT97e+7hfRMOTYIb94XW2hhn8QPEV+39wD1xOvaCKvyJog7S4
GTZ9vlviRRd1aEMi7z/vSxlpP1YZ8Ug0dFJaZiPGz3S0+yQb8p4ERW2GiNnx6yAFkAyvy21TST5A
q+1N97reNxIs1ouuzYSSLeHK/0Gb+gvIyVrtiwPvMXa1m9Y6soup4gHvB4uF+OVvhhDBzyb4x9KO
VRwLjFctaSsFsIErd9FIWbg3IUSTqdCHCZGl+DUC/JqVrWaZsH7GtPAUFLk4I0bZN1hb87yy5W00
NwyJ3Xv7iqFaadjsvHDMHPJ96JfIIuwWQU3x9rqrqhvObo0kIdE3aXmJ3a0lmBH0E5H2kH8GkcoD
fH6cewc5I+UxjSVSfLsKHt7S4LS5G6nuBYsQFVU2tx0OQLxT5ujDDXwkL0tUTGwXUB3t1CkVocki
LC6bzEh3cMieGvYj9wHzxL4tBvgRqiCHZrHowVSXbIEErDPdzRbjYcX0qIPSCZdKSfSkUS/0uD2P
IPlHpAGOaD5jTzzSReekBskqdo6v03W1HsN+4w+tWdi/2xK1ta6pKTSs6r0/HDfjPEB2oQK2zbOE
29HodknuaQGXY2kKw+mgjLV9EEDbIjdBN8fxaNhKmcxoduJvKiyYvHdrGkFshEZD8MtQBIhxw3G3
JkYKXhI4dC6oZo6eBjDqUeFF1v72vngqk9c12EZpPzbMeloshRVzh2EQngsLrLF+90XDx06Nmxp2
LcMJvFHeNM3+fpxC4OGFWpB5gJ3xdUtFbPfssEr5Tv7hmGFPn3GWmZ7FUgaBvplX9PihUf9V3lth
6X6Ptf8E/qqr/9wda2diEKxILVXrYgofabyo6eSnMtxJ/lo6KRH9ZwT0GAxG+VW9z8PDlc0eg2NO
Xy/psWOb44EAsj5dDeWosVhPkoP8yMLYD9lfuyHMrTxll0b3wuuc3qExptAwNkiKeOO0Iuc7eOiy
PlNWaDwmj5Onv6JOg5T+szQ/MIZr0U3BwRue5+fixpqtE+JK1OaXaCfhhrReqnb7IFK5LNBv5X+a
pb1iens88NoBJlt9vFHsmbiNLBLvdB0h+ghxJf9jWfzcesSQgPDyL1pSEY12TXZyJtZkBBuNTD/w
4chaAoiYB9BbUIir1/s0fzP/jWb2UHGBs9c+rmCmi20HnNiGMTkUbFkdP+Bf2pW9GXva4i/rp5tO
nUsceNZy3lc00jvLspETQEPxSdu49PZ6CMSa6VxCrdI1W4xJdViwlw8u35L/rR+OPSt4snxgzNal
eugs4ph+V2F1yYopfgETnKLPaYQ/aGaOaB01cMhNCSZ9pyfMODN2A8b9YF+wMXt3IU95IobMbxan
byaqPaf6LI9dzO/62q2ILsh/ZCK0PoLUS1ZqVH1cycHm33WwQrlWE/+u5H6cDuhOxZBgEDbDGkGL
uYk055nNrJ9kHnNw/kDsu9fFtdX0Q6w3rEOwgGCTCRYSjuOwJQUKuxu9gLdq+1mns/pCjhYxqqEr
HuV7jE41t6nkgxnS54XUYxhf04aUo2PbQ7rMI0fwYP+ECaKMCu80CbDGqkJ0Eqh/Olbs5EuCEGqS
XLHyCasllqCT68CtNZuSxXL4miHXSI2e3SSz6KREMveeLrNU0WE0N0zeXttlDB1+NmPVHoFbXo69
uSikfkoQqFwAFJlj8hDnIysKMxULTpbl06CbcHFCCQk1wDvTVsKSu243nd53zgCuuakNefsO0rhr
KTp+KFbkgAWXnqTgKfSWmkQhLPr/6gAg2+fNTIm4J5ssnDaHMbewCE+3NCndtwlrDde3U5zEVLZK
G0p93XCJcOOXn8jXB9e0p0KVlvcZrC65f6fiWmbwu4QIVySnut4FoQ1h95rypBmx8/twbz0L1v9l
wnr29EtYbImEB7mAY7mLKpMErHkomqx77i6dfzArt9Uf9KUXTo3nkn7dsHIYWWcRap/LSdn322W9
WPRQSDQn9j89btto00Ntmle5WdggKbKsnR+i6DfttHwLCYFzJ7AbkI/hgs4hIMIgOVW8zXn323L/
FwoKdTd5ZwarMB8zxKsWapTHGnc6BXVGACj/B+0nyvjhPaFTawFUrLGSShnEhcDiyVSz4iiucrjl
SBw9bKSgNm7hqHwAxI9k+eNzQJVbDu1tq/a8oPOL7hWUI0t88xKfiBthfRM5Q0NHYCGgSe34FjAW
TPjvcUWBQXf4iyCCadHMmiPUiCIyQiP9AbJVeTUR9EeZDtpxFUk2V+4tMmN/TLgYSrs72hm/0Rqd
fn8Zri8bX+ZNCnF3p5PGOG1s8UCDywYq9wtsjp7lF/sc6edQB3CPrn323+naTi2Z7XLGcUWlG3DX
kyAEr+lhLWjXHMgibr3c9g06GXs8f0EcZZkW3WWXSPLkrjAq6HbzAb98HOsEC4JuiImfeNBYKWOt
wGCeds/krIVJRLi3bgAlFBTZcxtOfFDnH/2nYxmZWghSdQyPX9P6pv8fZZCs/dEPZkHVKBt8yfGU
uuejFqx7J2tdDSi7D9pd+bDGDanXx8GKbJ8XPauXeRqc4ZdKeT9zMX51lA+ary1A1M5cHUjYZnMI
atfsFDSBzUN00sSkdq8nCeam+efGswiFyQ1AsZuEfQMQy40isCqepatfEuTBC4cL+97HId9KoCZk
3z8YTVJs0nsNGpzTNR9puaEjgj86AbKlqjZvYUnlCk0jcXwv5B7GT/XSCuBHqbf5CXvIDP8RVoza
Dn4qR/tJ70FLny4YXa8hzewGlItutZp9tZeUcKDnVkn/NNwgvH5ej0h6L6ieR8r/SIDfdQt1IYEw
i/Mj0QL5AlXqER4TF5nKKliaxZQRMczoARRmJ1IH05jJZjkY2/H/JhDqn/nX1Nn2l/F5TBOxY9+H
9PSgEfO5QgmwdW2IP8iK3NQjcGFnTH6tV+cfnVlyRiL2CXMeA2qQmKaNlcmvMoPaz2NJt15MZHAp
JSb6jvRyGJuCHd6Nf9wTmIFkkV0JHtN2L3Iu5ItpIGvpy3DB2A/CiC2mXs0SkzEClWKfCXlnFnb/
K7UlW5cc9ki/YoVLC9vFfRP9EWS9KmplqoEc8sRm4Q13828bnol/6x3i+puGluSM1Z3mIRo+YptP
fMmuMGiPQ1rBHGK6x1soOkOSw+ecd0mWWynwFqDf9r15iHTEcwRRSjgBqbCd1jnYoflWOvUfXra3
p9FzeXE0qQmdFTEHkFhw60EUmT4qLH5dzYuyGQw5xNy2ZGgylx+yWn1bnBy3iApsXVvk91pGBcKu
5j5VC+VMYFhK+RwT7FX307QfPpty7Xk3w3r8xwIkx+L8H6+rOilX1xYoyGTltAb7VBmnj+mXv+GH
rojBnpSD4Tn9RUlw2okC4exHdrAXFsWoL1+s2R1yElDwxmvU/B1hyXEi4BvSvfSMlW3Az6RohNFo
BRlTUOKRdqXMVDWEm2q9GYoGpbOfwFpEAQVVTUWT2wP/gq0wj8jpzSzyewifTO6XSkoR4RXpBqU3
SweIElN2vsLrfEco+J885o0qYOlz8Fa33BC0b0JculAYSTL6vu95Xov2FogbfTraIjtAWBSWRbxg
gWlJRTanrutZcwOzcL2iLxNfxQbU/NhFD3MqcG1Xzx8UXljM3uLH+kgFQ2mxdfZYswN2RGbbfd71
iyzdEZi5ycCinLL2+HyOcbHHXB7HmUOEqxQ829A7O0sabyfCID4/1gw6XhERthPXz2Ht3rYE92x5
aHRGcHJLeTjs1jz1gJQ9UKDbZ/Yy2WzWdNjRnBKd8nJ2bdCqZnV8dqxhaW8WfSKVUcykZ8jGePxq
Szm6TeDZy2/fi1tm83LQMueR2qygVjduv3sC8AyBkY70EbBSAKwqho2Bk7gImsvUary0Z2RdtqGx
Hx/nYxg9aBcP8qBHPHaOdVSqdlLGunc727f61/I1ZjiGkRljUOG9zC4NMzbETLUvykJPMXC8RKU8
/ScWIyTQncWJQW88yUHmW3GzZp0vzCQOJwCiEX8LiQXxf1YmXHIMSKqImtPkoDRwKVm+i3qHAHxm
Zlfy3qp+vv/s2PAXE9eaj16OssshHEMsJQAvFvmzFKzXF5gffyzaWlE6B9zF0Bck3NmumGxZZiRv
21OzbluG7YFMHCFiUJNmW9dYM7+GYK4bok4zF12HFLOlYgQvkg7c5Gy3DVpsVO1tXm5qka5+MYQu
HDqDMYEqxO7i+NBOh3Tp0kkONJ4BwTPiXXofytHeRMtA55N8Tv0jJDBtMsw3556yvKCEcsJzJcAW
hRhQ/S+vLTR+JOKYwrTIemJknQ7SbAHyIzpSUYkfcR5NmP75LaUaOjhkfz/CssQP5LLYs53G0pEZ
XVvCqfhFKSWyyYMt97LOpNqKZHpVf1affErmwXxkMkcypRSL9VXiaRfjEUhOqAz5D3BGrnbg0DHz
5iBy5rikj6CiFAOqvhR4crCXsPVAH4vvwQUlzoRs6yWx46OKFQsh4TXIVT/YACv9Hr2NMDtNG5d0
igvrzJ3aZUTClZ3yGlY7LidXcODvdFhhpTmsd+5ITDVbSNgXNvcdL/jRBu+yp0g39E9Mya7ZDRJx
bfVFholupHakYxapxYYNgrh1+O/olACx2l722QZZih4GB69OUsXqtJ8uAKWyMiEYnCVKaDPGXyIc
B750azmNDNJnjPxLElEzLvfRARirzVF+ZI3DGuN3k0tFKRpIFfes9IxJ/jjqWP4ZUivUd9+huJNk
/G2JzB1N/NQIhfu4MaWjqIY3TxV6vrx4C/wCg+rER7WpcJPT3204+b/bx/E5M1UGrhLsa6FeMSiC
ZN9eq2evcOwjUoBxing52sff09DdMcvUuuA5cMGHGvOc8wRuUEZWCIHVEAT2V2GgaIQjgAT9b6we
0qtnqw++UPxxNLYlkyi0QatjWz0zWQ2yvxuJ7uOmX0t9VhxtuKWw5CxsjfGPhjckXBKGW8KHv7uu
4TcNTbclk7/jq5ER7SU3TS8nLMmDy8ovQk7B4qDchsTcrTpF3nW00JxEOZQoPKdGlhlQp3958WQQ
A38sZ/U/Dg/rSf2AGqTwAdYhGNv4jgZ17RFr2916/0GYgH3+JMwwtPsx6DU5oL2+43Qbka5sO/Nk
PCcwrZh9Rs9SUaKjnz3plac01NezJlP+BmdEU8WqDhXMHzhXgr6uiB0OHlfgqdmA98L/QLp0h0PO
1/wfhu5JKxZWgyMK1j1kKyLW+ltAeNXYzl1Qgnbc8YZfiwCpH/QSrmqVg7x7woD+Rc0gQJT1jEsn
vnIWbJ5M/m44scLGL3Sxq4X2DX3JGxjtDOLuPq+iwYAMszdNOwm3LmLDUKE1NHixmORLtWW/4fI4
8PLFXUI2A3IvwnxHczNeDwYM9oQ3WAhaOzptMmlBqwMUCP/GiA9fSfdXXOr64ULhG9zAdirAW5Oc
D8SEBViz/MVostsKdEpZk9p4h511QX41nMwX8HGlFi5xMLKVMmn2o17fpjogNovpofg40RvngRMl
XJuXLxg+LCmzY7hycCMN4CFKLboX7JIz0NyFlZJW75knI5yrYQaVSaHlqqg5GmMXaWssnG1LBnTh
ja83vLvm1oLai/IHfyQMeoaJhFuSEyEcaBGboruHJshfpxAf/asSEbLnowYbMrDPnr4CLcflx0MU
+gUpl0/cSxn26Y7bJrTRtagasm/dslXPC8HzxAurqocIbbkgayfVdXiHj8oEpDPaKcfpU86TKMZw
DdtpKmlVZNOBFZLlTTG8yV2lHbaSAFgMKFmgu/K8rGVUYPtfm0XlZIvTqode5BIfx6eHwkI4CMoS
bmALS+ItX6WuSk+2B2w5P1To1SMtV+aIdukI6NL82iR5URn0Nm1cKnJ9FYZsxL8o8jxppu3hvveI
78ZgcgjamKK5M9aXMGc4lsd/gVDsgEavWHAX36oOHD1k/qJruEulu2vaFDKn5lsRspygS49tNHa2
+Tf43mTS1f6JevGHlGhTeOubXq7CKskzCNCRldQLAN0ZzRQg/HUI/19KTEM4vQO9IBbdg26qiQRI
s3PKaG/wfZO7Dxav5lRnpSVMX7GorHcNxhvBBxcCHHZsGtkObwLRSZR4fg7H1CpW0u+MvoPMWPT0
JO0mYJcL7l50oE7DqVTeY32BNQ7wWX8fAgjxKyj2ppf3IwVTRXhKtQrDSp+xxcJLpWwnsvfEJ+Qh
V3QAMWaEpIk1tbVCk03Wt4nKNRxzcaYwNoFJjeQiCjkF6W7zY1gMQ0XvVF2aKJvX4CZXXyQGWNr/
3jwsU8O00krdoV1ccpdSgWgCYj8qUKfOza6O+6Apqjk/u5LAQRBohcRiEKqT6c+OgMMV3UgMfqy7
3YrS0i8VotxRfMwJKFxk8oOaC+EKYfM3NSF/+uQEGHM+yHJT1DW7IQz60Q45lUXIwRqfkhH5+bAV
wk8j2Ktz0ks38M7KowMeACakcMbnkjbiApNyAZ1mupwjo0BsAwnr8cxpGCh55gMiXkGE8org85Ed
Mx57KpDSQxNmOXLWtk1l4gwQM70iFYzYNrbtvXOVRZTEzc2y2ZcVzxpmt5L1EmgH1Tq3PJ0HUEIV
aFN/A2Q0HjdzsAcD2/Qd6LikW5wcW2KhojAn7b4apXN96F3AXDCAWqE59Y483n8l8M3t61VeOrdV
fgC3tzIrqCJhj6tC5ye2+CZyrouUlP9E2XziCjtIblAgJeqDAINRpGpgses4Kfe9IrpgkVwgVpbr
gLxT/DHOWId4x8DM0CbfN/HzpdumgFNIwJE31YZdcTVRimve86HcGWuK+u+PeFwlOCbrh47zhOpX
3lMzoMviaaImE4uv2bD2QUozFO2f3A9jAzyT9xY/64OwczuzKHlm68yAxDjmQDpRm8MgCvCG472r
6CicZS6CUwA5112mcMth8Qe0WAAlGoO5om6OuoR0fAIlWReFrDmIK9EQr7/GM/8fGhu1WSax6dHK
u83IGNNWhuMs4P59QH1/3+RGj9x9fY0WHnw+dWfTMJIRfa3uioKkh8NjjXEkYBSlAJeN2wqTm5wK
+DReQPKxJ4KpvfKsecQ6c5DaGH7TZI4YyKauDqQyELzXvZdadP7yb50T8V1b9rPavWkx5kEbxxNU
WZoSk6X9g/CqA+YHJOJPUvE34WKyACHbYg09i+QcQu8fuf3TGgg6dQkS1jGt8sRT9tzyObcoMMan
8L54SwGmlLkTfa5fmryt6OuIr+1lpzKPrH8sq+B9TSTVkcYf2MNGscl9Fk5Dpd43eoox9OYfvRLG
L/9IZYQCyOfLxG1VzAuQrkuWuc1A/oLQ3K4nn72k9wekFBKRKUDX2AEHt9d9dZbotGTmwUPlKF6n
asuKb0efmkNhZsy6lKqFN8YZ0XVaI0dUKmUAzMzDk6sLBLvErk2yEPZmN0CFxnbHWwB28DuUk+1+
atfHTsXhOLFG9ewfNSoKn8Kj53D+ScYKkJYefXTd19f3cwAIPJIKM8aqFM21J4gWuQX/PmvoycVm
qZVKhVPUTVpHNHhmiH2c/x2+13S2Keuk0gKvZEZ/rlSeImHE+MtEXrIFjF+fUGV8oziqrz5ppSCt
4qx1d8zk2adnvmaYBBRhr2O8R4rKUyrcEtl8hAnMg094Rn3jufZUMhmdcuz2vUt47UNvR4PRCEvc
XH3kdaWtmkwKLSVDhUNtu8qV3uHopgNF+yk2fhiH5bt9Ae47YSs6AOB9Nrd1bg3B6Ilfhkngu09f
cJjYZQl3gs6k3wXraegNddl6avQy/SZt4qS2TTDINEUWxSWakOgHhQr72nvhvhrwzV6W5w2C7WY6
hQ2gqy+86LrRe8mmRQ8L3XGbetdaTkBWzqhCyyXXq1Da3nnIsafaiHtNvDcddQFyndJLy39gtWQB
Cyo4Dh49IECmwmvA0Grv3h7XPWZjO4SSuodOVUpmJtFxFiNrNX4Y5M7T1M6gNFv1CKa0sOVqcs2/
hGPzglKqE71B34VOxfD6jPV6BVGT346O2DekG6wwcyNAOtS6Uv0yOeCNsSrK/z2DXCS+WAcZn2z/
GY1WwIFbET6hxXxr+aHf/DAv3YGijuRmHGmbQ6WUDqqjFuRvRoCk6ny1p4ysietGczlEKy7bBMdG
weMkiW+XDoxAtUNdve1cpjtm7Qi9BhS27aaXSV/PXlaXV8CXutAOJaiLHPpoANtrxQe4/5J5bovh
BiYZcMO8CL+sJPt4rUaDrw1XVTsqM4maeNdyfP6rCl3mLP4MOS+LsL84FuwB5uiyomTsL8ZtgUh0
GL0DNEBnKEzBt/K7k+VLHC7Q92/dgdRpiT16thL0X/Bae0AvvHtu6QMhkS9KYOgP9VSJWQn+1wEf
znEYXg05VXkDofFv/pBq4Mou+f0sVy6RgxuLqq8kq5jsgqULNcIoz4SVqBIJ1V2we8HRAVat4aJB
JpuTcR79xVngb6ttNiR597/nHo1h335MYdrvt4cESpB+8cesh5NrEHkQPHUB1fR9GXyJNcwTzyde
P3fNVgfx7pVoA7FL2EqN71cbot/wTOLEwU29zDzIX28Y8lfSmLE+D63ICc/zXP22oQonGVAwdbZw
khciw3lD7iweeSG9WcBxLNualMmO5on0nXFVnAgkKCRxGZVmbteNBJCc6qExTeTEHoxL/JYNFA1V
ihLZgfVk9YJy74KW162pVn5zsGJPhDN+4OIIqOgn0N2WO++SG7NHjwUSY+MssVt15+Paqtn9UGL1
QEe9aE05UpdBkqc822AXF1Ic+gbK8YtigHtpm6fFn3EZjdlCb0YQUf+nPMVV6LSPGvgZO3l+ZXM3
98XWYpYLsvL4C4JGAcJDjMxgQlUEwneFMZtW/ipU0tQGB7T5LiH1nZPbLPf6DONRbEOfBHTjFzMs
HX+XR7Cl8Fe97dwucr0BB71cjiNdphpQq8kuVdVOPxqCh6YyGTofJFms8ETBObadTrG7B+LaYg5A
XvLcvpMOlvlwueAN3/WoT6jL7NASgIn1wvmWxDmVT7aZ2XAIh+04T3uNrk53fSOZarEyPzp/7BmP
RB7E8oDD4+zHOo5L+KFmLB86+Vba2wjI0xvRCZtnNCApIXHj1VlXblMSK2NS13ChSuN+GyAMJcbx
FS3IxUvEdVZ/FBqZLLb4Ccn7L54qYztNMXfayy9UMHckCT3/GFCSnYe7D3whXolmpVD70f8ksWKe
cuwsPLHFz2/wLIL6Fye9Li1FOlLFziKazVWxAUb8N4w9P3YltnFAuHEVIb80YxYUN0VS+kfNDmZK
irjPWGmxuu/0dZInO3OlBfA62tKUtwK8JU4xFbFIidNAMfZem5AAHmkaxXe3dR8zarNhHKow2Ejg
FV4x9mquWemhctDSQ1ebP48iXt6OEV8QxlIioHDCAxYzmZe+/yz1ObejZLM5aN2mzRsTfGU4Huic
3TRXggBDvBsciehs3oMIiP5OAdyetg7AOFgSF25dUs6Fen3gdryNWiwQ/9K50n8+Zo7w9w+bY8qj
CqfO+yZIsCaQvtgkrR+wYOx3owzrBDutOwmM77hPKN1o6sgG/K0RZHgx9Yx94wPy50AWwaePICzG
pBRmOAVJohvtabae7lfKqp77wFdKw62u1PBKUs1JGhB7zyepQPjqZPQ97DJdTEuxzGL7Sb4zg6kv
LRs7ECD3+EU9PKxrfJjXfJVZ3Xh0D3ii711GyVLNoygCMhSNppGm51zFu5W2ipEL/vxvf5FRDp+H
2WhW1XXHa38AL5aVd8T35zKnn57Uyf3+nzVBgB99Aqt227YQB6k2lIJf1FF+N+LaPWs1tel5d1z5
w+CWwJR1vRalepGTXB/EROWfReuPtKeJdQUJGRgdINqC3xPlyMACRPaqG46yt454+w482S7s3KF3
X6EsKAzZNUuifVQZ4hF0BwV7EuwuOUJN2EnzxQZwMZORwQgjMML7E21ss8IHIgryTxDTdtqBE961
+Q8+qYxtXHKxHEqOruI1f2Aw30gBL2ySWUYT/TzkgE7yzG9Rlqefe1CMTuXgSYA4RcXzTflBZZTs
1TbnSQPhKKSmZgqaTbucO9TKsUe1rv7WC7+/ZtE6+xzGXih6th46vpBz0tHUd/WAci2UAmNmSaED
rcnfalgtm1uHhCpdNvElyc2D1Zt2ScOKuSRpieRe4QiqDDB0lBvWTD/fgH+qZ7TSeuB3Xvext9DX
eYhmGrpy+ieoPdFAEv3jsv/IfyjHNeB6PE0XV33jWmIs0CTDhlAaKpwSuVtAC0rFuuPt4PrcDtzx
ZnNz3U55jQ4GgIUfDbq62XF121k8P/oHp56flj/n8URfOEyalrp9FyNPSYbi9n72e4HF8S/RPo/F
REXfGH2qq8Xw1dLYXHMxomuFI3W3Ky4vZHEuJFcCaMkv4vSBITeHTcLqs8z8v/zvXUqylm8huQLv
8+/dVOYspPU5i/XV5FsdZuXS07k04yATUSNJu/L27FCR9C4G5WgYtYez4rECD0s0MtoriLcUFj2D
sWRuZmIyQ6XoZ6zzUfhKjgMgItg8PCMi47Ddi5COdARxwBPqwYC61rZZ6/TSJP5wiSfjeGpWz5G/
zYtlZWIcagpiNLR4d6vSLBqo1e30eIxIPtJCjLU5zsXjEZQs8FwmsIKDjkHR59t6bOkVvSIBTt7M
5b1WxI6SGDGLbUrB9CmCpgZIFmp19axeiuQdPC6ctQZFhrIYKmACGnFZZEnvu80Cu31we+iWA0GI
TpLV4yooTlK32W0Vfx0d/kt5aWk/s3ybLmT/JUeaRPOAMe5Ecb6E1Q91PbzQyVShA0P/K++hJee6
I6UrVz/iwPgpj1Wc
`protect end_protected
