`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103856)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAOUJR+A5vTk/dL6QQdsRnb02yukpNuAQX5iWUpyHgnzVgJUZo2/dSoTb
d4QzzmM24kcLuKAdSAWVbsKqf3NSKJcwkGachkFbatKi0bSkABq80alh1lY/M1Cwwm2a7JhT6zFM
uaKrIBAoQ5AA/S/XA4tEoXJ/7mme3rX7M6IGfvHgOETsb2mVxmP4uSYTDZZiwnJ6tjZ3u9u40g9a
SJOYzQz72mOW3D9xtzfHSYJm1Rt+fp4odX7hC2zZ6EcXApHeAn51QGnYfnI2CMBRkKOtpN6XDF+b
V8i6/HKSELm8pplM569mOj14a7MUxDTGNkGBmMJ/VSedJz+wWDivTmGZzJtjyxR+9CPdaeuJ8TzU
QiDnhr0RO9I0uqcRZLg0N5wQXZ+3dRRy2stKMnMP26eVrn7cZ/bD40oxN8aLcXynrfzTB+yB6oX9
3wxp1q+z99fvPMXxSZba9EU/iM3M2N0y6tR0oZ/T5ro6OvUSDD5+luVpREhULfh4fc5TnjXNfasy
np4aENl/WDLl0oOCaFD/WWnf8HjwlVSnA+F0Btue//4XdiCm+nf+EypOXH0mZy+EyiFWVGgwjNcn
pCs7pnbKaB9CSCAzBcrhuEzgFEumYCVrUskQKWptOIjdJo0UPbOXeXdFLRRwIAaG8jM6vQOSd4yw
vxw3Cf/K7nEBghkmjDDa4oCWL0TOTsOGz6G2J4htECVHou+2EzxJouvJt72tvjuqDPxvlB1wztEE
JbTDYjFz5UPqFhG2aYzCKtik4DDNtRbDc6vu8liTGDtlkpSAZboRwNdGFeFXFI6Q+H53ed8ihzVp
8/8NV73kYhwW19MVIuG/ZaWwfjuWCeP1u2zIoNhWFhYntMer3V9vZR8Ph2Fel4U9qjOxPsvXIlLI
xkeC95KQnN9K1wot+RWfS+en2J6WDoXVFTt4XPXnRxWAcrLkGmv22qDpj3nNzMP8fQhhV51+ePGy
4FGvsH3DIwrg5iZV5GvyGYH/1VS2tHlcW1rePVOoKSQdlRC3U/4vvYYe4FH3IFNfjZWNrmI1IiPL
XVj781DH32MRa/O3tXxGCggt8CAitqpp3hvebLOcWFKfN9RFOh7NEA/HAeOQPToznXOpz9Phoi8Y
dcy1gHoT0Awh712UqnOSfOOqbiFwcF2g6niZAUdI56JCrn1YmFWgZ+fpafSAZpcMsUuSio4xW0zb
3Ge8n1A+3eDmcrflAUxDfebWcVJa+LCRwvGmN92y0/cJpWaOnXGbWByuW5fvh8xTzvxzguB2xD2U
WllpQK7aIOW4kmmDAh7gIgG9fyaODL3LfTXQWQlMk5nWA8EedRYjfEDE5EzaYN1NsuNPtwgVfbIn
nsgMyGVtTCel+JpVujZrf5ISdhmK8eGQCOff4axv1QE9HCgiinAO0ZXtlXxo2rC3Q7/I5n1Ny4g+
XC+iwlPBS7RSNL/fk8QETg5hAK2JFCUdmysoeVXEui16VWP9mexSc4ZLr1geH+75GUHJ0xAnYkNi
V0YT4m/YVW1lCrBqK1vr/M4is65ORp7PXl48NwTEMdklNee7B6VmcaEU+CtRIPLyb7bDLBIrohLW
bexGCufWK29kOnBi++NDQDwspvut5oyG1J+McxEaUd26M0veZ7lals1uuxa+j+Y/MshYMmIgoqjB
dDv93WXlZu6craUh3aFS7EUjnPbeN6aVa/x8SySmkEMyMqV9vBjFArx2/WRAmUfpAn3ybudq6RyY
mdQF1oTXmN2S3uoSajhSc5xyMYE3NU38Ltime3RVvkUql7H4LGeMZFHG7JuzJCNmsAxV8leL5nVq
gxLfj1N6n4r7sdHXWije/N9ksBBhuPaNPDF6b4NFhqo1iCvOJEg5wGFu8g4fxeYcdlurQ8SEbsIj
+1begC564x1sZNbqTNcpECcvHW9d7IXZUCpRsbzxrWa1eLgBKy3gq8aeY0jQeXoDo/LomN25er1F
/XbY0ty3Q0ZTJnImS367oz4MLf1SFlm97XCoVVQNPm/HRRCh+LIQ2alYCAhe9qCOBM1DnNsyFDCC
X+JTk70Q1+WKvkPdNixyqejKCmXeeJ1PIdMZ3SEY6gdACofGyHaZsiAqRSSnA/g/2P0uZRKGx3/4
Zbs3oNhf6M+0jfpRo8ttvHDFq5s8gfC2A8qv/wQ5eyuU9LKM15sWnOfkom7I+nGr81fUJS87uMcd
7a6INHiTzbrUmFkg76PvRSI2usjIrleXO077Kcy2y5oqf6f3e3rWkNgyi0JjmRGlN+Zyv2Z61iiM
afF35ill9AtzisI6ziKDW1FePRK9msvF2/1wg+vfM3o+P+1YDkJJ/D7IrKpblfvGauSRkgzwys0e
jvYPYzHD9deuRZDO6XF35GIK/x4qB9ZVDMHQShMvSCOMnJPNIRV4VobX0jkf+QWy/RE177TnpdAx
SxobQjjWkeNXEjmT5tnifP3q25zY99PlEz1/tsN3Rj25AwZQdfzAiCQ6fja6rFDfzchClblCVKEE
hIBy7bholktwyUsXcN2esoTRyMFWqnr55SMk+i+Bo/SdgNzlNEAwLHeciOUhhSASzuA/zyO3Uefs
5vBkOeVZv6vq/D0qfXkevKO2wiiMiwTsoWK8d91Y1rYk52Xr15u3TEZsO1xrXZucmUHNWIPbsA8O
cD2/0GXI5Xq7EurcgJE0yeIVcz2m+3KCLF7oGD8fhYVBPyAdSl75iaOm+rQrpNiO05hVWQHtnaVj
N4/1piSeNUPFdi6gu/Bq9RYhz8QoonDqn5MVhbG10PkRuNFchnQhNRqgk5371gUKBFW5MBEBGBTM
F/Va1MaSpnffiPBdGOFk3tDHL86/cpXisBLaiqdkVd3kW0QMj2QMKR2ItjXSPGsu7A17LLWZDMRo
hfOwxl/vgE0MAREWqu6BQaj3JZSasMSPJyEXy06tK7OzKqlsIwUwse6e7Gkscx9xPivOZRss81e3
Rc18hxbGXw+YabdEaY9Xftr5M6xRtMXGzDeCoihru6CT/5QWAyFS4Kz29PuzP2Sle02E9gV1/bLM
KS20ra2RiCPcUGz6qQCfJrGgPs4jhlmm0ssFoX3Oh9wvaYUZ9Hq0RFwNmHv3bn5ewf70oXsuEeVs
G1ThrwupUIubJOz/zppJw/dXutaDxf4vVBgC1lDfTjh4KZiU0Tp8oWAsYEsMnqrvw7YpouW2I33o
v8cUb5deLQcVYXtU1XgmAT+q0FIsS0oDpNeQqQttjbgm5MlyTpTLgL/qkzHmpB1uoNmfTeLLHXI8
4eVUIG65f7851fuesv1A5oApy/cF0DTQrD/9WH1V+aKO1pDtnCRg/ZSjPJ07qRbYkPbCKMxg+WCz
kFE+khYbWw+JWmiN1V8+z7Y7HnTr748t/NMi3NFJZfOHDxiPkVKou1GZsq1dVCSjnIPlzDkKADcL
Mkn0M/g2I27K+YIiGA05f1tr+KaRhIc3mJKwvc7FwEpMiAZmQBQ3btASGuIwgJsv1xkrTq+HpMlV
V7XrFw24GvBAQD0JjhB2tvATe+dPyY+0uC06KukmbYhHis0GuGbbvO8XvV8Mfur2F4k1VeYT80pz
31XFp9f9bnvCJlnErbr8Nw0H6VhfY0lb2DU3rfIA2YiFnLs2kbt8Eej1Q2WoO5BjZZiShMFntO0T
OuHK6G7YKaBCgGuMh1zHsCJd8jZ0l3Gx0M7kMe+6NeZSotMN501EK8GRx6mohHeBMKGH4tYw/way
W2Q2zB0EvpA5D202mPfssRGmrL/oxgUihxlEbC/2GxExJr2cObCMBEiWPI5VVKhH/2lDQ8StRkBF
AfH0dF4J6b8FPM0CFiJ9zxTU8Kuzt8H5h7OODfNn+hq9qFWnj0FXgthniWWyJK5YwZ4j9OIcy4MB
QjoibDXquljMUaqxbEXQuZYM7VRpxdRUSCCTQbrX4k2gpmBhgAMBz+PSBz1A64qwOi2Oy3yUdKJM
CJbRnNQo6zeSpB3T8u8iJx5Ecxb+di2l9UDkSKlL6slpviTB0mvX4XJyI2NmZx4MKpkC7DfGZl3r
DQnphirm0gP3b7Qc+NtDvBc5uxmYgg58f8l4KlZlGJRpN/Z3BRl4kNw2TmgWnhPROPkQoqAauri8
8zOUCeMM0I+SpywwWBPUqMmSAlgo2fIInPcaNZJr71if2CnaoaA7cLzgSeSMxvDg7nVW2TWH52Hl
z5Xu2zoVHplPkcpamgIRg+MoMQZj8jn8hkx6R7Hz8fHu4xLxC894ueqFE3cl2dtm1i1+AKMcTUMr
ykypgnvvbNKsRrjzWxDJbuPuln0+3WjLbR9uQtcOCdOKr/fCkvpJ80Hn0PPVmXu8hC+otoBVc+Rv
btLvT3EDCAF+nXJlsLUesUZWpf8rOCBb7g1OGCJ7Dai/ulz/N64ns/SOt7lcL5kyup3eyQ9dkgRx
hLUzy3YyjDgaMwXaqxujo4qlygF/1Zdoy5lFxy4tSBhXlH8xMWVVjDOrFk3vQ4Ker979n6Qapsvp
pCYpuyvaXfpjVyY47ynSkht6o2HOnUHtsU92CTI9p4HYM2bTBEyRFIovonu1Ok3SkaFkh0ji/AHq
Q5djTmbv/C6Gt3SmtkkPVwifQDTlWwICwJB0oUQJsCYJbIwWpO5C2GSosxlKlpQaUozvJcb/h5vU
vnHeBrG1pDbO97nziWLI0AlxhoBJDUKxPObUV72uTfeQsccXEBJ5SfZf7CJVwz547pOVoWKRmInI
WuBrYbaUvNdiLEF5mvswHIO2CCQwVwlvP24cTvEBKAR6dT9qMS0r0kq0/s8MSU57UnPrT+vKz8GK
4ug54ZV7bUN9p3/0ToKJInk6x8ZK/QPZN8yPaP3JPZWkwBqFxfVz275SIDCJqLl5b4gyTTKSDFwx
Nh05RCJazXN8Vw7SuJKbXCMuw6VVsZY1mICZsqwPKZMfLwrPmNPtQYfRy4tp5W8HrTLhtDXYzZ3k
vkCjnY+yJSyAGey4z6NMOE4iWdw07cI3EGjcDNuXFL9SyP/+aqiqNgmSYZy3O9AAG2jFREahg+sJ
IgHJbybGulHOmba90gJtn9pSMNFvyXt8oOwT+8zwTbsKMv/HyI2jrg6L42tOTN9M9OnbNryJtIqB
6vHbPbuGPhoR8Sys9jqn0XASSzv/u14ofknyXNweOkJje0Ui55yIWWK/+M9MwxU3CL5z19V6Mvrs
+T+wNusJzPA4eAu+znRUNjNNgK3chlUCfmBXQRP240b9GaEVZzPO9EMy90zINIdawj+YUI0i+8M8
yuweNZSaWLYmk7ievr8eTCmtgDwtRKv7kdeiLK7rBaW58BeqEN+2aTtSziOy9UjXyX5XIt39wou9
2Q4zf/VCVmOiiXjBRntqmZqbUuuPhmEWykvHpNbCXWO0jcxJkZ6MD1J83QPJ7spD18FT3KId84Nl
Dr4gpBuAbceAbQCbmEO6p/wjgPkLE2aa6CYHTcKUF95UX8ibCL2Qyf5xqsmhlmjScc9swCyABMbE
rpVZnEQB+xg8qSb2aYFvIStvLczvj9JIuUQCNu0IvPfQkiw13ke+6eg8+IBp1HdujeH7K61JED1h
I9i1gXsc8PyR5LwTdFhdmK9Ci+m+2GE4Jm4SxYICvudshyIRQD42s7JwQEpUaz64sH4iJhqsq2Ez
jYYJPvQYc3v+9/I40jvNZDdwivktqpXm+2SgtG1itvE71ZODFSCa2ezEDjHqgGE1EQbvZC/Ch7Mt
bjccjRz3SgktoDONBTZfUvkC3oNB+yTxFCBhjVqdJ76EBOB6gfDSWHYG1kkJH+8bwkjzGKwUrzp+
FynS5S+VgBvJ8iWvsyZCjoEdi9997M0yaEeQy1EWQ/3ako22ZOryUy4LyXo3J9klgxxs82+Bq1WP
JKa16LQaIPIzQ8mtuP065zAGzuKGBtCMLo79fB8yqnJ8CnBf3yhcxkk17s8v0pKVGLgNBzTPW7Ti
AbW6+n897I+nlJegUsoqtwpE0Z6buxmkSHQyeIFiEZ2Hij3JIDb+58ffvlfAKSD+gvjnasaVf9HQ
/0YIBmnBrnpBNblNMS8VFfpgP8TMFHfc0SJNq18+f8jTbV2IKz1vKFjStjcaybvxWpwC5YhEGdjH
hI60/RUlGW9ttW9TrpP+aKCucT31KlV4tI5K2XRpSkJAyRqh/+nJtOf9VPUGza1HDiKnsN8CwLTq
DehOXam/oqkL5WxA0ATZiCowx5wvPFsdiVs6xgt/y5GAEbfunIVKJXQyD+vGBydw76L8PI6HLDHZ
mWwVVELpZoyRmO5v7ZWwOvqanSq5S1SQ24Png64QxR/EKwOBsy17llmw4PeoqkxJ7xlu2aAb2GCj
ZypzLmgofnZr57LuJEA4iY1r+n6nZqa10n+su95q4gtnd7qjN4JqAyh8qtPSGjsQP5FDfKBMz5Io
r0eTi0FQdSVQ1rcHiD2vUto3ygN3UR7NqNrsizCgvE/z5kwkBjQlw7jBvSKkWKHRwuoBYsRQ7UsR
iL6u1IhvXrQx3dYDaKQFvnLk/VFFQBq8DBkxCRecIuaheJJoF3MoLxRP4eaF79fYtFhe5K6gb0ly
nFodkPmy7HyGY9pDI8OFMi/WG6h36PiOVjgFmL1TY9km9v1IY/cKRf5KqjdD3mwoB4/RFSxZ+dKS
cnXMRDgE2oGVcoi9aB6kYNNgtH9nAC4EooUjq2CE0lKMSflIc5sLwKfcP7PzoTCEt37wmfnLoEaF
LF2A1C2O+UMKoGHSH+ABNZkQ4eKXpYlIrwxU1M9MP3MNNvtKZserzvyHwb4Z1Mo2W6ZqOOTNRs8A
zown7RD/3U2CyBmG3CbR/0HI18XLLUbrQggCtse+FjykIt70GCtT/mdqJFuAPzPk/NVGhzkj4Vje
9f39b6aevkPZkM0HHWumdTGkduN2We1gUqLjOvSkinPc33zVvxq1LDeReP86Ho5HCUd8mViwKROC
iZh0LXk3SdAI9VFG9UeSwoLfY1hKSwmqA0kGd55L0wRfAHERJ+fTeMGS7/yvxbNIYmnPlNwuOnY6
vNaC4pi/Wip+sA0c5Myk7cIyiAlku6QadvxXckHgYytPMTTi1og6JVMg2ghW5sVD/wJHsjwzP0ly
3j1Rqa9dCOAjPdOa5+90/eOmuk66DHNhVbc3iCrRQAt0ZcWwT1nM4pT2PzbTa2MeuMCuXgEZrwgL
qf1nMnJn+7hhpybwjRmJ6Bi6JRYLP/VOJQosRk8E1UBEtMhEZnrp45JJ2EAQeemunSa0fAvT+duk
SNujiHrZ6+b74/MAWMgGgtVlrUaAFPVQCoNrK81EQytWXBTSur+hVsotuJ6XQFj6apUS6FqZY6Zo
kq1L85hP8QzeRTPbAITswmnFf0zgmxCdB4BJQNk6ju0cDDreoiBH71wR+GA9+PqK89MQl/4jDm30
brLA6fzsz5iiQtYb4piVIJvu8qFwK0/KNUFZSm7Mj6Tdar4VFlgaeDMv4tGKXzj8wMEolV8oXgj1
M/9FJLW+yR1SYK1cNbtBmG2VDpXUy0+FVaGzpEtFu9OFdMf6y+UK0Uxppqc96v/Fv0t9PG2XO5Ve
QYmYIobcmr6ARFkAtaaWdRnIV8mWVn7WsEMIJzSbGrnJynuMooGcUhfX8JFMeLowJGUGHzO/mBHi
aye5MZ5Czq4hoGGOmZp3xfROBXdcQuDjXL20P2nGQQ1r4+vCqsQ8mBemaMXkyCkjJIxZle/aY8bw
YG/DpVpHG0R30Irz2y10ARenTjXTJEsJfQKIg3s8ub8ntV/lDJjmMz8N03HTApFujQdpOjA8UchL
in6fCLWoK2k/ZHVirVU/hfixmbKBjP/3zfIqOpNyC6y3qVyzfyHU5EqSn9oyKf7iYhtcdNV1r9P0
aDlTNiEHzMJr3yobq4Up9Ej6GfVeNvvb5Y/tb46B0i6InQvBlafQHAXUFNVcDKINfmiDcOgnSHkq
k8Ro7N9kkL0YVJ6MSY7OnlAr5CctPEqm0/Dlsxio6vUqdiSyTXG+7q+Z6fJ9GQEmu9bWLWc1y4Lu
VnZ29VDPHSDf4Y1lW2YFh78LQgYBguyTwuqErrAHrjvGwRt7eXwTFzicQyZJRQGl+NmnlyYe26lF
6czh1qi2SlU9FtTzKtHWbA8yS74/o26qiX11WriF0XsQzKI1kMw6yE13nj6TBnNG+syzlXuD9AMo
UP/tU4d2oEB6OX/V8pFpPAGTT5tR29ySxOEKEZDm/CbO+/7t0CzHBd626s4UO7zk9Cy8WpkF+HgJ
m1qz8UV14V15N+MQ7M9a5990N2I+JwIVSwljSQWvUOViQubjt8RZr5x5/VYJMSy8yVcSlLF+nqIf
VlFksEPxfqQLPWFVwkryMX4gebqvuPpxVkuvsVnsF6G+VEZblJp6C0XKq9K1qkP/hKrRtm5NTbw7
Y42V2u1Z1zYvBZpMgCDbwP0hst1JwW+uZ56QjDCm5Qf6lIs7esYwXYKppIohzyOMi7iawKNyD4CC
PAL7MsSSJm+pyAYpKyGm92YdTEHIKDj31ALulJi453y+ZS3QFjQ+k+S67Iw3cen2B8x96mneatmX
2wn7yjxZsrTKJkwkKNz6pdBDOWAfd4LHJFS6k7cfu9V+suRCq2iHYsXatEkZvlX3wcD+EJ0K/R0T
NNDKGYDHoC/Epbfzl03J1QcRlatVDgz3DuvygCibhiISMHbQyk2571m+Yj6V/yvL0lD1+orDeb4H
rL2Mj/PpBo6VafyExGaCU6BOTUWHjw2DkRaRTDhvGs3UhP96o9wSAM+ln8BFqN8xUEXRB4AuwKv2
HBrXCIYQ6DnGe8zyCR7fKsxyNlYB/0tn5I/TPoa4GLX0ioYVf4z0nFl1AMted3shu2QEu23tLnxK
IXB5llmdVjOL/+FNyi+wXuEbpqX7Ih4KymYTTkVZy4rfkpqaxHvP3jtwqEnckPLlUaKcZ9nj6FBT
+A5bPpwA6lJ3IgfJgIjYC6RNRF3yFUYaPAW5eG23qJ4SRWzs0XdjVpEPu5Uqg7hYcsSGAgdtcV+A
6ShihZrutgFsMP5YLUX8tOkyCxIAvKbjmh3oET+bhMcdYCHktoG5G4oohGRwv9b5l+CIlWZRExm4
jOnBxM6wePj6drnSNbPnwccwdzT5xSqLgjmq6+s4b0TULU6YxkDlLN5PrnObA+sKamOm+u3J/9L1
02277uIBhXTcRQv1USfjVc3Rlk57alEOKwHQZTklGUqCY64s80QRl2ttmJXXfNcKwt612xlXmzfE
Kp6NfyyAzxGftnX/Wt/DfKwtdBCaZm3jR10ZoXdwVxIGO3Vg/JnIeOBE4kuj5j/xBQfuueXiHifq
r73Wuw6DPu0pi9e9EtiURfO/7i8Y/ApWdDVxI9EJzJ5TFopN31MTdQ124Yu/m4bFVaI4XD62+4rO
XXFBFzQBpLm/L5G9ZlPqKUfyI9cT+pqhSSn1vuwtocrz8YBkDvpcDroxLbLCsJ9fMM5deOhLcG4g
YG2WuFDXdTxqVZCBjHvssNtbHWrATLi976j4pRG198zH0ZN2PqynHGOejix3Cc7N+Y37WnXYjIiS
jMELtGTi+BpZjb578Krg0MuE9kcpwyDBZ/tyWREaLalzMp0iFQJhaI3AaIJexlcNRri/dK51UkBJ
1ZLfw0BXlPKShHx2I1FpejrsE4oGFWxJQHbeDjtHP5l8u3Kha146b5e51yPj54aYXPSuPnJqMmGW
ufanTufJFFwsYqA2NfFngJUozot7TQOg9qasN+nIpAoESITNx0V9gue/5Q6haCt4KL7v9W8s9gZ6
MCtQdh5YeRzFtzY2RbCGplXDpnEROvbgdHHWOMDY6JA9y7vb2aYmQf5TwIJJ36VA1mpkT+rq5jRk
9+hpvgqt2vR/TIjoxYjcS5Dzwbuvn8H8xc1PM/looHZtmk1tk09uMVlMGyG2/zc1IWG09t4qK1NT
NpZUuEmjYR83GXpdVKTfPbUm+sYXiN+6OUtIGOi9m2H0vUNeUuFfA3jfYW2bFVlzh9IyT71fdrNn
g36uHP5qv6i4PlvJtgH4F9hSesFiZ0iq+jhrmqT+LsfRLCXBHSxo5vc0r4mo4fMEm2iwg/786+hg
kd7G58CoMRIOAYpg4mU61L1yar+wU72xRBSCAa0izDaAejxH241AB/1KDICU+tK7yqP6OFSnPQ5l
Lbl54SpXy7sm7tvogc6fKDklf88j0CGOC5I57SxE6lDIHwxB/HB4D/HHZTapP5wk/s7TJD0HKaYP
Kee/8X3LPbeZnewxr8pE5q/+yi8BsyAVTQoYo5PTpWu45zU5RAYazacPj1Y8BdX30aWby1iNJlJG
vwQEHar95q3l2lbo+W9oHgHkZ2dCOWRATlQtWPHEDrRoYzSoatOuO87CFBT739mjjyaNMdf9hhTg
ikDp8aMNmLzVOSh8yF31zStNwfxDWsaokix+puyXbCeNRbYk52YXVYnzmpT8/Yvb7SzlHapYMBwz
sjbtHqfVRxxZqzavcew5wSGoqBPDHKFu366c/AJsgNitI2BrSdo2r+ilzRMsWi8hEsdvx7VYjjC+
qoIWosBNW2jiWoRLWPR76NWv5FAi4r+nHiSNbDWhJChlkYQT/0vBsRWmJWTPlaTzcR5KDea4hT/G
uemK1I6YFwGhdEuu6hNDsgzeyaJqmOjmShuxTQY0igIidLYT+NN0P3/8aRTJo5AksVaqoWmLmz58
FXR1SQYyr2boj5GPzdL0kPlg8imDcsoaKLiopbwlR6Tkz1Ox0OpPWkVhtQizYCQGD4oAGHOK4DaR
7nmmspDzpg3NeutME3ENokctrBaWXdY3NN5RXBHCWRkhLK0r7i3UWIR8C5yzlHBVBYyeY3rV+AnK
RtLJyvjMNZcqq4fh8lcwnAzqXT7w0s+2CJ/pxTJ1glU0fIJud3DrOgVofM6JobrVm9grxBdQNFUP
JRUBr+Nki1GS7aPsOZ2G07nxrnn3bTopXlwrFczueX3w57aBZEWczuZIBdX540ecU86a31MY8h3/
2lWdXUfWvMqx8RMS6xXGFSE4zQ09kH2iNKJU5e8vsP+4/cG2ky35wzWju/2EZM7w7cQkwOY/F/Zx
AjEWeDYSz+RD15WyNkbv8YtnTRgVHwwaP6CwJK0qkLJdpMSU5eWQN183TtkOJ6cq/pmQXUf0UDpw
yC9Ue7WmJ6VM9vNVUPsApm2o6zN5XgbBLqgiBku1wzIBZw6xKTH4o8U3O+3RctBKumxTKzmLw45C
0Hg3bHoHNSPLpEwb/CV54SMHJvrSAA5Lmm7dHNhy9YFDJRD1YxL7qmthPtJuH0E8zgUULM87Tdyi
iAzhFsAne751QlrVKuAXvIpsdKpgQnrxE7aD9zWr/nudb/ANS3XFLWfKqZsgRJ18eA6S21/GET+u
OU+ueviFPtCCrPXQZKkMsodrmUKHmmiL0oOji75+y7yJXTT5NPp2Z/gq6ms0WqJe9pD8lgMEq/Pj
VwCFmJgNpXjRg+pzNYUFidS3Y4YsmW5Uq1FjSXGLZr7IxDht1CHJagYfOO5v4fis1WPbnyY/R9mO
Bs+89xInpYOfWJvXKUI93iEqXrN3HEKMfU8rY35UrTPJTnQ2vYnXMlzxEC/bTqQder7sdhuz+gNh
M9j4HnCMiqS+qzwCZfGFPnDWCVJsgj8gCvn/rTsxrkCTr1rtKfugEZwAPZsrKKOcOD38Oya9lDgW
ilUgNdo7azV3JWaHV2+FJdaWHelNisQS8JH4gV/2odkgkPchXVYUPUd56nEHtU4D3aF4Z0akPgMA
UE8pRfPnloXsmaSmucbQ7O7/dVHMhfCbkfoq6tDM7yDCxc6vnrlkhrVgfNi1cW75ZWObgef2bF/C
FViKkfVS4gD5Pq+XS5GPTQiwyy4MKFzMONvhsNgd3bpQuGDh5XVVEY9YX2uo4Z+62SQIxrr9daTN
lc+kGPqMQUWc2/A4vXNkl+xdS6RE7+RxeCDIsiGEFuC/rTCCFPcjbbuAPYLY9+KeiIDP2qTTrMhH
tZ1NYPOOOy0fN/Ebl3QJki1GSMgNZLRNZY9cegXNT/Vrg2J+Dt0o6fx86tJ6XBWGcXdrd5HujHTx
OkMMrz17iKhFzGycfAAMHoGXW6+TICIoH4/MuuJM+l2wnjZnty4Hh9PGfGcn5EPW/TD/O4RmsFbk
bREKfh3QFB2bReicgtp4eMHeNmrjDIRTv9GVZIoRBo5z1uEbuBOeVPkheDZcnrs5JHK/MeThC5pX
Do5QNsttR9v+k2iUtoOCEqGUW0UKMISGMj0d5BoY3xNDP7Mw0LqxfHzm/WpdxnUfpmGbGCX2GcsL
urz5DwdDyCPOTTxUUucnRcEaqdFLC+IZr3S/P+yCPwEjKF/OSoy/WJFWPCSyMTttTXx2P0aI+pxC
ApYwep0Xt7Xe5uIMRi4IECmHi3a4xd3diMB2fymcyuykNoiEf/tFILLcpZlhKs8/kyxHwsQD8mjL
DhY8eaPHsgaJZjfZuehTALNNfGG9dsoodgC2ssW1kj8/kpL6xVWOwy+QdEdaPG+lWi3ZG9fs1JOG
vKeJgPK8nHyAb3fL1/SKmnzzWA2ycCsKwTNKWkkLf18Px4CCoZ47dU7C6zgYIhmO8lVZW6RVF76h
wuJH5sliTFCnbZy/j04yiwSjXszmZWWjcN8f2G/aoAFHqBT7DVy3V+K40vc/eoJiWxO7bEoA2ipK
NpopgaOrodBF313VJsPxe3z3DKzMR8MR59vvjlazoiQwYmJ1zCARQ8E/6XHZjE3UZz9QB1yUXNLS
bxn+lj/SusHE8zJ4NeSOha1iA65Mnx+dMQybxD8c12hoCSYHtmhWl1D9g3JsPTnWP3kFa1L8GneF
k6K3doFwS0NnRq/QehsRjxRd/e6sNfokjtGdSPNCR4kcFGVl7iVxBus+UNlgt5kcWdCC1WVDJYpV
u5QtyCFhlziRGyYoizRpDj3xpBEArzxkmXkpYMl+MXn3Rdsao0F8r0Be9glrUMxOvfiW9e6JqxzA
m8Qvp2Vu+Ar3ucDo5mC4VHUGb3M5wmDu9qvYV/PULTY6JYPyNqLrbbLlGd8kRjbiUzSIrzq3+G/D
sbLNjWmF/RbDo5LNx0Xf5JuWDoiTZlCJ062uDM1Vfn0fqZupv6pGir3i6jmBiVXPkAp9LJdnd6Ry
oPqrSpyTzH3Wz1elrxzxgMz2dlSkEPuPuhFXrbmxyfO0t5lrF+yUpBebKAqMaNrY67V0O/8e3ayA
++WjqRynPWbBeyEddZQqAx/Flhz/3dtI9RMxEoOKwLpm80GlGAhAaRson5WrGnOs5MfXWBjG+cUH
554ezKS4g4bnJTBnq/52uNydev+FaU1PzIpIWCcP2ZZNj1qiDNKgjSVGAjsk1EBg4IQHGL+PgbCf
Aknizd7SpMhrOtQf03I502Uj21ClsdlOt8mtHkJW+0+DCGV6mLHysDKMbqFzIjIIQsoNuDy3aRW2
LheUYIiISo2qw1KBP+jGNUaMhgFsyDBoEs3Lx+56MYt8P1Y0S3J4S/s8dH8utSRa98Qyt7Uz0EUR
5yqmj7L4Fb2+tCGNdmxJ7WWm0clc0LPUx7aMlQuWcRXlS3YuWEvO9GHPmd2S8X5pTGhmNsuOz54s
IF1KJ5AAMMGVh6jiNPrz8NxZxICUQfguMqjbaFly1NBcmD+h1iOQCS3Y31ojnc7aKVtAXJbK+uLY
HVLUcerhNOHOI0bG4rGquodcCAP12xO+pRoatT5bgCA1/QGbqgkWtQdBv4gv2UrsGOVmF0Xcl1sB
TOym/Z5p+6LoyJaRgPhA/lZv2RvIwsiAbKoGeQ+NFVpdcceEkx5WbXVgcPwNCxtydOaG/cKmFsCZ
yCIVTImcx3A68E6jyOLND5cKRGALfQDc6m8+EWEsrE8QXfxcbKUQjCqiWCBpkHEsoJGoNHDEm9vQ
xnNNs5iq5Gd3rnaDeghoCXVJSSha+Extd8Nmw5arIgV1KVNwonfFzhAsKbrR6XANFtIzP30a2AYy
IAaAhryoLNrZ0wmhnsXzeyBZwcECSX45ODe9zFXE2ozQrtZEZajBkCEQKquzsFaWVoPOcP4abDeX
v9e3tL+vmruNw1kdwc/iX23Zx3VHE8vfdjkpeiAUgwO9izYj3mVn7lVYqMBK0V7YORQha4j/+az6
xxU+0PA+329RwQzxVHcFWLibYFKCssEMp2Xmkfe/2qauAxq2enrDYfRagQbtTERk2dgUYOiWtzgU
mjTbQui3s3Q+48P5QyR3bMuaZTeEOwobLLDEsd/AkCFp+FSxijgXBnM0fFfN/yVxz1Tu0qrqa2N6
DGn9moyOMSZ4S/vvi7nFG1LWtTynbHUnAy458cUm89jZq0kX6gvvGwIDmBTZ1kQQP/htWNI/90Za
Ee18acgICGOp/8GblPOD9k/WK+HopRJXqfz312SWdfuK2V5jH9/zjRKfFhD9mHyrfxbKLglGEUYM
Hhz17YdnP0L0opObuAlr78vUC7vcuD3LirhZLIU7oeYrGgNpshxIVWqAi24v5HKBi0nnmOx2TTxg
3wVceBeEwRZ+KkmQY4Kv7uq7itPPy8z5MMSXN8ZKUbZBoIrS8IfH15h+0hKkzX+lxX8ifwdOsJcy
Ja8QYaivg6cYFNlnqxCMJfuZ0UTDEbiDJn2kT2NpSbm7hQmIE1rKsKzw3PXVN/90AhG4sQ/fq81v
sEE3iGo7GY05Dp7VGT2683glyF9LqnLEQViUX0KkkmIZoB+u8hhIHGQcZneTyMNSNYRhxkHs7x+o
O/Vkw4zXdzgOduuNroVVfu3X53ItC+fp2cZnExoVAdpT2DNH960GtbxwaeM2lIbQ8iE1ey2plPXh
P2mG/gODCjpk2QnAfGBoYvzGMm+rGrLp/GfmqQXUomo1NcdQ9rNw2yEDAd/wcD2+LLgJ/0YbjNc0
H5LobweGh5cAMax8GTFDg05EofXt0eDi+tt69qVkSkEQGVyNJNBjHU9LIDO5vWzwg4hfRBHLVtal
P2nF1X8Yh82d4aGfnAY9DcBFY/f4lYoMioO/KJ87c5mkbxNIrD+cf83TC3zZ1q7wE8ur+LLWMfL9
aBMy6ju3J6TXARwiJR4615+r8FhZuGnVhlqgE2niegGgJxkW2Yc/Zd+EM3Gz6RTnttUUoFYUvfg3
idkcfGtgcNGKu2iZ2cVV4FYs0nCq6tilczi6uYMn5vL3W7nrR6cX0QpiRLojpZIhUg3gqiNqANLs
+Uk8HAb0gsPTfCRSgTvHCKVqesBeQ48fThcO2LRgGXuFY7ZqFh/7VM1B030PqxYGq2WZBn0EjLtH
EZL9epjlknVUN8sMJezLHWvvl5ruyCS7gDPMjGghdl8o5z8JxXfAi5xjfOO69Fe6OZeEQQRhZX+S
YOCdcHEu+vLGJDVIoDq8W8HldrEK1KSvJwxh004n+8ns48nQ+iRv+MewULCuHVwukX3mvV8fhHjc
tBv79k8TKvcZ73LtRA7rzlaBbEZC39vdoRAOlbCWdTZb25jwPcJv2SxI+PbVFpZLZpqQ1v4oicsj
TE2z9YUh3xuKnTk/UCN4usSSlOWu8IC6zGbJyXpIq6PURBjgRh/yP2SQOsikaV7bwTI6tGCHyg8Z
9MExVM++tm4dQlvAWZ5sIgPBNBzP1bsyHSaFHN/E4YAx/UNk7BI2GgBynHOcPOnEB/tf8sgGQBSm
0Q/crDhMJQKZb+54RUMN108+Hhca5ME1tUaf6biJSCh29z2puFcrNrgpp7dE/vGI9CXXJM3l+KHs
B4nHk3Yz8TUQfi6BjQ+E5d+Uzkt+nukuB4c2bV0lrJmecwQ5XJBCucX6BfVeKlBQjiHsFyNfiaE7
tWDsBoBAF65cKbb7n8J8RLBHhkPUkO6HOYxM9rRmFgaqSAMsgQrfzb5Z9UYguvSOs/ZcNzVNhraN
e1emjLUqfbj/t/CLvEa8psSkuAPL6dIZLvCSrMEW1K+FVhBc+m6tWkXk8BTVOe4f8g/8HZ3aBBQ6
2HldqfmzTvcsnhSoaEWqE4mlwCmME3CbyHf+OzUSrXJUl1oB3/2iPcTGy7frABLadYeWZVrsMxD6
FWB/GBhjeb91OjO/yH9nI/AqEdYwCs03VV8nc6w2HkhM+gYLwD6o0Np60HvVZ8wyVZ7FwRrMVuDT
h4k5Uirt9WjPcd254AokFeg+jP6tYeI3O3r6tCR5Hp7JVFp3HTqfOZ8nvlwp/vBNnXizxpEss6Nf
NXZAAjt1A3ToMccpvcuaWB9ox6ZQYQfhA+0rxXvXKvyf1m+uA+jbRPRy3Bl/RPfSPDRobFqlAGwC
gQI+P1MMFrBjOXQl6bxv7RaZ1aTLoE3aOHoqZ8YsA52l6+fwwNx67MfvNHFONwrCPaMFJ1iWCZht
cCbFjEU3ducPnRdlW19JxqdcBqBLnIXxaiA2jeoehihCSB4T6Bs2lGvKcI3R3ekNBiiBQ9nt9CcL
yAYWKhBr5hz+9Cgg4wwH5w/grNBy5C7ZorsMSc8TlXawyjJNr0D18UkzSlOCYzVIwxHKP9F9WCJ8
B78jlyqs8hx8feQ6R3wIhJltiIN9++eu6Jx5AXop/0uFSdHLEXkx4YIcq0LcixID7zblisr9GUYm
MKoRL4ZnWD2zW+D7SGhTeE6xYNeOUTGJ26UUw01eW6KNSQEUBdHKSzePpW7gK8hXSLP8R1Mc5oWk
HvWC/cfJkHodrxRmfbnL3Qr/KssXh9H5ejzyNjgWiA9KxDP27atzF68Iuq6KVQMzkYUbrrlo0K4Y
JhYeCTlsnKnIpBIIP+/IFaNL594EMTRdmeIqXT9YaoLYpWvMxIYS0AIimQuVDdgwy+L6zpUvvYwC
hLutIgFDY6O9Rt2OgtJ+seJ6P9RzqQ05ABbpgkKOS6WglemuMzfGF1QILSWlhqiRauOuyPJcWCTy
tZ8DZ/L7VdV0BnNYn8BqZF1YspsJHeHUED84DW3L8EjVfDN94E+xV9T+ZeCyEv5cxkI2hE1C2Qke
ma30r++V/D/L60IHs9JkG6NYs+NuELEFtm7gk3pOYoyaGAyUbbbG/btsbbx+q6WO7qNYPzRQdzeS
/1TCgfCDeV97iHfvIt1cXqs2xTmhe1aP8VEHF4PHE5uWtls4Lms5WunwWQBYI/4dw7yBoa9Q1X5n
h5cHJD45XXpjnad7kzCu94zDVxFyx+YnY3HvCXxwTcOnmXO8216vn1chca10cVCjON1fx3WMbQqx
m1DZto54pswwszZRjIBqIGAhTQIhsudzgsOxDVPGcYPB4oZXBCRTo8GZohCtZPd9O8/4e2YooT6m
h0Tlo8/jjXCJAGyXzYLCT5EDfCt+ob7ds8lRjo0I8Vka8HN28FgnIiEphEinCVe2MUNhpyrARown
GE5hGlStMNP3GvDr6s1FndmQRtoSb+tMhdqfT8+215fcY+sTVSR26/z6cl6S+5nzbFbZDAlKFH8A
QdSCw7p1K6RJ0FdWnLGMR95CA+WuOnK47qXq78KCZ2uzsFyINrGJlVyJTVyFHpxxbWEsDuIWrQdD
iraLWD+8gcqQ5HDoLPUisb4+QKJ2FYzX0OuU3jbeHRzNTI5+nRx4jL+LrJO35BHvlTUwt3NKOnvX
39p/ZUUDr69j1Nj9zq0jEwUx+Iwj/NNIdSpFwpnEmwf3tRNANGZvn6+BdlDO3plyZ8CVNoJVMNAr
VdciMrHh0gBQbQF4mZrzzE/Yg3QH1wRgflOHYqP55aVcT8YlVFEg2DBfoiWgVaflK7I4qkmUtHGj
xoyTxsuxReMqnRcmdxx13FI63qEvPbUSKE+XHJmJiBYAXnyUp1nH4zNvQELyyyArWo+eRbj9/VJT
c4liSY6TwR1J4mkQWwEh046cx9/q01LcWcPn9n1qEHRvnbTutZmF3C3Lys1WfN6q6yo8OXo974y7
3Yr2/lhNbVWS4nbfCdeZ6hbLtrh3hO0//S5Rmvs8kQgxwTUE6D5oRKfIoINKzBGyJDcGVlOKhZOT
5I5ImT89emkswr6699hroecZHi+qLWPJtZj2Om530V48GTgEEO3LxqwgXnKwJiW/o0XgKgp7xfqU
Y/AxNShhPfC+wdZXSSuqgv18C1celM9yH3dPFQ3eFb+xmnPFednv5sf1lyfgWU8OYH8PDmx0kJj4
DrcarG/cjimKOr3o6DTNowKAEmsYSPDWv+WkCNsQJUf/6qAApj1eR9vTcuVai1TE0efy/0kcdsRk
h4VQscb60FcygGF/Y4qinDBfwTReEbkpCv1aaKKRoIKhDq03kyvSngKVlV7vlpTG38IlWp87z6/I
HFn8zq74K0+YmElgvS0D/w9XdVwFilNFRGM6hriA0FoMa2sqN+hd7/XlEd+lLrgUj5gCy+t0NNlw
8L3T+jRVaEOnvOdLL8dd1TBnyrYaES+OoL4QXJcKvb/+bZkyI3IJnfHo8v0rK+2qEe5IXF5eVQmh
tZKPwZFxNyoke4L+30Nt10sXuRj3q82JLYQQRVIXEWQJBk37LQiG5YBYDp3ZApFpEBd2eXpVMb0J
h8pc8nRtym9bc0kOqh2ib4KXj3o/KS7ZvyfMoGXm7b18qAxonCYlicBc2i1uVDlqtNM4TKUeOnTG
eWlR/5oJ3HBolPIGHT84bTfbbsuCJkamzau7IkArDl/5Liv8VTIX7yA9EPJJAfKNSNbzBvibEfCU
UwovE13/y1xb6/B0z+yjcO513krP/JUu12kPKpfuimhToUmV0b8xjikuglzldDtuLehNa86EcGUD
XlxLVxqvjINBojA8LAT/LrBeuTRkf8x8ScAw8nIRHW6/IrMk71kNWCg463YAY4fwrnoppJHbqvuH
zNqEv1PXn1TZDdS5v5bA8qqt7vA3OxiqGewWZ+uXAMiswwrKJYswyMOZ8eigiQeRSCOkvtM5ZY8X
wR0no14uefDK/LfkSf28ECpwgBTQluO1pPDN1Oj4atjRHHfVwbtrkTvgTOj4FDTewdzMma4eEMt5
zX49kNE8whtigwXe/74ROhUo+SQZ0wR975HV8GnA7EZBZXlyeKPWN0DoQudRrS8CVfb759y1bkkL
8HK8VUCH4bbysuK0w3US4kW5/AQpIZ+I7Y0YtKRdAvFaZSxWLQlmXCkJApj2Ga56ruoyTYFoZREv
rr77Mmpr2vPEM8pbhD8ZMBX9xJ+wIPHZc2cNRrG8S0DeomimP408A7BrK6/Suaoc/gUjAUGHGLaU
LPLsR5X0iJ6FiDbT9nl6WV3tOn2dL0APYXdCzSZq9vWcGXg+CNpgV36OUeB0gsVGS3uzsLvFQ+93
n8iXMXS2ERjzI9dHDhOCBJrFCm36rGAGTKwoXJ72h03ixgS2Nox2xyVXzN2VEPuR2swIhC5pJLj5
rmRvxM6STBC7VNMAiXE7XA8qOZK4tDQtI4l7vRR/olRbqYYXklmyea64xm2/53I+XNFcq07E5F+Q
riNh7um8cM5UzrvoYY3r5PV+sEEKkaAZqm8Za7StcgY3GJMoENxi0ajc/HHMtQzsnkO8qoKDAFWd
NFBwO54uP0LehzllVDUEMOAmM+BS47i5hbCtFcu3yV3jaY1uE17f3wq4BlgmEDWuMQKKAOEZHTMv
BJv8jNoz1Qzjeb4BVW7eARCyoavXZuFpOTvnPtMTrP8rX0CS8S20SqJOutjLDLurHyp2NJMehRsn
XZuAaeBJrPhpBkX+I5ESP5q08dcnhxR7qviKtDthuZxYTjYi05d7Gf0HIWTMtP35G0GnBYzd8kke
4+55RkALxBYIs8HoQruAofsnKNMS/oNKQsTAkTZ3GR4aOo6jXtZeDsj4pGXRPUsACcT8NyZ4o7Cb
3bZNPxIuWS3VC5MdvyYgDBdIw5oFBAl42mVyj937730gMlAnp1566WROC7SQB7wYJNDlDlhODnoP
a4cPTEEtzci2H+FVDYLwatga6Vd0FcgJi6ubUZH7EcETEpkKx9ErDTP0RGKZFTPBKNW30KZ0Qzgd
19am9lF5JyxIRGPKXy+tlMjb2h6o/0OjJuVdtCZY5WdTqN+lNsV+7o+QqfMuCudZd3VfbQAgt/iy
iW+iyi/0MjOhp9vHrNQAE6gIYQUKMRg1d/2Ma2Mlz81x+ue/tsuX0RD04ybERE/ZNgIaRhCnw4eg
8ZfgHmpUKro1pxzf5HyyC4koy/1IqCsxJIYeGIjpVWVUikGOfpdyshAxfUTOe8zkWp1Mc655p1wD
sPt1LQ3i6WdhDjancQXiqTce11T28LpapQrYLHodQ6uKQpWmcAk71Dtj6sp12FWioCOp7CYtF+MD
FTQIlobXRwqEwnSOLVZNGnMVB5VGqG1tGyAEasgf7WcXETNGv681xKK3Tn8D1J3ogYsZpjCXSK+C
QpU0M1sAcSPHfNYM3dEzh4Io69yle4W+pr3aNA4dhSizP1q0xRaSi7NI7Rfch8sd7e04S57rCxcK
TjPy54aNHGsyYUcao0qE5fvgi98jvylcHP58KHIAKQ945yRYrqR12PRruUpPyT6c6tVmm/oc8aoO
R1yymySOGS9IbHYe5Xn3SOr/hZ2woQuLLvBr+dl9aXinV1uJSPOF241G9k6h+5E8WKOrmzz2P34c
Ch3Zd3mbqvhWPHmj4pbFHxxmJSIoeFZ85W8KfmSFDG957H8adKt32HWw2rXNJvyqmeyQyN0FR/s1
AceC3/ImB6u3sNjzFHhxcgHoH5miWv+WN+v8esBS2M0JYWFUDNmGd5JwkZ0XGTRlsTpoO9MRi2I9
fO8vFF7wxA5C/iBddM9hnHCL9+eyAqR3lkXZSzRgpJImL5gK/p4yUFVLxdWGU81VaA5mDbJfBosZ
v33hoYLJ24hPLhSKfXNplojA5FN8+dpmar0oiPQNqmb1dv+GffcreC9JwstdzDsKmj99a42Mbg+e
wmDqNMMlEVHsGdEZtO58tpoUBwND1JXLNjBaaKDlaMTSuuZqArielzEdSsEWhwlkz3bBArYBN4/8
Qx5Y04SZSc5iDSAgwbC6t2xf3KXMMol4KRFrBi/qh90JiQmb79XpyD3n6gvZZwrjeCa+igGn6zp4
jt113yl1HUN7UV9jjjgVUZpncWcRo1l/LSwyzft2Kya/fc+OuQ1dLkyAAkVUUg3z3b/Ol/abCsRX
uZgK3SIjn8W3z650B377CNIrkvOEjD93CwuJTZFLTult3HwTykr1/NNdpkIbMIHKqjSeGMqz6xPl
BcZ7S0Wk/HrHq8V9yqAczyGEF+mlGdDpxc2Zmw3YwU9coiH09aMfHdWgAZJFoWcs45fYBRxoXxn8
YsECFBSoDrFm0fWtLAyQBz0bz8fRa2gSL727acOesfpt0syP02ebCIEy5N/7+BArWSEyv3xCG0nD
N+4BNXeWifes/bsdZ8mS0lJmnF7sN+EYw6LP6GesPv1JaDnjnTalqCQYDMpg3b/bH3e1hAeivH1Q
JSeoxQOpawqD1qvuQ+CU0f3RNX9eOrgz44fBosKxrWbscH3SIzbswZvWudSp8zwL9RBbuv1dKP+i
A2+Ds4jK+PqC0AVNlJalQf7Nqd5Axn3Zcjhr9h6MdDRnVFpbzi3kmoHrSWzPtYFaL+CuXia9+mgj
vUAmi149dtxuA2V1nGy3CCYnqaMEmguusDZDcp09aFvE7sslZ9FQcpjeicgPHex9LzVN8PeeO0FC
G2yyc5GwLhdeh6rTEk0xayDuHks2KQDbmiMmJXhr7gocAfJ7fXlkDaiW70JSNSE6yGosy22s5dhO
lXrbbXDqN43pNa5g/kAKGq5p2CzwCGwkGN8qwgAo1Z09946j8U4yA+1YyVc3rTYqNis1gHG0jqjb
ia68VcNw3m6SE3lDyODzWA+CSGCiEdCZ1WFe0MAtg9hYH+ldYEbpuPTsQsEQP0zVDOBXmn2Sk+Ph
O7jziIungjeHG+cNmUuhy7WUfmrotx0X0MlQKQfWMcvWJH/1iAq8pQi5lbsGST1//qw1RAdBoxe+
L8VIck/tRQWc7xN5un84BZ0Bv6+cxSA9WkbZfzOB+zdeF4rxjuswdxBGpEk09pFEtHA/mTZgsGa9
apy0DaBVzcotUTiao/7yKVg7sIMmVRBxnbmY07m8qUWK3gL879u/uuJurZOMVZNfvH7mFbZypWYS
7YF2aQRxZ2foYYkRXcFKvqbh5NeC4G2y6dneDlrF6cDuEQNEWakD+4XlqNjItFRgKbnBF/kwRf+G
uta2eUctVFV/Rkd1ucvTRW7btDLS0H7UBcpaZsx0oa9c7fOy9hwN9kMg354dusEsx4V5LbaZgal5
na7aooZpY5bBQGwU0XmA1xsuzWXDe0oETbZmv5mKn+1bRmc9Cr6VtHnJ7pZ32vooTlkprWCEQOxd
LZ/3ucSCrDX9Skan6GUvPgUhjd7eNjPSWxWH34sQ6boe57JbI7n1IdFKpBZgXjqFnbFPVbWizlpg
2xbxTLNGUe0nt9hQ2k2hX8lvrZo8GBhdFF14SR2N7eiuS0NEB8qteiv0iXySdPq7M0XHOZmrWa25
2RojZnfAj9rDrZXLUV2NqxwgmFs23lIZRcKhHAlEq2UIjpMC43etVDnhE8HZnVuwk9mjB6SDalSH
9oYPvN03pckv0KgyRbI3+0fO/hEZKmjnOSws/GBBN7e/Y3sp2w49vJxQRZVuGEZQdYVeCx1LL/00
B4HfHtOgz0CocsEQpyJ/odeX9ARs02xoeWysoXo7aPRrArEj0idN1YA8IGu7GyShuTY+RPxt59EO
BwmM0awLrsoR64K4es1i39Z3XdwYZEWpqRb+Ey0kqzaaAWM5oxJwuiNHfk6xhjBEwhrUSU2hzDSn
MZj1OJsPP6FuMa4nqIbLv4ZBy/aA9VG9dtFJwaObYkquv6/qV8+YNae7c5cv5kZwHTEpHTdjRAPR
PNn0db1RvMG0qTCVW4vBWMkU67EBcaSjzF6fdX1U/acLEKN4FgZzgjkuQjaUWHwcNB4VQXRAdJ0R
Aj56nOembWuWZuElv1gOgn6vof0uHnDKuoBauL3sk1gx+KZ6JXHY5zD64FYJxrZzPRkFSIn337ul
B/q8ovp+HZxXRr2paghvCBkwAvL6cXpxVD+JIo4R8+6xSPh7MIY3AwkAx2r1zAo/Buwf9+QgEika
i1tpNQtDmvX8zfXE+nHivXdcYA+syAoNk8N5o6c9PYj1XNhXcxe0QOGarwT/u60tvopd/YQKa2mU
ow36WaNbKPN+knxRCxKCybpSbbYrSU0TQIwanyoHqQaORFr3McRgeV1Tc3WJgtG5BP0prCtTCGeD
d5lZuQwixKIdUi8Vt99Nyw3SnBSW88gi7JypV06nA5YyzZwiBTzb/OXcTprR93WOE6KMxVuhEzk+
RJ0V4Lt/Vjb/IfrQybXEpU/k3RJfdPJ8Zg9eR1MLun99wCieJkirPT1SrMR62xceP3bUNvf5ywGt
EhPfYj6XA31sPFrk3D+5wAsPL8r9HSqX+HBkkSSqlZnjURhyJAmQ9GXXclY3Y6rLxXQQ8K5cX3SA
Elj4k7sWInM8GaZlWAfqISc8Bf5McO1v3za/0VBuswGQBbLmCKROqI4vA6qp/KI4QF7h1Do9VPnI
YraFDLFcV9GpK+jwgOOVUthH2o4Vha5gSS1iODncc2HvFM8Af4VYGUCKSPUilFLwDbtqu+1/tLil
wcPmzy1V8FzMfShrIavIb1bgQV3QX+ckLkoQ8T19ksr6WJmRswCsTbdRUdjvkND3gbGSfPDPuXpu
1GWGJV8ud2m1tc8fm96bGKUUxhDJl37N3Abk/kLDGc0xTBUaqbTFLVxTNHVLbQB07igRDZRaOmfs
iKCU6og6krvMP0utsBxFYQw9RDKV3m5qMPFNNk5o+m/HAUW8dOZhIoFsIPozN1A8LDP6wT/hjXuC
Uxgs/vlSdW/E8dGbkfUh1Z6wYJokXqcj5d5uxGx3boHHU6o47Y16St/iUr5G3vzJd5yAS5qgi9CT
7bVS9rKKo5s+knt4Lzq/1eRs7cK01UkVdHvq58XHWRMoFfMQzwEh1Kchb1IA0lWqTMA05+Ff6RSU
Y8GmsRdyttrgqKw8NvYJyLfBs3q1cq+IRbQgddrmJ/fgNPfjDdi5Kw6ZqSapdVKWhhXe9POOjtsB
3GFr4NRCqrF69MPOMKCKfDikxbAt57E+namp2z/7+KhldulLHo9qp+MDKUNrrFIfNfREPAylUZ6y
jOyXJZJQlPOJJoTZUpbwo8GgdAKER+zQOiF7pmWmc1MpDJC1/p3JpE3SAqbT32NutCG2vu93SgV5
U09+kwRl2QG2yNT8HBowrna+6scmInttexn6srSG0QoAjTnXyblQDeL2fOlBlp4sTVC5Vw+9k3Vy
IqLdOpTqko14WtpufbBqCmGHfYg4QQTjxVy8vQCD9oOCYMnMAiTuHiQTFO4YqH/dJ7gI82OhWc41
WuPBeYVaek1fY5ErV+V58kEbXVulTwQ9lveF5kwoMOs+Pidwz+re0NlctL5mdfqZ9XOcx2iD5kg3
MJapX8iG8pAW2WOkZwbpl3TgHAVx59lzvJVuOWrivooLo9784g2V7mfU5bJ+slbAzMwscZzT55s0
ElMvCmUii2OFjYrkqxL70Xq95cKb/fygSkoyaSefpYDp5QlTjgacdMbpnGN1dJ2vZqhS2hpsuttB
T9uZMTR1pOQPFeUInsfSL+yF3C8snobHyT6RyfE6SDWmeZSrVIo1V4Ev7WTLHWE39kxFSdLgNG8O
Aq+lvTJ797PjaaFVKA6dYB/EF/K+EbjDAVgjDs09Uzn/I43sAY0p9N+D4EoS4RqN8ulkGiVlGhpU
Vko36v886HE8hWy9cQlVmtp+qlmXsCmBgzVYYvQUjq7qUJipyfTBDMraJJTcyrW12x8E9T04GL4s
OJwX7B3LAL10cR+pPbRDy8OK+/bnUabmeUuFVv4xBJG62prdKaaQGvDKA6ajFkE0ahBqfM8cDfGq
y33FxoGNCpEn/4W+sMrI5JUiReOls30EsyLwk5bbV9l2ZFfyoke/gxtHrMosBF4uJSzyhewxnS/r
GG6PRkm+Feg7xLxrI3zBzMOSz6thWIqYfoVAxixUuZyWwqo7vjL2oxranVXEZeB5GFujSkpRdsnE
nNuV3bJJgbBEq009pSBlSWm3IVw9dK4SM4rX+f7fOoi72zbKc/hgv0CxLznJrrkQHusef4cWd1D2
1rWEgIPO+jQfIg0vk5yp/i2fdNrZumfxZpM5at91Wrneur3A+8QKmAO//GS7b+Ui7HwRVcMzHD1p
UIKc92PooCW1heiYMDgkVznx4dbpYxGW6sqY3rT84Bc/rgF7HRMS9267Ne5Xr60hnkYCtg65k8KC
uEiurlWqvhdS0MfJtOEFrx+7jnJoY3/xp9okzGfNIEPz7QMUR0niaLQ3+lOUUw6hWPvj7Rd1cYl3
loEuFwZcBC6w9W9oEYlBo22kTcWMyWhcKeWuJpnNpWA2WdCQBxEJBsli/W8bRbm1UWD+1M/cqI4I
t1Qfiz0uyk2Apt35waUN8a6Upo9ws6mOE31M9622D8mARH77jkJ8SiH8HcoUi+MBumGFrXF+rx1g
J0M8LK9D7lcykeZGbeGlm959Jr1ngObaJ7kasKAWS6q1xFiSb1T069NZsXJMHVoUkWqgAvTr7PK2
FqXjgnTyRysIl+Kk/xFl2hK6GKJD2a1Jes0oKeO5XNRHDYrOxPO+pOo6zYY0h/Osz9LHsUZqtD50
nsN1N6mYpbvxf+qQf4tQVm3iD+6euJTUH/pUC1l1CFe/v6mSUQqXiOh7lBcz0hXbWAzpUxXw0577
VfEDCHv7OEysH6B0NObz2l92N1gHpJ2pZxRmnCtBd4MAqT91iDClHWc/Gwu5XpLBW54iB/V4Oq9X
yFX5+ZwzqZ/rDeTwlMOx2/ckeHUp6HTo3IhJ+103MkM3OxizfkLY33slq3AKDPqo08SEjZzLZEIM
016qxW1RnJ78eYjO6H5zXAtIoIqpuSk1tWM1GztCxO+v1y//ZPrMoqjSL5ofPoDEPn8oFiYsw/lg
JqOL8owZgTGaiKwiq1Rn5zXgJHv2gweJwtL84gXfAOsOhsiJZ2tdO4vVJ1GIZnwZZyCokHGq/xfY
hN74yNA3adcgFGGKOqc9usyvR8sGbkkU497im7GT4zTMLzflzX0OIYP7bleb52LKi+JHSrq6xGuS
prfgMgAj17hc38NyfBjw3vIIUKzgWvZq1U/7MVuOa25Q6mPJP8GuK8OHnNHoZfxr49VArWudScws
Wt5eLCacfZszO/Hco8b2jy304yHFoAKBPYmnD/5KAhbKcL/ZNpGMlXXTqO9tSu3A9O+RTEfS+zaL
4oC5wVZ2LMAt+UOni61S2C4abNJplw7CogKguyLJN+MtMikE+pcXulpHB7PjpBmAurC2TfcJy6TU
DsY088P6mqiKs8DTjc5twjvP5i411gU3hg4/srfcsPaEHH3Kv/YJRD7bF1X6/PYrK0O/JC3KgDwW
HppQp6fI2x2acJKrM75kRl/hWecwlrlu/Y4Lp5wCZ+l8zQPQudpiKVQPjgqNFnE4a4fNn2IC2aEd
cvJ+DB81sP0f8R9vhC6j3Z2pAxQAKL/0UWgai1ysFZCNzf2sS8ykb6lZdyDIl2C8K4oUCXDl4ovs
gDZybawP8LJrmL5xYKD/sA1Yo/qzdLQk1AnUp1LO0lWo9FEvhwEHoMmenuNKi9M2wtQlu198qocy
V8WNTjZz8X7kGi+9q2vsi4CrHjW6BEVqQFUfJUpr3lQhzg/MXivyUpnDF13llIbmFhPkZYkFhmV9
IrQOmh71qO8TYJ94n0mAqJ/0GRIK/t8q9jVsMzhv4ouAQbyJa50xMpxmitikMq+XTUNavaYRKByW
+wfFwp2SWd5B2hsWhpnoEfs/zitVlV2cXa36u/NHurudzOQTUd8hyT05PIKNkuWBnLq0JGSCMabh
EzopCeWhZ/YMFA+mFBRDQ8Er23YGWpy/vFYk/CdO7b9VHn8ibciSTDvYxnnNDhyMs/yWT2g5sh+q
+HNnxktyKQ4wF0O25bgkBgoWL7OWpOd7fmS2X8r9WAJ4XoUCglnUYdO34qHx7GJA+gMe7/V1HqjC
X3ttSOPlyZ6AF5S6MoYWA/95ZnKHLdDHsEI/iHfx9HK3AMxyZ4KTUGVLc4++DNtKvE0QivW1TR0K
1AcRHfCqacSvIsuB15LZmpqqZQZR0/VFvJlkrrEWhYdVfiElImUDyu+bWOM41JZz5pDpVKYdBuzm
UMh2NeHaQ7dP+c0LbGOELZihyWwgr+QkRFQXGWlwyIaR7WhXljjsnWBX0KdR+ZTuJNMqndWsD6F/
THjVSChPu3S6g1BHz/mkHd6cVMGqiXD67bkSyDI3AdX0x1jdH8Y/VLPvwR2DP4ocYS+1o6R3+Mwx
llp21qP+LNAgi6221K2gazMdwL66Yoc4CGDKeOiMSpm0S7I2jUSGNcLLh913w1mkV2L27gkPdCzn
qOiHf7ylN6kGr8AoOoETY+Gy0c6ODQs5CsVd2A9Ul+Q5n8L5B3PQzTuP+F2sk5izzYLn6BiXmmxO
RLGbumhvI5Hd64Dkuyezri783Vl06R7QGCSllfTkqPc/w1aAdGRSgkHI9GbHKrbcagtCeGdNhnPW
OpwhMzQLqyIHJTNuTvDQlj4uoIXMenUlPa2WmTjo+2r7Pstqj2bbyj1u5pfFj81AN5XmaV8c3Bnj
oDBUBmLEmAg+o0Pgz2WE7f+ImQoc8hxWdK+pPlDa67ocgTAK6cymwQqKykTXG3gyhSgz2LrjiUqP
ynTiOYPnsigjLq0f4qWUZjMYlzglb/PoGOw8qp/BkBqTwvs8f32TFJWfte4k8M33pii5H7Lb6wwG
R6EXhaymKKo8kYSoUCwQ3XjW6giJuc9aDPaMmy3Yh0MlX3VeoXcreR+g5MYPPjuCri347XjYc3ox
vmutOrDgM3dPUKxTfk5NdncbHcfhhg+LKrEIOHUlkYgAVK8crANfye6KXkdBSyitjuVhNuwAmVzX
8Ol1O2zKIf32pwIOeBS6Vt0Dkg5qzwEAJRrqEX1eUNnCzhs/Xo9tk6n4GjECUbshcrnxTqpQfJBM
yJti+WCLc4DavhX9PyjHaD/ZJuGY1HxvW9prJUZ5KoeefXbDZq092L9djTMiq5YXJBLIZKV3Kd80
8s++YJ7fOADdevtDlEsj7iLgKMIgqUmg0XiIBuTTmqfKUZUt4jDdcaMpFB88OuRFGMXioBCo9mNE
mb4mebLQCMCfaHlzDXC98g19tpGOlOVYojGZ0TJZGcjWHgX2nG3AoszchbZeYHyF5GMHwNlSKoIY
tWHpo45rBmHeLR5VgEItbLIFZVN87hcb03J1BYanEqNiPBVlYZ9gbTufM+C9CBsLfdMTh9+f5jAj
ogKJp9cxp1TVhbcCsqATbx2XGSpBzFfxBvlo2KsOMpewAJf+NoQkAUjbCqw4rkdfJ7XTbbF4BlKN
mKvVu1d9OxhVYtA53Vg4tDLFh0iPu5rDssV6t4RVKbSgMkAWZg/dtjV8M6A5SJ9t6eUc3gkZVOf0
Qog8qnJNexg+nF7SO/DMGUYuV9J/HHSeG00ONuGMQPUOu/EkOfVXhV1dTBcEusPkA7a0IUug68qy
y8RA2NvyMI7SSAFyngZczPdnUl1yPB+EWfZl6eWylnQy19wa8+DYVJMjeLKTs5r9rRvPHGjaYl1T
yjVtA3CNiLscF8ONg0kABx8M1R9BYaxUMqq9Kf8P7tamUemYNfXcd1PuPuWOAiIktmfzTfJk0V66
EgpG8f39qD2FotjPCEYQCtFMFBTJ+z9kXwZceuvW9qTET2TUB3Ge4BD6NhIaeV8tHkkkQA0cUgZl
kJRQCXN/QTkwooYSy0yx5LBFfNSsIki9AyJrS5o5cK6AJZQogOsmUCPK6/N0QSS+IgsZcwPDyjhe
25O+diy49lLAPiAfemCfOsTfP/nDFFCR8QjNKS7s5zlT3i4up5wmmLXySeGvXHBjw1vsyN48JbRu
qd0Ns2JKDVmdwDFhxILshagd6XKGsgFdORk11t5BdP6CtpkrF59y1h+wio5SnOGmGnkUX3xQzK9i
c81m/1DdSom4GpUWjh2PTW5K73WZBseYbbbML4KBbi6/Dt9ghc6RWqDHJs2DmFGV8deO0kvKrXSU
ZJAOYlPaj54oXT1ngc7ZEiZxllzHhtmCLJFSGRMFHomul3QgVc3HkfDrPh//XV658pCpFtoGeJ2W
f0iy3WxH+2sCDH3SIImzVD/GtOw8IxSimlKZYgZVP2qFrFAXEKF//SGOSFZkOPElXkEFmVEwkw56
B47fgT03dSc2WJMQnaKtC+lBpDdmpvH1vD3ndogLu/7Z90p0TGdTjGmVFMEAwC3+DLUGRPzuuf3M
yTOXivPvqlPb3bRhoTkvkdCVpVupt9n5dUYTSWd0zXkYfI8aBv8iREAOYL5WsucnjP+feeFcm1gF
s4jRkzy0xIUfv3nR1+Rn5VnsS0JViUv3bj4cx02caXN02YSY4jHrqXshpb4+0fwBuecuKimln+ql
6W1xY6fLxseLnD/hsXOO5HCNacf6FvIx8/pQik+Bc6bYITkwLakIyLAxq5+ZS6QVkQGjlJVKnEcn
GLXN7b/+zphsHQ7ls9JfKYNS2UpNsmyjqdJ3IGocVSX1UmJ5nDhDZBUwY5PMgueyFSI6aAbgAeO/
Kj0krZXNSq0oEdmj2rwijIrCz7dswgABkYBF0bxfwA7OWs4l7Lmz4tvOPJpkN7obAbKit3SRxCjG
d4rqEdk8ZHMy/jlrHvweDVvuNSQoEsPmbfubrtLLyzxBa4vfVC9ZRediq/fjZ83Qrd3UuGIeL8/S
eXyPrOodIJxzLCUHa4sYMl2d+eUssLala61A+ucB2rvScSdY9jvF6MTjN67mwAbcoWtNy2F2JuYs
SgEDPJ3jxGJto+3p+G70eNK7lE5y6HN3qhHv+VGbW9ORE2TIbyxHJ1gI2Du+rBN30OsOeHgcaXdX
M4vNH4Iki8GtGrvGolCc6tsPfDPJKst6qbzgvMcrRlc0/lzR3qyL7/sqQBIcOqQnnzPUkPZWxKfY
8x0O8Rv8wJd96SwwVLYLcKHc9aIAAB6r7ATsZU/acMB1GmrnRTOlD3ztGezQfdruSEnu96UXCpX8
2ur5pGT7kCAb9Tt+dvJxlNi54fMj7lxtw86jA7q0nFfZZjs/CY/Ph5MhDGQelxoe+2leUfhkzBJg
z/+jscq1KGcl47NN4hxk4oh0pHc+kqFk2NmvfOJGVrxPM+S76wRfTlxAfxGTor7XVhUH98g6ZI+I
j398dO03QoO6xPdz057xx1j4I8i1N/jp8ZMIv33PtTykTQfxCa5BEYW/aqdvuacPilR/c+CMlN/R
r3jrzqXQz/eyvM6vCpt1A4yd6qNFMKb8SBo00SjDOm6tfwJk5sAqOnvyb7GqFr3VLGMP4OGDn1tI
4a3s60cpEeVnbw4X86j+a3IjmbytxbFVqLfoeyrr4tivePD9Rno/WOSXu5kuyx1lbFoWGC7HIy6b
97K8uy6eVsmwDpqkzHShuIHfp7dhL8vXyZvHTyZJZhlSnNRCeLFqCJeVllaI27ELx7ouLYdd1sSC
HxY3ca1h1fmCFkT4ZiB3xeaTZHBmgEZo+HQ3HaWzNk9dA3EpldozY6kSqrodERHTm/LpXtJOFP42
/Nn1eneKpbi0fyS2FR1oEcORi3hY+YLCYo+jcbuzTdncsHb0i0m7D0Ax2oAgJRsL+G2m3HEnyR/+
qLTITGtVqA7e9C0uZCQ45f2k4Ze3upl7fzknwESsjD4cCeUQ4JR+qpGMX0S5kCKlTQILN43NE2rj
GP2YnEXh1cryPeTpuyA0kNI3NonNUta/JRetiNJnJyCM9N4OpAdsh4tmSqJVfd+JVXOHxPDo3QMm
1mmReUQbN4WSL+TM+IDHubnAlnD2rtLD6bGwbWrt6jg/T9ilDY5NJqVzZIZpI1mfoqUsF+eSQCRS
cb9ItPBWNfUvBQe68TdeF9fGho6S/7S+a54oqlG1hFbFDW2XWGWUDAQTRwxov/DEIVbDn1svmQur
oD9wNXZs5FZ2KuRURVKpVFO91fi4tLWh1frCGw0L31vw5bHAHBxRry/Vq9zJfQhCgOK8jmTSOUkZ
8nlaVGV0R+2PwBqZFuHbCOTKIAF3UGCTE7+U6CTlEWgu0mPKDjUSCsX2OPZ7V/KgrzmLjrXmqmdV
+X0h2hfmqUfleYLfbl64R9SZvm+A4UYeFx7ii9zf9MVsmcGQDRv1yfdn4QMDOjWq++v1lV8YRiT4
DBBcGQLq1kFS+15u+8wUppxGn0lW7R9MJs7p96QfoH6uEZGWJ9Ae2uNJW+QTMIwrbkpgNLAjgqbR
H1OELJqx82Rdh+35kzGdnqIE5Mw8oaBvbGicl8H2lDeIP4cRjV8azn9u1la8Khnq0Tdli4/VrtZ+
3tJUDH9EZvhmB5f92HlcjWAdx2+pQgtA8LNeKw8O9Ouy2pk9wIvABzdUegbFFxHMr/9BHAtx5Fma
U4WYab0zJTFKWjDhovD341InZwr7d0vGTpX7SqtytDovsZuK6OjsiUZrpPosaCuhAh4UuPZgS5Uc
yZFZnWEx47qGeb/fnRTeae0lN71Cn4N+uUELpizy2c7LK7TCGAV+zEOkb8/EDXMd6uUHXLG1caLc
Ip+gge/o2rk7W++hSZbf4l/3y8Vai9a0d+6Pfhodn3diPDD6t/5KCiqN7sKD8hfeSIpOb1JkBs2o
eE9jYtCtsvnD5ntGIOt1902GW5yKA2JjPnsdouErGNVcZAyjN/lv+IUc6oO2tu0P3yM6D/WsdiGs
RfaSdgkCvsD9ipT3hI80h0j7u9709rcSjBgCgf7IdbUVY6eZhP5/+MW7SAfGY2Lb8cUDpBEqJdM/
gzOdSjSW6zkc+4YxQJ7P1eQtbYXOASgadZrtkJGvPuCybLdLo2RaUVk5n9R1BoQkWekvnrb5T8hQ
3c6+POXvsorLgUDTiMIEVg/blL8WMyNlRSUiLqVdL2PCYhZxEeS+vdK9U2jyv8A8muYVUo8RnFH/
WuM+ElEusgGZTX8hutwAe+PZrfxOtk/h47gNCBbhdAi8qk6UKqpCifHGJF3/OrVGRwqW2IMoXAdb
FY6PtSwPbIOGSa9mr5ebevZjEhog6Xu5EK3s6FzKb2J11Hs6ts/bo/NQGAthkhuXC7x1/rF8IzXh
z9kzfGywtZ5ksDzQw/p1IFl0x7C0l+ZsG1SrZxJKYxhImUl0gbkJeg+Bq5JUBTiNKL8qka0QNhUP
5BUVPMmMwTezvZb9sM+6c8FxPf+djy/+1zqy87mr3ow67tCuIf3a8McowBUNy/kyzOUdA38Ofhjn
7x0Z4oQN0R8MHaXWiZjm7SuXO/hudhfTdMt5cKAjmoWr6EZmR0pkB4kGJBEVX33KSfXwZkfTeAL4
lwI9hkgkXzfPFH9jDuzxXvDeHQKvsb9OMK/hAigereBUW8tG6XTU3jwTNHdaQOH93ffu2ZQtkPAp
k42+bifOakSeOJgCxsXzBdPyS2OZkmNKLY6IeHOd2z8p3eYfqaHhQQ5lMg2c9zC4vfZl/VaRZ81i
lZ/c0dlvnSEMkKjL3abDUlNHvLCDbcf70YzVXNSovqeNu/dTeg2aIvjZMvhC+id/gn+dBDNLHmH+
tEPfSqdfTJbTV5DBCf+I/z8kLGTfiE6nlxPb1Iqeo4xh21ndesBuCC556n+xfz2nRVjujwf5bDTB
YotAYCFZ8SP8qnqFec1xQQN0Y6k8D09I2TM17WWxtcMhde9JmTazLenkZ0Ip6nyR/pgo9vEzBZgO
2eNwfMHX/n64rb046uK7UMu/yiwJ++NX9NQ+jsp0xkfux8/oV/TJyThe0AM4qjq4vmhAAqFT+7Pc
RqTUuEJIBOkzk1JhriuSzlxDPuCAcOSxt9XNuF3Jj2eV6/gXs0PntF4m35a8F4A+vb/DZSvu5VBi
y6x5s974weM3BQOZVmqoCkwwIJPVLjpOzxnOyVkN1KABOqCzdAxtSotA/aXxFrHWDEy/0FU4j8NU
XO1gbFgOuBr/AvxNTvV0ZTtF3461JZyK+Vj3Ptp6oWTDD1I1tQin2TlM/+0ULO1AiQpe9MawChn3
NnEudv50wAVPeJ0Yp3ghkJfnJYgqwhP16hMksx5w2UCeZpta+fq5G2vA3V7y0SFadURK8FBcmb15
puUCD+vcpc31LMnKXi2dxU/OPpRRMfqurUR5W+lw/omeyH6AsRlMFf7tUZe6lndqbzAtEfGgYQQP
rnhAtXhFzZ14rrFF7yQi8v1dMK6Btp7bMp852jCwDeaIUtT4R33t4qZl9MOCf3L3CzY2+s5O5qyP
J7at9OkkxHbl1JxdmLGZNYqPybdWo5BefWHf0gCY1by9ynsKmp4J8Vh+YW745d+O1Tq7zlPTWIBT
hJ5HS3igRg+xGuYRuGEh1HbE+ZUSZwLSeT18ZvkYxpkQ4ml1OZAcYd1dHg8O3SAKEnsqeqodKHTl
a1lR2YB9JXkGS3GQoPioVE7Rsuf2UrsOWFJBoU3yIb/bZJxeTHn/vmYUY60yws3H9k+blpqP4Ruh
vNUvaWEbs//dk73qfyPHBpqa6sMxYGDhm9pCvSoK6OeZObQ2K1+u3lVohS27h2Xm6ZqPFUFWFF01
w6AGOaNTxIcasST1rrehPH3R6vFe1ey9jShl5QgptEoCI+wJy35tasFvKGBqjfgcXeUaB9fMpDqT
8anYQjY5J4X39P5XNNA9PnBZRuUnnZEoVRBrHSkje8KxXR/6gbMiPHVh+L3jEO4UrqAY2Nz0WSAk
7+2WLClcDv0P213+8oat/k1ruzbSJt9kQzN9yEBXE5gSfPVaqCQcexRJ91uI4HhO3Yqxc2GKlGtn
iPmkQKXpN/IIxHiEE+OWj1inyibDGkf4q2RryKsrF0ipAznDUU9dGzw4zYFwB5qUZSaKnz+cYqYR
LYHox7hDbdjd+/XZtxGlTIdvWI4CFsJ1D1zNjBTQPiK1UwS1hs/feAHfveDzv5BEe6x0a+cYyMBR
4LwbT8x2PW4fydA5WubbdGh0jkrnr5VvN/kxpoA9Ga+pt+gN1zD1PBtEXwE0/0EORSFCBeITrxFO
LnMVQuA1Wbj4fUGPg+SaLUhA1zDbDNTxI7kmUjug1x6NVPfse0DBJfqcYc4Uv1nVaGnaG674yz1w
hw3zC9OKsukKsy472U8qN+gJgO4Xpi72D3EgbHWMK1z/ny9fkKTROl4tQfY1XQ2pSOpA4mzeUSDn
mnIi4Hem1l03PY9ANgX2CAybKi0RXErtFYftNHMccUo+aKlov1jPOc8r1aQcW0ueS85kXrg7JWbQ
1m4Pt2O+tlyZlSHNbKNceLB8kuZbZ4/U/pzzeppkCtVFl/F/P4XtnNmf501CkKC2MYoi8u641H/O
Y5Wikvl1WdOmIQZmfWB8LCpN+1zppe3i3TR2vDJt47fXsqONC3Zvic1EJCexoZrE4Y6Curyeeii4
3mMXASybx7f34znbirRCxlIi8qwdx7IKNi1OgyoXrvAbmyWvd0pURScKpzqu+s38iYcih1m4dfVb
2uUG19zhrUf1V9HnHCiUd2sg/fKax+zcLHO99/Zu8cwIT7ObUErWRB5Us64x12+1ABPbYxAcG0vb
OiwjF+wRft+XNuYgfgXE5pXw0+/bSV50ZlN5K7QlrNb7qpRbL4Khcmw/56f/OGY8htrQkkWsy1Hn
7/8EtA4EYONSilbRY/TYYVfer39XHUd73I5gqBGRNuzt70/b56wD/5/CjNt2iwmAaYZgZZhvDCCp
UZuCQjPQyXXMctetL+5rNxr8SEWR4yFwPcJDzX+7vU8Sc+AZOvMheveDMzZZIhvm/nTH8ANhywVh
iva/ZF3TEoFLWypUjyqtuGhqfAbj3jQtvRfC6ASxCdmSurvIbvDWOPThW/vzENMZfB3P5pYtmwuO
j5rQSWOPgsX77qs/3rKSB9+1baVEAzU4OAjwu2dos9PP9npbxRCEPE8oZwBGPJA9M5POGJauV14e
Wqz1pWu83kwVBAkWHqDLs+x7ly+Ai2AtOVKEnfkU0WZM3SY16WnXi7auLr51W9ms6GEcsz3jBfUJ
i5iN+V/r14CBE6fcg3rjX8w/G5Vm9HPOmCjOUjLE26c1hnhPFHVBlhkAax11zAwwRc9lRuWR4Nfw
TBfTpqjfceS59oPJNkZ8wyqavixWVM8pEh0GEjW8z88rrYcmyLJOX/43MriFgBo6Q+YtTiZJvLiQ
yBK9daENkIndVLivapAoSRstJTiM3HyTFct8khqzlOrRT8mTcLdczikp/f6nLAUQmKJdUmdzQmZP
5+GCrZ4DHseCwmOLeDp/7XA/sdzE2A/Bo53NUB1TpFDBw9S7TZBoYPwRqqi1HZAUGwoiZfkgC72k
9kp6fbnry8Hmb2LRJl4TWL/JewWGMZx5wXGpgLW3gOB69Or6bCKhJe+6CCMAP3aW62W31letmbKK
qqgNJkkFLu4tSH/YkUU0ZlNEI91uvhidockvjyOF3vAsCiXV8YDLbCjqx0pq9vpASqoib9fL0PGz
/YIWfUW9BlEaC7wfL2JUsXtnxMwOpp+7OzBy9UGHB7694r3RTCMbr8kik+OV2sR1WAKTwRd1/3M/
OTAkKpVZs30S/JTTsbERtU0QtgDpZ3+k1zRYzuwf9+3O9/f3FYteKnHSinVgstcaXBKNKX4Qe6BN
m2XzXQwXXfZia4NYnJiF5LCCaZgA/DfdCnnk8NOkiaJK8iIM37CJhmEMglJZACTWeO+xL3piY1kD
rOyVoZCPvIGU7mLD3ND6r35WvVTtGNp4wh1FU49Vb03HwaAHIiBeTZncPz23mC7snU/89W6oPRXd
UGjspBvvoH3gG8Ki70ZLz+RNvINcTj43ePzYws954JvhKX57M99SZI074RBF6pTvzlo0coxpJCbF
qvTRYEGWdlkTweVZby/IY4tgoJJo+OgFy6kfyNte/2zpLDDpNkAGxcgskuK1gXTn2/eM6fq9AF+E
qkgrTP3WHn1H7huUL/FZ7W4lQpx9yDsa2mnGX2v3wC4Sl8Xy7QrbJ5k/jgvaCQHs34hw+wZzvEGp
V+SSjk3vgj9j69WvOoVWrh7EkGxiaLnpnEvqEAJrEfKAkdpcN9nVKTes05++a3FTvMBZM7LMdevr
1K8F0ClbhErnfWJQ0OpAp4PMr2+A75MXd9k2MD9EAa41XOAtaQg+CplqSdos3kl0Z/imSDAGZ49R
8frokVjy3ieo1NZNYU9GIJ2EWezZhmAGeEWouPZH5FvwyFQ/fQiDxuOfxkNO6uV/gzcoHLNXLIg1
7UJTrNKuPmgxTQzvqF3P4subB47OSC6xmQRtw56BfaxsjQiD0yImOIkYjXIvBFH8FmLZCnAeafhv
WZuGhB2ckckqhBytOyFXFAPElHOGGJr7eoe99T9ysUT6hxm+fYm/XBI9K7XXi7qXwwFoXGkGnt4A
wsV+PqnjrJxsvIm8dv+QwkLKUaGPGyDWiPHysWUf0sfjkTo96sMIXanzwapSyejIcySlB12S5n61
UVfEDCqLbcTKirALBpqY5LA7KPdH+mezQozbV0zOiAN7l7ozQmL3qg2/5yMTLbMXDhdvwsRRn/fs
KTCmujEebASm0Ob4RYooNNAggr+9GHBiwNtoB+8BTs4sx9sLZDXKCAA1+wzeyWbL5RNZFB0IY6PF
utYGTWd1EqF0sS0anGQ0it3Ja/Sj0bm2H3//nF7sOOeenjabqUVsPUmaDYoJ2QDhN4RmtD1WvYgD
3JBqa4tojiQstNk/ATPsDMPmejy6UbLD0VB9fcfghdIfwleNkl6XaxvkUi3bsJsF48w1cTOyITH4
3vCol/WjvQ5rJsqYVrxIzu/6C6TMvwvH+wnLg4jkVBpsJJrViShOpHGfzpofHZ5IJxaR3WGG86tv
GoIOlyhZLDDuYBFtH/Y+spOxJHDT3dGiEPCTb+oAABqSYxlvFfhyLESVkDfn1DJLV/ACe6Q3hPpr
/afUAWdEd6K1OyKiZR+eX3kg+TBLjrmo1pkJNIdHeD3ddA2x0ev1QTzt5yLcBeQDxO8NshNzLYXO
3ASsvQrJtjrdcBrnTiGG46D5PQeJHrxjyfdKaUZCHBLyGY5B9jOfLPrj155H8C7FRv0pvW6ZzOj+
Jh7SCZokcMzBHJyIQBZM8jVHAZCaEsiQ95JulezlLA2bqEeahHCiJ+BLVGtUeKCQI/3A+hytNZu8
+OESNoDMU8TRNxHVdndrr+QdiL2OBA5GY+CtVD6XLxpyxPrgOzhbUjse+C+mzLCj07fgJygwsNOI
GFOF6PnlI7ZbwfchxxSJpoZSlhYx0iPA7eJONy0/22qKBdSzMSsZQFrK0DfiEUe2My6KkSEjULnQ
MadBasYsKZ0Xoa3ZEikBsmZjmtmIzcGrAjJagkVxInbR8f6RqEbA836AKLOzCdq4/RlOMF0uiGti
curMLkpRg8MYPW6VRSmOaBenq9mdTIBsV/iFhaVXXf00exhINW/AKa+x+4qyOC7uyEgluiLdILUC
YupcPmI0p+68KVRtXsgg9UvBLAvWmo/AKWAcLVznt5hWmJIcZR+PZr4EcRrYRlb5R4OlgMUHv2Zy
pVDhLKWi095N/YPKXAOWvlPG8wiKZLFYfP1UEsvIp7eOonmGIyMwdRzy/AisPFEDS8r0bS7fcktF
mNK4IV+9Y4HZfdYov6lsDI7ya9WrADt1ftQAkI7MfBZEeGz2xyyzoi4bQzwyG/2zEaKTA094nf4E
vanbryw39f1KoI8EPmXlBTI/Y79I3fR6jFX0qvRQscbg8BuCWYk681h2eo1yOhvuWzXlpMYiZIto
E46Tk8OztnKSOqnfuJOmnjh2+qFhFV4G6PQt6X+2nk8wQsvE7HPCyLQ+iOd/7jcFkEG0UrmlKMgW
z5kTZwBc4NxiMo5g0BUCsWGDPPL85HtRGABw96oAmK3gKSr+8GcaYLOP0I3MJQay06Z3c70tpbaZ
VAgMl6zi4vH+IUk1Ki5BvnIptKjTwkpPRU2dwCu7xYfzd107CPF0JX21ECS4DZkPnlWx1FpbO2kp
a7wFzgbZ27ebrW90V/UZ4tzDneHjvP655Zck+dSCo7xMfBN3eQLbluhrtCRaf1IL8gnHh1cnUoE2
IDnzGVAD5UI6EKff8I3XK6KNb/oR+JGDA97tziSHhj1Y/u9yKrUyhKSnUOdk/BMO+MnMveERpwFF
faJT3qY3fMqBhY7f07uZ+D04/kM/h1/9/280pdlkS4b+2rHZZtch2tSkHjqFLpTNT0S9FMji7u91
+0vMZ6DKr0++uv5AsyZ65/bfnUoKIuFoMuYxiXMcwzN4KHdyOuOfI2vOyQX1g3TQ8Y6sB/Ha4n2m
AMMNU31GsyE8jwausWftHQEgQ4piMQajcZsKe3AbNmDb4tTjwu6lHaEbRBFGCcwZ2dPfLHJKMgeI
g/W+0l0L7U08/EhpqpxxTp5iSro6JGvzb1cQm/2v7bK83p8GapVr3JbQkppHcuYLygcrUcKPJ/Zm
fl3hdBXFFMhm4vn5hCvXsOko42+Wbsj/UWBkrBT/ZCImpx+xLT//NfzEhyp90Nof7dbRzCq18f/d
MKk/hpQsggmZOC67d83cIQLiynjncUjJwPuaW01faLpOz5CSrhr9Jt9gbc5NFtlHDgzknNqktOIa
zS+T6sFO/k+YxhtaiUrDQrp4pH6MLDU/z6I4LuvKBInrIbe6+2ixC0/PWtEWERF2cKcV5ZlaQLFO
N48ArQMRmwBMlgsbbNViqY9KyJCx1qtB9a9+iNWvhd76HIgOL/YV4aErtIIfTDX6boHT6E1gGDpI
oZqdxgPYOoTkgo6RgXlTi0RopBRVacJlBXHxUAtASvOSrqCo0b32ltT+Fuoc9M3IY8mOiO3OQsic
qTVIJrwKBldxRtnN7E52RtB3hmyerMhNhT2u0OaHPjK+m0GRB88pefwu6rEruSCBqo+pi5hFD//b
nHO5D01pxJqAO1eaczV1HhEiIm9CSpkr95ijSXl38lcvzST957Di+XGoDzD/4Z+Wvy8aXZP2fBxg
xXzNuLDxRtJw7BA4gQQpzza0+DllFeAWaxVlDmp1Gya/0W0CUpFLKYshnnBUwmqpv9Ib5lnZJAPW
gdYXO3y0iMLSE0vjWNZh8/Dquivg0NP2M9/nvCk3IqB5GdPNjVOZv85TzenEetkUVBwgdMIvWUFA
XKUG75GgIrilJZn/5/RwaqQ5OCO8KnjtcZYOG+Uqd9SaEwdWoqOvJvXV/SXBgxYWAGxErZKQ4OSN
yD99Ce7pwTLrOzIFIIWjvC2LtRnhQrzlFny7mgy1omYoyhH2vxWy50y0kTAd2hVURbj/NjoFtSjg
L5yUm7/rS6wPMINgQPQbuKQL1pvFCzHM+FfhePuy5sB48SD6W+j+RzR5PfkmLGj+kXWDRtaeI3co
AS05BQ0JRUB5UOZOmAWPm1sfrWePQ7/owyDKDVRc9y1sjlBbSvqgmnjjAKQzAWt8x2JdDSZfwvGd
tXDYrCDOwD00QarHANCqCrDSF7Eq9dQGOsB0MVmJolrQC/vcoHcST1/Wxmg1+yJ3mJIHi2oa22wQ
yCmuqrV4I+rTPvU+rbLa1fClU3aatn5x1lUyib7qyrTemEavyAJo1uAgTtJIR9mlRjFpzCTRf6K6
phmogtJ/WMvSoPjQDIKq0Q/Uo4yiE2wrlH/oVjbYmHSP4mPu4L7z9u/Y5iTNitiZXU3VBuhMGFqq
Iu/4Y0HlFlCBKspjQjmool5T+UFeHt9jV8FpHWyy8+s7btlcY0CV04PSpZTildoWhoGjp9vOunz+
W7E/BxuLUgMvZAIvm5o5cvoaWb+qXDg7tM0WeFOZYGS/ekYX+BioDNLpAmmYoJZ+bp6JUjbYixkT
N53bbX+QuMH2XR70nqY1F1NqvAEX2P0iNbSoX8RA0sT1+kFlZtgVdimgPbWIbbaQ6O658ngRCMoG
kcbMX1RWxi6YSpHUqw0Xaf1wysWyse6dPWrMM58pRudZKtFSmmXjeMgaj4oRrO0bREHtU/yljsEw
8AbT7gW9SR/y1FUVlgWDTVGftNfRJ4UOCL/U4IBuNI9CrOGS1518M83xZH6fVKzjLhGgGM7WHcwA
If92wcbxkR+vOsJ8YUKvDpbUY0XmvzpXTFgIjG7m7//sg0rXGDjWR8vm9wdklh8jpgatWbchiXpo
4ef/k0Hd4RHDqO+XwajX+GByRVAfv2/XTRKlgW/cp6PTr/IpxP6/DneQSjuNPeN0UgBEJnVwMErp
agySMy+j2AE1HJWKrYKxOEUI75jsIWXBP5kGxNMAve2NGTKWxevarleszrlHv7Jj1fIwWcORu519
WH4pGykGSXAqjA+oIDAOxZT6X4jBgU1+Hczymse/XH4H6nD9xDGSu2FQIa8AkOFRw9hzRrH93Y/g
O3VfoRq/di3+ywuQiuAoxexuCntVp+zCzKfZAmXE0QoE5o3Ntx94Q4XOca3LqgdQ/4O31podwspN
6UQVXE2tSARLye7U+elGyyZG573d8p6vbmEhEScz90VdHyOxqwFwPZ8sGkONdgUB/BaFMf15R7jj
pZxtnGr7L5dpM4tCF9DROm4DWTl1bQ62EBB5Kygez1FcKRdvLDlQOrq+kfwZPTCIgItiynzwbZoC
SVTLwmulQ9IPW8WiWdRGZo26EXxRqwc7yutzw4/LdXYhPzI1a2T0KthVqcClZ4FzsOFvQslyEfFq
hMNGNHspJeoyQ6IvA7RPeYouItwslvst/Q5ck3zR/MLN1huhrS16LXjY9vdx4MIqiD995G9drQwL
Eqi8iuC+XbjAunPHFoDn2zZRHGAr+h84IQAJt5UCODNuvlzI4g3+/IAXLEmR8b0xWAdV3p8/D535
UZGvpTJhFF2+9oE47XN79DL8rSlq4pNi+nG3g5tEVp9yDmyV7X4umXTk9xtgUSWZy+L3EXnZ2jvB
NQWnIXaUjC7lvVSZjY4h4PbKb5ti9vPhR8sG94mnXoODHVYiaGmCEsjPzTyEB2NpWL1uXAZwFQ5Z
cDLltlWL3YVfoUUDpKJL1B2WTatZJy547ESu09NcF3JRF0u2Y7vci/D9WZVMSpiwGSrQkUMe7DRF
/+9cuJTXRjPhQ0tIsBppgkVXx3eslpi9jLIFK8jM+e8VhNR/B1CZCrrXmMYYSfOMft6z8oK8gwCs
CH27rfMI3rayVqdiGvntnzStvbexU29KXLkNC4hbSd3/HIoLelJbEwcn1hGVc58MKQh9n0nbqNo0
B7Ha9U9mpDgiv5mA6Cgwn0bJlob6I5EB96UFfo3mctQdAZyag8IGrefOnWkFOq3DeSqnb5pjyPAU
rYgwgcYkRfMBg+Z+8M2OgYX5zBGVK/QiB+CLNdc1G8Qgyl1tTzLPvxLR1PSezT57q9lTxw1hk7EY
vqAnN42Q4fbiYGCOrejzjIAHAJycJUtXXlvmyjyhoKT2FS6ryyf8LbDm2fVTWFL86Hen61TJNv+8
e9zzq2L2LCTtuYyuR/Sn3lUzYz4jP9VOCUDcFOMRbKnS2t8f4PM88a4ffxuLh/72e7uWLRVe5mW8
hfFzJh9HvGSMopoB6hbmwESyy/BWyFKlKVvQ/4dkklEng0Ht04iyq+TmErO033dMZfwrBo7TO9b0
7w+frg48eQhEm/vGWXAo9yTnJCUWw1YhEep5W3293Yd1Y8w0RFrhoxnyARzewAss113wWyLAYc3E
Ca0QXoWgMlaT03A2py8/WxTh4iEkEJwbb49Xec8fCHbYskdshk+jbEuMGdewAxU5U69rtENYGEQV
FF8PyjgLD7fgoBjF5Fx8Q1boK+zuKRtMqRZR7HBqtPe8TVpwKVJF9VvIHpTD7tQKk7J9rr954oFO
kjSaRE861/3T/IiW8e7SKgT+uoYGAkWcZa5WHAR/uxKOubZkiYps0+ne7yahsoi5LzdGBJaBt3s4
ErlOkwrVV4Avqob0jRcMRG9nvl89lGV9IoLp8M3cad+l+ujkHXK3MLhkyG3/l2QFS4i8o9U4GeH7
jtcmwKW6oWnhLq8yiXH88Omx1joYCW4d6fOnSSi5o3H8UTerSv0pSZte3PSs4kzisj6afSJbm5Nr
tsigsWR/96kUbXm6lJu00RSydMZk2fWXYxjD8JD+8+bWhxmzhCCPuZaMPT7tNh5r95Pm4Wv+qUT3
KO8NRZdHSxvnB3LROqAfie2b90+ucKV0c3zuWNltpJsHAD7s3N4DnkzN7ixY5qbU/DNOZ3qNkBaE
eDGxtsR3bVYCIZd4jlEa/xqFR2DBM8h29U5IS3pzNPW/b2C4HcH3aUlj9pD0JlC4evcpFjKUPSZj
x7rdJH/GmLZDtV8XO4CS+Y9Dfsu804DL+rS67IzcSd4VdZJT+qMf34ZMFkLnXu+nlR8P68Hn01Gx
acBeCkufWsY2ZyBKu6sHaCQBl1ErFCtdQTDrJjh1izLv9ubeEDiWiCBEH5a4gzHkBbjTMk3Tkzgm
gYnsNDsUG/wbADLh3dOMDlBLMp433iXPDFjGCS/WFLpcYdFXXn42gkRzS934Vtag5hxxzFfJcoLD
2JT85mkc99F2KuUGzHeZE/t+T/4RRfBYo804VbKCrN8nSQaOb4doZWuyWFdpuBY7Qp/evUfcjmWK
/r5706xr1ilSZ0Tztvz7mH+q0a1zKBKQks48BaAaqAIVTD3NIQj24e917czHy/YCZykFT8ygrAeG
vX6k3ResfcGTUGAvdixtdM/nch3OdGu2ots/GcC803PD+QZNFd7ILKXwjBb7RCANiTz1fv6hI0nP
b/bZIR4Y3hLs2WP5yESBP9eciFGWCypBRTVyvj783mIHdT9iorKsfcdmfME/PrNjews3Q/18BQ9H
u+mA6pCVys6efN0KWN8IIy9K8LFwn2/XTQziZwXYqZIvyPDi7PdOBF8LnXYmH1wfWXGmvLbucgl9
HAJCKsUO3xcIvl5S6EvhXlS/Wi+R9/wm0MxX8XOKYR+Fl78YP7tYkTXsQoL1gpQ71cHTFNHFkJqO
qqfy5G/mmkCUYRnpFk3g79Nrn3P81Wep2dSthMNeJg2LgOOi/Jqtg4/7K/pVJH/kMtJc7fR8o6sf
irlKKCBj0lnGMCbdgRN0+D/2ZhqlSoLel+I3VKxBalQfRAM3Skr3b9A6g/5IU2wSSmUp0CU8zCKp
wftgzB8FljolG75v28KXEyhi26EygSrMDeqV/O3tujqBqK4gxMGA/mo+PQLus4hakwP9nUpUYhwB
2U8VK7ix/aVs+8q/MNsVVWYpgYobPaO51By/91nr36W+5JoHhW5shXVM9+7Zn6QLNgtAwKHNxI6n
6AoMzbx71sVPczt+KjkziJMOr5xMP9Rfw5LC4M+DGYtTxWVMtaPNv6CJKVWnoFIs7LhaFvKkMzQ5
7RBXe9uySAOYW6tS9PTJuue67LiFSsYJBYB6LIyLzGmSsFmYZoD94Gpl4hVYgtbuqlG3fJOnrfyF
nRVfKhTzTGyqavTD4OwNhWebn/MDudqEtqR+m6SwH1/JWoCvTWbTx51FcsdcP9+ZB6FWTWiUpGNS
yfXJ8p3nlDjTNoLSfXozkmd5IYfuYPmyiO6cyawIaldPTaB2+BXEDc9V+IjRykdnRUR63T0r8YN2
Koq4LJP1L1WwXWReBt+CC/PhS72c019ZijX/Lrgxvi+I0bs7w21X4nNxbPM+QUZGV5+fi+MBTxmo
/oMDR5yU77jcVoIuJGnVvYrmmMc/Ho8QWrjm5xlrO9WPAk0qTENTU3iSyBHZ7dFrWPbXmzvT8HPA
+z9Cr964cyo19pl8EQEqWa3lIrP7fBdhCRBTvD2EeZn40TppHLgMRvYqMwNwg9TM8yNlBZ+wBhNP
fyIvJt4tn5ZY1GBnc/FZdTzIEIEKjnqbQKduaPQ673z9KNFtHyPSIFPF+G+iPbshSx9bfwedTNIp
5zeu5jcVrOYNKYrVDVn07e/q/vxRFtRExCf5hxBo+MwuwFilbI1QwKYb+lUDflAg6lLkZUG54MQ2
P8gwUFVoTRQuFthplGGjP7xVTbke5Wjwe0yeyjYaEy6wUOTeN8CWs1yFSesG840lvY/SX0gvG7gB
F0AI/s6TUkOK0WdzgizPXpHSf770JXlGWRwL9SqgktwdRDeRqB2ZuQ5lRhDOaKtToLAnbtmUcpmu
StDL+6hpyi1C1cVXl/cIiABkyk6RpbijT14tLQxtPHIV0sQkQA9Ti+XPDBNr1eCjSDsUgaddWGrd
M6omhM7mwtt9oYdIC/LzAAVgzS9qXjalrhtC1EonIESV2/j2nqxIlP8X8XlBVT7m1mQQ/NTmn5+a
DkZNIaygcXFfK7qA4J+X74FazWkY4IGw/3Vl+XzB2Cm8YCcz1/ofTznuV5h/LLskAgxSsfUeMTsu
szlQKq9sybHEJ9bSlHTPuS4/XnAY9CKoNQ0BjIN6UIKfQDlSmN4X+mvSphHu9PWnpyJE2qv96mXS
peiUjaN/NthkaA6PlrkaDVREc7YNJagpgZL4JZ4kcMaF5vttQ5mfdTO05nushiBpchUmouxMBuC2
1XDp/OJ2DYqdN1LBSb/hi3Z8LQ3hxCcmZD5hVM342GF9Q7jC/ccbYOdjtDXxUncNGOzXAULwgXAT
m7q96ZR79GXaV6e0F1OaRYkd8raJGuRoCJq16kf9EHdjXRRKkVepxPV5HawNYPsqI+V+l4qbapn2
0wTDTmQMlPhAWH8sQTRX1Cx125lI8AchnjKj7VwiN9pR8sCIAbttg6jAqjHNv0kT75M2TfbOU7x1
xlnewigLlcsf3/TkJQ/JLZ8Zxz8hUCa+8aHMLXgeuDbnkeOsAS5DaW+foSB6q0Svl8vyrzMbYpnu
/F2adp1Fg6avKpQB+40rmVJV+uCo1bm5gHPZBfVGVeaPk1E3LI1RNYbp1xEEecaLzeBmdmYNRYpb
uPxY/DdztjO+6Crxywg/4J8o2niq+K+DCLrtIyecEVOs1Z9mJ8q7tgWBG3ZQ8FZueFClT/r4H4jH
nYyF68Ej4fUY0dJ/rexmv6Gp4wVovqOGvn9DFk51rot0N4UbgG/UTMixpCJePqsRVrAY7bqZX2KE
fYOqC1oAFP5dobHk1BIMKJQ/CUsTfFhasVIOexxnS+z+2Hm9qa35aSx2JIPde8LIcZ0J0e2P6uLp
o9u7b2oN7xUZ2t6vsX2XpQhUI3C965xkQBiVD+PvyRuWbE3pIrEZ6guGnN8dm5JPRYF5ZS9RzmLp
6Iv4c/cNzG/uwPlDgFM5aZyTPBvTTcJc6Ftbh5DtY+sqCNO54rLhhTF+AmNsJXzT3k2e6tzX8wsz
oylOxjKYWRJ/zT+N7wf879f32k65ldjVXCuCQISEM6XkUxrfrZYaa9i5RCE3tF324qZQyPBVaGES
DVNeLBoAZRj/uJTNWP7V9zvp96JT56h1RBZbqJoq+1e0ltnBYgZ9FGcfgg0H7/NsXCmKYpxZNXQ5
t57WaH8UFGlcIf9nFWRScZMUZvPrPQTAlAUf1KPDjGCrp1tNIT9QDH15IHP83MMBTFGCPntcQ/Kp
CdwyKnw7u1oLRK8f9MZ9Faijv5+Ifx7r9iq7OcHg0aqPHfRr1D4OFINFcZe3HK8g4UTzZXBFLDpk
78/bKenBx3Aq0b6T3soWsf7ZTi37mhFPujqw8oNM8UcZ7DZiZGB8I+c0cp9C8rZlFW5/KZkJVmir
8hMy1q/06gyv5gYG24i8K+Q08jNgSJioac3uDtf4oVxFaUyXaV6rgUdY9LtSH3gTJ6uonQsuv2lX
HmE9f5NIVooh4GJGIBqc8ItIGuAgbiASE912QhVx31ZPnFGYBBubpMkEmmUo2TV5CRZR7Ic2fCHP
57j7p60OAKp9oCv/x7opHRHNpJXi6+827cPRu3mD9GY+8lNmTX2eO19KEGMpmBBV274uBLCr2Yqw
Tk6hl+mFF0M1ay+VmPgaoInyNKL05Cv8vx8h1THTfceaUtunwpNhNRw/ts6U054SVGXePQvc8gHc
QqsVu5uBxU9MOARZ/r+l0R2dafok3qUQ2Xk8z/3xuQL8sHTI4w6fCyAcvB7K4O5QNCF6nYbNqQNs
Gm2SoOtMdYGth1eU5oIxM4PoCJVrYcupLPJQY3b9tChoWvRgMq6pUiomF7Mg6sHREoo0kle8GIXT
N6o3TDRuRXFY0Qb0r5Bg+usNcvltORam+CYzRhlONZSckrRW2yM0gp8hmzFKlrqb+uDtZ9uPPE6v
wnFTVTXV7W6FfcLZfg4guvFNNsceBMq7hg2fHqfFP/qblaFxl6iKhql5+CNPxWTKSdU3b/ylTWG3
Pw2VmTKZ13BUvkU3sftBv3q8VtJwuRUyJO0wOCb7DwPKnfHPmUvg3deRW6YuJFIaWHtXym4VONDB
5lmBWD2FS9u9sY8QvM4dL8yES787H+mUliSwBw3owTlIBd9AJtu2UdGfSilGHZ2iDrtEgWseAWKc
mmqLdNzAbyo1nFsSYro3cPnsv9a6BEzlqFbbOf6ur9/9xep+1u3EXYdPUD2cBdFKRjGjQAdsF0cH
DlhufyuMYmrs/1NVMmwMubMFGtf/qKiYRDzxR/Rj3jYBFJg3Qh8TwVPO23Zd1LBPe3egl7J89LQS
HOS1dOvyZHJyW9Dell1LPWCd5XddJRiuDJTyMjwpHq7RBP7A4peu5hl0J3Obwar73+wHDBetmKEw
WDQnZRM+dVdbrx5Htbp/DiEYZOPw+33x3r61TnbivLc/5Nss35LJ0cyJOqWJHkcAYlIVfJ6pHvdG
GVDguSLpGWhMycirO7vflwpHZYQ05O0syzH302FyHFwCaQdxMuWDlNWeC03GoMzdnlWSl2mQsTYx
d2aLJrO+BiiPHrOqV6EVvfFmb5YaGO1IgZvw7rrt8aSz2qBD9clT//GfneoKVK4kueCgJ9YGXT2S
i/jEtgFY9S6muPXEFKMFSI2BfkSN9kcdsd816e5+gIPxANWRHca3dDSt9AaUJ36FzvQbb7b/ktJZ
SVXvJYF5UmVgRxXNqlANqneINLaErBx07BkPW5bRusjL/zASOmVKR6ie18rX20QZKdRovQJ4fzq8
PuhTKug3h24c/t3bkH37pbDFUOcIi//ECNjh5npNdYWjlCefPbTVBWLk9MujNLlUMuQFPb06NCfH
TJ/LMgKu6pOYs3ndtoZYMLcs+JGiitxUO2WwGwCIC1NI4MUcsF9h1LucQM4mYYhqCDzVccjnFJip
1u43m7xzOjyeIFWXDdjY9yDJ8XJYYgc8p4ryvCZfp8PGplsR5JOyO34bSIk3zIAvYrXGEPBHZA54
5hOTW5JFOIzz3eJMAggP3DnBxZFmUW/bHbsyUg4zb5J8dvpQYu/eESuxodcNNNrX8kj0iYxZJgAH
np0MK3WzOAVfh/lS8JUh2DCRyOzcoBlUcAXEnrS+D/tq8W3n3xCL7eDODsBrtxD1BkLsQrcfr1d7
HbSwPYZGBIk7JX6byjOhbyxQ8on5k7/P5hpq1jzieAQnqfhD5uvwwmnwLhgZ3ZQQJqLwqnv3krp9
lJkTF1tGrpF0t9RSLOoCBD4wx4XDOVHkPKobiO8J/8XT2wXJz6e11ElR9k8z/jDQnLQWD1xHhROL
ThC1xaHMoJcHy5G/S7eHRuZwNSh2K9FQY80roxIlG6Pp2mDQeNhW6TnXdezntlgWOEBXDqpL5esS
ygDji/2zyePbx1oscUC1Ka2ZfeU24KJRFENyFMBxLOITbobf0OO/pk8dM8AD84mIdPy7LB+0UCNW
++Fy9HZ++y3jkDYlueXkPuFhW4vMxA7X3TcFZoRImx2+m4dGGpM9AMt8djfKXhMgzh331aZDflY4
6/7zSSo53ihVQ2om1jPcsozKo6gbFEBRZu+VdJ/fgq9IiOVRkB2IWlH7/rhWnAYzeQ5gv9q15Sxm
2iOEJ8roE0+f5MQwt8pqAmw+aSvS0eSeMyRUkYbBn1xJgbOZ1HkG6J0WPn+yb3tuKCEVsM8xesC6
S6zzRFGLiR0xRCir22OtkNlkFznDi0IO9tNEKktadasF4ozM84kWVTfCDLsVEO2Hg3A0cZQufBpt
Xo3thawtCtGV+8kq+ZU/roGbn5g+7Zt0ppJbbujfU1QQcX0Vr9f/spcZyKx+VYh/bI903QZBdNHW
ZFd4kEgrCEdjZqIBMxmG8oezxyR3/PmLi2oCr6X5rOPpXQ5IOCdUym7qw8vOhpczteefgBu2lqwY
EEFhEJNtk2U2quW9cDk3FdeWRoqcdpsjxOgqZdZ1QNR6SmkIB/SUUHzEVzYF5gC3tNdek3tLNKx0
cBrIxxxt0EndD9IlA5OmgAUWSMocqOw+9qssIapRd6FLoQRYzwwwXFR/yo557bh+kego/v06/65R
rNiLBsBiaim2hEeNq/1Ke5QsaHhKLwaHclUAXMUU0cADOzt14i7752xzAWTEzd7VdurKVYVHgsko
P6PRMj6Xu45rvbS9aPygD+csEBVbgRec+JywKM91ZAOy+q8uUaoM9XnTrg+zE4v+U1a/MC8oKQj2
Rlx0GNmgq08m2Fw+pwQmfz0Smer6bWPBUcShpT9vEI7fsc6hxTT0fYQ3SpeRu8lb/y4ZlSYV6xaR
ni/cbNQyuNjsMMuDx6WpfbBr5BWS4sD/z2rYeOTlV5MIXwkE8DQ8WdpuFuTOacXzfOmuvMz6ElF0
0K1hIw80/wi1HxiZp2DJRdoLAG3A0with7bxD0Q850QU2uCasBZBqwRei0dmmzxd+I34pzhHSp5v
vhh8aQhAXOcuw72AEiC8k/ZqYMR1zHBuwG2l8E00uT0W1q5SJKV67f3xQfbgjFQqB6XekxsXbZrH
vtxYGOi5+e759xGlavZ/gnklV93eF06ku5NNhiIoLAsfvl0WGVmkPhk8TCA66gU5JFfWkfg1+bZe
fCYNM9ANLQydnjYuoC7pkdB0vamVefss1XmWOx1GpV2UiURxawW0UzYoyy2kTo1pVJgvJCufcErN
/HZNaB51hDKnE6dbnOEGJQ5+fXuFkWflCF0oIIZNwOAc5Ue5A99OPpqMSzmH7tvXvDpj6pmNo/0X
yTDmGT/9MjNGwA1/rC5jRAuqAJtLAPSi00dZ1Gd0B0V0rnb9CmrdmbliI8lQIzeUWfu+HOjP37cu
9ML40LA9MtZ7Qjklb0U9So7BIXJ2nIkFLH5ixvktgIj/SsJ/XB879DBMk8cc5LrmD6zMI77pD8nY
EahsUyL71pluhYuuh3O1wvHyTX0l89S9mseQJ44FdjSzGjdZPmkTQkXzZpXYvwrlHdgCuf+AzdiY
g1roZhabmSs5W/LIjS4ADX7LqCDux0xJ4kQH17mqggGcKjn5dAS+BnGUvaI+ldHe6J63lgNDZuld
B1CuRb3CdkMTxrRJWfvDFxza5HDB+b1ALp6lGZdOlGoCxrvFbtQzFORCHem8bnJWkQdEEBABVfCp
41Nwb9yLc3cMzwc4arYLiU3xql83aJq9sfFndeuN7V+8d4pZTJNELl8eE47H/2BSitzFaU5xbwVh
TsrTnw5w6aTECI+Sx8dUsl+jfIbQjGoQfhccMcgevwZbxSrhdFdrI2BCB/0jbsNB36w9Ty/lbJJO
2f0Vy9Cmz6SrKTVp1yReA4IUfWOhI2L0fWUU0M9J+67kpXkSvPgEZGX3NRb55+Cnp3tf0sEtutHQ
aefFXpRsoxAmlzEE7OGTj/zPlR/8xAoToycY9gis5vZm9P5QEbTvDD1VeWuTBrzNBhQiZZ+NvH6b
/oUpKIs76cm+rqAvhDg0MXysCDm8wpM728sRG6/EVRqZtZE6Gz6xrpHoZHyyHkMvQKRPdM40MlZH
G2W4+4PgKRl1w0WVFVRR7rjvH/nxEmB+U80GauRDal8ZhpPLBWhuZBvgi3AFdSd3f01iIaAUNace
vThMIUeibKo7Csth6R+1Dtu7E7Dx2jYxyZmd52vzcGfUCgISn8yMTzpr0LJN/GTjDjSH9GSDPjnD
saj3M90d3Ma7xMy/Mzym0QavLSIvuZNR2YVPIFx1AXS1mDB84GDTZNnedVEEJ1VNxAfvVPYbaQFn
j4tf7VQyE6XXOcNtwE/sr+hHLRDSyrue6Mnbp/Shpz8oU5ZQusst1oh6vncC69MeBtjv+5Z5iTpV
f7eG2lsEQSm4YFBElsFqfHlQvHsnaEhGETkjdSbCO+44B68LVEWlSo7pSms2g1cwfOsiGTPR00Dm
cQSGC8sE3omM2zldCozTWWslZGQWxSvH/n44vjmzR/dSC4FK0pns+ex4dXI7QNGDUPDB/VXPI12G
GrS7awWiPDt9ka6aWUTj/yU2UmD+/DSRHCdHMljiY8QwSVnWxHCJI5FV/5zpFhDojui+kn2CYsXT
sbhhqyAa6glv1KEhLdlL63fXTFygMSyzqaM054V36UMqRYiOo17A/a3SrfhsFPS+xscfw0aNpUEj
/M/UhZ257VmhdgKXN/E7G8qqetvWohlmK1kwVkMr55p2FS8UMb6y2OOe2PCn6lDpq2K3y5T7M0fv
VKJXXz9oMLjArA5Iqn7oyzHFali/xULxluIOYTB2JGHXBRv4IWpvsN5pE48m9jkjXcqQfEM9DAtB
6JxpPFhGZq/WT2xAVJCiBn1sGSp2paLuvx2/QOwFFIMyQdYWx1kAupIs1V4UIi9GDv9ci8AssJeo
r814Ou2MnELdhM5Dqt2yxVgUg7H5NpEyS0uRZWdKsi10MiS7dYhv+5RWbPQIXERZFBBFiG48F5Ze
2R83mdQYr+36gfrAh3upe7WJynLPl6rdhceL9KStOTK7s/nmwfrTvPHFwQTnANxfHt4ZXOSVgNob
xqj0TY5RzeAF4rOGvSsWrD7Idyh2IgT6TQl0h48sKkKYr1NWV2v9UD4uZ0ZS1ON+MJFRUW/dsFHf
7TVIfTi44v4gsTU6XLa/kaV+Qu+aQHyQCVxXcrEsb01mfAX20/Kx6LtLmzeLqmIaqaR33yiOB4H8
cXafosd1Sklp1EJVtbaDUiGjQWNysc8OMGMlB3KzY/V5RDu27WDqCBmTr2wKNAgiv51AI/pAWsN8
n76R9GaqDuSDPUJMOFzBQRnez0HZiKICNMveSXUJJSEeQglVklT3o+m/vRSTZYDP+lL2ANW89bn8
l580ZutIDMFIiq/QJeJfuavYZvpQmYTWt0ZSeAUHvBL04twzS7WJSCOr2+uCp+WGOIqr+YM9HO9q
tZmuU65zGAGKX2ecsVSTIvppIjDT1K+zBgPjN0BbVaq8ZiFKvQAUKiFtAFOyv+uoJG423hWuVzmj
UovC96dvVNAJN4Z9ivKa9BK+/gXmTnKItdPm4fhq1Fm6kOwrd1meNmuqy4MvFSDd2ZuL2SWUYIoD
oSm5JfBcuIOfdvprsGXvBcqt8nYxXnE8fnTUkKTOso1pG84QWYAPjtTi8A+/R2tFSCCM1uPyrv+n
bltNYyhWTbplj8xZGKUCuZdPedfyy/gCX0dlqMhgAUpS1i3lFjz+5XaU2jHcqz1EzPZizN4s668O
lJQZo692yC+/1HCuGxSfqjKGofgUYPHMj+3hI4iMAeaUu74Y830kkXF1esCBU/pcp78NO12Ch5yi
6n7t3xTYgSLe0W3DLzU8UwupESjKa3mKrdQGvXjt0UjUTAch9DUYA2+wsSLftDc+LNbHdFdKiq+Q
GYoyQvbKvFzI/JgTLsw8RAlZXsJvsbeOr+LgcIvkCYp0JlkBWPBbbg7B9ptykhXr9L1rpORbAv5B
EoxMhufivm4ZHCSBrnNOM9JeHy1f9Qk6WvhGGYYfrFK0udCA+k6rhmv9Nav3P/lepS9SkuG5WPCF
i7zfoKG4ifbI2Zhetk6kJh9pW41Xwzyhddrilw0xhY9vZX0C5sBcd0GHgl4oAT5d3i7TF1Rxe/yU
I1NUn35zipZSNS/A9M+CxKarGFYeoyLxITarP8rkidefIsya8x7A3TI/YY+yUu8k9fziXeOQQ5An
kXnK6slCV7ocPk2+IsqykuYhrW/ZD2J/nDmUIt0Y5HtqfvbUC5+KQWExwzlSfHtFn9atlzcNBQPL
CtGCNpWwUBLCuDdmw4lEoxQ8cKPmUUWOHK9jIP9fGTFXdXhffiwOH0n9bU2ifGB+UoGDGhf9H7JM
kaXjZ9fdfZDs5XZieWak5MS2UuGzqPXm3zoS2JcX0JjcHnn9YbOQhSK3S3LRC2a2AzUJhIFIuKl9
lvZ8+te5lFWP4HDTDQpAeVUu28NxrzIYACNEBhk1/89hbnXKLqIA0YLz8lqzf0s1+1+iPCXGYPcg
q+tUGkkdzfNTXCZAk3hyzcKpNyi+FIsdK4fyPx+6Vd7RV7ciedcqeTjLUsJNONBP61MXZ4GwsMhS
ZJ4YeVQzJWm/HVrGwEMbTJIh162CP9k1LK8EyWU0BC1hswgm1hDeUTvJvbL8TIPWvfZjErk7y32s
Pc5lOX/QsxyDIU0vLFcJQXFgVZcS03CT9uo/yPqXpVDsf/OD7Ov7s4WAcoLG8kxLw5/zMIkHOhl6
EYvkyPJ1lmezERV6q4P8wfZ5beGGj2DGRhyUhJdA584oiDoBqYryW+U0zCI2myHIudausyo3yBgo
fynvIqg4HboL1+auOvZh1ykZukM6LJMxyoRM0Fb/jnT84P8xXWlguKE4NqEfRJqqn0qONmARDFSQ
FErYPhOfZor/fDjgWtStkSMCz379t66X61unpGmYwY14jJuKTpeeASqsV+l28axcli05j/6XC/Tx
OIIFKRA9vcW0yl1Xt5gi8cc+n8co+J9exN4e/BBBYaA7Q8iWVXOuZ5AGcOaykQ/RPsqshTGoCyLq
b9xoD5x40KNfSBIM0mSfCArSE6Jgd3snx7oGqZCADYsxhoZibo1wZ+vOl95eFxHLflkNW7ySqVvD
uhYzQgaNEJ+kc3UZZOKiswZnGov6Sg9JpABFkzSb7NvTexzFE8gpLNR5cmnX5F6fzizT2AG5QWHL
sfRIFFHRVz4ymHcH6Gi9qBzOfgQ3kqL0nd2fZC4QcTmSzA7+V/x6IZ5gRRHK7jbA4Ae4MDtW1nRx
MiuB3xTykT5pWqky05bPMEtq0wMfdS9SDmbIqIXpbqdAz8tZYx5kqF/yRFqrBVt35WNt/Bky2QvW
t1xW6UQ2kUigDUgijleJnauqeIw8OK0FFfXYktFhhwKmMFelC6r3nr/DPNSjbQb6hytDXIUE6QoA
7T4dWQi7JypdUJ+E0PdDR7m28K0ScZZ7c4dcnvxYdMpX6pOqAoTt/jsOBTvZE7FZYsQwxqYXSWcQ
yJva/EC0C9ZBuspoxBfML6ovahrtstEJqE55LiK7IIAfgyvJCH2CtNSVNG2iuaEPbKVLkiS6t10p
UhB+KYxYVV6wQ/7RugsbfXfm3dMcShYAjMNOLwekZkCPnguWeKFXt/2zdfjDNgYmqtQvLLB4Yjnc
gWIN/hUEnY4/mMa+F5/GZuHhUbS1jGNcIEWxINn4g1ewInTUt48ZZza+V07VA8M/paZkCghINAhs
iqyvrgL8IEdJri9noNNW6Uit36my+tZjt1Ju+5U/aGjJ2maaco6dx0LIN+H5XkiNOLbBZCfr9/4F
WT92i8AOdyQBGsYmN3V0of7/TI1nAbkVzKgTbhKjjNQec214fiy/Go4VvWq26h7g6iRvAW0HFuyL
9l8XFAkZ2EneFIcsH6Fo9u97kkm4FV50Uvsud7yP51DO9gE2dH/HF1cMahLpvOPRViX8p3OA45nA
Lgom31Yj0QFDEnFQlTnWZB7/725uspEcR+8LRWic1hSnJ0H6HW+xD6xnxk8z86EbgwEIN8q32bLl
8qSHdT9pHB4vj9ndKwu0gZMwup0QjAMfAOP8btQmH3r9viNAhpCJHkTMJOurvZ/yF4y9wY0nyWJb
slz92NhO743HDo1fvu4iejb4UYelIMXDAodeNznRRrqEsnRuu8NRnQDRHN6NVlbGLgIXFodvRxk+
lwuhNEnJx0mpNlzPqFfCRuTeOl+3g0FR0WkpzMGICbkHgZlA4eNVJZBjZ8tzw3WvxIji2qVj31VF
/LSoAgSvqBWJpe2smbHjsSd4I6ubvLISLGAF3tuzwkEiQpmJXXTFHSHFo4cTkCTC0ngj5q9NpLPT
AsgUC/iPPI9ok8CoMqxMQDT13w2jDQSNGV4KKE1x1KC/IyeWrrxXeAvwhTtSWv0l64pz0ZnXZJOf
EEuqsNJkJMaj6zfdzqE6bTiGMezhXwdsDinBDFg4Tz3Kv4o5jUEf5K5RpRKt/fw9rMeVsNNDhLL5
q+qoYS4+W3b1qwRRfndPBEVQMgzk0LPL0k4ASsrOONBhTvuJ8Pbd/+xo7ijd4ZGmzAt9Z/kmr6b7
YWWYO92DjozOLAWqCeyh0NeUkNblGZaVlhYgdGiNWkqHNO8Na76YaDvY+JmdDzjlVLEo0dh6XgdE
2aS4chTpvgQqK7FcyZNQdcifPV5w28WR1RY/rctvNYdnOdr4hXvf8S/tPQcIBCUaz/7DjcAkegli
S8jIcGQdbOp78qMBQ3tuB2Re+n9i4qNWwSSYcRov1T3OeBQDEm/gUSWldJXqc4naQwuu8pwGfe74
YCYvtfCqvqjcY62/GipqDsAQnwjWin4p6W5p7uHCy0mWW+sypCzkZTXPpY+xtkzzcETi7g9HIDfq
lL//hTzvVHtcHrW9HXGJL7vONukLKK6QEzV6TmCdjBUs9/RWu3oCorQ9encfy5SKphpwqZSm77Tb
mceaD1Dzzh/Q4p7rNhOaYqnnvAtWqOqYK6c3j0rgMQUj7KDj1QaROKHjYQrsUv8Yzdv5X/oTgrd4
81OX2vGnBrRAswb5G+CvjhCCJfP5Bn2SD7/oM+urC3DWGrZPzavF31QtVltCZhTuEdX+iFIZ7wCE
1WK18WwXahdMO2Mwbsu1O3qXr3igCvGx1GRMZnr1p2yqFTSbik+XCHtp2+7h9TB/hoogVaWs/38V
zXSvovPrfbxUzkUvMslIRFFyPtUXb21VE/WUbAoIXsFnnYBrHyUCbcE92M3mEkPFqQZC4vH3v2op
JZebdxqeexB5sB5aDHxWosSUs7+YLDQxkc7H0PtW5bFnAk9+P4eW+c8Eyn1JdsI33JS3zqcVHtQt
tUgtiS8rqmk8VedVtR/dRMrcFsRuuP3GWQFF3zpQAGmQg64AXSKMmybjg5Lv6M+1UHHzrAbGKehP
kZd/LjF73DImAMrTVT43wF+cL5vZHEVa77p90y9yXTREeud8nGigqRJFaItK6+uf3fb4JrPR0Q9/
f8mhXqvu8ml+n+5DusrPoSERLTdShTvjc8HEIrWivezbJ0VGYi4f3tfNxxTS6pxrskVCr7ZnOtiz
LcztFpjHgHUycXtcmVumEQqeZ8ywsc+IkTA+zx/4na1AXVGOIueo8jeUhZFOnALx7tPVOb5IPrDC
bxPKHB12jXWsShkdDo6RfmWOflBfkBoR/UcWV4cApDJzQnCEyC94jLikDy2xpjHeLFpvkUDRMbg2
1Cu9Yb5S3QUUDZG2CG6pWxHVtXRMQT0bTOlmr6SHuHwlO61ut8nCv0y4wMDo3U33uHSpx3csbjFV
W6Z+mo7yTYaakgy7HIRu2VQ6eE6kir7OP5mXntZkXrUyUQD/Kv+TIwzSiOS86LkxzkEaOVbJBInP
d0Bgc3Yx95IUGtQzNfskB8y1gH4LpYxygOWzoaxPOGJFWWnhJijNvaj9+BIuzlkfTCuPIU3nyLyF
m7k5+jLBG0t5I/8vxkJ+4sjqzQc8SaI61mJJ0szolrujsVp1guqnd4b8KnuIDJibwmyc2GCoKH1D
LggBvANrN6dFit8ZBzRMbtaNaZldCMto3HnC9lqSuf5LldDjKfYUVlUxPhN49ljFWGG4imsqCFYQ
z1d8yQxqLwV3RRzqk2WK2/0H0WUD6lNZZ9aTBxDeY+ESC8NoiHFUfw7r7nvbnGPx/sxZrA27sbQ6
wuSAH1LWhR6kWpIcbRrcJMepseWCPY7csIQ9T/Rm3QZ29MXlxZxQFqVVu9MIUcfL1Fdb8OF9hGY2
rsnMYSvjNi0FPphgPEG7g5KMo+1jLgosHLXbIh3e2T+2OpUYYo/KYcQoPyPk53X7aG35IoKU23U/
f1D25dEUq2S442d4Xctu0jIL0y0x3h69PfmEtdg7cAQUmjI6S66Yh57mTRs1VRjBEZlbEU39ST7V
3LlSwyNJ1b97nKjQQCEWJ/j3/MtiAc8HGOVnR1Tb2wjhDx/gG711XZQ33oYmlhWwc031rljB2E+W
rgCBkeHvnoEsmNUNizKVzZsMTyQwOAZHJG2ytZumvV3Tjh6bwTf1kJfpw1TnA4avMaEAKa2SWZeJ
XMegr5NzLGlvTZ+lktjHJVJ49xtpGtSIsH4FbH8F1JWnEnvkcSAYI0k3FASat2/BZQ7+YBALWY02
xwLfDpWvbIYalSr1m80rLt2MWU4w3WQg9XDItgs1YO5Qud+ISySTGtzbFl2yD//UhRhNdEBP/BTo
fg+4AY+WXvKAKY5nOwY1f9SlVXlj+6z0LQn1Q0GL8bENyH238Lw4l6qBJ+6Q7OmNIAoBL3HmiyKv
iH1/0Lvd+EQEE+KA3DhZEkFnWID8WSraQkOz4fqCx3rEBwiSBAWs1yiEwkyHpo1HWYAVz9nN/xmT
iWfAT80Rsy6s+iBPAG1U5KrBjHLv/nNE2pndJcLkYoYZ1uo1DI7a3NxGnUBIi+OqxTVw3OAHX1hm
MEvbrFyHVcXnusGIcDHkrKjozaMIIcrFiBWkTIvFKwPfomBUDly96EaGBtcMM1xabWrd48niHvBA
QcIbVC0dFhJZ36Rh/QJd4I/Xjd7gEz2WSmCryRSwZZddVBxlLozNZHMg7bGfmOC3hZ5ssCYw6cjX
D8m7cFcBx3aSbmT1dyKKepdWLiPZxXdjLVDee1DFz3GQUsFTnyaq392caxxcwGvcFjfogkLzF82q
l0IXHvMGak0Bxr9D2x3SGFOdh6TxylK6jrUbunLy1WszsiAjebcKcLUGuEVPfwgqsJmLKo3yqW4/
0nYXc1BytXF9xNAutSkSbKYeEvKlbwdOmc1i1HQHMhOg6nakj5WyaUh/lKr8YKzJfsiAHppXHR3Z
mHo3nNnoJPLiN3qNfs6QPHHvFjQmH47l4mxestsEKkzEerlNZaaL8KJImpQQTRBQtLftWe9NhWdW
IBqfCLE8ttXFaAh5jQfNb4DiVl+Doi8Ts4W5zo8AZH9Ob2hlbYkaOUrBkgWb8h/GLMnT+iH81iVH
FXSMGFg4U0TOkzN9feDC9shxFcxl/Q1ynZDu17t34TS9Iym8m+prmudI7lNuehFfnwdgIV/IEE6O
WwiU4eQDAL7FLEe4samufflDzwMRke0ZfXka9FRNOZd0LFKJgEoRIplzriWRy0DiCiQdBPIjrvN2
MawblLNUWEKsHgmQqX9S3hgXFielGmnTLR1RN16xAV1OEpm3IZG6/XG3Jju6JBHF/UrrSe7WKNBU
F/J1alJ61A11Dc0eJ56ETNwK3LyzMn61sXSPgdLPw53MzEsG4NoemJxbue2MAqbbS9rI30UBaMT6
vVyOFbakaE1mj6OgFRE/Vwq+J/m0DjOHoDkU0FFhoRjiBcZKdJgK7TkKEQ9RNhsFXTgE9cNC2R3V
91vksbNlHX0joiC/exX+tGv9ahinByN7lBqrMh9aZYUb0ibPNwBHPLU5M60qBZGN7Sdp3o5oC1YV
NVerbIC/Bmhb2XE1r//ieoPJv8TQDJ454oglXa2Nsd3iI8QvSV6MGPXzvLywq8C8a6QNrr+Z5Ljy
SfITvLv2rKB+GOHNdRKOZYwWUwLRpSutwWEKjPoOEWcma2iV7GZCUqTYOLmO/Bya4+7tXzCL/6cX
Ks5dbN76Kg3FZ0VoiX8/IC6gH+0Cz8B2VhX5mnMsKr2OxxPVVPvF3LtqjK8D4Bjt6d4KXaZ5xUhp
Xt/3CexUXZ3omYFnJyYArYHhVtWyUPTxaRdTbN79IvA5U9N1mGx6fTBk1LpevBYXSsSDn9HNcMV4
F6g1Djtn0anQqvjdPtouiQ3/4vxg95XM0v3KlARkn5HguW0WuKaTpg+4AgidXLjfzeWZOAqP+CgU
/hcZECYallGjQ2WW5JlCvn/JBpvwlpZ5Q0CAge+LwKT20RGY9JolCHexaQRG8VohOKzmUKdwula7
ro31SFXNa+UXm5R1zFx2MyA78SB/Imjft8tbZqErK+vW1rJ6DQmoAw17jVe+FTSt2gtewKRUX35U
3ffsQ4ZLfrEiFcGGhOMYvo+J+eAIv53KwF6ixg9HQt1IfNweWEG3RTx91EGq0LSJH/jtMjQwLdot
6AjyfR6oARYRzhdbt9JyyKFx1iOvrwU8Rww4s7laig7uGq0ESu2q6a6QjTbDiijRYiQLFELZqURR
qY/ELP/eQ1XjIEOgkVTNrF586tztvnNKerve+PTBv6mcVk9R0yOYHsIi0VJ5sFaQJI/MK24aEPaN
Q05V2LGSDRrrNIxzHQaO932HUyt/4ouF6nasdRy7FLsjeAsM1DuwSMcirMPWombSadE8bgawdmsk
sHGn0wX1rt1lApZUZYptEVdxmtDGKFTEKCokHuBtRO4+u2Wj010iOsDXi059vENsL7n2DWBT8jye
TXfxeOSnjxU/fezZRMhFgzzfuDXiFK/jTTzlJHEXOXuQ9jWPrl+jj9KK4USEd07y2DVgIVN0/3M3
2BOWzdvjRnQAffAkrRb/iQ85GmECWlG8qb5xY65vZ6yZyBpeR4wqkfXZbZIyCzTUbOp3sm7dYSaA
58WCqDSo4jj2zJkZBiTFwOmHajm44Jg2WSt5rb+2vzg0kfF3XT3Kzh6I/cIEu1KHZqlX4VG51e7w
978UWmDP9B+576NQQdSZbgslj+MSnU2uWcngSX59fFVhzcWTbLmoxd0OQFFZRZZKPPkeNt1keFLN
H01qyLEieX31mQI5tJYk+n0kiGMWoHAR35WvBpkJtxF6doomrOABA/PVcibUKZ/dS+gXQWBcFFU6
HNvKe5x7O3mfr0YDT7o5r3b83DIrawgFIMryY1VaGyB5vBe2NbDS/OfLujOEX24A03ZHnJdZDra6
Vk2csUfcnRwTy1/LANXL0TK25IDHu2Da/s2Ht+km3FRhLjcJA+7QIecQvXB0LmuPfEHmfAHURpwD
rIwRt0XSMIe0d6R7wXy02WYCNLSW2spSX9vqIoOIufgdNSam6XwW1RoDhhWYpi8bIQpdeoV4yuR6
o1lO3SNbxQduFT4zMkOcuCLaqtki5bKttD1GMTWvQ755Kht2CThCpuJgrr+tu/tU/YCnJpOZ9ISj
83BJNhRYkd5F/ZsT39wjkZ7B8rkK1I8dURD1ueDc9j9pCk2i1pncjHl6GvXlkeCgIO3lHx47b3rM
MzXcFDu9eA3/nhItXmkWc9BvgNned7WsrBSPwad2SoajpUCKTvIu6DakEWMsPNIx7d3+brTABFrw
gZ1+y7TNShMREVWBvPRdEprFVtnHCCRVsrJqHjSuC6nRWlJQytQjH/fvBMLWVPW8IFAA2klmUXj3
gw4kbEYJoYCHsuxf2qSuLWZjeWe4HMtrFATFqZ9zUe5PZ7y3n8emSV/qY0pFDu9j6oZVcc0g/vlr
xJHqudSuNmP3SyRfvnDmhw6027rP+SQLpDd3cMEHUNOXLKqGHPC+5CsVGaPWHsAOnzMan1MeP9Dd
kbQIk8Lx3aeUq4Yq7RfRm7WQlCJmXHftRI1xM0pGxYkhmJHHz/2eYKyr8YEHI9XBIt9Wzk7zdCsO
DE5eJ6AFyIIFx/tEiPBbdfJuwz7Ez59WdykqKbeMntMo9Jw5oSo8vLXTVtnMpwIj1LdOIBlAtUu+
WTK+WsS7rPMo2pmeixhFEefwtW2+ZTRr4kmJuBYmU86mtGZfB4mmiSb2ZonAFcgimai2VcEei65Q
WuJATc9Hr2Da3ibsnQlhDf4aw5Vpa8AUlMDWBT0pW4VGVZpiw6uJujLVSVboTVyMHpDlnbJGTCso
95WPHLMDDeSKafmYbnPKdlhTHikXTP8dcbGAPvQZ88t411fYNpfrgtFJv727OW31+PdX4WhsbCwd
h3gacvfiNcw2/hIW0aR2SJRSHf3kWkjrvzYWDIbzIQI1HifW4O5J2uTzVG2V+x40ZiKMFhJN92tv
77wD5iIl5KEt/vFuMw7kM9pI9OlbnNLBSUJePiOgUCp+iTysjSMTsdKRgC+XtfXzkagiHCnMzIP0
TxIUNGXQkeCWVnju4Xny6BCP/NZBsUz0oyZNVegz8XnIdkGub6ie30PQR07pQdI2XfA+PwFmMWvj
9xfd57S27D6bonH5ma8dR+t1kZX4OKvS+pbyiRkd4ftjM6bP5kzIgmyq+idwPdfZgflhv0m4bZoV
Oq7Y6lSzl5NeKICjk8VGrBS2n6+PwzwjyWyukyAuYWbgiRDmcfI5VpZCOP+uB7wtR1sIq6Y49OJQ
5l/hFW9ody9AH+KRckZ6gYJpXZePPj4yBSygbEnRRjGKsP1OujccvY1k75wREBgfTFmdGX7uExqY
9krv8phA5xRqjdLxaaPZYcfteFYizbvO5nEffpV7eS2BgbZonR7SmZin1MZLsBT+heBBFBaHvpl5
xOkasqKyfuMFdM3a2GwasO5HGnKxgP4HCRrUy6N/68yK85RRHDHZ670M23PSdT4xwuNI81/EaMRA
RPfaRh/TPyC3J8EHiGFL8p+phE73H/yI/rzTc0qhfZs14O0TAEKMtrJrakD6Ua0cn83Ccr2hjX1X
XTXeNjVT7D1hP/qhdTZ3g4DixrGEexW8SfqXpE8l2UMG9AP6QNR5yybe4qY6shgbEfWnTrsmasTg
nABcbk+Y9YNyAtWnfckhS0MbYBq9EEd6EzU0MQbjEuU9dqQFg5dn+Hs8ff8DwMxoAyW22J1im945
rM0x8G7zgv5iZg0ZGmSfZohRjIRi3g0qtIY3MQCFKwvHgG9w1pz1tD72XPX+OoWAuk+Ost7u+ZTl
ZWJByP3xUH7NudZQYxfCTnUPfMcwNC9pICJw0td3g8818FOEWBvZhwKeJB04OXDchFGGh7HpXCQw
a2bVYy7WiNRsFBiSzPruXIaVf9MnB6cUaSyFeWH+mWNRM5MReLAl7SPLBg0+O2rAijc/P+0hy2A0
6Quj43t7OnS7zMh+lPCIbnRJzXZ3pkxaGQ/qTlGsZ0trrqXVB+OuilRziH2NtcqfSaDMnngeZgNm
AaTmBvSnwuX7GQXZrMkL78N2su6HJD5uAmXFKjJQx23FYx84yk3jaCHntrEmAIbeCu/jqzxwziJr
zE8ciTmXDQL1EiT7sBz4WmupKoNvh/VsPo3RuekaNZbmqJkNRubrfIs01udSuy1Ty4Et+FKDLTyh
Vp+kfQJbJcJkdRDkjkBKdVUfo9ephzfRJi1YQUqt8XBIyL/w5jEhqBQVpRf561oytqTnVgJrxt3z
wZudTkCnA3hXL3takPOFnJRIMAJ0FVGDiJAj/U+srmsllsTnOownJpp/phqZHAVG4TkFZnP7ZHPX
JNqN277t2dM8ciZ3qYBlIKR++hv4+RGMr6acg2u/yncYWPqdA6KdJrmjW2e6xpE5j25fsAYjgfuU
fbGxiryEe55h6MlxMNgAqD0MgdypZZyhipGMlOzb2Oc0LGptbgv1fCfXfZdFRR0hmT5OpyUMsOPt
IXbhkggYVxGZU++Q+A1vM0hD1rfFP3Wp0BjeEZiTDAMH8BTcZLSRgzByjatLMsxQ+/GFXDQeF32S
YEu9L64ec+Z1RrTC+q+uYgsHWOIn8SQDPcG2EcsSy0BCZZ17lo/7J1COZBvHd0fklrY7l5WUmbyC
zxteVP8pHP1jeTiuDuQZDAYWSwCeWD/iuMgblXgN5Evaj+FxXm2j5lpNrUWwkdhFSBkmcFhlziSp
ezeTQeLcg8naFmS2faDxqg77gerX5AKR2UOi9A1NPcTMJkoGoAPU51PPX34LvYkrvIp+c1fxB2sD
5/a2vptOV5yGeVSiVVaBvmQxVhA6JwDEOKnYKZYekidHd+P81QUdHvJNNY5Do9Bo5QnCf5TVRVr7
lbO4c87pjmxbPQSDJg5aydRadT6zZQEhGP4I9BVo5/h05z1nuRbySm1Xl/axWqpfLtT+7721Kw0H
WlKEupR1oI+7C0XLIYwN9GGwgMa7MwPbm+BJP8JzO/CwAwzbkPupkzxgwf2rudTqVuSc4MFMY6FP
L9g4RPRbcN3jjg6g4qPQbvC+d9NJ0mA3MH9JHr0GQx1NhxvHyi+AxiZT+WckbatEkBqw3lYgl3/Y
JuFlGuWK5CcwIiWotmnRboPGHglli5wgnCBrXW3KAsm+Liyo6VVLKVDQZlp/svJL7SQDDanqcmhF
zQPel9i7XEMSKwjUyvv2L40tGEcYCcV6GAS7zC46WyIMefLvmCZTyYJm1NpxMTPBnmpdBjGKzV7M
ivKsSl7dwJGODSf3U2FDHEbqYSGA2R1DBVqYtWrT/evAGUEd7eafiU1QOMc+DLMruLB9i+NHzOHS
GpXpUjQiBkOAfX6EkOvTU7lmKp5BhJEJeuIAVn/Tq2OTjnVO06xvMpqzM7MZRPBKoYaLhafpaMus
+pgShnae8SBF7PQHPds9HOuVUHVp2daj6BSCEkFd+6cTkzwvu1ZLAdCnBHR/85b2Jq/TiReyNOGt
SYYNeeIWweizqCFf29sUMRC6xYGn/u4vM/2re0jt4WRFWmYbcFNo87bz+WxmI4yb98Hjw1I3VXXG
ru1YLkq2tJBLKe2eEe5IIWq/0Rwq8UN3s8DH0ZGjCRLMlAUOIz0Dd15iHSQEccRJv2M0qc+DiDeo
W+Ds1PDICnV6Rs5zKSvrCN6nq10U3TFbO8MkHRB4DxuRK7TnrgBoc2nMHEekLUhGYdhwE9uNw0bZ
aq+D202Zc96EeQdFXDrBdyesJDRHEDqTPcp0juwAOgL2IzBq2gLsp4Mz5ivpTLOKGaoAy9faKue8
U77KCAD9zRlrOZwnkZfZFUkj2CovS7JIWM6xS1RZnAPty/66spyn6PMjtU/CPvxMFvFVIEq/i6ug
+cg4BO9vg6AmeePQxN3zQss/EVapT740tWAes7Ima0mgcwhQmPSTGZJWOdGYLvOLwXB8HAl1pP9C
dGmsg1Dfusur5Tj9fXIzPaa6WcdyMcNte3UVa/CzWumvHtHUFNPoyRNFCzPJCZqXeVX1A5cuNV3l
/eqZ/cyCRgxshYeR0YP6MHdEpYYEN6jXKUBiUWHvmff1z6aS5ABiLNVS1kSBH8Xxqu1bltHzxKL4
rE0ccBxlvHogSijPnAZMdaM/3p3If/xA9YVzIalLJkGA7UU+NyS0PnvSH2xLeQyav4YKc0Uqez6n
bfPpkjrZC92+nXufmVpN8KGvUfAqScVmTp0qBtruFszjp2sXaM6Vd1gPx8SlS0yfHTiz8+t6sQ86
eQRqyQxuVXYJ/zhbiC6zU4oMZ1U6u/HW/kR2QsSWAgKLZMttcz/SUPvKmZIM2g9hS/DUy6mC7z+u
8dsx61S+A6N9xTougpnRM/b4/QMSggbMpk8kjK8VFfJom2Na2ZwyiW2dCRsLjO9qxqSrRMWlTIT/
aLIbji+WfDNs2Lz+X+1iFm/+gSTfc0dW8xkKKzT9vU8aD5PDAtwo7m2W36drq9sBb5RugF/IfXWB
Fv7gFP1lMdEEZXbMYbPykAEd4UGMToM8r3Cm9pgd5l0iXs5fEAm06ojhZrYFj+zM7LwiQLXhaP3k
Lb/V41elG+5dhBs0ILff29Y9lbBBlnW/fuUcUTBu8JQfdhJBGhj/aR7ZLqrF/b6NndbT4D6S8cZT
ZPuxSqh8Qr6ezIQ94G6n2ag0/0vW2UYCpV4l+NUL1Ks2cYY6Y79tewtxrLWkIAGug/p2CbR1iy7s
SEL+q9QANrNK9G3RKnJW0zoQhAxudWp2Io7ePvz9MLeOx+qOHYn5RSu22C3X16IQwQp/tti/8i41
JuUqmlFU+X/5hGm6VqsKAJHonHohVAmgmHBiue+OUXXwf/ZeWfowwcZ510ppI2ODsXHktjWT3coh
uCnl6Ihhwkp4YqHECALKnpp+OgFtRi6BTP6prGVKra79fiDqSpcO6AlJtnJKnjR828coM2pDJfP4
FiWF8ETh+g6VqMuOiuw6lyw8CB4f/CYeLDDC8X5YbhXCLy66S6V04Opiu2tJerlApwTZI0N63s0j
r79agLH/1KYeszabAkWaR2fhmRc9VsiSDdiGNWe6VLsAP1qvvhDtJ02/fAL4apYxJP+I+zxNHvK5
WyXMxU6FSTFl+BuS2uPMUnaIo63PCiDlRcFgz0yH4rgr9AAQyicXjx2WLEVv6QremrCFvCOG1p5x
T6kfXq8BRDNJDcnbCUu/Cis7SjE2TEl9G3luV/2TSgxq778/FsczfPhVfhKrE4DQJ6IA0NuZjrYM
qRFG8ntqtQROgVID592+1bbrsIsN17k3IuUr3Tf+7RW4XhiMtT+6+yY17OPgjXQlosEXmvwtN8Yb
5dtSvTtrdGYddwB6IKwOTSLhIjaKa+aQhYWemGdtK1wRzZo1I7viFPvWdMQI3mecXYONqNIXPHX4
YfZ0xOWyMPK5bWBoPVqqbGooUHPeeZ87Wr7FBWYBWZOIN9qAwUspVyEJQhSojIR9VYd0/9K3Bk6Z
C5Z80AQOycASzuDfXJJHcl9739ByG2Vk3uEZlsIsQvNNra+XqvAIPEMRKKqAZTHsX4cNUjAW2rzA
YcLluLvA/lx537/MVaZWAP38prNtbT1zAXqCQfyrLce5Y1b0D/pCtMQib6IkUn1LGHwCdLRCwgm5
XZ0KGh10STO9ayyupCMBFY3zYAOStylJs6Tjpn+uIOWY+5HQMnYF3pveHg9RHXZKeJRUU8t5TzXz
H16ga3fPrspHUduzW8xoVoNUaLL6fZwN1buiUPY2spSDfCSdddVeNOFNFgjy7uAXZTgpDC+6pkvQ
pxq6kyy+9XXwRQj6gQmIBlzDV8kc93g6JgNrKe7a2Vx7+LogUxuL+qxwvsBb9IUPN/hSpP5CtBWW
Xa87mZgJ/IHLcUA2AZa8J8bUvcbC+LA80eEEunQZzPFdTbSE61EqbNZoeBrJHrwU8DSy1ZhmBERI
PfDboxs0iHNKJP5G0BFdA5hApjP90O1pEI91VwO8eC+tOlBnxq+MpYTQE1hMl9BxxSsdEHfrbBAf
/E8Z3DXYDl0zkkX5f8jIQfMydfwzwnpjFIh0CIl+08roETgADWweXt68kom2zIqZUmArkV7ZVsE9
XqjkVidccoNb//LrCT4pTSPrbTY2BlE2EH8aLTJ4f51cZIFeSDzdB1AwP+dlS/PitXetyD0FyPis
b0kTOmlxmYF3+1amHFXug5mWqv4tZ9OjH2U5CtGm7bLJxmXFcgJKaekiQvfqFq5rbiqb0xMmyLiS
pCR2VLx2cVc2iWaRhhaiGILx72VqPOnuf7mwukTKooBuQJMGoUHCKlql5GmtIPFRMAiBy8DOxtOX
94PLzT3E4vVrmE/KglGipYXYtVvioOMbhkYg46BqZtxcw8UEGRz82R863OH7JIdkcA+OjNMrwvgR
Q/g5aXclaz9bFzIFsvI012hCF1sOL3aGo5tLESJYkjgxUlSU/ZUEQDe5cflUJdW2G2ny1HVG0Bz0
JWh0Wvj1BsrDQRvUP9yL/N3CAPJftCJmZ9H6Yu6ZfdEiZdt7tpcyAGtX5GRA+Q1TbJ4NoxUXMVLB
BCuC0mFqfH8D7D1zuaNsGtQD5LgDeJlwvvMizRduIoueXRnLoPqfKpqjrXI7sLEZGXkzB3960Jrp
/ojl/yS6TTVSNmCXiTwnkj2IjBUwbWqeQQOriDUiEQ7Xc5fuTOjl5AP7mH2R4TrgyrthMVJcwoHT
krGj7FDiczi9MyfdpLDyBAl6P/3DjRIXms7Mtd9o710qn2fIOuJ4kx8CvcXVzH81QW9mhRbXo4Qi
FFRHKTROhTLWwdklkGwgbxT2+7yRxndF1z0zku9YJXAEc5c2R+hFnR6fgwukh+mUwtP7ySI6x/JH
vuqJ4oGh6pGTLuH4gAHzPVCtnS7AflkhKyLEa8rchBXv1BLdx2szbi+UqJ76MiiCLMSq7np+vEjT
hDWWTzKOGoGyN/9jzBYDF1z0sWMTeiZJxkJCjrwQEclbOUVJseE5/uYRKK/u5H4gd3X82bz3khtR
a656u2gsZc1YTAjmzEtdAKbqGmAXqO3Yt3KKqIl4YPdpgo8Rrg+1Ledqg/N2gpWpSFdLoQeDYCHL
OqZcnloHK+JcAE+f6HJKtj+criSt4w9nLwZYBRavH0YQI//aYfrJwFDR2ZmuvVIAygxV17ED3KWe
FOp6X0CGYwSwMLNS8YGkOTStwiqEQyUrhdl/UBc6J3MYrCypFee6Gg5P02qHGouIKKCUi/4lQVq2
teGBPD8VvHFDYLcG2PMU4cR7PROLv15LPgrH78aMNk+nFJME5qcc9bjqVcpt5OpTi43oMAhTK87Z
ETMU0JptDOqaj5c5tDZQlKpbtQfgKfYY8PysROtyhJ0Tt90H+3YR3yBLiBrpxwBokNLKlEpfiyEi
DoTGnM2Gx1aIW1b0laXeBZPjBBz3Rg8IWN0o5YrPWkmH1xknXbC9UG3b9i++g3qtFcwWI7L9Rv4E
xWwK+zeYq282xo/RcAsTXoatRH+5KijYmGNqZ1GpvEOOEdUUbNISiB5pKr9+YQWg4DqhG3XgixEh
QnV6HAXuSP20zZnwLNbQR28WrkggAvpeGB2Rc4mHCSazIp0faPEaLQ1BlzUiTDVgEg0zX/WItqRl
FZknEFM6g9NJRLangN57lMtGdZduVBUHQV1Uwae4593E1pL8Okihz9wLLUWOsXnwK/OOjF2zcDnG
pxfcTsyVb5pRpzu/9kc4TUWNfmqESdqKucyCiplJKVrUemRvEoNgW2cBPjHaSsaabOYMoV1tJrC2
GeBHTKB3cDGQVc6+edx82B1NfqHg2SX28ROR198RjgfYwfNQWv5ceO7sAwGuErmTZ8GassVgxjN9
Y4yCT4fDcSakZWZ7l8Cmd8E5dRd5Y3Q/qe2YMnC39e3ix7j7SecEuoljrJFpkQ0KzAkruTP71Ipk
5KeX+IWJnetiHeNLFMeA7vMjZ2TmrsroLJNj6K8eReEgXmInKvaiRG1wMjQ17Ug9DW4aNEGCQwWi
/mvkvtJUJH1bK7yxk46TnGBK+MdTjb/9Rv0QTca5ik8JAwno7DSQL6kBBO2Q7cogigjdAs7eBoid
5thEou2sBUt9DxBqowXU+2qW50FI8MbixoStI9d5XOuoi5n3EpUHH0SM23bu/zb4CksQfvYi4sDp
uo0bNQT4rk9I+Nh73Yxqlt4t/SoW2aMQTgfyfpIoOL9geYGEiJ1dyNGn0o9zkqH3CfBCJUXSGUuS
FI1XbNht/hgM3iU9v2m9dDJ4NKOcQ+dt6R5T5/sg1M2fGwbPodnf6BbhUMfzSU4hntNDwk6/jrCP
GROw+jAk9a4P/S3rg0uxq7tRr10Be0LUOPNWKiffVPbhUQVVmNsnc2484gSTlEZVruN7IlOFz4mH
iubVWBQKj9uprjfd9rS/h1/uuy9Djr4+8CNlPm/aLp3Ujh+Js7+gRGV24C1gLGs5yCTYleJAQMnp
c9qwTKVWFWkuDceOoCU0V9tUoYZFxLNZOp19UGWPGkxIa9LllYNsTZILUDZTupNHmwcdr1oB8ddp
b0Q8tkcFLQRoBIY6wvgGJiHBb70UPYD1LFloEvU++cn2ol3zs4u3ZVa14QQeW+aktE0SoO/R5Y+3
K+CmNEDcOy3xCMSmvo6usaAWEijelovr0Wb+olD6bD661G4ecaFxP4s/NoQlUomXzWYterPvKa7Z
/ZcN/aX7VLdr3wuNNf7we7esT11TUS+9yreHLTRqj2qp8A8zBP9lmGl5ZD03AloV0fC6v5M85tSF
Q841x1g1sYEGV5A3onGfwrGbzSTkJquvQC4UWOhLSQTlmDCBOLEUonP0n8opXWoyMKaDVIRu5S5S
adymO6MSUCqs8/OIrnCojauI0SClnDvrsqwKHRnxqEGms1ne6NNpOE+TXAfsI4rgDhNYrvR65jXo
KsagkCrGPNLzbCKONgeyVnGwI3BKAbgvSxLeKa0YM7g0b2R72OuVrMeKoslOehaPG3nQV32hMON+
Ck2Njfdcx8lYAAvcE2j3tR6nRc6BYHbP4aH7vcCh1j04Dq4OjDdf9Flj4mc4ageKDSYGDewOGM6f
jy/zDpZZTqb7wM4+OBxsz7WhukFAJOHUlqSUKOEK1QgUKjsHTC1O9Ic/yzgyyRBVZ72y/IKy0iWg
3r7Jsjv3ck4bLYaZc0ofxh9UAEXZYi/17nrG6f1cHpe7nE3o+w0zLEREsUeE9neRUmlqUFuLSUwH
TQU/gtFlpr/80T4HLQNoQUXZcynVMcaT9/ry/tkRVb2Oc99Urwv+zdeToOILRGsWEEKjayEwXo9I
BdGsNcvmCKSoM+7Eki5RPktkbymULGBgxqNIWmFf9uA/0MJpp9A+Hb7QUbluHo60NRzE1JP5zMrX
E0Kd0wvRxaBoepwwmzoLJxIdjPUuX6CA/H9MRvE4opYzhrtR3O9l2hPSFJrGspQM7ixF0NBgHzBq
JEPP3DDKeqT/nR81iFyB8eawuY+csjzT6nvqTDI2CtslLsErmNi3ilJ8PNEVmGZy7Ad9UWpmA5ug
x+Wt6BEUjPMnXE6H0M4n7RnzPkWL04ynIFjqcQFrIyoj1r7sfvFG3SbtO+77vg7GnohLUq2AkH+1
zdPkBdmKyWBsgiJN/W/fRSMo0Kj+R1bpVhtgcrk6szn1cvNDHuHWKmoiJKA44jaFJrPE6APKoqAj
Fx+fWvyakhKun2zNVCD2Kn3VihhymxpegU2attek7zMqur3xYf0AkOUn9P+ratZjLgyYASdZ7MPI
pslUcNcSqKAvF5DouYD3xkHDft6B9CqPK/AwxUcwQ/OGtYMbRcfHS60c2pouUcz+Ra32WxlreiEu
HLjQv5KGKYPGB58P3bGs4Qg1IVf0g3DkQWZ88LkwaJB6Fm5rk85ket1N1FroMgNFDDD+bVzD5DrJ
cbimhPuw3BwWC5pYHeyPmVwWiLnkb/6/Q7mb381a83wzoJiuINnhcuTI1lRsGvSlCSD64lewHSfb
iYlfA7CgG+OOg+dbpAJ63WNGFUHUj8T3Z3NmMcPPCPon6rJ25YWz+J0kseIL+6ZisIsxaLjbWOj0
abWU/dJxdcJK/1cL2onNsozVcRKkIDq31Gi7/9zjVSlP4XsBqeOZww9VTXYtf4UKSfZBBg5Brndw
wrYUGMuHANqv0Wl1b760tFxNN6uwf0nfoyKerU+wvcENljrVb3lXmfK0dIasA0b5qxLEXc4DjjNk
uhEvYUFNPPEZbE6bM7Lv064fbeBthE3rAuP/xvBQN+EHlPWm3B1V6R7yE48G/tvikD5OjAkHvBIO
/pLB5KebFJ8ReajaDBDBd0e9z8hCKjxmWZwcPuQaGMfi5uqwe/0DXXWL4t9T8IaWcbhy3PTgGrfl
A3OvHlH3bZZy+/huVlbG4J8GATtKRQKr9zdHEcIoZVJrdu1FFxkNGIEtBdzLrXg7VBu8wLJFhJpS
GnqZvo5W8PExng+ETBpU+/pfx3g/l/Py4nusYbgG3L4kAyPh9psJdXpS3vDnjW/lQTgaqdXMZnxu
NjvjY1fB4Nx1TNcM55aRnDjqWPWDZPUV+QuGuG6InRZtY3C6a5HdtTO7DHOYVvIIm0/PoenJubuu
Ll//2QkwtIZwnfK7cutIb7gcyviM9DpIq/X7a/AdP5aoPxBiWRcX987tOr+Qc4mJfh0hQ46wO4mT
Z8NN0p44bssvRd7Q2qp7MXpvCThUrWpNJ/aQsDT7YSuYGqCmvT9fQSajaSZVJaGMjsfLs+PSgz68
dtVL/EEFPz17TPLI90hHP6UinV90RWeNtcb37yvue2/FFI5k5ae0CBGQhmEvuQKfgCHn7x5xu4a2
IgnGCu98gJgp+WXaLrvnJAPKAObBNIVDZr53wlUbli6S7AruD5DzYKBP2HNpKeVTAv4MWsJgOG11
T6iyg0LNNZ5fkZx4OJylxQtCtnPm2dkb82IWwpyB4UlMIW3XerYTvtyXQxVmtNGg2Om1NEJWAqsy
ND9Hck1RCQz4jQ24OBWuAZfePRlFBKKW0c47ybov/cOjAZZwVgP4j3lknJXMFExurF9nx/t1+e9B
I2HJGH+ApbPB6Ep40ScUYcGUhRFWvzrsE7mirsAP+ScPrbifZgh/yeL0Pg6Fe08NF/qeHm/ngRWV
E81NhBDD7C5Qw8b/rRneB3cauy/06ovbfvNDpkMCyaaRsrSAiXjWUvZ1CTuQPx/3hW4Uq1aetHMl
Qo7w32sZLtWYoScZKdVgE9/19/C/32/0pUvCSXbEbI6IEr5lY5sx/ghs3sI1UPZqt5F6XcjKqcyn
EMIWyociYX0U50M0PE7Tg0Mg65LIQl9PB1BZqQbUvryKDnWN0MWjwd5HC11cmedZs7fElZeCSs1u
9V3Bg84fGyEkWu4CA5XFRToWsKdcLSL9XCDreU4ifJP3dMaCCIstuJ89F5OI27gXFDfpHl+1Tcoh
GI1BpEI+Rts+fBFV1VwVMwtmXQSfP/5/zyVN78SQ7Pi2K1dranbuxtYAsyyXuvcyBtxngK3DqTaj
BRM1M8XnsuBK8MBa9iGfvy7xOoiHwJJeHolq6wfoaBWWV2x9qUWOJVyxg3qhJyBfgg2vB/TjCp8S
w1gL4eoK3J7I0GgJ5tKRN3TJllrACWVmFvUEn7BS9xQE9Yj9MzQKKfLtzLKH/pC0OJPHn4UsTQM/
/lUexqLMTGAlaurpMMJ6ViesQG8iExO2CyWbEHbytuikFznJSlMS2EaW+KXRt7qqSD3yNXE/u9qo
gB4iEcszZo6GD4WkHd9dTuWlFO5SzvWDTUWwLKNIxB2UI73p6rdQt4Y+9P8Vj+9E+8h5UiFD9Wc7
ozYWecMxMpYf0eH1po9K4Jyt0k+bJPA7Z92+MGbrYylHuyBGOiXqpcn/DO/ewA7CEYrxxWTBhONv
QpnEqxPfkFrxUuDVEW6TpVUCXFLfW94eD0tGYwU6x5818DFo4gRVainsZXGbT6eWXidgqXcuHbvb
cyJyku8jSWTUNxKtpgZz2zT/uSyS2z4jWiOg+ig+h+pU0bF5GozLn2kacJdLGH+VgKh/F/w8/+L1
UXxBTtkBgl+1BrJAYNbITObBL/KM7grgblgRcyAhodNHg4Ucqm8Xn8ZVO894WY8002FvUnrihXTu
UwI2VLtsQ70I5BhiyullvR83WNq79PGeOU+fczADvtQcmkPYNPhuN6gJaoUAvjzqH9MV1Mw2M0tr
uw0U4U2NYPpFtAAerrrFjkR7X6CLFUuvpCNCevIdW0QM2zdAjcE8Lf2eZvqh0np398Bc/ALpISAr
NRPDqCRmSOMtJ7e8PRkNUGC7vCMR9ccndpbw9Jv8exRq43nag/goVGFGK7O8iNYPgP5B2dH47KoV
DKFX3NvFa+UfshNVhDniA2I2xbJZeleJWlHeX0CmZsgLNGPEH7u1+als26yoP5GykBwzRhbPI1G6
/Pj41KkE0hVUilDyTxi3f4YGly6kO4fGhGYKwyH+plpazPMCuESlKH4bO3bQDYvLWw+y8tdMzVj6
PWcHh7tfw1K59v45W31J5XtrJJYSvuGnbhtL+RchsifIOhelHFfT0d0DsblYERIuCBE5emECSOfI
klYKCVOVagLo3ilJPE3Uc/QWKgbbo5MEywfr1DAk5zr1D/XQbK1I+l+2ZJqGjgFE+YvaFk3Dh2+p
RRDYUZSnrXsvR8juKHp2t+/NqIJrx4p2AI3+UzqD/aRFLLwnd1DbpPKHnf9OVwk3Ri1EYdJK1hmL
Ky30ucWyvpD0papWrH83DLG5450fVY65OKmNYoOppRdK/EE4ssyYI8W6PpxkeX8O9/hSg5y8eK2b
LBk3u2mmUkw+VJ1aTmw10V4N5bBxbmfnrVw9+o6YSqK4wyzgjIBQgGXwLpGYdCCA+/aHXvs9zoEL
nsYlemmrcskv4tzrYNbdjdzGrArjrsHIMs89VUyevMYzY6JNJr+ho4qHEQQLXY+YNJOodk9jmMT+
wd+Dc/z+tmpcwG49ineievYOatQox/m5SX7jAzglvQKfRLTPfxUhH/ZoH8iPOd0NakxYeGKlk5NZ
aPChz/JkJ+npBNnzLO9lbN7YYt+yOJUNWA3OmckabD0pdJYwT+JEuXKsjdFE4+Qh7jKLOYlpWn9a
NdlCzx+4Iu01JVdGp7lKrtJjlK7V+q99bqhiGH2fpRDHSARcqmzfnwzSQQXllS8tqFwaTIT8mHBK
ofyRuaIOSkVQNF0fJKXwA6UmATBv5OkO6EFPmtB+dAlUoOswQzUIzNJ0LqN+1xyfICOWWrOXDzTV
+DjH0JLpkyV61OG32ZRm9G1YErPH7aCw7PVyTyUz9Zuf0GLu+fe/bpkzAX1+7w/Nc2Dl/nWMsCb5
bvC0HShb0TTMT/QIZNvELUhZEuNSVLMxNtJ0sW3YOFSXzqUx7wnfSBGcFiNqSDBBzG8maZ0QVD7Y
3lbPLh6pdTra/XOgrX602Dd/uQShuT2CZphMihfu3ZFrBbgkY+HblRQuNbKqS1qCppM9PEdpWLvh
2Yz5aCYGsT6qM36Xs1RSPAJOdFsqjpgmhn5o4/Nx5CCqK/2fqUQ5mg2yS61517b7+9Lxqfwtun2t
kpmQPwWf41/fcIDgk/AKgiVAReXpfJ93KeyJo5neM64M/SYtRMydrgZT7a74BDA8aQ8Ye7mCg8OS
3TlOpv3mYcQtOORDUoou82s89pXFsoO2kOjh2xLVoC+ORkU91icbzlnIk34Km3dq9TPmo1Jdb5O+
n8D0wQiEaYgNiLIqfJx5Q8CxbcgKBaPa1QOkqx0/1dwNNmsVqDDBTsrX6S8N5PPu/510ggMJyFAP
XUU2HWzWftOJ4dA1TohxORs6aulQMNL5jjhrRoASp9/YH4LH7PBswGT2zxAo8wQ+zOHyBfd2aWc+
s+V9Omnofe0OcIg4sJTNAQxCcALBPKsyEOfDOEpmCtV5niwRv3sXQJs1pQU6yEKb2G4BR2cX+P+k
pfYNjAOrHWpF/Xx7kYjFEh4pcsy8OJQZHWAYTMiKBOGQCmvg2fLsGwgskinKVYaELRgESv5IYFvZ
/BROHVe4hko2KZhZL19RKbH7E60sJMnTT9uRCBFakZJfiIHfilDCb+m0SH5O5WVXe2Xogm/Aq6/A
IT8NkjjPvgFy8l0FLMsui4NBvXn5WXPBWsxDsS9wNgj4B0NcNY2iRufnsNTgHJaM8NUmsnA5tlHh
N5gXI7GZQAl33PwxWOr+R5GyEJNmo5qOPHFhuj8irzHe5VG8OC5ROC2/ONDgyChcFLnt41oKsyNm
vvFHFY9mN4H1bID8ZBxymYVGYVj2NCwr5mIvMFcoQ0eIAbCJf5x2qXog0n1xJNEr+4yf83ECn/+W
Al5Ea2nHEDAYAkL4LQfAyZRl4v2JCUvk0jURJcSAoayPxOjUjGVLKqHP3LQH7QRuN1Tz2+fbNoGY
48etNsGrAht+xwgT8rP91iic4QHeUsCSx8XMEN0fYCDmqVpAtc6Vdi9hN4rQY1AkzaOSxOletBn5
HeHe5goqq2Mf50KmyPyc0T5/vbgdLYNxAkLRxDWE0S7FPGq4J7oDi39Cq90Mc3n+3d5RD9rdDR2Y
c2PUM0SXCMRgAfDYWCXTaxFVuFiIhtSEaDMPsZ/sTiKqrvPO+72E/sMKZOSWS0gvpww8qcrnLXYp
INqjToqf0SiWngDLlzMGwdkXTl2aHW59i7FNiUqRuLTc2dfxNXdsYwz5xoYpewRjfUFQwQtfSeaT
qfwz6TPC+2PVwzytLYXerHvnQEEuqv57hlavRLjCzFMYYcfVLYT+8kXevH0yAPzEtzjlGi1FpG1v
yrObci1UlN2D5FsPK2hlHtBoAxL/1UD/OpeIdMds2JWW65csB33IqTj5QhJvKr35879lfTbNFuXl
1m9SPxXaFq2XYusKCJJ2BR5jbI89HYtQWqa2Fxtl9DnZ//ehQwe3ir8BflsIQ/UT3y1JJFLGhoxT
3pNjxTyUUnz1Bb+3Wsffyk92KBdYr6YIiyRngVGmEa0bvWWsEYhRUO3P/x3UUUdEn5hUeylynHlf
pNklYHxvDcA5LQqJOhfACMU6juKRnr0Eg/P8CwIsYClA4BzziQT7a3aF8dncUvd/XPD8sk4y1dvu
QpCQBDcIXaNy4K6NvBaSrCj0wV9wI9A5ZwD4uxntjJXiHJRXXZ1GeteUv6TCP7cSMGhZF9Ux353Y
pBU4qgwpYRTjru4h1hrjRuFpZwaQgHJh6hOw+nXOx01rIiwxPXph/WWC169nJFb/NesN7Dkb8fRI
ErMfCHYCseLIZjyjQlyDCOLV4wDrVZxUcNRY0SYpvYW6TzIoinxW+FMSLBhBumy4KnzHBJtxwGOD
Xhwj9ciZU7J4ij9qRfH6pFEquk2imkdA3JkgU9yX/e7MF2oCCoAEUHo/BceBCGi8FZSLfbTJE8iQ
+BKa+GCHv5oRXd78L+4caRUCUoZuiGSeNCtoEs2FdlbhZN1XAN1LCxTC6iWmr5rggIP/L+SbXHI+
FmNu0m7R9NkeVV5q5Aac6ROt2/weGLM1AQ6E9Tw8Kw41b3lmuv6Nbj5Vve9yreXIg3sChERYmpRE
Uf33lxp5ufpK7Mtc7q4mKItSLQfu6LlXxfoJG2IkNGoWaFT+WoFNkAcYGOQWHzIQWli44X+QgaC3
eoUg9LvE3Z8f+1JPGtj/FsLzuEYukPzxO0rdVbwqWHgYmLDD6zzm3EIBXK003adfUs0iAwQd6e4o
i+MCkHfNh7mAkixA1p2H7NBFnCPI+yEQnW25tnEnHqsvIdzoevOir6NGTKjhd3guJqIig/Z64xIa
KcNVCqitrzLhZdiM1MkV4NMeIqauuNqcaAlsDXrpQ4CAxIr0p97D8h6WAkGzBaLAnPPSuI/dlj7i
cc/IkQpKv8oI7MT7T76/9uiddsReQ/CgoIZE4Lhn2Q5BjuerCIcPUR8r6rBAslQp5olQWDsHLjto
Cg8xFQDWsxOH0ZkraXdcabeH6k6Z6GUjOe6QpBJFBd9KPe8jrHTmv35VLVC1ntEssoez+9zzp44Z
gbUECs4QNJ/MuuzTIQuhjFG1YPw1LT2/pXoBwu5hLp+L8CaAsnhFKV8S6536KF8gPE+nrEOflWZS
YP5vbjLUVvYh7RNocNkEtF3zb0Non9h+j6H0Pk9bCiYtgsQdVqksyC2r4bJ1CBU9PSsfjejO9k/y
3WaqWyVWlK/Cm4iJgWgRdm0SDuWDgqSF9zw0h8JY1XmdM3yKbYtW8Udkwv8SHnGDK715UEfoLF7J
q/Ja3pq5EZQuBZRw6Wb9QiyJU9qBXrKENJvHfPjjzYD/6wUiU0qokYlKYnf9rvxJ1G4aOJXXu9o0
y1owi9WMy09zX9ITfB5aM/d1u2ozkWs1W4DdtkdYBEUE0O0ACuxS4OlpHyvJr55fliuimsqJADaR
RZFn2+hOKjgDVoT5WhYzJqMVkDrruUAzDgcVlgmnMsPMwKV507ggFFqqkZ87p0rIG1ss3bFnO0PZ
7SBP0hDRXva0C0e21BB7aDgIjj98atUI2iEjofFzB1yDkOvzJU4lwQFWDEEOHsfUoVVGmqCDB7Fn
moyxxqx3QBHuMZNcPQnk9DB1NF9PCe19mvhcQu+va5awkvPGNkWw74NckqAb9BO6hdodrW5lKMcA
8/gy5gSR/FCcttlTq9Zh5z2hMbuczS/wBynxadZw0X/zj/KRG3XN12F77x50bvqk3xFCQ1M/2Fm2
hqjYjoKdjB1Y51iuVjp5MupcOqizASNMEKP4CIDuEcJSPiiEGWzKj5RwiHuAckyHHkNQgf892fS/
myIsr1cnwQkRGBOqZBrt2JiBIMOOHmDgiZz4p6JgUQ6QfSI/gNGZOcEu/nSjV6xCxhJxSz90A7BQ
g9FE7Gs8BRT4ayhi8eN2/1U1nJflkIVncB8khDbdJH8H4UagMVt3fRT3/9tabiweIWueQna64n5H
NlLF+Qg59vlFqA9+cqVIKfnBIdMxmYNM8UYo8wJrWsrdg1EqDOYmH9O5l7ePeVw43IA2mfHEarJ1
gHIJOUhS1tdcNkbqO8/0xwQXrbES/gWxQAiYAqVYyL+YmPkZgUHhaFnMRQG1m5P6SooctV5wLIOc
0IVuZElZHBNPHAX2nInWc3cx0KBF5vD4Yj23V6h+kHTFCfoGCpcDfiB6FQXAYF+6Z7K8S60tri4S
MOKPldwoLZ9ELmXEBxYiicE56vDb7KG+OT5EwNkn0VZzqRuDStqRGteP+OWulJr+mRBgDoAKeHSp
r9pbcqlvlCNVXLvop82EmM0gKyVwKLMB4IZPVvnIogLSkzlLAscvhTu5HmSQmFcBq0oXX9+psEit
osGkzNrThBanmEjOFU8CVeaAM5xSYHF0s1d1cjMfcCqrNzfCxajSz+OXEPMZuCe/JZgKCW8W0yKV
huMHAzYyDgHWYqL2L9l8XJeAJzpEpsz2lAwV7I3D9u/AY37Akvgv1P54mDefhIJsz+KcR3GgtXjH
1EE9V1GfqF+Vz3siWe9XCGfxGbdtZsROJgH/TVk0dyZnYiDwI0BehniDubSF+SmrRooXDyJVYroU
EHQenxszuLfW0mMkODIKmYS/N6dbfTV6NplJLjm2d/O5jkJsDG7BS/rLqi0IeqSGBTwxvQxbKqcC
/Gr4Rijuym++VhL31kNuhdj7F4N9gsJrIAE9aVc/Dtg+SPGgLlFRRZzByGeEGTX/mueQP7Jl7qqO
WCV+lLRPjdEPTgAPRQePgA9gYovJl0TTZKlqNyBtWS4nH4Bio1akB/0EFUja3Z6d7qaftgSlUPS5
lUeThVQVIuq+0CWszPCFvp76oPOhaM1ItMPNiAeDZlfF4/Gzb7PPzExWkSI7eCPdJIN+OpymIv4x
WpulOd3sb4oBZ8vrMTThfcxK9t0V+n/yuZthPTRQfQAbR0UqoXf9JBkV1lc2yqC2I98WsTaFT66Q
4I3DAFnKX5+pl9N4UL0A6E1Bqs6lsenKHt6tn/Qm0C2yYgmPb1N5TNXYlK/mquvEvb6e0YLkCau6
dSU1VgZGMnhqb5e4sPW2XqneZvSg3AfmB8Q+qQsZ4AGZ9i9J4YTWxOXjNtl4lrkISTbjOvDCVm1Y
uof5DexAApzbXaOU7C/owWx3jIFiv0VwpeDwqAfP1vbKC24MW76kPiVxXpAIEjyoBKUscbf2/kxk
TISaQLD2flKnLX7PMHiqGRoi+IEaWZsmh0Qk0sKh22dI6kznExTCw68q3mZBv6DoUWHUPAEPUN6r
TIHb+PD5G04GYJopITHZ3N86CLnDxPvGchJf1UYDMNpCdCugv95cwS0NgFfciOUAqam7wVEark0e
suCMgoNzR+tm8RKHLEiDzlqhTSk5XJLS1i73yp/PkoHDO/H24OOehqUDwGHjBEVtIMqGszwPzBu3
qSap3PqZgHWmg+w1RVuYp3OPTF069bTVgh1ipwAaQlF2DWcfL/TmyYopHPFrBkzHN+TvyGSDMAMF
umgu1T4aFM3L6P/C+2BUV5MpMxEae+6BExX10BodE65Gqqeq8XshuNKiCh30ZzmfjraiGXtJJVtb
XHbVqiiZSnULWx/J82WqZHW/YZGQ1G54wAIDAZN6qMbC/M3b2F9OB14rug6+kaNlL7EtG2rG+AYK
PaEPAt/s8J8fpjSHU1aYAr29BqmAH5juXbNNGjxFVrzccvtcxAdsxUm5QdfdXEErlRj5/hnqgG7D
HI1DhD57Or89LPqheztXIcV2BC/OyU4QpvXr9V2w2Fiba3nzE/IXxN2Fr0JaUmZt3Y1Aa9dw9gII
3nSuBxTIk1Os0PCIso3o8FAPX8nXEKc+epWEb1Gov2zfOYqRgJtcGXBVhNl6WJn8is++zxDZgmRF
mYjHZp3zuQoJV9OwrYinoNQdF7+sxtoPv3U1VOoAQEtNQEmIiEDbYbDT9TlxSOiwDp8RCLyvev9F
w+0ACztH1K91SilGdTDgPkyfaseGicwmClXZFklkVhwWiHKsrzTpKBwwXM2L/ZhxPVKvXOZPMK2B
AOWLAfbnBAhLY28QF3p1boLFPBH3OpU2BscIANc4lkwBRRbnftTit1Vcb2ds2UHG/7qjOOA+8x61
O6bQbNCucN9Lo+dXPtS1xSutkR7Hhku2oFKJx2B9sfuVXvIZRs1hMla2khds5nOgknsBKf9WyvUc
rLyGBH/7oDUxhj23LlcL/jnP1gpkpd3Qyq6k51D7IQ8O8zp0XSGhSQySFn55CKmQDILXyZ5Tzv+X
DIoTI0OLf81OCp8UlUUKu8tIN3odZf5gWJsPX4ksm2a+ckGx+NXuPOEHqM2osmUk6yJ96sdVLd8v
IYOWW0aR14mcdqXLrIwSN1MEikMfcMMDinf9k/QpSI81hkfA37+Z3ute/nceYIH0YSUf3IKKudj6
eUocyEvwPw4PdSlhr3u4Aw71cA0JPivynXfboZpMK6zsKr+aoqpG60ML+ujmJmXpxmib49tzh3dJ
iJYl4dNt97/dWBr2pDEvPGWmi30g5nAUloahb804sSOD7SkeTuZjUqswaioZAjqiwlCXfbz8gCb/
CYyDwOj/c4c9ZAg6qtgrfH6Hj8wqHwiNYwspuu3EfBSb+QVMu596JAXZStV578oWxchcdMv7RVjx
uAQXastiww1LzeqnM502kYhRgLCKEbJrXw98GRXNDJvqzEr0jsJ5y5ImXzIK2zYX9TYjfb0BpNoW
QKRFyh0S9v6Y1obkugpu9YYGlHOmam0D/fZZMsovcJ1ZV9BMhNdCDHLD54amsJ0AXaNVFBgEvjNd
yCqF4sQKFNQbGpN1cR/xSj6LJ8nswHRv0M5Io5RzH9bBWZYCU46S4P36kGG006fcctJp4bjKudVQ
QiS+cHiPQG1nlNieuyKoQ9mU2O77xitVKJsKG6UQm0BBJA6NGoGD2kSWDvU4OOSVj1QWmOz4OcnE
l2dhWuLoAQeVWu7JYegfo9HpeIN6H8NXOUDUKzfI7J7FdQjWRk5WtK88Sn4VW05W9wkwL7QjNxux
8QgG3HVTv0T66Ny4AID4KRIxK6qwvZCLIEmcQ9w12XCBsjwQoR/4bJPemWZAePPdWcgxMuGYOOGP
crlXSwvaJws4nff+a/oR0JOpaBu4FlD7oetbp/5CC7q96H+62gWVBpGffBW6lZf9vKwZesBmLstr
qggcmZz4HdzXj6uOZrWDh1wZaRTxfqTf0s+G9iL+8VSuGqgHPskmpQKcP09eFPq4byLmBs9TONU4
cVMXkY8n4uUbCNgOpRrrP7vwFhCoD2XpRFWzdUG954aKoUC5Pefz5KAeW7EwzftrPra7sKssso2w
Rao/w28wwK9+nroURXkWrQ4Ya4IVP0rZsEeWiwvzVM0L/ARqf5qKMlwAz+a0c1YoLxonGxNkwOt+
1y6g0o7tRVwF6RCvj0i8+FTzlBSDMnbS6lgkcREC4jcPPB18fMowjFZlXWaRM9FIMOBLYORccEaS
ZNhpzuZ+zu++kf//EdQz6D1nUVbI3GJLqcHQ1yCoppVyZYswrT3FV6Vt4qkXWvEkGpU2BLCo8iWj
YLztt6n5grB+XHu2PhNnm6T4xMSuSQg4f0yDAbaZmOouYslMY2CwPKTbEz66WmT1nxRA//NNTm4Y
ncLEDffS1VYClhEcl+rvxYRQh2tkFNO1GW8ppdd5tnemnZBsOJtFnzayGfYhz2qqtU1qqJcJjTZj
hIi5Z21IbYGUii3L2Ti+LdHE9HUTcQSPnHDIAuMIw14CI1fqz3dtmeI80KPG4+6GRXuZeLBZ4H3a
j9RuuqcJ+j0EORNdRNHDu12I3e26G/Uz4BgUVv4LPa65tpLzVL3I50zHo8kg8sL5h9DzGiM/eL5h
h/WnLjkpKN8WrL+tbr6XDZPpi5Wk5DXscOQ6x2nCHCgWoAAKqwJfS4RXSosTPFLYzQQy4F+uI0+Z
tEV1MgLZYv8L8ZohrLJThd//VVP/pVetsJ9dLG2KVnwZ5cU2kTJUFeCbHVyaK+pod4QfnkyrSSlu
VpCh/6LEtuDuEFwsbGh5J5mEauRcghsrvqbq+CE0m+j9OaFQCIYWtgvZoC4naxZdXzB+lUXc7OTU
sl7Suvqw0XFF/QMUVW1LSnI64Thr94dzWP9And08pxRmJHeKXGxRvbYOADyDalvbralHpDyLLgZ7
L2KjJxHeFkQeAqItqfvDHHKSwVQl5fLz472mRwcImpidM/lp00v/8uJujt0I5TGJM1O4/M8zUgpZ
dvxFht4kCnMLsiTSTVGFwVsA94MxOW6D1m7cugzFMdSsrcxJ7/ZoCeJjTtGqjRv56muR45EoqEG/
yJvj2rjo1TqK11tUi25wYxwdJZ2CoN2rmnRBYDKNqDsLJVW4F4+QJfcakheobdhwxkVi0jzvOzxn
/viF7a7lBYPsZvQxWOnW97W+mflgSPFCwzzCkIhTEn6tZ6B0MJXAYyNujwjso27Zmp/y4oASx7Qd
Ull2zb4bKBE5v5GIEpmgxkZb09TT7gxfyBGaiYMayz8EWLERCdZIpjGT+p0Z58T+0f5mfu7R7Mxv
NNbJJcxzNXAGJr1VxROQwFUO7HY4JZuwHLQx1XUnmglGYN48DdSvgbjyfXA+Q2x6SRi/kP20zl6P
eLie6PgPPOr6So+dvfn/WDTMD5avSzeUHzNolgR0ClAkESiK1uFXGWlR4OD4bCLhi7F9ks0cWfBz
/x8e+DYPoMVFenBRensv4//72Y5gAodwWCb+lkRJFiw8nrS9ffs4xNKhRR3a21o8p3PpnHo2kIY1
QO+VBp3neqHGX0ac4q4p4Kec/RO4N2PQ1sJ7gCiOBT5OrIbIcDi9tBxkDA5DiqMi9/iRcvRip6QK
u5XwI57BiA7jw3yoFwOvQ68hpB8+4SnDY+J3CsMdyvMsmlJjHd9bkZyyNaWflKsDaRudejqh40bv
YpIxjCM9/HFS1C5KUxvBooemWQyTd8FiUsPPs9YMQWs5vB+JqEYoJyn8Ga2t9ta3PciAh3X6wxxt
iyRrnSWRPvweTOuBpOcMcdEa31siHufXJ6oRWkDqzRQa7lx/8pFd05ULi/iNIE3k6UfLDh7tStqc
MUz/9uBm1xA6y9tfM//hhPH8nKyl2KHYnVVeth0tJ4gYaXLZEnjGIX2dhrzyQ5qt1kkLpe/+OlH6
QnQMOkpn36LWpycs0ahTpiGu6WMhaWBCZj6bJqO2QUCHi/nYQwHo6kO3WuwZ3VqMhNH6z+7YN04w
IOv5R1IRXvw7AbW/pYs5VjQDjEc2nuO2iKyCXGeE1ef8JV97r/42ih39pfoxF+l5wN/gPyYx6OxW
+n+wNHaptcXvRP9lk3XSE6glZjVOhKTz5ypipi2XzGTMmqss99z6ueV8I3m3pikE0BiubcDPsP9s
JOUsq6TaZKrbrIsKxxGYt2TC9qNU6OCcUJYC55n6xRltV2W+4MNyiyoFlgu3JLSwB83zaZwO8C2L
LawUC2acazy6LhRTAch3t+Bedi37zXHvhQCKIX+tW22TxM66zlUGfvBlXSp1ILuaJnh/IjhJgkNR
uhsmGn5ksK0Op6yHkqpmPp9Bpg3xNID23p8NJhETN6ukzECsImBVxO7OYD/aCdX2YaGCtyRWldvB
eJh4c36GHKxX8qrNezFRj537miPm2dtEEdgQ01Gb4mPFPoGt/HzmfdtC7qgocmi1/s/TDcLB/ByC
2n2x2A3Fg7GBdWpdGMmRh4cKgg9HBts9UM1GjU80wMPoeGm60LyS6rUvxKK7OL9bPO+0GzA50369
1F97idIbCMSIZT9hwP/vNCQGYJa/JYnBy7UmqCUvnRR1EQpakk23Ahj39ufWDiCffBuRkNfoACHT
ozuNOgDgVVrJkGwjGg83xVQKy4zfJIu107X572KmWlTP0qdaXMQ38nu391AntHI08J8KHm7fT//T
LYB9CDxdwH/I2stGzW68G9uWiSv41Cw6JiFEF89oDxgA6PuiKwPvk7RC7rvFxzTsaTuARZB8FyhU
KgqdmbPeqp19RKg3fvX9D058zBH/9BpyYTcEV8cReUc8UQfUIG/RrH077yb1iMJTQc/RRNM8dDeg
q04n0+WOYYVNum6lJBaUC19dk0TDXFgCiLn/LXWJM0AeIXDTWU7VGGt+ZiDYm9JZuuM5uo4y+tyy
m46d9/ICYIIJW3StJ6geA8VkbOuNnONJiqPQXwqxX4QFhY7ELF1hvdj07VufqZjd8RthJFJyM7ff
tN8HVjV/y7vbWbGW2xD6z588H5ub2JOOeGZuQbYaKCHsn6puA/1HlEqGP42VgNmqfV3jxUd+LZ34
Kd1CiqQwnstYp3kl+DmC9sl0Uk01EaCOb7QemqLToucrSCn2XcKz9xumGUZWnbMS9ztjG76AUb1o
UnI6GM1zPR5t631kZeh3VJQdkDZ3Ef0r+9ELnX4DtJdpwW8CmzeW8Pj89ta2ZyRpTVenYGGtECTA
4Gf6hEDe9hq9XGbgm95Ert3vaMnQ5MZxPLawPt8sOOpckr00Vx/dqiz2nocl1Oct1AMtIPzeVkQK
Ov1SKyjeQiNp115y9BAQG4HBZ4ir2wsClbNd42qDlSQf3rjkHgU8hsWSfkVDQUqQP24J/7PTHK6k
jl/iSJfaPPmJgpiHHRSp5TFL7hay9GXW7N0MFJIrxEAtHJ1aaRkiDIR40nOidClPBoqM6mWXgKgn
oAFLwyBH46pbcJJi/BSP6gakJBHtLCiZ8o8gWcoFqoheRwMff8XCIJxLs6FIH6fQJq1qYWegiSpT
k3E32uuyt1wEkMMuUw3XgtoLJhDiN+t8B+aqYl7D/azLaP/fQlV+UKw1bJm5fgWIAbafQG44hY5S
92W4JfXbQMXTVketFzAC4IgNKP84hG4BRGYg45imRV4GXuTHq3Wu1OLVprMETdcJOPYs9HO4+tt+
/9dorLi7XaxW8JvepXKrsNThLItjmhJhoZ1T3o17/U5K7syHq+Oy/UdXoFyeZ+MqLsAzAWCglGGo
8Dc7W4ecSZ+/DR+LoiJghiIOo+W3krn2a/+TbD3YcsjXjMCBNXDiPVMO9YOlZhMVn4wC69oOcF4m
Pz+Wr1oj8QP7Aa05CZcksLRwscBWG5XBu7K9oMRCkHg4VnNL/QKUMypEji11Zu3UtvVWidVUBCkO
4cj1iHxLXLgTlg0q0D9e+txpP3qpnzuBVWz4yrRMDn0PMjbVPq2NNh/Lqi2XbbEjCRNrlWFZazV1
I4z0n7FcKkpXM8Hlkp1g7HCjBvTq8Uj9r3+NI/T/fdH9qty02hb28n3cxg2frEBnGO3eYSAgvmhS
m48YpVyv6Mk51yuUIVuudLanzbsbGW44Zq6TwSmyNghvcKJWoFJRtpAdE/rJSV+aplaYq+rt+dwb
7DxN5rGJMu22Q984bJ82rtf65ytXqr8cKqmMDEMUWvGL6X9LY2hhLva14NXKP4CPXMq3VPjbND1y
G4YuG+ImLU6zO+4DEhCMI8E68bfWtT+MS0mz5nMV6zPQ9ZD7q9q/A00tyeTvnTY4cnx8xG+QUSpM
qIr1qNm+gRpDNuSK+ITAE3DlzAMmjV8cD4xO/U3T7ZCTV7xJ9rVaEqpavkTG82JM7Xbz4mChsa/m
KoP9z9KBrtTleFwGLiXvqNWOfSvA2zOENapbNnOseZb3BUiYhBG+H5kRJ3JGioWwd+GR7czAeAIq
FJEHNW7awFZwbkYOWkK5qB990Ab0vwR1fR5EPN99LjJPtkk/T1axT94H0ifW1D1nC+MlUPoe/tyE
KZ5nJPfRcksHSinMotgnVb6OP3Iz5htO1I/YIBJsvobHItuxEtGAXaLGwI55AVrpGypqbEmSXvf/
GwBEnVwECqYXxPSOZ8STvUb9WEmBZE8L7H/EnFfeaKtFslikqx5rP8YJ+RQI2LDkr/uzkT8KR6RC
YLTiKUqHVMJOlMnzGHnJKm2gNkI+43N5LiRVtXcRPnFHIHOur0dS6ekbkd9fq0+BKjcoWpqHJZkS
VyvLyuPM7sZtK1U+TiFxyx7BbXmxPx7Im6nabJuqnbrDt55BTj2tvomMaiPW2LKksBx71yMe5uXB
8loXNv9siU0/Lwq/dVg1YwZBuNfa2YB3Kh9Nl694E5vIPhkoO9KuZ7bCcd7FyEXpxABAzlduYI1d
qJlm9UyE1YRm1q++nefhEPAZKLyvllWcVaSyBhwyBzMINf8MYP4rTXwOeZgWTfzl6dtiXE20t9M+
feExfDhE7NkVHazjlDCkXgHFxL69JDI2SuN4UyQLUGUR0kmIZKEhoi5aZkxIL2J6q/I9gvO8CVvP
+zyNfolvyk5WUZ8Y7Q7upKfZjVKFlwX6CdhUmAUrjtTjrG2X8mi2bZZ5zAiU8N7ZZ4Esp4aIvJeT
BRrXY1GTUIZpH5n68+6RPF1fwEnVuZqL3PhPdnyQ1XsXtVDl3Crk+mYdK9DssGN2Nsj79NoP2ZVe
8JJ7HDOiZx9TnMhDRLuKPWMrcprSVS6DzMWQEi9FZTPUYbmPmjCir+lCwiJq9tKPnK24DfOC5LEB
09yjTX7JVYCC957ZHibTdOkTf4L6Jg4SLBnPa+xQ15Xp8rWbSkenLIK07pnfIysQr0HuKJqLEOMG
LaSsgBz4NBurX2Dfeinwq+EOCPHrNX13bc5F8Yo4Iv2MqdHaNos1SHajPgIYYJufDFJUSGfR249C
SUUEHJ5Gl7s9WQyY2yXUZ8zb5oC/F5ApfUDQ4CXOmoDvCuzNshpjCkt/pKTGlPiEskM5qi2zz8mc
ZnrsyAoZ45gShOCi9H9KOB+9iiY7qNM61LU0x16YwPIoKxQxH2LddJO5HFDGl0hU1eLcAkcWICUY
LxmMUEskJ0rbl0X3xiJALTOlKWM/0kv6Rf3z40HvkR3ohynJwtIsL/lRuU4MFDg81mwadPiflQah
HD4f/OXe34Daz0tOjukqm48zOMmWI82H8ZDNZJzxn2Uo+gZT0F4mzD7U1v5ePMejGfstMoBuCqPg
IVSkcjQHa+UBi6a2cRno+lNtmA3hwv62ZY+6LSDiNnLoCG4iTwJkZm7SyropZg3S/380kO286QIS
PbAZumVUwbAFddy/qK5Nz/HoaxMgYGd9Oi0uZc7eaeXPXaCHn4dDiMOFdXJ2ag1GPyfAY66o8axI
hBTLDZQifzFEHJaTyEY2pk074xF2LJ3gEOunarrJPZT5p+zU/nfp2S4xev0rk5e+qEXs6XYuPv0Y
c5BEaFONoSqUIB/FvgYqjDFC8LN1t5rkEszTgKkgx7OgejMhvD+j4+TE4H5Fy3kT72979hnWW6ts
aQ8QC5BjYkbrwAsnL24Y4CdbmCNediSTYKKJ4xQw6br+Tv6lamktp5UHKxRrtW84S87a/RKYsQkM
Q0JKrB/ACcS6K37rRNSZOXrdRyQ7VHVK6fCZPdboQ4BL4jjKIe0tdKGkIzm4lnD8N6SlQB4JHrWt
JYsvLDMp4O8lpeo2eYV1HCzoq+4CgvQxQdxMFYHUm0HmDFdS6an2n14Pkms4VXAE/TGupSzqi4Ab
x5tlPUnzh7Eg8MIlW9tjAHefPm3z0UFaCU5UQT3EsR/iJ+1yRZm+WcDc8aPGTrDnUs8wf7I6all4
HJJKyediWBw5VIxIl4zi32NikZDNH1HEdiHw0YarQ22GSnmahFD8SNrq9Qa9O0Izo5L76LGOqSwE
T0sM0+xkfz9+qQ2gUg0Dg4xkzH407lCMI8KrXtGeXS6i4LU5X8H5NNDOe8e4khwYtTrettA4CAPI
juUcaZUoLRIcTg7UCY/ZuMzD7AK/UiYaXIEnmuisaRCC/51tMt1fHLH9C7oi5KUb4zfSsQFbv9xu
PRj9zPRwPEwibHWp6ev8FOPoOPUjSiOX2YddMal/VHBUJJjjXYS4Hg3CPQRFtlTnstmSbIyYvtMJ
hFH9PU+nUtFK/BqmZ8XAhTiRbMpEbNjOsuhKTXlSZ4jYZ6dny6AzdPA7BTbPDAASSdRzj8Z4M5Qy
JqkmkQr792p2hmw9eegvNhE1EaM+xgkc52dEcttDIx4fTtaV4ZfglaUCOG0TqNvJR6DbA+DIHCT0
JNY3YGoqoRnZAFdpceea7HLfEX9mcqr1BnmXVn0eeskuApy8nEXlKfuZPay99ySOR2nfu3Py386W
SH+XjQWYoFDdbmcOv9cD7VUuL2FQiq9Qo/T4Sw9ST3LqPW8nlG45XrJ9cCac7QMgZv9Jr5akuEE1
KsedOmdCZppJLovlnBPgPsD+2Eg8BqaC5UTJtUeEHg9BWq8YsJXSXX5riwwHpLkErxTcvP9k0Rv3
gK2wZtqK/3KygmsK8WI9G5EpDBV4B4/bX12lDJDrVP/FS3NrK/u6UeDf4ie3bO04OpKFWSr6JNrB
zsyabZ4p7J5x+VIsyWJ5GUZBaW+HwmlFl/4lZnyHjZlr2mWFYWkxUxE0nhHD4kd/mkECpHKHiVfj
WN5fuc9WCMdk1O1hnGAt1diwbtUZ59jif0zetuj8ZG0DduB35bYdNwL6kYQPVfEYq6WZn9dA7o4O
Ni/Mc2Lbec6aoqqO1+rSZoC6FB3mCCpKbzpMyhqLMW8dic1ICm3nKbwqROO+JdWAKjsnW9AemaLE
YPkPPAx5R2+Fx8pGqirR25j6q7AU91RxA6J0ggTIXIPPRYNZ3LITVm+qUxU6avDyrJAv1/BgZS60
icrkJKnco0sY5FIiH9EOpxdJAIhQLtc3qZ9j1g2WDJrjtms93m+iXw4tmawTE/O0v8O1vB61ElNE
BAygIbIJ/jgyMnRAA3CRZrPr+IR+3IabGG55gVpFZRcOKO10JAh++jkH+sxwZYKWG+K70utOUJAI
3p7Vb6bWWTnHkp8Da3kIqGbPvBOFF/nrVPAR/Aih+ILRISnttMr+xFO/U9MSvHh0rh4CYquNwq9s
XwV3W/N96RpLGJxhAZdnkzm/4+JmoxoNOnS91ssgfFk8eAO8Urp7SLmboX4o70tRtbIi6IVHsz5w
EnVLBEfh01X3b2i2+okMJjJhxE8yBT6hTY2s87VIifVgLYXA5zeFqPxdv4V3cSQEdYjXwSD8jdE4
er0IyTLS4o1LKdN6oOP7AewiCnUIPxtns/YleJqPc7Yksyechh93gTxPDcgRBI/cdNKYH8GO4nVQ
1o4xNBbE++tSDPrlplD1lvK37zsggbNc8zP6E24nv72Afbl/ZKeQ1xpQIX7wqVffJ1akt5NuaUBe
8R62g6/vAIdcyWWwEQ+qeu0XVktN+XfPo8qM49dT7VSHZ37Yyy5Q2pI3rE9+ha+UomQ272ys/yuf
zWVhaSsMiDgwEHisbr7Ldz4NbJzhtv/LJtPpheKVapeWMxhRr603zQ9orpJ3zBeS1oOO4rpaNZqg
6oIMitptb1AIaW0M7D5//UvpwCGbEHZbgswMfPixh1kSnLqQOGXdZiD77utq0OB0tRk+tNrfJSzU
N4rL+2SzuJPz77xuD+TR00vRaaTNjg5BWVHtlXjMUp14Sr2/0zMKJ0ni4is3+qhdQPn0CV1QAogc
pSzIDJV9dsgYDKyjQkp++uRI0erP+PkGUzq9JGErbpbIOJCYEC+5Ce+j+EWOqbbdf4VXtl/TeHTC
MLfSs0BLeGXTANMVJ9IPcMABSgbivfLUbhuhYR6K8roSTZaX5VdznvqWroNyaeHwukcP7nas9Dzt
PxOTkdczMlqKorkrYe7lNB6nzj1TDKUjR/GNmXOgbYEuQ7wSzQWtH+0MHyp+WXzwrrbpSWt3HivQ
tq1kuUVpSkrrBxWyyhLunzifgoyAVPMRLH9v6nRvmDEgkEoCwwvTXhZknTH9owOZXEzlV0PrDLOP
yVmEPjexaNTDiwke2eqAUfWh7thCYOGepOnSHqNBvQdPICosFUfe6lD/ormmuiK2lVgXQl+2xw+5
xVe8F6sgSMSfWvVY+QyJ+wPe7QdJtStFuSlbDjyKsjedgjBN1+cX0YvB1q8Ps1fqeJr2RWlMtiYq
2IJSo3qiNykwhffIJJVdg7cv8NSe08qpB3CTvPUGyCYBBVKbMJTMWu0FQvDDgaG9ggZR9F30kqnA
ACriND2VmO9F5V9Hu3QWIoj6LivZcfhysgv2xeFir2BxM5Snt3fx4MdUgTfAesmWQSTUbDiGAlWY
l1x2OuGExGmZEUVZtIhZHYK9kg/3NAb3pbidtAI/tJC+mAG6RURO2MQlB62VNa1Vg4HSTp/uVq/V
ZjM9X+0F43UZdk3OHiXQ4puInTaHdpeZ6m/hiw4BOcim7WQS3BKIqGOFssM8LoyR+tt2W6ljwrD7
Je5pTCcGmfbiTOZcKLYJf7x+9GpA0yZ4qFdhd4UUDhnfgO7moyXjujKUzi37zeES4kPugchWoNoy
JouEsCjkRymQ0Xe55KP+iPwEksXfbVoLWG7WWTrZMcaKCm6jCETBYCYwIEUaCDAG84k408TqWVg+
mwwtlhwq0y8G7hSIIrUxYmuOaSOalhgqwWPTw4lpdo31w6Ll/xqoYrDju0WFWXt/hh9iDWPZezmk
IEtoJh1XWvKUhGWYW1DVUee1VGF4UUN/SVNl9c5RiPQdz5908k8YhB58g17AXh5kxOSCIhrG3rZH
4M423fEjyMHExhQaSomV5CmOKRpIBtS+u1Z+eQxsVIwOax5CYV/XNe1xU5jwORE3ggKqUhuqE+nW
PvVB6DBLj1Q0Ge7O3iXZle/bnVUcRGVD2h/RzOwLZQLG6ZXU6fsZ/EoJJ4sSy2OhzTHlbxIbwn76
EKOOZTJ76Jaf+srNF2Gcf3m2UB5W5fZbhsQQTu1oOiywiQshfUlsiaCTw52ekP6HeDi1npBk8W6f
BiFDzelZopK7WMtPmqUfyDH/s0QifY1iW6/Js8vCdDnKgkJE2IEUBO+Xge+A4+P/6hJY52fEgERr
V1nh3k2COA/2CLztj5nycWpZWglPFVAOndSmnY6cdD1GJBX8tTr3sjVxclaKWBFLdHzCKlfVRED5
s+MfuxXkiVikLomPaJXHCYN4qTLo0ndYstej6OAkCjswzXX1gRBKOW4A12jV4titBeOd4j3eUIyw
tJYv+sHdQfaNw/jmFhS2+vSJMm5x6f56POxmXYl92yXhPCzEVRapZE+5NYfTqAQxTPKdCVvnS4S3
ayjtRRF5wNYyizg5UaGDhK7KzMv5CcLY4SSPLM8bNA2Mw+nh0gEoN/yxNlU/+27EFXvk0KIf9uCe
9t0qcakdOuqKsPgv82LpkldOBQyo3jUD+5Wtw9uDpwPItp+pxYiAFvHSnL/B6+eY8Gcbfl/UUBPY
GWYtKmOYAje1Uj+UI5EYy2W0qI8M6gDmcu8jGU4NSpjWi4lDEOpkWEsaNBrx3/1fdcxE628TNXCN
M5VWZTz6lFWr42OG3N4/DfkABPEuJOmuW+N4NGzCusgvGcASU0GAhlI9lsqUIZPJoSXckYZMpKdA
b94tOlTALDCwHHbwyGhXt969bfPUeNCtOur1sYiPLFF2liZkdwhb8nzZh0iGQv+QtHNjNC+BFiNz
Yj5PXQQb0AqQMPk+7PNq2g+gYko+sdXnyqoZ8lA2NaC+G4yZgYBzYmD9qRwLabRo8VQ5LxZndyVp
bXFyVkLyGZemeUTOqMb97BQ9oXNXBROahfswD45MXbWuXahD/mtB7hglv8BIlO+pnr1b+TWaWREB
lraROAGTzazcRY4oJWDzdRqOs0fjIUtasHr+nml9NZkw9A3JtgSmuEyGbMeHYfIGpgEYZXnQk+AI
d82oo7M56Isf6IhcF1j4m6zQbyS0VEkT2WU0JQu369EzFQXyh6ni4W9xFtfIXPJQrDaiLscTW78j
BIRMbYkl8oFnX32XCv7acXopoXP+AkmhRuXWJnrO4WEQ6dt1VdHXptFw4ePvHSBV8OYq5cHwZFC+
7sB1lNN0cm8B8Vt8An6dP4rgAyW5PdeLG7GF7aB9Q9XZvzn5rWERMQTJ2d8zWKeOtHXwVXm+49ym
KUk0P/PnNUaPr0nZLX/BaKuybP/0DyCh6vy3k9Om0+YINFnhXA5NmJEIUU7Blh417+Ip+PInfQzZ
bcmU7dpY+Cift4vQxiteKKWOGNYu6DHwWuB6dK+IveWdRvnzMXr88qr7P0GAUetAk5m7P5McInNy
4UJGYqWgdRFym5DtjckGUBs0zqJ+ErSA4zKVvgeorJ7eRwTygCC6S6LTTVhga7uXGyK5cieQFHZm
8KXzIKgvJeS4WWUEoUHHgH7KuriVV6r2PS85yxFyC2FDh0XjynxTC7bi+S60vYfOx2PVczHEwnwA
sbyzEMyTUjcSTniLtnJQib5GrW84uZFKkDUfSfWiQSv/vKDJcRHbWmAwii4g2jRWtpWyM8c+Tw4A
gQ1qXkp/IUEKySWgkxlsQwd2EA9d/9HEuOIaaQK7bnMbADN7zmBVPgSZ+vk5AmQInt4Zh1Z9Zq+5
/hql5P8fQnyOh4KmGiGqkQRkoi95EH8GcDl+ITMOZBvm52nYvqCXggq+gjJKP3bvJjm1VgbiO6Nz
Ry98N+T0Q1zK4cbyEh9/g4o0KBb0YE9//iK/N4R+sCOkz9vlQujPufJFGBxixdaNQ2dbKCZdpJKE
3ktPXtRoa23WL9mEER9wbVYGAgGFzL4sKlUQ5ik/so4qleKbmF7jUCoA1X+uN8XBCqCY6gzhZFt/
KgR/xRH+dwdl6ZMWzXCXbSQYv1t3SqIb4dgnoselk1WeVLvx/Sh8ggQTeo5qCrxaFVl/1Rv9rpQx
7J5hqYyiHPr+0dwqXH6+MR1Te1CwhWPxeuMOr6nKWnnrKV2ouzJUgDL0N2yp//EGDAJV5B5POl5c
kLKeDVja3SSRCV4laiUa8xi0NbW5B2LA5juaZn+k15R0N9w/vGN/UuVfY5tocWgffdDSUoQ6/PAM
+KilKJBSc2IcCapBRSRCJzSjwsKRcp4MZkuPXNN7sEzuaYZefx5TvRjuKMKzpuGh/09fEbbZgkT/
kOyr2fvCH1VdfyxmOj4Rae4I8W00+elhAwKqYls1nXXd8O5PltjbWrTeX6RhCSuUsSNmmia0YDvB
F9K4Nc4imN66UG1Ng7TK6RjNGNAY2NBKYv7dM/9NU/O8fachAtgzVnJSOQ2YPnod/YIrPgHKWruO
21Xnue0kbgoTQ0ZvIa2TEEU/l00qAFYh+x3lJ2gvIgzT/oPs6BnSS04zulP6ixTHe1Cz92S8c45l
MXElK7BN4Ngq02aNEqNmFWziz1kJhCw8uF34ihLK/aWpVfCG1mGBcLikIMsdGx9grP4RcErlKyB8
A080NkIiJ0H7Zn7kusSORgYOiFjpzX0rfoOmfebnyd6Sjee3nCRrzziDJyl/EpQGOOSSCyFpJyMt
9ySp/9vHEBBhXl6XYhVSPDbH4usjft8KjxXvjg0ZrjaxRgyk5fGenzXX/wE4v/TQCJ84OEF5H9pS
OqkTy1UGqoZ6QYFGci8GeKBIqUProN0MrqwvJZ2WZ4etjWiF9N4mSJ0NSljgWDktVIjij0SbUgFI
hjRE4akEiLtffxZZxshTVXEJTZkzWaOscZMzJPL6y3548xa+41gxB9tCvRO0hRy6Aeqx9L2arKds
Q03lrfYfCi+Y4cfNcGarVqJGotpNcGaecjQaqhwLtR0V463CvZx3M87LSB23xY9o3YeGrhJBaMMW
9uT58Ma7OHjiydbrU8TDbnJ+7+7Ja7B2TtINYoapz3FKWNjoBJtT+ao9FMCc92EWOap80BbBDdPj
GSoC+pWaRdUiAziOYp3hk4cK1a/+aD8ImXKL0Eaa9fEtY/3BUlwiBAIIdHbw+L29fIe4O5rWTTp2
CL/1+wQv7EMtKMCM8mJZTe27OKC/60XILLc+20G2OA71PsV5mbe7eQWiq+htWC7AW01WeNsxlbuZ
ZOM4yelWgX1Uvj8YvugTnWVzr4qHoLVGzqkVnk0fraey/He2FUa9I+ZLHlHBe3+7RJ0rSlkaius0
QObjoThBSf7TRAn5lsAHC/2W06EM/e2utcKDLZfkcmXeLqCuZPB893Nd393RxuOE+3VYPs7Ajfu5
+vhcC/Kuia1vKhX3/K2cn4hFYOSbZ6W87Fm6FE446wAWklDcj9hYtMtPhtnroArjUHUjWG8ODh7w
WJg3SF2F+NObE8+slaBpqZriaBGuaRojNx8e7udcTf3sT/wjV/WSsoLcP3Hob6bcAIaM4dyS172F
NPdOX8RV7vP4131scMh9FafjHB+F4Gt3UPtAPFsaNuPomwl91OMMjf1cPFbaj4jWwCYE9VDSal0H
/lHD895JYX0NZP+M2sMydPI56ZKOSt5h1sczXCiuk6NGmBrxFD8kRqm/IqV79T7H2tseqR/luiHE
SVboopCx93V1tuGDrfcf59q9OtFkVtx9etIT80lSOfwzISTzPps5eNnvgKjX4FbCLmAlspYhiUOe
X2JBd1hxnjvhiUNT7Qh8U1BbfiH0sBno10JKk7JFfE+G/Tl6zFsn0i0t49flmqRNi4qOA7C0Kv3U
ov2xVn/bvdS6vJKD5ovxZ2OOYnCxvVBMh+DsfOXq5bSfOknlLFFCYgipgQYSCXeEUP72tUGQqc1X
ur2WXeSWunuMxFA32/NEyOpYwsFE/U9U8C/utpPNRwak5CnESmYh0XNu7Vl9cXmuL3cfq/rgzhdc
253y0AW3z3DSPNhY98llft5ZSjNEQo43zxbjsrddxG3NELWjG9/+ukUggCoF0um54iOQK46PaMQP
IDGr3i0f5GYGZ+8EuoCD/I79FHWf/G7pIbhTAFjRF9g0oVr0CMnKFCTODtPSycKPBlaAQ7nd+IK7
fW8O1vazuid7F88rkU0OxfPwwV9YssRJR6hoGKyuPSiS3xELs/OEhNA1jj2a0ISgha+ucZeC6jt1
I4Nz98QrU1yKvIdpPoVwDZLS97sNXOiiRcvlAOZj79eY8sxHvscvRpLv0/1cmSO9hfGcGRrguWHg
bkzTzoQbgRAJ9bxAlU+A4OYlrLJkTtN2K91d0l1RAOobyy/mt+5CnCxTgpmC19hmP0ZbxahMG/+K
TfJQbZwLYmaqdGxIkBsacrRCWbUibFrSAIAO4woOh3SqNXdcIzbzpML09bG1xqpBxUT7XE1MzVhv
JCXo8rffcqjpiXlF9iFtjjc63RGrvudkUiJ35ht3FkBk4DvoywhuiNcrhjtr7GY7c90Q7uPUn2JZ
HnfKTQ/wlpDZQRZ2Nloh5+mF+nwfuLkzx/9VO3bgeFKhTbOuAu1OdPS25vZNTW6rgsSLNJa64tME
2+Zux02quganMcQF8fDUSKbaLEaFVhwdnmqqFYvZfnVxxdq4wdNCaXa6s9Y0xHWpMc34hhnOQ0ek
QBnei6ck6BuTPNdafTD5VJ1DrLx4ollfxKc0LvSwSMJ9b19C5SKrBHrTYlH6Xn1EJF7e6RwX7cy4
C4Gk7ERSHNdAnOpebC9P3nC91Pn4R/7R1zOPa9aj/AuWv6GxFWkXARKVm5cB125WQ45Wg5qBdbAI
XkowqL7hksIVzQfqG7Vow3TvhrlhkeuqX34wLYfcOLFKPv072/nyPPMQgIYqcj+T6Qm+9jPFcw53
j6x+qavIwSJNoeK2+0RHDe5Y3Wnk3Yx3bTIEn7RLy+ZQVKiyOyMyQZsjKdMtPTDsGP78HyMF8LVT
ZtE9Ah7z0c4yjQ97zr7pwJpNzSdNGnt0qQeB1P50MoLqdQee9lu4MqewZ3ZdXvcEaUtw/GrG3xK4
MButCzmvzU988FYx2zUbGKgADerZggbz6tKebbb+bGRdf1jNtgNBtREX2BF71hlb6f+Q/+rS9W+G
4EP5Vr8ZI6ULu4RR4f/3ghgi206y7bp40mSb8rQwJ6/9MM+9Ict6L5Brr+244E8cAH8Kv7bMPz0h
qCGa7UiZUV+i7odfsGJkm7MxJqinDZbqOBDFJCApfVxOhULTDC+wfQ5oixzjxGa/KPvUy2A92fKE
Xl5FQTug7EAw1uQ3LG0Ud+Xa7sDR659KWRQ4TD/OVNpxPd4R9O1I5zUYwCm1AuvOELZ7VIxDlvWB
oXfPizojFXQ27+rb92RI2TGBo9Zx7v7l+mSBbYRUXuaMGpDoxWnWTj5Tdyu3DBjaHuu9RXmEDL2d
tq+xK+MkMmfYAdgFdjxW9LzhU9yeMqhDegwOoKEVLfIXd8QejGW1KeKBFnIBPB2vLhnsM6ruWxJX
GgTW85Kycnz9cQXn0nDQ44Fr01u4kjxWZpcTLIQkl4j4i2fxBM13d8vNzT9y5KCT8G0wI8iPoRKA
1hcpKWfwh5D9hXUVZOBkCcDfvhC5slIZCADNUzAYv+xbO7/hvNAZ5KM0oP8zUNS+DobkUmhhqzZt
KJkQigrOmrjk6rRVlisN4o3dWryFWABzYnkk3q2PlpI3CHoJ/da30+ur2UHBTZb34gsp+bztDGP3
xb6FD06v+cTkA+GtTEtGHw9P31wt8xis8e9MW1eHfoFz5Qpfbtft2gLFHXF49qQi8742aH2OqUnp
UJksfWKUmrhHe94o8HY0Rvs4GBAbFsMGWmPEqnUBE28P3956GoxMV94V85wAM/r6ezvOXXMCMgxp
5J69Vl/xAQv4samZWD6oGI2eDkrhKw5mapjpNt51dDuQ0I+k4KOFFyInjDoGWBKuXtuECpmFp1vG
t+10V23jr3fhAWnUPbN5MB0LzRrZCv9etZiMm+S729CVvOGWxQfv4Bj7vjbxEPZAO0ERulmhoJ3u
sZYna26JmmHEYKVzUdcFcHniQNvQQV2USsoSV1VkfSipk/KpJ8Wbpkvl/G0PgUxVkhAedI7OGsIB
GuoNdnMQsA4RToj9fLTymIcoC1v0lKf1SXmpi9wmYkaH51N0xVQoBps2bxxPCgF0kaMQl4+4gGVh
Cm/Cg7IEThyFVG2exTSuu8KGSxkx1WIIJh3J8U/OafvyaxmXWd0O17eECugzkZ3M9PSeRxGlcAI5
miMXmM1Jb00oIr6bj9jD+k5JfZdIpAGS7yI3pKT3DQ1FdP2Ng42pG82AxQ6veWz8LwYJRJs1fegK
Kox575PPV8cvD1hz5L8/fb6IRVO+TpnruY5aMGGvaXvE48SHA9Q0zttkC+5lJAYMjo4ZJ5WKyegw
B5cQt7yComoLTgbRkSZkZ2nMGqzLqCsOQtCE+ExQMcMbEXR0bry3hxViL7BRlQwLG5IUXMXx3XBV
PB9w7O6FiZWS+2nMLkPO/Y/sSnXRe443SQV2BemuiEt/Bk0FvzSoZo+Y/0R1VK4w9u/32hpH0/49
PNPJ8S0qGXzdGCIiEG2uaoI4okIXfjWFKb/53VEbh6qW/wIDU45s4Oc4qQ9uvxxtRk4gux1N4ng3
TTi/y8acZfE3dud3yLIIZTp9V9Yzw1ji52HOKrAAJp94K6RDKo3wj5YVY91t7ZPc6BuQ3CBqMW+T
b4fQg9HpI3BCDi2yvPXb3ieL2VAXuNeyjA5mAlHDAmIofNnO1dp6kXLYc4cl+kt5fji1XoFlhf3b
NgXOZDe+7vFyPp2OUy6qt/jEp6v13B6BHtkcay3atIAAZHO32+eGCR+HgsJ9uO3nJrorIuVB1tzt
Gk5lYtBF6U3M2VSs9N7qVsOChqHmZQPHRinz6xLUUABhwT6KtVZGpvcAFPAUMT1Fv375bHOUhPVL
v83S0uVPyR1xRRHPgX7aN4qyZ8xv2L3V1kEilcfus5c/fYbZqZKV/yigC52i8lgtfAdC20clWW2w
FqE0UkuZjNlf/PbKT6b7h9xPNpElVZeRbKS9VhLIO5CVqXXmU8P3LtjkOKu2BD/PHr+oHhuZLHul
k9NhZ5ypm7JYH+T3yPjrtEEENf5CHprLhlcxxTqRlFPvPHbrPmqmss0rd1v1hGCDEUO9ciuLuvKm
PqNf9tWnEENhlkPMMFxX9nZJqBB0QLeaQTWFEaRDQAlk36/yiTQJGgX1Vks7/vZyTtVW4XRoKV2I
dhlLpMhuDHJwCZuI2KxksWCGm/OhuDc3MRFIXKzUdxC6K4INKcDktVGN2TG6H2N+abe/O4jCXjML
PiK2LCSgD/mUwCJicjCOyfAE/QfIkujik40h32g40gfqVn6CFakRTFgz0fj0pQlH2HkPQ7sM1ee9
WXG/fc9jnEhtpjybsqvFszFILa3cQlsfhn7Wh3CCiqPJDYGpiKUke32pSMjAABedc+OLFHCJJYnE
5K/uXjCSOcx3cTOBgeLv9bnQNwRquIZ7iBwc09U1W7ZRFhAB6ieHALncNqTC+ltvwZWeyh/CUBOU
tAA1Pj9f263iyNiiFO5py0RsB5/HpeWwhQ/WDC6FPI2RySPwxkAyDY+nZ/UeSJwpZNqHBWmJi/+Y
iYdIjGmTB1Mdmpbdk5DHtl0pQ8mdp8dgO0ej3Wc6xGTN94Rd/aPcmT3SfxbeVLZ4MPizbnbj4T1b
aY5k0bcjbwKJdTYnjwShL+B2+O5qLlLA4cg7Ait05y3bZKCrInscrcdjP+ll8dnWBFpLzzR5zu0F
lI++azBjqxJEMEIGoII3edig00ywdj7G+E1bPZ+XKqdK3ieuNUey1/8NLs4oePvyCnuh4WuLbbp1
prI+i/gL+5fg4yTmT3B1M3C6xDq+Nv+4E8BbyH4tyflFheVbCTk4EkBQtadtVOmhp2HiO4rMzb/j
HwSSg9UikDeocgKo/mZNymLEeJUBYO/kuWuctZmctyRNJsRSsj4IQRKfgZPhi47MqL27qHu9nlaY
dH/ABeXtkeZjvl5afrYapFEPuaTXu3ntm8oPXJ6hS4T2hLhHzSRi1oBXFYDVeAvFe368LRbl/CfC
3NQbeYKse2tFGaGfWYTXwBc+KkYfO1tvcN3vj+2drcr11XQ1pjtMcKIcaMrZ2y374qANoD2iNyG5
bJmM4Htqm5XiqI6OyzjIdR+c4CceABX7iuH4c1Sd8XuNx/IhGnxqwMix8oU5bMA+GLoyd5cuClcv
JLbaYOx9mfn8Udzw526PHDlVLarcyXbcrpFy1FBGjWGluQA74HS7xJ4YJid8m73S0F1Kfa1A6maw
tlGFRnaKsDVgkOxKuU5UkDKuTPfO+jvMdXXWaerAnhoqki2EwKzSwF50vMWQfaja474TXPE1alWM
2buyRca9cdfmqq/fu9SjTLCRSZTbRr8v6c0gjskYYUVRiXHZBvca1Rs+lBm2jHcVxg944QSCeMA/
zmOE2dmEqW8GyN4e+jAzIowH8cH6mtwaE0xVsx2Nyp8JV7ysygS1GS7IskcMD7YLXSmxvAGi7Ltg
9Z4Sd+tZSFHXXSVMcc/fIj/ZQkQGwMbn4CyS/2QF0VgeFio8mlBiuUYiOtGziE7jLipLuz3jPbKN
yMsOYmctRPJZAIS9aE1p7COSiRMJAWYfFCtrYxFY7dtQA72kL/7fO8nmxZY5D0ealSo1xkPsv3ll
4A0MB3nY9/fsseDvmk9ozL6jsexeQU41M2GKvzW94vTjGnuUdujnLpXFoT9vLZFNTxFrlwMKOFJA
BsVSFPc15iqnnm4BjdwrRxAEZxvkz4hUeh2vetWGqvTUyoCCM9AcY8ugORHogq4XtwY58Oe/q20/
NeAhI46KSOwUDeNBEe7IxLO7hhswI3Yn+ESeIFVUNyv0r3dhuzkbxFmEwDu9DyFDScCvv6e1chd7
4X+es37Hld7O2pNRy1AbB1ZGnSzUmPzQWyy2WejKN8qTSIzTYYtBC4vr2F8xtbp4KDPbUp5t37Zt
nbSoW8yrhZS0gk8qFU/m9pp1WVuCfu6wOByi4wrzTr4qZ+6aIU+wjxxZHq94YqfY+mC1MQ7U81fJ
qh1mNUE2+7Vmy8nTG/Yx1ybWTG47x5TUDLaOx4RqcVUQ9+YgsYJRQm0+gxB4CO5dzBWFc/FHZJFW
N7l/r50pZ2xOifqgneO62pVPZ/FEFW2/b0B0evb81hsW9fJbvZgThTUQ3C/6bbpngukXKtr0p8sR
UbvEMN2ce2rYsVy03nKGj8usBe7ttzeWecE9xegCVTRQ+majNS85BMYRwSmdnEdxV4iAtHYJY6XI
Bo1yei31JnQByhLYxW8nG08I2GSDILWRXFZUOLe8ZPCNcOqKgZ9u3GhpJLHq2HPLQMzRs20bFZhr
Edsqc/mGsLPPtVTvbnNQdBVfx/tbMYPXGOZB4htzJDkkoVPEMGWXb3D74iguzv9DMH+2u8622xP7
V4SZjNykY24fyEO4X52rrxeAo5LgiKkO6OVcRtmEQZ6by3PPmhWGvkcpmD0Ra0XZAAgZuAwL6Khx
rEzyruu8Nw2nrWJVr6WvVrXJy6hWYbEIW/6x4zlkgHON5o6nHxHXdjOUerMzfwR/gKJt8XXAa0G7
eDwafm2h97VvNgWAd4q9bqKnD9p+QwfvPXvPjYXJPQeTfNfk5YAgwP/1NymDfNU+VqNz4v5rqXbg
IyPAzMVoBCcS502o8k2Wl48I21XYS4ZiC93Z9vqtN6DBOxdHXHPVueEQNjGUUXYT9d9hW1Jvu/TO
ym2PBhtIXXUT7OIQYL0J+bdb42g+dTpRIuQAXYbWQebTb9QDKmclCFRpQjId/6uRlu8bEbSK7IJM
C6Xp1h/4Fyzqq8/QjE4Aldlx5aBUfCiMBFh5OpZ6TivXoDa0EhyTagib4abs9EpIClSW9n02QfTj
bN9NTGDNtH5g+e4z3AWIpw8seNSR0QzvY2sPlDEnq1PvFaeQ3oBbV432X+r7wTot7N7CNZtLTWCd
cYov/hwWe1tPVKC+oVS8/t0Mw0mbkbCog9cEPQ0O4JsSIoH/IbbUxUukJ5Orkaqc0vg70iwHKCDL
6780k14BAKN/er55zrV/YyZCXbAVE0wEgFblRlKHNEebbp6f8s7jrh/KNp3NXdOwNmcVW3nO838Q
eh1HcLjbbqwjoZ2IAIhFmUy/kG8j6Q3LjVC/RR2vujj5plAq8A1/KQ6h6Aw3twDc5O9QIKLUzpTt
F+bRjGByE+ncuEyyIXmAhPz35k2SmkVMYYz8/oOQfY1WGrcwJJXO5NJIaT0LRahmaakXtGfl9ynE
sCe6XowjvEhg9rooxaUXxoI9UJjfUEvIeLmRZWTbvD5Yj4NN2LcW1AkggYsYG1afuIRZSN20ww0x
3o0bLkLsPt158D3SziFDVkdALYFvNzvjaiJHI9OQHHTmY9023GqVXE1wFydy3BcRlt1X4Jb20/NQ
Ip6TY+pehcSA91Og3Nt3lotkcD6x+1J0lVfBUwCdzbn5JhjJVHUQBVGti60JRy2NAC5mbaG1OGUv
XZZNbzwJek7bsT60xkZT5kvhwJKVi8ETQ68cUUmM6p6v0dBa1B9HnIgD34daJ8Np5T0l/3CNLCGV
MfoGHW4LHaTVo7jIJjPIeWx57vhTAWQw5AiZRs5X9HfNwHQ6XCMhdGu9M8wJ2kq4Xe95n8K0LcLW
k/v+H1tJlU+1d9LTKgbaH3SFECifu5//Pz8bup0OK5i2qo00Rbjl+sKPvSWMEn2W4VK3AeWSyTh4
Wfgsm6mfKlasmP+BAmMQO4OW92HZcwE7ZV9WdcOzHUCwe7oREMSDoRdKDYv087TRi//cBQykC4sQ
ltflaq87VGNEkWw+8Ao4xdtgCYqsqBqOb6d1PcBhLkC8kiCpzTCUYc1KxQRIqO5sei4p8YGU6ywV
bFuhPFuXoN0hkYuTHCIdr7wgSGoX6aHvydHG3RTITOnEuBnuJP63OCWLjRPBZjVkY7OH1gaC+TeA
te4UQJQBOl9M1UtaxY/1ls58RQ6ziBCqgv1rm//0a9+0WnWQlJOXpPhSyrRsi5+svU453fVx2Kep
ZRng5YokpbF0/JcGczVJ3/9Bi2EM4whOaCTqjx5BdwrNl5nCxMUItx5k67rB8k2iQf4vRhrDJxhV
xEi8k0tMQDluPnl+cnALcuAsL4GkrjrWTZm5ziVnw455YvJpgM3O5jMOEu2OHPzHSho/rcWZ8iCR
YpvQFpXuOyPYZ/R7jRSHJLt/cYAGILjRXBFP8aLo9nhDGrfYG0GQxS89MgraHBhe1cWc1GG7fm+v
Lzt6d6jeT019ND4s54aWEizmQS+gm6smb69cKF9WJ1wUrW4qqtsagaZb7BH8xgzFTd7WunpvMI6d
/w6XxlvjnOy0EOtBYYNDXw5rpSC5Wue5IOj3H2+PA4GsYCvAMYKn2k4bYOwGZKWi/f7HWh3CMC5c
qdLjMu81iz8OH2V9+rAKhA/VoaSli3cc/w+FvRRH/3cCcEKGMTT9+CsWgoTe98jmljHCjbYwX1Ep
X0lpguJy3eyyv2mEzOkuzKrgAafgwgKjOUxt3vuQjT9O/8reniTTaiN8xLqzUPMMpq1qOKrDBZcg
uel1bFuszZY6JX6A0DZgF+nFynAbJbXMjmK+ZlL9eK2J5TW8+mFLlmsNhL8og0wfV10XCi7yCW3J
Hrc6AhCKxjU6Y/0DqR3Eri8gdkux18Io5hmjbeHUiuApg4uJU2SChjlaUlOMSkfROdu6/BcvGIuF
7qINgcVxvBWn2GTj+nJtrGtJ0yoPAkph/htT4FzRRYoIrz4wdW151tO4SUzvMvpnLE22mnzuPc/j
M+hpRcWKveOqgD9MsRw46nuUL/KnMIjdUnAyb+YC+PJiky2QFs0zdUF43E0B7AZ5kLH6CKWX4A/o
RZiRiwznZ/4+A6T16HOVunVzRR+U6Vl6sTCnJR3OkO3sd662bIta0WR59nWqwPmwoofyKt76+SIU
AQxgx6Wq5grD3JxS4Zojz/UR/TIuSs+mZqbuCNH/Lk8foWUY2R1bz/zMJ0h1xIjO6vsyx5ZsXVdJ
SclQdFYPmkeYw5bztaShqry64h2SvMwH+GO8e8zsA4oQ8ziqsZvP3oMbbi/qPGffr33nuzkHkE6O
Zb8v/ttYMHWOl2Hs5Cv9Urte4yML5z1oM/XIaPgqvjRdFasZnp7s2xb70UVLUjqiupBsTJn2yLCo
LIZQiwX4YEg2umalxlMYsv6uWGM2Lskb+Uch0giA9a3p4OJ0VNSyAepUeCY+IYHyGmg93svTC/Eo
jzy12yerC4JVYCgWGa8L5On9a2uxz8ZS1785/qUV9di0qYWbrkWpjJoQ9aPTd2MAAzdIHKptq/ZQ
DRHsEd9sHuCXuRfFSAr8rT6rD02+i8eWmAu28z6xFgOwCB/1jbZUmWUQEK9Um0Uye3Pmmt7k8P8A
1hQB6vz23cny0L2a/PB1GogTw2Hx/1byuMRZdeCczcDoFkAUavTQLBhmFMZHl4tdEtxxQdsJ9iqe
RJjB3T8dNYR8ixa7VaYeHOsAputDaLTWmCOmScLJrn84HIeIRvmrbFKvHcg8Ho+52uOWskGk6IiT
nOSL+b1l1GCw0sc0IYikwymYQOvJKqjtw5muoso+HZA/HXzqFSpGR1LpEFXO+Y5qkpc1NUu1y2gn
t//LoIOim541wvtRRpEtYtCj3sJM8DaF1NoJ6sB+XBc8i7lYoQ8Ia9/c5JawbHJhf4YL8H/AGYCm
sQ9yV5dg1vkHqYX2EQMjIkP8BFkGkpsL70ILaVP2Ek27Cf0jRSvz/r8IrjxiIJnvc0X2nuzQRTKM
VDNvuj+17FCxZroLNehsdLDCPFsWAgliTF6Rp/oGZqmV1oVE6tP64rkt063vwJxK38NjJmKmRfut
z3f+smiKR0dmVcIeX17Xam/x9khDuq4kEnAfUDZ9ISZRvTx+wIFRQ4e0H/IwfWRot4hmJMq+tcPI
OVjD11mWr/oKHeyU+wdp9Qagft61s1OiVHruoLFUcGhjY03SBm7OInOqOZTH5SQDRHSVF5iLOHcQ
pskrDg8EhYuTBesLnsu/7l6+qp+DpxZtFxgIQm6IJ8z1Er1D0zfZr1rpRJNiI8sMFHasE+v52lWA
Ugc/iJpp5PSWnPbJaiAectMEwEmNDSxPb7P9c1f1Xm0j5blsFw5gTeOkLhAz6wDXtSVTTUxM9Y07
FnVBVHYttecyOsvKO3i4OaXcimNMb2JdzTwgpEFhPi+6hYCM+KOrxxahgx0hc/w6O8PF25NjMR/r
EtbBP8Y0ka4Jr0nudDhIHiN+oOYl7B0qUeifLf7m6y1rcy44Iy9O3LNpA5Q8F5DrIWqqMVjBbO5j
RLw+kE0CzKc1HPY/+NBtAguykQpZYXyuyE7t5IbCxZYgK90tfw90qAKf612evnZKlBxt5/yNc8bm
MZyvYLyXtW2Hj2msgUSzoDq6ynd9Q6NiF0QLFDTMp7yiUHr1xoaqkP+NGN6TATsF/Y25lRSVVL7o
KiNeMdW0lLW4PvLEaC/9QxOXhaCVb07917YFINcqM9mvYSKtzH3DLPTN8PQHkGCLdBL5V0VUXKwN
+mBVAnDxP76/MrQpKskfg0s89d3+svPOaWqpe8wi9ivcLofMcYPYj+QG3MuYkmp+nnuxkjLxb2v+
HAakQH01bi/rqtYmjFUfynMzCk9x/U/UD3KTzU0gMieYiVsWvqjyCcXtKpAjPnZN7YJOwQgcJr6e
DVvbh8Tj9vf5vA7ONmLo+QFM0qh66yH1Yq2Xy1oe5O6e65JCVfYMcCc3+bCe63wZAiGJG2Opmgs8
A6iocjyzz9O165MH0VzFNgD4AkNloTENvKk+mfusFhmDp4V6HifJaIyHKICF2cmizDdI+9/1h0iF
dtoe9z5dpzKfIWjTIJp0lVE9I6nuqUMKqquijc6rArUlDOF9TOOn0cD+Pwp0IWwiECXRMwQLvR1I
LPB+qEJ9TQXhMk4sUAaQ8Sb2/zQhjMa9y6KRdX5LFSXQX0nD7QPA2f0pK9UtKXT6ScqjKHhc5YTi
Ge5ywFMqrl/G0wuvPFlVIjG6kNTow5Cp/GkjH6gZpIWG6Xcr9jN62dLBu8ir5I3xRO9C7ZJwIlqE
6Nf/tCrx2ssrLLai+0/clj4kLalngDb3w8gblcYue2VjobM2V+7/wRNDSfCxenBAtdzoX75vSoGr
ndhSmLIODNJeg7aWkjnqBjqFoMtwVN/BuBhFysUNo2hiUQNYGtP8uCGkhYFLSqkk8k4IBaRuzo3F
klzZnqOgDe74kAXZpYbg0aRG4rGAfJjWzJ1nnVydkBosqn9Vk3FAMrjjbdmlyf6yv/+piFsfpoiK
MmeIr3AJEvHXm1+1RxqOFTEXmSZnOnUA8LWu8xmqHRG+o/P7jjaRPrtm6C/QQLZqGJSy6w47Kf46
BRLmECrfqTEWlXez7/fjx/axoBqWnFdwW/07UP/Sk0GLrz9GgqN547i1wFECjjPUuNXwTMF4WXcO
zMUTABNkQl/g1OEzfUbYS9TSYvVtFCt5AgNeQPEuEesQChZh8smFb+AtvORLVc78NtfJrf+S8Weg
W0xK2lnZozU1ScQqDNZvPnRrMALdneqQNbQB8w2q5dvcI5ys1feTOdGL9jFY33xghcDKx91y7gpD
sP+fqfAJLj99un3WObdU/+PpJrfJRxpTp1APjvWrxWybMxf3/FCAvEWKQjZXKWYNln2oJVDrse6Z
5YKUDzPEAzrM/ISb2q78P6j+mFJRSH+3Odt/+pODF9Fn3Pa7pG6n5L+frbkH5r/Y1fpVhu5i8Sia
sDE11qYqja9gyzfgl4l+LxNUBolr9eEUObDrZMA+A+m4gEROVm6oCExkMKEzX7X1PHSX4YnODslO
m4ZbqhTcyV1HzjGKAj9d8HN29OHAIIxw0wwhZK5fTnpKko133tA9ocv+9k8zHs0f3QAYFmn+VjIe
vM0byLG24AK1iQ0ybsBcFKorvdlguq7onRkwleX6Q0KssP5aYX4rGuwYnw8iVoqRJgBVZxrpreji
EIei8zTGPtQjHitqV/rsaf8SPkDTL80LrhaXmj5ZtLr77qYjn1C8X03yunJdfvVQavzipO0hHead
Tgmg5WHkMDdnW4qIm8kW2IjchGV9km0oN8PNTw4MsocJZ675UKne7rOSj7W5Lf9XZvM1dYN/DjQ2
QrEzM7LoSMPHtC3U94uuCuIVq/83VCFo/CXxT9XlSLzBbSRro3L5IWcVM5JmbggUHnZgRD590oHo
mRz6aL3TSOISOMGAQxpTcFTZ1H7Zfa1yS9CS7LCSTpcxq4QnaFBJYwKvJBhDY9mgJ4x53gmTtBFn
MfQvxtBU4hNEmzbYJ7w+o6MRiEnMn6IQK6VwK2Rh7Hy8d/xxF5ALO0lDdaELga8bCYdPZ1u9hDp1
yJqCIBkUPDPX9RgyP1FlpMqcV3XU5pdeNIB+UeloT11MSHdVa+70fVgabkBCLijqu5jrU6rR1ldd
5Xjs0DIgFSJJ8Y0ArpkM50NFp+2/vUClfmrMCCWO10tSiXrxtXrUFpcTkbIRivSuWYiuqtA62R6s
qyyDfaBIIibVUE7ONxFe/LgB7olRWd1UPPqoMa0eB+norBG5Law/OBZCWEimeDxIzpG4BPYg0VzC
bSW2Wgl9uTt8W/gxhyYv7PIjJPKweFNbS6Hoke+Gjr1j6R/1GmaejGvBac9zsRMxHHhWV9irEpMC
mAlgYtrt5e14WPhwhQBV/Q0/V6BXuG46cfS/Yp/jz/FBsFop7xvkyNGMVfuJgfofk7INgBWwhYWL
CLfwgfTy0VzjPUrMVrJqzyNMwKIdKf/xhXA79irbPyX5qoYW/wPC/J3w9z2WoI95We1kYrroCORc
WH48d0Wd35gzBNiF7PprMyabjQk5qTPRXflHai8sWGgy4blBzqH/rz99b6ao8E4gsfHQUTlM1x0y
Vd7/FBRGIhYpJq7aXaqwJgc0E2H8UN1N+IbEdKkrOO/ps4LqjJDI3g00TfJrERU0FoARjZAkfoLT
j6MHa1kfY3SANGQkrLo+SuzcusfqHWDh7On1uKCX9SCJaZBXhk4qfp4ZYS1b7gEfUtwYYXGugjpb
q+UsfeknfhCKHRvwnYkUQGofSmdwIfselbq92DEMan+2HQcYDaiefXyC5N2qdk1xXHmdFBba/Kfn
ToWaRNsLrxjCWwxhkeL8w26c8boHynypUVsa7iOKysphlQackQZMg1lmzdRGFX61355TbhkyQ6nG
jBWaYlQiaL97rhuZgq69Lv4RGHcZ4ChCyeyIHA4PzsdLyk2fU6hymQtlaLXrAi/QwIV4JU03MFzf
zGRe1zVczlSituogMB/jgRc/CmQ7wB6fGnMrmIwGyb/ynfop6zfaGCvNkn6z3NBBXZOgfHYAb87k
ExFCxmMFuLR5w9XsdPv7+py7PtE7LVOVytMfXST1WF2pwaDIk52HJJGIgp5pnkNXS6+cteE9WlZk
Vt+3cx8A58zK1hH03h2lj44ZjWAjKUHpaYuqQsYqAMCE33fV4kWctu8Fs0mGOtrxDU/w8OvV/N9N
fstCkPZ8bjBWrtNBBH6WzYT/vIfoh94bsDoeI3igRynNyfsTRpNoNTzp4CrgduDBQ1Puc3TvvPDe
DgSZd6SUNaTx3S3sOvb/vwxCQxmrL3I5auleWdAF2ecrclp/9M4ncCFKHZie4HDXS5WOxo4gEnI1
JIhY0QfwE5cPqMRHyPpDKmclJID/Ruo5lSc6Hfg4iWlPDYdnwlK0zJg740lomAJRKCFjhwEJJnif
iTn5nabbZa1TOXJRojOJI+FtxGAdNSlzYVy2tuql6yUwF3XChJgQUv8kQmOFdyXd3V5Db9vdq9NX
DKv1xoVup9PqBbPRCjCM/fGHVskolpMHft9JWcCAS87Cz5tV7sXi0qlvn32EeaudCGjkxfcu1aXr
ZscO/WdrrxXgAQdKJ6gTk82B+1f9fka10mExYl4/PZYW7kFVASvxtNSZwPAryXH9/TBaeMtpXhva
7rQHTQQOJo4SWaq8GxxBH19FWFvnxYddryI+tW9nacWH0chbIw/Nw5SxZDXLGCzEMmHT6b2mp0Fi
ZX3jNk/afZMBL7qckLt+rQsIaZfwct+WvGJOIdDFP0RbtHGP62f+n+wyvm3SSwQwFKO7JOxjMrtR
tZGVNaYJIVfuTWk2F1MG7HSR38X9zVixjFCBL9tEcgBtF2ehc2STb0u23SLUaK0FRsvE40HHTcfD
t3tN4PhNFkgJKvtqIw1yCVw37fQhzI8RgKeCBPZejS5B6b7j40KWfR90CXgG6oxEe24jRTmlgFB5
o1jYHcjrfYfr2en7R5kgtQ9BNegw4P+mKZfAMkyjCfN1WRdUJVnfH/vGII+odv6JUW/lKAHMLgiL
dY3c1Gp3qGZPP4ntqmEY+qCny38gHV9FiZKydesxWlLf73yymAr9KHOyAx65r5/WA20F39fvby6K
F0/E3euf/ofklGsqbHM3xUJltfA5bqM29C1qE3B0doGvjXbwIqwok+2eAMwq40QyzIw2hCHu5NCJ
WLw6oIZ4oEirstN8pbyhMcDvDY3WMqx1Io/2dv5Yv5rrntGOWq6VebWgTh0zIqD7ipVKaS6HPDqy
DpBMdcCwxgPaA6VcyWPncMmHbaBvhLdXe8GViqFzdbRVJuunOQjc8bxM88tNyDLWANXylFwRTYQm
08TQhOvRDllduQOxP98wjELYOBQf+j8eqI4S/4GwxhacLRZvaFjD8JLwpUl7LMz9yV0gO0gVMqsX
D/UlZ9IOZ582C8rhbXgspSsHmAwIzPeihJJVinRuJqs1a+zXmzrYAydglJCDGrCyEHA9BIdDm84O
9vRVnJBDqExgjtysd8+f+Yd5jhP6PHBi/jAM4CJR1AF0voSOLe9LLJCjapqeN8V0Ztbn8CTrnGNd
02jXIxb+96Sm1p+uYP16DmSamGDuhJDrJvGslV2MCK/Y2yAwjlgZ2fzoTMtNpaNgW12qY84JXKhy
xrc+0RjGvGgnXDmh5JZ6zrWd6Qw26KDGhHvtXOlvQSsvpdekwBd64uYznJD0c78qMsp5wyn0l44Y
z5ZGVZWjBOWdvNOfOI2wStTL0DiFB6uIdnEgHo/rawY4kN1BVUljdgCoFr+k7iQmQE72HRscmrql
r9HmV7kW6lr565tnfvPjiw5btDAEc1MV09KyaclG4D9+NHXHNmKB1cj2rAvdhL13P+rLlD+91Nis
GNyDqrNF3uEDFW8JeMmxUddDH4Ws2LjzTtMOHVWhi4ukIL/vrioXxR/g04ne4ug3c0bP3mIxG+KR
x3bQx7bbj6oXgsV3xRbLWQd8gc+YrEH5KjnvlStSjjk62fwb57BQ5U25fTk/pAMN5kssZGhQjAy9
4bPT2yg1Mm3YNMuTyFOAVP1QfAsFPr4tNbbfO81GrJuoX957IELd5MFUn/8EfmHuhW0U/EfDU+Zo
+smoiiF6uQklb5fT7VriqHfm7v24zBvtTHFjckvxaUm6f0D7eglPYGwdz7sMqhDrXvJbjhgrKc3E
EZ7+xUHEeJg3Ph/dPwALhJcD5qBW6SL8V71wlZPfVN8D1XbuqS9O0AI8jWojd9yOYFcjYDb+3wNZ
vDgNUrziwssvaWT5+TiFCgnM319MvWQqVbCaX/l3+DnUcTwEzn5jtiXLcqzskIzpGP7JBTnrjkVT
Uf46hMtdaXscYd6khyaEMCYOz9CAKYgM0H0NUcwR2vVhGc00pnNx0hmpERFoF863Pl1GrTB7cPQK
WuXpdbpwaU0D/iaIQsMK/rcZQvBFQSOm+h82ZvIMTiCEYiRiNBkBGrR29TMibwXFD+2jbwRz8sXs
arTCDA0ADk5B8tidLvNv1caGhslqIIZjD4y89RlYdtQMymvf1ZeN2pgPT4+qqUv1r+3nr5qPf1bK
0ZvpP/YxlFCd4MJ9nT5B5wmQrU6aurCeNQIuRtAydyzLRartpwbs4EMGmbK8o51mRPnL8Fsy5/Xc
AXTgZ1K8LW+y9V5ZEiL0Z0KJupt8rJF3ruTFLLVhXhmRlChlWDNK7djHhy4b/41VxYrStDfVnZMS
ViAR9MVT/gmROwGPKnsjlF8odzEVSh2kMxVnoRoA19CMHWWYN9iUcqhffdvJDySSDorU1YKgQnCn
F3PC/b/wUfdl4kZpyQeEdc1DguhJ4aY6N7g3RcZxv9b7oDpacI0fYcankeYzdh5g1QeN6xowBQek
F5389a5yNdCPMXZHDfOKNuPozyZbaMnhVSfHA/1JRJst7yYRbb5Jd8UrOw6VVXo7cvsfVeqsO8Ky
3P8rYDb46Sa0x3478mfotZQXS6c2EdEqgHQiZwDrWwM/M9l472Fkr8A5YuIDnOPkWdAlqDDswQUO
aia2iC3QA2o8WwvhI/eNomtUCsHhsIvOvn+YSWx+4uztgXDA9TBVs8A/TjET9QQr9qEEknY8P9zb
bJrgr/yW+ozEs1+haqZHEy6by7ZZdLLUXfAMs56JxV2KkEqBQbrlEjfoo/RfnJQpjZVSQwVYJXQS
xgsGFHEAd8G5LGHbNku4T7pZmS+bjM4a+dwcXN6k7Dun2LpnYMz1NUNgk2RdbsbD9yLO9AwNJfIr
OyRbk6Vn0RXPpnu1S+klmcBysMh/PPWPF/1/7LCqes0WUalD6pqAMM27aFC+6wkwvAFCPqvh5xOk
sgNQem6uVpFBK/1Ch/jQW6vb0pLGbXT6RMqnHLTLcoTIRhEnWpHavXuqj3RA/6agLTUzlBeknV01
HzziKaxBnvYm7sqnRZRDB9rirnJJQnkm8l1/hwf0XGhRhAvjxAJkPMai9gmTXuansMqDALqVlhRu
98BhlLimTNedGJFgYkIp8C9kIfge9lYGWQijLhdr+8HIl8SAj0LHfRysCuuCkUJE3bfBWvrXvxpV
iCH659zS8M7O/+hE0hs1NuvPL7a1si7smM9znu2P3HRIrZ37/iBscIDLqyQHLzD4uGXRtvG8JrFF
tDrdfyE64V6q/h8JYkeQ2LRAJ64WOpIxQ2LMwTUkYXs2e+sfMJow+X4tjdUzEhg7OlTxFcS0dSaq
pz7VKxpuLfew9ATdjvfVkYqeK9DQJ0zA/BRTdd+IabUij+ZkqxD/nJq6UEehqefSCHHS+CzFQkxA
E0ec8CS6ogC73pex9IM3AtMyn3SAKIrOtexiSd/4OLaiGiQxoWYX8KZLWQjGfIt2HIVF+/EV3iRa
k7IoujDRMn8V3Sng8NsS6KmlUzoAm3vIYde9PxIqSozzzDTQl/efPXkAHjr+h6+4dmWbjpoZ3uID
AaywLnKXl3uxZZga4MkeQhUW5XCKz3Fg1NFlPxVFNGXz496Oe3HTQ2gpi1QF9rEZKan61MODqOZW
+/j93srWwwfjNiu8BmXh5wF87TX0m/PyNMK5Zeskwwer82CZSDVOS9gxS6gCcpQskI1WcefgRZgE
Sj9oxj88y+im/zpROXXo+DaS58biz/+8CvQbp0L9841LKMFY+sAzY/7Ndt7yhk1jNFANvOwVl4/H
gP2kLOMGeDaWXZStZ/zDnxPOkDoVcT4HSFgXKXeX7E65n6X/h6X9kCm9WTQF0SsrLi1L1eVJsZyB
CLW8VyMPh8snhxr20rM5Ms7lnhinhFZLYfzSfUOBrjQGn8VomTdvUdiwWbCFpwpFUqLHY5png7gl
4//27TZrJENwla7h1PKWiHDS12bBUrWZHCauFrmHzpw12DcwpYpQwqHLi07ly5f6l72uKePbc6er
Smb2qSqRvfyYlQmkr1m5fPCRfsSTn8HKYLH7lqRTparUDJgTpeZ4+rTXqIuiJbHV5NENYTQotoiC
Fxm3vE+Fp6KihmMnWExMFNSHjkqonnNt9vTeEOhwrEDrNkSHHLaeG3llAi+Uezj19/7q+BreElhv
jBvTlYLFLo187HFEZjxUzYcWQaskvQY/vIEit0umzksNwScRDH9vdnjzQujI/+sNIZPmapaFptJF
YB656ao8kaCuVgyFAJffa3Uax3BHBoyYTT25dgD/qYTHDeG5ZK7cPzHSWpXUu+qaH/DK4pU2iHID
AMaolVGE2BfUUSgZ3mfVeJfuTMgu1m1m36a5HaE3doRanXs8a37iDR+4iasxlBMxPsgdg4CaRh/d
k0ARtP4PbTWk8ULW9mrWYf5R9WIai+I6J5iWgPhCSECP3sAH/LI1vgvhZb3x6YBhHPl7Kga2gYeX
25q0PFb/SnzDvHty8r2wzVio8wWUhl9Ln+4g1ppZZC9A473emxWOl4ZCvA9C/xXfNCOnSkhUK1a3
ieep4Dp9+ujIzWdoFQT7EIrX4uiVJgIlKi0L9TBk/zVOaD5KYiVi0tL30+eTC5NO2zNhMsLvwkBt
wPVNuDSpOQs0dmdM3w91WqJ0BP3j7MLl6apQf0lmLcWWq9AIS2BQ/Awjj77+MKMo7sADgo9hW/qx
osJxW3smhwQGQekn/2Y8nnwYopvD7qbMetsCnvA9CaghcYYSbsFh1NJTAHrHEXhzelRIofmuFpnj
byFGZDh1JW76nmaFk9T43O7ZXPnJOweYuTPW+/R6sN7ELWU86BQ+K/RxPARDm1bxQ65j4S34b92g
seWGbKC87PXcjwYX/eGR7DcliPnhaENpKtijlNHpwbSX7tBHKveU/BKBFk5ricACyA/rrAJLEUGW
X39ggX0NxbeSEEaIsu5MIoAZgzom2Hr9oQEztSQ+spgTT/rHC0PalMHNjMB53s4D28IyR9q+sJsE
Fo+aVfghQMPU/qT233aXjD5WngkM7d4Pr/B3Susn7L79OpDUY5ISrnWqxbMqzdWSEhpVjq9ncyEn
EFccOBEPbjOX9wy59qm/HnBXGPSYWOmNM46HcxyyDRNSTp2jkPyih/SQSa95P2+iyV+ctOPKtWRP
qfYO0CpxilbTU0tw3Ws9JSxL6HZ4NohNFmqns3geTcAhuqrTVthBjxgV8qSCZR3kYi1uNSpw7qIy
m76WCRwQGXUqOkhLeFJacUT4y0I7tAwskWmzRcWTZ6fjt4Z3UWq6C3qcPWPN4N7hW4yTVNIfTVJY
7P9ukEjGHXJ4sMtr8zTNPiqkruLgMPgQ7nEFK9xjBIKw6O/LgwmFzcZPx0/CIkqfW+mo+RNWmx+Z
pDy8ZYw13TXXlTlPYsuW9bHi/Kq/NCU1hpPm3dUehoyt7a5BjVPstNtU56xHc7RLD9MXQn+fhoyq
VBjmkNqYkfVGhpYFtAyDJqdjSfwAm+5xDcAq7k9cnaJ6oj1E8Y8y5zhhq9Jyl3ltUbF6YIfW90BN
QW1emHVG4FlAG1GUwJxTXhQxS3f9ZFzLFO7fYmg8mxls56neKL6OKGPZPZspkRNDkKaJncQLZ646
AdoIBKpMrd6aSq/HUmStgnPRE6bhQA+p+kkKcT1S2E6J5RoU66yoHkptu8FaQPppqKLBpAQCfrep
naK7mHluaqXdATCCOQHPVAOZSGby30glpACfHv1QSUCOX7X0hSpB0za8rpjJKnzmLXl+9KnyhcDB
Q/XEtUcvL1L1mEDIbYaE1rkRmZcVE89gqLzqdb/Qib4d3ATwPon67+cp4jQ43w2Eu2FVYxUhVSD4
Pp92AVeWpU+qA6Qkn3sT2X/api/87TVpctwaDjIAmJTLzKlhw2TmkX9cZXbM2h6Ynn86nM77emsS
mEisjYx+UJlS9AxX4hkQawBBnPXl16SMTka0jEXUNnIjhQWve40edgyZJcjq9iblVYsU01FlScEt
AaQOdh7iwi3CvqC0oN6n/g1u8tanO1kxGv/l9BgSFsrASmyKTT9GNunJKB7l7NxZxOwzVctmFKK4
Gaz75cjrgeIeInLk8G/vCg24TmC53ayDOf1LmFCQe25RAbPOGFzs6RO29DuZiBZHSpDtdxCF6rKQ
WdgqgckCv3mJtztVndYcA8PGc7D7JiX+pVO9jscNOadlfxi986KPwgLta86l8o/ZZ6FfjpyBhLhd
Xe9PrKD/hKTdCSpg2dbbq5sFjmXTBfAvyUfe0kC1jKfMpwic6nvfzMhbDR6qavKAxF6+pLOXPzOX
hbuz2MRQ/s46dvxD0EK0XH+eD6i8YetnG8dYwSTSIKQo2AIr2AliuSIx364hZnIScscPLnhOM7Go
Qs5A+raIOSMcjxwLhd2OJfFHgZ84O0rphxYaWUpP71dFyh1hNeHOBCEiz/c5pGbIy/jkxXjbltmZ
v109v3zeeXFJCyT9FlwaCtm/mCrf/8fkzFCzw1Vi9FtRCxOm29F45LnINNPbb45AbZreUAu1TBBl
8WE4ollzA+qHxfmX39iSKgpQ12ISHMKVIaRTrqgQ0ADzgihhSyh6CWQ7DwsMmSusDTGucIJQ1huK
MoiTqPS+fvLl9nkeKrW2MC63Smgw5cJmdezh6jvX0Jdthzdu4uxfPogdF+20jq/n7njthcJz3XYg
87hbCUJdYfCoXZRzuG+/qatLhHrq18ueVtUd5z2/r4o/KyYanwmAmw5ynbMGv1RoU8bHRnK2WRsG
EfrHpJ2UsM1KlkU2O8OwiogEwGS2ms7sA34eAeZJNxR5VJDmDlEmNbrvcoQ+JO9UHXMaWFie2zzb
31cS1bJu6tiROWM1tN7Kp3ziO0bHGeac1pxTYDYfmwjiGSCXwkJxCjbsgdWwIQPn3hpMrekUQedq
k1JU92f3AiR0R3OLZPs6sj2LBfGKjmH+gQsn5/f1kfGt8i1YKugsWxnroH3vmTWmF6pyEGGv6KV+
qglG0gw13VkckdUrz+PIeKtdHaakxQXbkNsY95nkyFQjBd2br4KLFzTPe9qjufGMr7DeB+eleR+y
K0/RYLhlBSDL1m2G/7Jicr79j+8T2gQoswcd1OUbIII4cxMYnyGgWq3BD09tqKp8IdBO3SvcNLV8
ACKOzYRJXcFQVUlfp4hD41Y4wXb4KU8ttTWlMLm0hDj8zOROVwMeZoMA+UVS4cHrco1zpMHCCzyS
G+AWxWKpuYzCzSRBaHWC6fmogi/YFGeROaz+UUJgOQ5dXDOmPEBjKo3L+jMnHlLhgnC84f/9m+yD
yte4YlnJn+NoavK0uHEMrXd15TEUiAfj8CENs5iB6nbGdIt0s3DdjN/uKfh2m/Zyurkgwlrcexds
Jsey3LpBOHrLosBUxsmcxQDQXZXZOc19YkEwWvdY3oqrXBIyEK1912OMLTSoY8AxjfOlM3UswSoz
n6Ah9J2a7jsiE2jLNhgG8O0ue6EIcCzSQJcWdaOBwTgOOQkKc/atD0rRc3/I+yQksY2qN71ieD8i
4jxBREc7DgamjdGwwN9RWPC1ujLuTR4O5jQ4beFKIn+2N14hqwNLKNgS8Fx5b0wov4dLHMYF5vwx
2T9uUICPdSnaxFhlz9DSnY2MX4N8Pe6PyCCpLKzJZ8Rhh2YaTXdyyKPa2WQGzHK2apsWzezwAtQv
8c6X58AYR/yTs6x5wN+8mrhX/m3ps2oYeioKc0jkyeGKUCzY84x/L9R73kAylMrZAAugmT8Ezzwt
S+HVc49Kc4jofcvQo9cRmxWZI5o02BYIB258OfUJJuBhMt1MyUILRjp4Fb9gzSkuyZ1jiLraJ6Qd
Qz71dCWuUGaNExwyjy2jBTEHo7ON0nPPpA7ShIgRKmy0F6QOE8GXkZuEA+oLVjIaB6iFd/UbIpwQ
GEsfoeWEvuWtUF1fw23DJ2DVDg6FAZiVrcSpueu5lV/gMcfsdTt1fZtc7nHlB0l+F9lDKWPRKogz
cHj7+828PupxG/Sjmj6ZQx1O8qjiGVnVLnu8NftVNCZtVlIRsfUPfIx8iPx4Kgk30En77I6DxmBo
SdXnTiXkL+E1O58iodYlAARIlHJieB6bWWGOy4N2Pj1EtXLSHCHXh/1Rv6X4OvyN2YXTpFRgeVA6
6sB22nAIm+Iw87C1NfCJ18dnLV+ag6RlbBB0SmqrkZPerncaXk6qEtVA4D/DzGJ6NvQVsC/WjGrh
hvjA4lhq6/shUkLn8IFNTkxzDnjkmHlL6/LYCog7bzcLcVPy54h3pvnF9wJ9XLHL50EK0JVZwpha
vWB7WKslsEdRqYd7p74MyUR2Hh+n0Gg/O7espwUXCnUAHl10reIyJfVufEQpEKtEmJJF0HCpfrfF
W8F1cNC/3XAN2UtEuyLD22ryy7ZwLXXGwVTSUAJqJTL0gWpulv+JiY1tzAprSvWTSUVFEgPwJ4PD
1NSrfm6BYpbal6RZw+6PQHHsRuvEJjvzpaZU7J9/4hPY2ox6qtOU9ijPv7Hsr8xVFvAfTqWIWBDW
GOj63h9R5JEBEVfllsQbHlpWOCJ0WPshR7iiJfaOExcCfg+kvfWii3KBHNTUdFrRcMltKMupdiCG
63t9sDaZ15erNf2qpYkJ8ZOWxcI5hT1F7jA3nhbNNrP30tyDyUoc6VA3cz9rRl2N0WlXb3SbQUdB
BSAcobfcqzT/h2lGKoK9Zix8tYxY0PY2CKhVes1q8EWHIXP8BHqXnjk0yKoZC5jNLe+NzLznGWvW
6C/vxsAH0JYnE9+lsxx26SJS5EdCGtoALzSLJMB0sqgR+5RRUx5cfBw9AwIJvOGVFf69+WEjWp8Q
qAVWIldiafsh21guTC2iZhDXyrD7DcD5Stj2YC/3CeDC5eZpVNssUPoryH24+VaKrt53a20HGyU2
EK6C9allvrO7ki7h9P0XXYTRZNeka9bDc5erqXTIQXgMCqka14fQRAE49gYv9Lf99+wNT0VRGNwt
3qZJzj9cFtXzCF48G30Ms6mtshNSNJp1FhbYAYPm9cUR+D3aR3TF9SWsW4HcKLZvvxloXg7+PyUA
QC76351bIMWmwecMNQTaxVpdrxOz09xxomUeUWh/UfJIsj9nU6DxqZEF4JUzkdTdQaJxkSM42iiB
3MZwPLwj30uVIv6N8b56CtHGQEej1wHvauzbuesqS6rZEIMspjHzdv94nrUB2EPlY6ICOVTKlTss
5eUAjHLW+jpt6j5oQq0K4/qEt2YQAKRe9g8Leye+BaTHgoVmHiMkg/H2ZYE43In0u2h/dprvDaYB
CpzzQNsWTVSBVtqNPAjd4+KyBZMTBppqg23eLFCAlVtKms9dLvNrQhvEY6KPgI2s9ZBN8x3auZHu
1M+AES5rz0meAbWJEfvZlFTl1sgE8OTieJTaIDmB6ngpijD8vkNPm7Ozscduf9oUxRO3qkhiV+QN
FC+6XMdFrue9f8T5bLZJVJLRAx/x4s1Jgl41eYn+uMaOHS1eMYP/c4YPFpgcFiWGkxufVkMNxuld
wa/hfHE4voHsr/1WXjwAWOHADhRTOl28xYEUdjGzsC0GjOG9HNF82vjobu7QSLv5x5S93aHjRP5H
qs82x3aWS7pRdn8QN8otdhgcqrrZXb7URdRjdIMtpDLX6miavsY527zXbnVbeWoTs2glGm0uPK7f
xQkVRP8y0Ml0i9Prtl6VWF/dUmWXLXhYlEo9sA6zBm1+52FectUOCJMbCXalr2KcCcxTaAMtoN1O
LO/16oQPUF7PMa/xiFw+RvQGrxtIKOjQas00agSwFLCv+oFtLhGCmWhOEWfhADRtsuUqk5bA6mUC
7DitWxktSLQvpze07Gf0E7ZDHrvrQKKgmcKJ/2I+2fd/TtSwUWVwW6KYNHckj1GJ/NFaNJrHYtDu
ekWZq52F2Ci3tFkPUw3SOnmSnJYgpkzIOdZ/CcQ70xc1DPvQwkedRV5q49hVPW3iF3LgP/3KnVVP
8S7j6lD0k3ayvP7+yvt2jdWwtQRoyM3sF9YJCIGZXZ2ePhf1w3Sjn5Ix0MzTAquoIJ8BUVpyeHDR
5pnEzEJY11W1HP/AOwWAWMB2Tg8UQ+2GSKuF8Q5jwMbL1s3RrwAjIuQWeBmCq2jtCpdOAIFqY49e
WRLxH8ileBsWptIV6bz8CwC3/JChVoZ7DoAo17IDBLNrbtEGsbMUduZPZi1Z86ndHhiw6WwaZhNe
ToBnem6lNGrAp5t7Zc4EvzlPyiK2oSmG7YvadC9B5cjzJNIH2/s2nOqDeq9mDkm5XtiGMTdtz1yP
bwfCj5iXyFwuqpt1JKIlNisE2OMHS/Lk6C4BlkZXPuykT8DIyCwx4u8ElFyKHh4vd0l/JnWD9Uuq
FW1+k4DDr7kxGdxdXB0oKTwsuC5Bljgyho3NQS+4Dnt0KrV38WjtBuj5QK81PIS+jUtKcVSo+ybZ
ZS36jtSzYr7YV5Y7M3VE2XwqOWY4TIfGo/52rt3eQzvE3YrIFaCxNZ2hfspwCF9UqX7GFw4MO+yP
cy0I3dQXK6MVjLAB/yHCWUcQ8NKLxOPxGYDOtb/WV8XkYsCjasYgwmy6aHq30Bld63iH1jtOti2P
26h+XCFJY0yj7oWUoWmUD3Bxj4vlji64TcK14jSWXZXlcbFm8kCkUwwn4GGfUr0dI927HOphyNig
AKzdvkTotQ1y+AyXYZVjAkJ6ki2rVnSg+CFukjciIY8ZSLuuSYUAONvgDgi0nmXFBAiWGbBz84Ek
BciI+MTnZp3buecn/NZuLNSan+2MPAVtwHqEcWkG/Wf4FPrKYMaUguiu3koUHDXNZUUpgJQZ/4Z6
bsYtF40c4RqlNdw/bXq556tNWb3y3v6fcNJPuKF2ggvYGld/p8JWtbXirZL/ZE73II9lSF38B0qI
jNimy8Uw5p1QFPGXbCXNTTE6faGLnV+4UcLb2cmwnSXnstFCS59XVGjWz/3o5j/Oruio8Iy5aLfL
4TdfjdXh4Nlqgbc0vB+m5qzgN6/LKH/BvCNlYfURYP4Z5A00EIKHz6HgYPQpyUJ1jCtC2Fc1r2bS
BgP7wifOu8jKhX66mWwdh4pJlilX3Ldj1HJnQLEJVBA4qnJz723owWoXIv6qa0OadDZgb+XM7UwB
ZDlTpB85tOjyNors3/dhsbvc1a5dzufRUASzyNkuLqUVmgRnqM06f3aRlOqvlRGYl9/SLzAhDhOo
SHsrvXljH/3N2XU3EehIu6VoCx128YGGIm71S4qVwtamiRnuYPVIWZ0BAr7/b6bpFzjDnHAsg+HW
4hU7MhR2MBogguwPpWzXxTQZ5GJBVKStB4uhccC30CH07JfPYUbtWkjloZzIs59QcvA2b+CTgwQW
KBgJmSEbBxw901zYvthx/1xJ6VgoV+IEs++fMZG7QxpY3H0MCmwYjbSOMFOVsF67ZYbofaDypTKq
a6+kmPe6EZ242Y/gd36HipL1VVu6erY4uIiF/zQFmQay01gikZnzLnTG4Jhm7KPDLQGvicCqYxeV
B7T3CRNoqE75rugKmvnQRB1b9N1G22GbYoS/ML9bnt4dY6KdePONHUKR0fd8F3MudA/AJMX1ps5U
EXryX9VDNHoIPv6J7dcx+DHHgIs2+nKs4aZEZ7N76E/E/0JmHVfp+xV84+RoOnadple1CBt3QvlA
04PsI72W5nzHyK1e9ZkySPg2ndebbLa7o7dgu25fpbaEls+XOs0q1+gldS0gkcAQQN0IzSeVpAK5
N6N7D8tYM1JPZdGkWs7+buOOD3atIJlotWRaVEEvLUtt1OtmmuADqgOUUWusi6XNANRaB35F0noq
qHx/tc89f8zGV4aog5FeqT6oJULE7/ZRO4htmeeiWQ87EOj//YbJBdZglD3X3zYZfwCQ30CC0Ah4
MhZ+Eg487DXP5Z/rq9CGHhNUV3nrPI3qyjjOI5sjxEk2qYBrSyteYee/rd6XmwghRgZzbn2lwdwB
UuMrEbL1ZbVsfz8VQ9ILB6gopIowQFUPuE2JX+wH/fe66Rg3Efy4IYICoPNLK/0cOwS0+Q/0Vp7+
dRZ+MsRNZT3gAAMGLCJCUxa4FzTIePFX/z6rdoBvNv+WToM/nLPm8yMovsOmHQjRqUiUfM6Hz2+o
YaQ7cvyLxHSvPm+ih/9BRmug3upm+AimAJghKuRh3+eLWhxP9KH5pwp7rvKgYRZxQDU6F1cptNAV
CRvnpP58A/olqaMVSxBVNywK0JXZLdW4/Qr2TnQkFD9dZQeobsS1JuCIIL8o9huOEWtniBR7LfL6
1zkeYpDAc/k/5EMXB1DBd1Hi+YGvlGktR4rgl9Z1+lkiv0Zon4U+Tp5aMHv1Z8n19QkOzN0ceMjc
6yRrXCxkQFbNy8ah63ZvcqoX9cLMBpcYOYbNb63rOgPpxW/f1oZEb90XDuVu9Iu+kU2n/5uGxg9E
tUFDt+MQi6XMAdvFuxps3c/F889scmJVCtxn02TlWpj8PG/ufh70ni4Xu6VFSFCZs6aiZwXavO+i
UqPvzLAzr1XEOOFARoDMaXT6TJD6353vPnowN/WvMWoVvB8RqfHGLOuDfk3zu8UthsvqA+mrpWEx
86hqFbhgcZ6H4q32r8MhPc0w4tDhH0I48BBK185sRLQxVZEsb7tpQqX188gafEFz6wdEGJ/ZFhfy
E1JWT6jyuH/Hzu+enRQBmAP3WLp79sgozgn/YSev3CKtvKLKR2t8UZriT2p6NizgKvx5DnCK3eBM
FkEiXuPFdAPaFfoNCELQVgQjLty2UDLOZymbNqvVGkZW4HahGGbOeXALgT/qrGZNHu9/yGUj/s/Z
8H1BUUJxXrKL40AibXOuEWW8eCSdPkwYGrEjN7vHOegGURP94oeA7QDJKYAz6ACKLFvCIYLBX6nW
N+FRpWNdfTxfNpOvkj7zHqxQxCfgxQAiBI5BRHUdhVcXC8bGtRU0iAdQ7AkQD3HmdJ/B+xH6lyBU
KhWt12SWC3xU2jWNC5P/pld9tw2NtEg4zk0EMWkn/6o2gKBHiA6y1TSBfyumNsWgGBvEs2264Z+b
nFn0UVP6wh5SMcty27onPRmAn9oADqd3SRDK2KXaxzNRZbMzcspKYyPEOPUyjVDKvNeLfQkBvKlT
y24WPsIEmM9TjPqM6UHfTOlMnjWrVHCWwyjqNeTiBP8ETVNirZfkDQ6i1eYxzQw22Ni/u7NidxON
W3QxQ95t7eCTo+/xMqJVGCTjo5wTO8uy90ljxF2b1QiiWUpKtBe+ihsWICLSHWptykCCUaZdQf8q
1HRIQapEzYHrS9joa3Wycq0ZKb8P5botI2hoYDQ2XXLN2Sqf81FMqYIHBuOMqqB+Eb/EZSTIczPl
6JGZmRlCM02zncBHcDEBo8j/yEN266cI7TiIWS257kuLRPNpCReuGs4j4Yaqm2J65yvfdDN48PsW
V6Vd7L2ecXw5b8Ltd7r3by+SlI9PjLGKpUrwDsYMbjORWAgOT6DB8eh1axGquuoCtmYpFy2i5liJ
kyVyRtdRgJT58/Lu3aT904AuPH6ADYV1UspULpVVa0HjVOiX4TZcsNPmBfU27GzgKfqlR4E583Qk
YTki5m2GzmHyxtjfXzRjLivXBL1LCZCZQA73bzRBxtLOqb2aVR3oEagTgRPO92mkZGmRiiZfifbp
tUtuZvPlf9PGcPGLqZr25lMVPxmS+Hb7vfoVHcjMsKaeVEwHx2W7Lbw0tUkM2lCoZO9ens0aQ9YD
fhN+jCHBuXWI00MvMa6gLsDdVEaNwnZhFcRHKfz3MUI3KmdZQr/hxuhQkhuMqzqa6bNE7QiO5lN/
NO1+tihnGjh1699uiklZyf1kzYxT8aqpzEleptE4VkRt/CehmPsyd204agYjCEHo6G5bNhYQvtY2
0eITxhExNmKn1wxs/5TENGSFCuyObS9EDiTxp8L2psmqkSzv3M8cAwh+4t+y7i9OEdM7Ndr6MbtZ
90cXn9KYSvNBJJ1fi6A8tJhpuvgpYKSI95k3UJ8167sUaESeZ3BQZf5cMYozATDXqzsJNbVwH9Fd
5IRsMIuRBP0E0R9loQwhkhW27Rkkn8dp2xncaWGXjS2fZxI6MoyeJfUbWBizVXcdhC9DO9M6Rz1r
0zFApfg+exgmh4Zu/fXX/lfLKo7xfUKtdt1odhKNVDy7inX2ihkPl0aqBis8vC7fl42BM4JwzNWR
5we5TOEzIWnjNBGdvVUap9jd6J8mji5v2umBxEUK95T8Zy06CbGxEgYfFGekpmMo5kEqwL++lmRr
c/VUkdOjjHTN6f2OxxtPeTfMNnXQjw/hxmRKvwgrgUm+ZwKPgkctif3XyqtyQyxaU/q+6TcmGjXy
pvHd0sdu5z73nE5ckXvehsJOGTnsaxHFSBjWxY0aPWLkhSihbARaNuhVwUnc0J3wuWTnZMxOkiRV
8P6hGfsIMGVObd7nqC4dO8tbo62W6pNR/zBr/Oq1wawK4Oc6P8enP8x7zS7LVapjxdCAzVqq1EZO
TIy39KqmGCocLlk0SABR1KSdwAGsUbzLl5+P5pF5E62NbttcNbutJOZGnZkfa302SC4bFdvznnW+
MGn3quq+UscEAyC76fk93jVpiyOko03pOu2Af2H9hjjwN37O5j7vh/FoIe8MtyNjEGSr7m/1WQr0
cNMi9K8gQte4omDyqSu4TVi8zsQ4o+CKvD6O64W+Q+PyqZFcZOylghlUi15ttDxwty+6yftnjdXl
hjEVsGRrYxcYjcfWO1iDVqNzfHzxPCpOVDBf4mJjJrFMKn4Motd7mUSToxCK4Shud5bS3nWgm/ql
ZQGNP9tmI58NZmZctnSmDFz+cL6LhFmQrXh2FJAZa2ZPjB3oCyC0I56iwKMxCgoThdrfKAI9devP
6BQhWJQSQ4YAN93ZE14Rg6/M0ITMXQYrFnCO2augIMzB+2CkB3JMRZtKE0wwMxYZFVu0TYOntskU
IA97gjNfhUT5u+mehlgpck1/lT9pLad8AOPRkEqTalh9TjGPBAvfL5kJ3uQ327YDlYUOvZVKOCjP
AawA0L9+IPsMuwfgdbCV0+s4pH6v+q1PaKjsYL1u0J7JmUS4nhDnL89xzeHUEjstYlb8sgrj63WV
nlW7Ei8mN+0mu3ee3viI3Xb2t7bVHmgHy1wa+r60J9NkwAElr/ErjwnMFz/UOE1LMZWixJH618jH
0AfbiTPe3wmBFe4JBFkKma7lEptX3MUF89oUvr1er9pLITlF6Lwm/Vjn3cwCJ/dnykruCdsMK04V
r3NLH/8+Fg2PAF/0W2lt/9F4t1gIh+TjTsig9is8UCadpY9VZVP8xduzrqd3f2mF/h3R7Sb1Oryo
JKSAPXeoQCy1KsY5j4h8fkBAoK4roP1YIA0lfjSDN6zyF/y9uaglLwtBluXDGg/QNQC7qab87SGY
lvQI3KtOIOiRrDpaJNz/yCLMrlihXd/Ft00Qxko5PkLohxcD5a0kRyvFDac9trcTGHPii7o8fiCz
Za1KETVwetgeRhlosqZzzUtq0yzmOX1FERHX9lM0XFR4y1SfT7n/oSN9eeYYxzdPZo+/h10WBJSE
HaeAWHz2Ct8Mhr0uBRETkvUuklnWIPOk2AAC7rwP/YKqnCYRJLImxyBjKkC+VXFsY2glLpWTOJH4
MF0vI13abrZVuKZ5M3Af/L62BGEkAgPEk/Dabf8Z2uNufyRAL6jDZKNgcvp/FRxVpHVQegKFMIHI
yHIdMgnP7kvb4eSyqXcwmGn6UIkiEw7bK2FkI+JQwES8/V5AtArnBO1BSkJQWeblnW9FqkevMZHR
JIylo0EsP+OqVxLw+iUQXFjkceleaZ1Dpys16L7No3sXIDAsviOa+bjHNcPo/ONGB0d9Ft0qPi06
XeU5NAFZCIDCzPZRj7Z5UnBWZGUIbEwHAEbXOSMq7I2usrAaTla7nzjhpTu/4o54x6KxMX8RLpKR
u0cOO3MVmB9NS1PNc1Erc1rKD+f/SKPAJKfLrzmX5Ld2LuJuamhhgAoB5szcxtcymm2dAVwja0/x
Yut4OOf6G3QhHwLTfDiPvYnbI8IeCtyJstoZNUDYsRU6dJ6Ud/cJS8SQ9UHF3HL2w7lg8s2tQ6A1
B1m+16Re7Zcq6aF7kxwgnZ9i45qDuBauXBjl01XBMQ9O9/3aG2GRD7Hq5oKYUiBXzKEMpaqf6FbT
qnAHCFxHVS9zcSaapT/b5rFAU/+sHoBWT8LMiKRG/TXdEcifnBKowFFpxaFZ9y801z8S+bEHuUXT
i3OUcIJv8xced5LahMlvf9r+6CA7jLbQKtX4Yu0NEh+lKG8D64NqgxBLiPmOPhSDrcyC68YdFBIf
3CBXhIA8imXdG96k0Ysc7htZObgVonTffgCKwyTZgVLc0OPI/gGqf2iV5iCfqDVVf14GWjOarugn
84obiZuEf8H55P2GNZ6m0IrXsgoWGAAO7iFuQoCbF5Eg/NpSQGKd4X3oW9QzjdNgu4+w1KUOHhXS
O7kZfmFOweCEhHDe+7cnhJvCWdbmDtUZozG5SmpLAksYSgLyHUz+so3laP/LK7pp+KKOIPsIXBiq
Z0YHJLIc+kWip/y9rh9Yn/0TQLufxdxLsxbK7NO39iaxUbNCx0lQS4R0TMQCr4/hD9p45pHGhtLn
OR3HeST9iNNpp8QiKfstzMYwNUSG/ssZIOUM98bMonSb7MvDIeAN0Gg4CSbIz5KuTxfpWxtJFHbP
jox0qWRy83OruR4G0/JHiGEXk7P8edpoI1Xfxj5tiAPENCBxXG2fo1W/KGUvsL1TmTZ+njiSy68+
97QQmW6GVynN7r9OtZeKqsMgb3drkVFDX6oKoUP1z5lluC1/Seh3Cjjo4i0LdgQ8hiyR4rLGO3qd
GdCD9I1ytGEqlD5MEzQPruDU4NaNonQ3Ia0Gj/Nf6s2bzVeDrhnIbEOU4LgFv5AfB9xmRrpfqiWk
AVWVrQDOtYmy4/Iv0TG4bRxp4G05e0Vph6OSW2j9Jw27lh9ePt1soNILX8SWYyvD5iviKX3giRu+
SghXVOEXoICTb8Su7YlcaacFQuHBEFQiC/DloCvrl9Aesl+7xAVyG4DoeQVIgnxs6C3gJIWzV9RF
1/G47ViKcD/bTwuCQNf0aSUrg0LS7z+sq3JWQwqOMmWY3tn4hGOoHNo71a9siU/JyHB0PA0200He
jiq+kyXr/vvZsAuojfgOSlkJ+kgwMm/Tq06SoOK2tuetf5NEv0bqTFhdxrQJcF0v1n3rRWKJJKJW
/EgrewL9hthIgfXyz0hR3Wq3MeCaFa+YEnLbfaaksIS/QFcJCAGT2/T5tiIDy/f1QQjb6fRyPkX3
lC0Yyw5g/LySayfsr6Rh9qlsOocVJ4b8xsH3tTSlcGti8EMldh6kdnprrcoKCzW2uKGiGgx9ebev
4XYzv9/w7/BAsn52RuNSqx60Mjxk4+D0MUSF3gvAx5MjDHfhDYk56siiAwVn7/OBxdCJxS+1wsl/
VUAxlbTWB0MF7BOVC0USc4NBvqLKoSWw2T7+8Ql4IZspDM/Fm0f45LxG4yFbombbGY1QursCU3k4
UM+qgKjGLzqDVnkoLLscONqmVbn3dNJ72kJRDXCeAaBgdmUu38riymxnLw0oORCH/gi85R41TRZK
lN4CnzI3FhmQb7RYyz7f6KfoB8ni3VaKFOmuhGV5yKMqljOH3VGl9o5rSB3WCtQyjF4u3iTGjy0X
qFQILBJcZhYT/pGA9ZC/NiTU9hgtJlRth11X2lr2zHI/O3XN0xBNDvoku9WiYIrrASZ8jNLfVjDX
vK8MK2xxaQuIPjE886h2yP343kWfyCxOpGCfsmvk74yMD0jrkeU5ORi+/5ST1UreLOIkewukciSB
9VyKtmZ5uj81UemR2j20D4qL/e0FZZP4L5xl44jJQBZqQ2lNrCybu9YyEhO7AFKGdb31QhTGjFfm
eocOPZ5bmMXMJfGWw6yPbhEWaT0SzYSwxqDadOwUkY3xKvi6IkDmK5Uvi1zGxbCrYVltUY01dQc3
4o8k6w6SeI2tapNwnpVMzmI4vqcdlrk8HxyQeNJlW5rP5BRjvB/wUcpe2ekT6vPRtKIIxE0Ch6dP
u1d9iKftKiDRJ6gMQBm+k4TayPMTzHVQuBGL7yYx7a1duPylqrD5DTdQGeTCwGR/5LaJCFI6rfPt
2dsNhwADw9r4FglBHapbPCACJS2+LtfyV8KI3EB63aO5kJ/J9tlJvG7AuAM9UABxVtAYGotI4/kM
R1rGfNCUCxgLUb/OrzUGb2wxKpJRxE10PDGhx7bbRcu2EyDEp8fLHamnXL5H8WJJkpGo4osRLB4R
55SQKkLS7JKwYGDYCd+MRhuAmIk2bHNMBQ3vIOM37DOlg3uhJiLufIoTnBctXo0r0UBw25i3Gsm9
LGWO2GqMijOypD54GcUkrmFdzGgJ3XZr6po6mwSkSFRaOonATzle3mQ+pWYg1jRDeLTXmnYQ8BU+
RGfJ2I8zjat/9EnGVUfDsklEJfp/suUcKNqhBm7NhZDWLU0aZatnc/1ScmtWNzSeFi//hl2XYXJW
6x+FJE8TtEKuSQ56UX1MOegf95j0udz2Rgg7ZR9H1NLtN1UfLUb4EFRAlrcKUjkeOLDq694mXV2l
DtdwEOk1jLGpMXM5ya+4oP577VonfPmGQkKcRll9ZEwhGdRj5l6dzS975OzlsAKE9ed/Dhdpc7F1
Eq7t9+TQOMVkeA4DJiCELKnBwH/rb3LxtVuro8xGj8BzleYFz/yNE9Thpwcmm4UptV/0bhZU87x/
7jzVsDr/fgL3l2+LxBmCX1QkoD65trBwphwPX3+ElnikOnM675pGzZGzZwRvqJRw4qqUxU9s8nox
CzG79Wo4lWLoW11z57bwfocZD1dg82t+tcvaBAUegZ2hJp5oJz0S/Un6/dApMBa6UmDcXuM/6061
LeXkXCRilEITLTqo7JOXmBPmjzGNBQiPffq6L54KMnB9W8WY/kp0FWCeoOz4V0mfdNTg7gfX0lhI
8qeEHaHIkZzcNFp6r0ZQDSDWoOtZoTRXHYq25uo/7acLQDLp3S4zRsKEQfYyLMgAsSNV9BvqFiDk
9CH6YY9WSbbE3JqAjBneTZvw7kW2Y6Q4RJAsYiV2pUqJqPglHDuwkgt7dRt7oxMrgL9LxEPd+Gkt
453ZCa3Z5cABG2oxtLFL/Gst16GYUDix0W27ro4oERwGBWGnoSzmLOoBg56qlHW0c9dtp/7/z1gt
adomkDd/NGdKkKLNiItZUB/wRZLrDAfiTaeSlJ2IxURfFy77k+7lCH/jCdTUJ2YO9Uqxx3gIstuQ
2ESfTl+fyuLBIYSrMyezCLw0bu50tJiqEqiauLVPgYqq9Iof1UgRPYVUSoiIy1eek9lMYx2AzegU
U9IYrKBMHuDxlmXXHkGDLV/TdejNFLE2VR1gJ9A9dIoZ/WnAKqYeqdcTSsUjbJXeJMXtU2wtMt0j
QeU6VKcdFNDHS3vweJ8wL/2avGRUgVM8R/AcLB8j2qY7sbVFVnI1tudbsyfzv4vvFJIMLUHirlq7
EVme5Byl3p3UG6PrCmpsuRJspnzf9uxOV2twWA4RHLhM5dwHNW9PRcCNLFaIgS463gRQW88yYAKO
A4CbDVdCt6A5QLU3MJvQRyDqk/uny19N/ENQhn95krVgae/o+B0FxBZ9oK2BDQo/zb1NFMp8qfQ/
U7fGm2H6kIePHShTBRbw1BbeH86sE/lcNcPvt8Uc+vazuYTdI73wBlF/JfNu8ycA7lpqHOX05vv5
r4wqPz11ItGzuhM1+ZF0CK/rj78VjPQp4ccjasLllMTt23KtBY6j/32eSjE5sj+oNN9EAzi71vtu
4Tc2cZtnjjRSKTrPEjLrnoE8V7bglzQfLCDBeTvxLec5T5peCSGQYm9xazOvE5N+LCzUBLUkNGhD
+Fv3K27LzXhiqbaqs7grOSaEtm17uE6u5kxsNruEluLVAlgdOYJmESK2V9O4qmZqpaHWI7qP2JTi
Jc7Ai66CDOFKOOQVisCboo4SGc88oCpDnfRukKYkn01Vq+6Wo/yftAUP2ZuHCnS8aJ5LCgtZrpBj
5VdbgqR2AMamXqGFEJayiB2xEjCA0en6wS1TPfuqEGZAVmLyyBOe7GtbB0pGxxfXcPnxL6hyg4vy
x5Sg+zsh/b8ks/C9Gpcnppk6iU1tdG7hYsNEC3HJizcb6nP5+prqfczt52fsuUyZFdWqoCiZ06b/
Bpuei+JlxyU/0Yu8k5E44PcGKEG9WYmOdJ8Mmr5+7TxzOP6LxRlIs4/qOUKacwc5ji+4vs6Rh3dd
RC12ydEC8YZAXshJnkbTQci+y9fykJemJu+B+dakowEZgnMxPsNKtf63rHN5Ccokwj3fpyBE5w6o
VNGlRakmWqYmhPVw7+9VkqJqEeVMDXBxzk43FAw3rK4wVyntSUyuKZHSpBnGncquEU4g1RReUpCn
XrVS/GGTa9ucduZpMQDU75LK3dH+dSRvW/YhSLRiyu7YeDTOJ+CGAFz5X2yhLGcuh/OAOjFnw/th
8lggIA+8SwXc/PDuG2QQNKwQ530CnoN3IB/UoqgEdoQOYlyhUtNpRm346rA2Ry2pvLpayv+OLLSF
3mBqTBHPi5gWLH6YkCUVeP8rcd6zwTrRSK3xyf/ya8sO4QTk+Y0Fqq6cXhiAjTrL6WZIKUs2fLuj
VxvNO4i6tODf7IxtZs9/JzzgtwH8TJ9aTnmq3RrtaLnZjdlU0vIz5F1RKhVjwcxWe7k18icPdIWt
oqYTUHWskycsg3USQFeOLONgEWJxS0th6gChzLJn7XbzLY++eyX7agoiHPY7dyrnpGUZLzh6awTh
9iLfW2vyx7+5eg4SdcbhhhKaw8ffdNhKOUBsc/RFvsALUuL2CXHAi1LxpYJg3nTarjrtmE56xD3U
yemjGU8CrmM5STsBLFc1la1CvNZ+pXTMsTN7ggYXGMlavph4sohHHJBZJ/YporMQGpXkZ1ddiMGe
xuEjpXAQTeIIhl0RdonQp5kPMi3iGsYSoa78iRJONP9Qi9sjUnd/1Ow0Ru3xU/mfny3V0pEtlZNa
00O9vj9it3EVyKk9Iom/OPwCUS307fzvl+WHSYv8Fvvj9nXSl83VNHDTWyQL849TPeohIGOgj/FY
ReySZaHqKaqALzulDsK8KPDmApZGTKByHG+rNMyWPeb441PfUG6KPut10pavppQK4SUf7QGOiIuc
7PeysKdl+n5f96GqzBJfIvGzfmGzbfcDVV+IsSe+xh215W5duKnXR/jbjymh+nHJOjXWVL204C2K
x2QurY5T4Fgarm6i8PlPgaQZNzxonLQ2ZjFjutuGo3KOslwh3fhGPYrgpxJEz5B8miB/MMi8gFSV
3CGQDhLo/O0uufBeZefjASXppXlPCIeHp1ar35qyrU9yf41qbnU77ScgH8kEvQrGYNEcT449oX/d
EsiOx3b4sRQAt/lWpjppOPWFbzfmZa0y2WAKSmCT8BVcTLbD7e6mep/TV4Eaja0tF1t+2msEoy7e
XRT90+VLHHPNZaDanDP/bo3CcHmVBqQW065v1hwVVU9F8VkqvQ3o4fPVTwAnzIdnbSP8CIldzLnF
WmiVocpGizdDfmp+2YpDix9/WVN8XRTVQB1EDgqo5P8NLRHqJdFSgXgXtyRwRJJkc2stsLySGR0E
vdpZUy4QtpVAAxK+o08nuO49yuKuhezOAtj/trbK8dJw5pfAAJMjWqXXqk+ZwIN+NKpb1+QoIJ93
DnbwEQWSi7RYfRbeUUrOqXyAEGP59l+GiV6eKv+LDgXkr5Ua8XFKGt0DO0zPQQDsnaPeNt5jsCw8
r7zqgxxyjCaBUlUcyBIeIM2ALV5IgcAUns3eayxKMm/1e27TBmN1nXnZGXBaQU3KwkiGB3JTgLIb
Sc5bFiIbd3h8ALC/aPIeJ6gHDqCY6fUtTQVBlDRpi55izvhLa1mZI8ggBV6HmgnxZCvlCfhVQD8j
VHD8PxmlVwchDokRq85cVcMsA9in17qP8KFw2P5ckqolNEiJv8X2yXcLqfb5Jc/BkotuYyqs9P49
eUXkfk/qzwE49LSzSbw6CXyaE1/ZmnIFzeK5LJcJsD6oDKVGb2ijkO3oAyKMp9N5EOQs6Qpwetn+
mm8Bdl/utiy+Psi2ixSUrTCm+VsdwYHStMCGGkKFVm0bbzSEj6x0WjEvuQKZG7YzCrSrad7xlmUq
w21We/8ONiGbP9lAFxwyvgwH3XbWjMW07uCWwFTS6eLyybMV5ixj9stmUFesGKQwrGaW0rvpw+2M
BE18nI9jpEziYBasACUTeXqAYJWji3GonDxZ6dsyRBiZ0X5NW9Cby6Vok80kRI0V9MBD7NDW6eR9
lzVTqJdPpHT+vCP06pmOOvlmBO12zDKVYgFj15de6+1lEZRYgHV9x+t2bTww45wkh2P9wD73MBi4
LfkJcrstWO+YokEEF4Lmylodkq2pR1Iy3vzAFmIkn/CoagQh+9RFk3SF33hn3JYl8AZ7cxp70G7i
zYPLCrTorAQRpyi9WUMFTsqx9TzMsdJFX9Vek6e5K0b3MTfmDRHet6fcQYnxgdl5NCNY/A2JNKS9
17TvUasUWOWFIp+kwkkJveM8L/ND9ybucer00xRYS+UVd1hu2TP9mfVyYNadkfZap81A5GJ9jqwd
c4flgWYVffTmiWIs+7caDMX0eaTJg3MKZfbN3keKwF42rhup/wJHNfir+BRHAAPjMyc2O7wkWeg8
zhTIrU+vH9sd601gKtMgWWt4O85pryHLnvmLad55sRi085VNlP+c4bP/4Ndn1/APnztVCP4WSY4/
QWziXhhBIMyk6HBWuhMUPtkXAjGKu/ykix0RJTLuMXWSEJkn87eM3+05lBxGFewpnLHNIwxFnl9S
hOTNxAJKKTjqTddWak4MB6FuVCG9jTzNB5PnwWlbQor1tyqhR2xY2aBv5dkVF1/mKlexSHRfZ714
mxiXwg+3Bc2jzsMG7U9rOgRF9V4zdH8JLWfVlFZw7QMteIf/B+9MZBVzRHizq0sLSnrgO/Ipw5PZ
gShZ7xIaZmFMpMWr2pj+cV3rUKyzLyrSiRmeJmknojukoGzCAZoYbQLomsNIo+kCCrLkL9/wr8e9
VDf6UUrrCSBAW7Gecmc/zqrDTJstmHDedAxy3p/5ba3XaljWd43H7qtnNXvJryy2JqXtyqDy8kT6
nNx2V6vw596mHpWWEnBavF/fMJpZoqatmw71MRDfBpVGXv5IzrlPd3NKJLe3uhPR6GL55gC6P/1Y
xNNUqZp1fo7NsbgkeETu2pmGD2fzSAtIDfGnVgF/pE/8vBjXe5xtNoBTBDOHSEnM4YnlOQhVgjVa
ERrBIItF0G7TKIvKMqsG+ywZ86JXRLixi2fAySrtgcKNpeS4Vm6FGpYc90tm5vc1cqMrMKaT1ijZ
xdQI6Ny0tlFy2SZpfVH125aoPRm6I3Pjg+Sv34VWo58NFuvkxUphYC8BcuOdGJrIihhboVk/xFrC
8MI/N51bsNCfvMHVZ16u3g5C5lWihu61j50sN4MHwUco7sSOO48w0SeIC4JSBzdZf+COuzuOeKh+
bkxuAIeF4/f+eSBij/7qJGr2IlifPxBzpVi3eHlt+GnXVtpjeYoOQR5Rub1iwMLbgyxitU6MOuJF
Lba8kDSB4Lskbl8Lg9QDjDy4hTk81jIeAUHt5Aa6pd1D2Tq2LSEeAFy/yuzxntZtjRMCc+CuvvTt
aoZb4+xPdzudCJC5mnARDT4wnFCsCw9EiRn7NPo9AniXEGjon6L6GPtAsZyqMTlHSnQxFo3dSJZ7
2WL9GzHvV8Yv5EjZJZDTyPWeHU6BBQj7RqNkFS5Tp7Y1TQWjBYhGHf/ol/KL8/ihssv+M6YNXe9i
/oibkBPy/FFaMzs0ww6XXgombFVDH9wwhmFe/ggqQl40wOU7l+WwkGQEArRFFPnEddUC0L35tj1K
qfIlZsExPTeFT7zamrInhrS+aInJ5s1fPjLyZInTxbLWctZzRL9CGECjzpRMJ9SxuRmljHPlYqt4
9a7AhCjDCev/suYFtCju1vGTdFiO4ALXQ1JqUGE+wJeQsB6Oiu8lXKrccI7cZv+R7Oaru19T8Jj1
tjsd8DZWvwU1VHJVTMieLWWu9g2M+RrZm11V/xHqQazk+cRU1lcLolT62nAgtbnqIUfub4jY3kn5
n1T5wrqiuWRPS6s0ugPZizd46OIcHfnK+MvaHAe4lQdIHcGNTd/FGE7Jffc6XNgTOoJdpocZcFCF
B7QQd2LICmLQ9b9lBhfp1dMP9apy/gKpLx8ni50IMY7ftTctOoycCXzwIGEHlMQ6Ngw7b2TMAg2P
87AShO/lHmbUXDqQJLxL1ihtboXxGiEDT3BWdJsKmxicSO0k2fMehl4OkpsGqDKJNzdLu7d49+oR
o+mxsGJAZ4rSZL9JOTDXXOXdZk1iXn1kYi6h7xPR8AzJ3OYGKZyjoYERcNu0jZWeOAnyk61EYqup
myfj+iQr9w4qUZYFbX3K9rMRRKL+hAvqR14ewTN1uyLYs3WiZx6sIfXproPLualXTihwgOWBTnTK
NEASgeiaVnshgfcFKw1WwQx83EP6oujKf1GIVikm6tC4PT9Dmx3YHZ0sA3faiUI2mYFZdm0SNhkX
B23eQ+QyKkvfQj8/ClpFqvm4mdDEivsRW/IiWotd53Mo4LGqupwgrVENJX96DlKSAeAJQzX4lMdJ
ls6XGWML4z9KZS/vyI9vQJfgQLjL74SP3qxlcaF2nTbLEuis7mdtH6dBy4FXXUdS9e0aAcYNm6qB
2+Q0EFDOO5bj+DDbhpkUW0C1XuhyqKmZuUN+U+4WJh7ZnCy3g8kzN3nGGMjKozPZ8ookq+LJktQf
vxzMcC9cZyFZKr+aEl672+wtDy8MRNJYc1LbPRhpCv2ztqUaFkqnfWplcdkEauuf9JHcsG9+tWy1
CgEHPLGiV2sO3aU+oyABFVjfTATtcOiZwp9w/DoKDJbiHlG3R6PWIAeHfLdSiEw2CbDam3ZH0LA0
SV82vata2gsKQ/rYScfkiDLdvOYROC2QB3DX/TG6czxAfmu5dAjgODK5MNESAHD9Wjgg4i8ktZa/
cSLjdNkm6sJLt+Bka4gxHzbqNZFOto6aDqmu8ri9QXyuLSSllmLQXw31sNCrzXlMEi4im7Zawj1M
TKMB4P+itgMt5DYlYfRhu+1vy8WqYYnwAf4M5cFUKxAMRCGHHhzqhblKJ2Ah/b529++6RUrykycv
8PKWdXx41sJryE6djTOtMtByALTOAucsL2fk724bBqFwrCwqA8NbWdrd5DKzRY4LFdSPaC/LoAdY
L99+9uMD8UUXIVazfhfk6T2vSeDWpBxd7rZvQFihHdwJwDubpjAX7teFdgyCVekCTdbuLjU22lhV
5ICxPQmqZFuC++J5XLzQJUIa80lB2PoL4H3AFc9ECePkG8Kae7hCFCS3+sNpow8fhuKc4eYcgTpf
4b4brFfM1oYuFdOjU7/ifFkcrh9lfCZ7zYZAruYV3QJF3kxikJcdugw/SePoh0jKqoC8OsCquMsl
SYnn/nlXy91OjXuMT60WQqdQ3uYPGCTL2INobQWpxAvubuDuLs36Gw4xcfhK/hQUPY/zIs9oDlyB
CzISKzyGbfOKYrdhpjp/FUgfdjZOioiP+m5IAft6RjBNEcvzUbuV9+N/6nMv5m5SR52KBg6Nqeav
9uW8t3dS5EJJb5/31M+WQT2Ta8HvN67IoqBclV5lvAhaI1K1w8N56GYNB1/JZ/u0CKaJ5FRdJGBh
qJ7TFnKDwy0SjOJXQyJq2tOWpV6R+eZNSy4LUCJt0PVw2P95MGuznjg6Aiqej8sFroPrCiD+SHYr
SY6O6hibsApmjjFNMPLQ7VKeztShW37WB+XgRpC6+70hIhrkumgXC2EOXnmRmfWDXAEEhy34GgxZ
i/eRyHUz/o2G9/ReGivcQJQgLLmVi2NEbrom5wiu7+jsYrVaNvl+izQcybR0ff9s1f0QIm5kxWgG
BCITAbS78zlQ3A8TPXUt7+3AdpbCZ5kML2KJSTbuopSUT+uP4M6uY8i9+zkv2KuomI57RdN6Hu/P
mXg+qq6lmnYpNEdeaxEojsdGC+tn7ZE4/rEVgxdJCBbRdCJWyK5cFJ1fSMPglKHPEHEq+Q5uKtvt
C7xpz3nCSpalwU04EjCV79ltS+bIViRm4E7RH/7RQTHtKtcHeV3nK63NhmL45GFKvz/UssF3TCHy
IU9bWHlIueufFXC3HTj1Ha2PgOrg0q3XnSVhe0Wz28GqZvzsL0O5DP21a7dlY4oqUesHtrNhzlwN
qcXuFBrG6f2cxGj6y5eqAVVcFuqoMvzVK90ASIMOj+j206Vt/b3/F+CTDhL2TVIl26fJcsjKAo+P
d7uvbzu4+UNi2FkY5g/vurASEbWDuZfiPgTITe/MSKMHzwLz6LJcgKQtJFF2oWwQKsPRN3fKAG8n
twIctiJnOWtoJk9HZFwLMFpySjbqa+6AzyJW1Eea5Ul7NA91DJU4nbA9H2lAXTZXQGa9R7xTXP5G
fHT+pNKZoNWCUPa54fSQ/IAtHBGzWLwLSqF4kT4BbBUyn1e78j1qcaJ6lAPdv1P445lWG3pF6INH
F6vaEmzH4zBsZutPOmsg/qjoj8QcVyy0krqEycj8JK4PvN+21IAqgeLZ5ZyyxRU1WFlCdhNspQ57
6Zb9JlFqYdM971Hp8YhZz4u6qILMtI5LgLKzsiUlneNhT/fiEM3khmLSQwDuhPiTLqSYSQ8TlnaD
j22GLzTS8QccHjevB7GeyWNEwxEniSZvd4/uUhaVtN4bdpnm/ymLxeVklwbodnbhVokge0c9eZQX
keJHGip/21fRPndhr40YhxuL3m51xg1S/CktcRU0GQ2fJut6G5rorAKuvAaJb3zXxZBIzbx7QB8A
/RQMubvm0KEOYpWvsEW44oH/9GHa0X7GfMTB8OVwOuo6JgT9y2NsowlE2My/MK8db6y/53M+rqME
17eMwkALWwU0iEJ1bfoF5S/+V4yacIZf860/RiK9TX90fZzBfv7566eM5eIP2Wk5fdRs/j5avuwc
oxBuACm6bxuCWQM9v5qzw8IoPC223mSxW3W1D/8Mayiy1v7Ls/TCZxtZN000XwK+UoHdQfQ0VC1y
nCUFwT+G8SI6dLdmfp9TKMi2iIENzEans9iXroDWnfh1T9Uoft+uWAusSb2eGq35HurO71v24dzm
0anMeAB1rfz6nG9z9xMvf4Uu+S/CWPDeEPGlZFZ9QyfXi1z5BpilXBHTT/4OHn4R9DtA7/m/Wv2D
VWWX6AO2OO7f3WsMPVwu/OW/WswMmMGPLBdhk0aS7pPq/56tRuqxOeFJNHKcbQ4H3K248uMMQIH0
S8FZC4ZOYF5qhnx9OkGKURph4a+znLe8vLazGf5d9Vv1dHgmBBTnoQbSpxHV/6i5B2iXk5wN5s/T
7t0ktKubsq0XcrOHIUZoPWxqK38vTdogqFWEiCLxcxTuofnte7l/owGuiXxuPMZKvebA4KxmJZDj
6OWIAGyxdxLvAD8kTzMGvc40uaqbsA/UFI73IDfC5RYBs+EPqXNSBEBUsmvUQe7tmXsT4kf91b6Y
//Ir7wS6uJFEKL5TtPnkYW1WTe/W4eL+leWCxiUcHkYYgoDlZZKG9YaxT0Vi5HKpeGYBZiSRSvny
t85ozW2XBJYnSI3bLyS+pRm3vcttPgg06jiDmr8ZIJeFfWnQXriezOBPilFnvQhKD+9plvUe1YCO
TjN3spgnZXiGZc5CseshunFJ0ZLV/m9x+23Izfe8VAMyAS1G5qdz3+6jU45O9Z5wT11EcOzsi70F
Ay+YL94RpM4/A5Sv35X8YKyPWH0gl9zxRLCx32P+gCXYNm5mzEytOttmg8B8/N6F7nXaSPCMMBX1
sDo0zZEMXR7HsjWEcCMjnXmscr2kX+nQSeTQ8mWEz98Hpg8GSUMWpz9E3mzRnkpf6hYD1QnSHoS/
3JobpxnK8Xhci1m589/asr5f57bPfs6ZinNJo4Dr49efSMu+kbO+TAYubfKZo9N8Xj+t4mLQ1oLI
0KIjsAhwaHz6fJA097kRFiw12MBDizxEfrD77G1nO4YWB+elUnL8Bc04FN7ZNe+MR4hD9nONdYO3
xkX00jIHTScfI37qkmC8MFBLiCEv1TRGJOpmsdRxbc1kp8Qh4Cuz15ezCYyfRX600D4cGI29Yqxl
GkoxujZ2MpH11ZzKXUz2g2tOGqCsRiKdLS8sh/AVi5j8/qxhtsHDu8UZrUyUsRT66rHh+gZjrYj0
P3ZQT/0M0TAl/1lQFTSgUDQdUIC5fbct8s2eTDj5tvgibsXQPiK4vtRr0S1kQ9yzHdyawfp0Jpak
6cwiV7zjp8AYOnE5xqrFW3GvA14mfrWCyuRNIbg407qNdzDMCBtkt8/tpoSNw6RBTiZ5W2Ccc7yv
f+VXGeJ5onsfJ2XedmQecyABF/Pw2f7KnE3kIIsC+dr0NEBY8rKY5NKvUum/OT/9XbpXYP0F8Yja
ly5D6GjZeYewbglY7+7LGQJ01SXRF3HrxJXoTBe+T8dPIAd8ybJH9oLNZNjIadBLy3H5yeZ9+C+4
xG9wgpOYrMItuTP10s8pLVbsKy0COGI45tzAoRhV4Nq/JQ1fnq9tK/FevD0C3LNySk3v1Eec4v52
4OSwEI1wvCHxZcBP+n7vgmquOAbr6HJuBdfAxTknvUZr4PXyruvXWwolPFXBrffRkXjWfWsXkwKL
lRzORKWe5XRAY8gWG9Y8kUB2cpQ+aly/fseoL2P8fA2XCev+2qqoZoi3sye2QYBObn6u4c5HuY1e
j9wSP6MGuzb3uVfZ5S8L+OlK/eZ3Ec+OndTeLO4cj9EJQaeSLuDN8KeLW25fFgQlFSD03WLKS7Xm
mKBEtGdqJLadoEFgZxlODQkHjCj9tZUEaLuRbcRqUQOBMi/hmmjn7C3e2N6slM6QcP713pd8/C2A
mgb9qgtecN/hr7EbxBSgO1U+19IO/srU+xgUGbE5J8zj0CKHAF0d4Rhu3KXsiEKDwMke+bpPlSy2
c6NZKXaErix4pP5AvY5WprGnFvBPlRgpjbAlTbDthas2uRreUA788m8ZXwByOj+i8nnuJPp5aOKk
XeL4UozvH6RccDJjTn2lS61/ZLpC0H0S/phrOavd3fKd0bSu5ehtv4VY3qZcSdLdGva/VQ/AdOvh
1F90DoWi2z12Zbs/nAtL8iC3H6D0RoPYvG9M+iZckjjK5f/B73Nb5Dz5+i0nH3xlA26uiFcWuUh5
/+Tj3wgldVAWJIT57OSKDw+dANHFFmP5L5g4o2dFssd08FE40WaXotpZLeb+iZRanCeAzQvVSLix
mv+YWkn5s9iW1NjYWLVZalPznCKxC3+Zur+iaIxatLt//gpY6b1/zdDYHknooYPDRhb+LDfV4TnM
6xApqMTKTfqSgqysUfclQ4PRQXSUih5gypsTy3FDW/mNpYlomVwlIFh+IrI5QBO4mpDEWLrBZ/Ye
4ziu5AbMvxa1XVChggzYgg3FjCpTIOxiNuUCVu+IG+SiEqC7J2ppvFMFBBi5VBjL8K3L5nqKiYpR
X+JscA07gD2oFTDb6OkyfiAH1LqCUHv0OpDvIojQECuMJeUKSA7uyRgE6wx7kUdPxInvhFfD+Hlu
8lprn+DPNNP7xm2A/HL71MSAC4TGd9LedUrkSpPgTtUf1lZT7x57rQqU0HQOmCNPx4Ru/9Uhlkmo
G1Icqf3MtKTNYgRJ0e+deR4Y4Vi279SQ6LIqAVPYMwh+EZkWxBzt1+s2MCdf0/RR8L4TYSAVDEBs
Yj+S9g2I0IjJOoQsyMkyqR9FbOvdLm2jpeJL8y1jBEPaXhpink2nTlQr1YhurnYYLPFYs34NUi3D
rVECtZ358GQ1f6+kdEa+uYK1tPqy6p+Yj7iH51lkiFORjXHJd2WFSwxjtM+CEYOFO/o6Oe4VpIuL
fSwVQooQvZHXpsF94TVcORjuSYqazzHrFUS2pQghTevleZWLznUG8vofYdh7YsYLmE3VTLXH8mCv
8pUHBLTgi1z24fgCjvUojq5CAHVPN6r4fXVvd357eNQMPEVzNeOltIZ1mwAKE3usXad3Ew1GnlvM
L1ZV0APvWLcVZ2J/rPU9EaKo0oXVAN11qSIyuLFk8dBNIFLnPV2MiaTpVVWYtqBm5jhW3eadDyec
TGjCVc4xKoYni0J6MNTeayAMVJ3S5uOZZ+Q2E/bnbIWx98vqpT7LegeBId+tNIMP0pAy6x4qQ0X2
A26VYvsIcRLbEsrpLQzEJRAcFHPPZKCKbubetC16YezHxNAnf4HGSn8S2LOn8A1iT9DjqdlNOCU8
bt6iuV9RtiNjBbEgeO/kPDCmcQaWgo77YaOWB0xe0Fe1CS1b5NkeRTTvVhjEltblmf2C6eI14sIO
tOaInjV2FWd6j+MkTktCIPS3tVU9XjU15lSKusJBNKNcOwwVjJipnnUM7PIhSEidOiTTGIpbZ3IP
YsvO5zOpjaLHPVASzMHq9uEA1Jzd/88v/tXW4buSGcwXkIejX34thuz+/9ztSlhhXYH8XbJVaAEt
SiB+niwnZRJ1ale9wIl04thLGhTMtN0AcdQcjPlDPyRB3IKaG9cRAzubRUhI3NA8Kn9Uf6OMAcKI
jk/NKSI/sIdwnUs6y9WETX7QjUEeUM7QA8O6zEuqqS+3DJFDTH/N7ub1B7Bn+HCkNaD25nz40sVu
MzKpu574QqvSee1l2nBC/94AKWc9ekaINLLfS/HMR1szVssi+tuN9jwefNRpFmpFbNCa7edd8l9B
y3fjYf5tTpNMkcmlVVLIHAFO+uXqS9r92BPDZsGSVinvLrz/rFDbcrKRCowlnzQWMN6DUx7H08fn
mRoOOo3RnTYWODhgeWOttKVOttTnwOIykwdO3ly7EkbG6LaewRs9/KGHnfg3eeDEkwOyTGjIpseq
oh565YT5pFq12nXhTC35O2CUk3LwVY8/QaBwhT9Ze4v7PC7EDcRye6oiBsAMcLz4kgxiE+tIhXWo
Phd0tBcJCI8MeT119/NOyJi+kYqEbAqyCopUQuAH14H2UT4D51xw2mFSA8whNR4kLZO7oUp52ozs
FO9QPTkv4IDpoBSQ2m/kkb21YVhExeNrtZ/RcjwnHFAZsBB9pcNtG32VyuAXmC9Ty7bT25hRzDfX
sGqmI93k1HxzLP+avwQZgg//e1Io8hEAGrQK+AfbvQZ6zbgVfQkHG1roi83avashmROMZkFLvOMk
SoJWoHqZ9hB5ucerdb12VCU8gdLQ5sOZ5vZUWLJRaQsqb6GfAii7ksSE82zyTm1fE3Z4AGJdnZke
WQOWUO918NaG9T4RgBrbbWw7I3b4+c4+OYbkXrgWKWDGZxtX7iUSdZpY+Mgo8y5O0P29Vd8EGwws
yuqbJ2QHQXK9TdjGlZ3a4DHnVsv5HbDYCzobSbdjMGL0AGD+L/32hTMXA3PlYX76ScCT9jWbp2Dj
cCQuqCIfv8rf3cjoEJ+RtJuOKdF4mQuhv5JRmZXKpHTSolmLSnZmYjO2Pu4gnaopkGPW2smwlWj6
7qN+1bAQsJGyKymOg7FVCRGR+2opa6qUBxVUrYu7mhxPFUz8Kgp7rRJQLZhVkrBrkPYvvjonaWnt
ZfG9gHHe5waTDQd2cqxaG4azaM7yQb3GTBMm+Aplo5vUrDJRee54stAzo1YRsab2EB0A5gpRVKLl
nWCB1MxCjChxmIIlNp8+Pr8B9OSO7JXV9zCDOAbio5HpH/tUGiq4ecb7imhI+KZ1ZrBHRgc/TA6e
mLPYen7xHGnHH7HwJVd9IAOQ3PDmxX9b+KXjZ5eyqvGSqW0z4MOKdqmlhuP7WE+FpsUxUzeq7Y8W
QBqYcP6P2+OMaVIZ88TFNXWkmGfq2Y+Fkcq/oHvrQZ/+h2VCl6nJvdWCYZi5ZxBlWFxl2YLiFNq/
9jzQAJuUqHjKB6r16MCak4SWcmI1WcclDznFJHo93BpMnCYhsHgSBewEElE7t5vdJt4ysaI9VNJ1
MixSzVRjuI7msjlN+HG1/E1WBqdSBluQAgFZ0YrW66eSh3brqOJnKinRqQUcATU3ylIIm1IVYMce
HaliFo0Jf1jv9a+ZSltkq+SqSjaCD+PxUdM6y7Szp8oeiyJAqvzmZndJ2kuyCdg68vaPoM5GwsRc
Iw5TxkSgzeo/bjTJ7fFzPjRdMfMUOFIbwpnrZhzycv+nQsrupeha1tI59q0FPMfvkNfbY6x48scB
tg3eVkf17012JcitkfFB+U1G/vjM8UN/q5ZxArIyS3rSiJuiSmP1BgLSPC9nB2xj0Gr6hdUTDZZb
qwM44KjpYJ5nWz/tmzUD+D3tDYhG4XyPLFS9UIVIaURF62beiaEWf5mKuf3oV6qg8T9S8pVWN9gO
HY94yP/NLJp3Gezpa3Cm73yZvrieUjvCbkNeOU3cNq9RjNJd3HDwboq1TaXuxICpmnA5EajKILnQ
rqsqqZ5hkMh0wg1RvpOXawOOGOboH0b4d2l2i3CHMHp6hATBd4SPL3eydMHEmphD2u0yLcBJZ9lv
AVzfylrRYVmAvYzXdKd6/I8uCzTtmwO9ydIGr1Mt1AKqhQHeC3sDx74CDbWVvLYdB0Xrm/sWAmIh
0yBdYPqSi/k5Dlm0ivyQwMsFmHCRjNpcSLxFteh0neK5UR2irS7qn8BIj/d+1csnmLjLW+wEoE+5
oXtLkI521864n2WUgwdDBzu9/NtlmwbxyjLVZtS8kYZDsRKTnrCl21iMDqy0j2etMYIsJSARFWls
lUaaurQxrncrGywtn9DPmrKV+s0MN5jkPOCm1b8odddmJm8hPbf2PHLmalryxKiu6UO1Mx+Xox1W
qMK2TpYAh6QyZL1VUXlysP0HYoJsCj28xyrrBKonUvj2NBw75rnN8sZiItTyBSZhj9qrifOL5z57
3/4YyrVIQi9fIdWSQzRX3teSue0BfQquUBE3OP1arKeAEER4l5aR1oTSBv8eVaw3CVLBWoq3lcto
LWiVxAFhMEwL4L2dt751AnaS6FUOMUr5Ht3iRcVNF8WJE+AyGEqmUQTrpH453KFbUXA+ug+HPvG6
CM+BI8GgQTzNE4vJ4t3FxIwfQXNhRAvJbW/5Ed7+1Igmap/upSyNUP/F+KHG53yGrrm9o3/Bkou6
cbALlSF2DZzdnr9uEgexlw2icFdlp6eTjtxdwghwYfEV/7Gxy+V24WNVecAHS4LxVD2WLjXJKVdw
GWn3Oh40dtMDjySR6LFvz8OyewMMlJbNZVAFa1YoEYyvn6SEXV1Z2iTonFdDopBdfW/Dncc9cb/F
jvGZUB14s3ArGupbI7fLtuK8LRwNpqiIMzkE/Eopd3SFOraDm1o8DaEfG8WGBUo2AYnOI8y+t+Or
pIib7pfhps/6pm09pyM8qYXJmGZZzBWLFxze3bQidNtVQiYBqzUVb4zdelq4v38aiCNiOuPfW5pF
T4rjp3PR798VeQ9TUbVM6SUozhCEiz+zMlsbbhYsMqGWDK8xjRA/mLPiWbhNX9g0vBH9U2a0Rtpd
2t+kLhnwVpJFwi87lzyfyd5MeRUFnuVnJIoqU2EyyVcdZSVjLBN9UevCfNaEqeMW9Q1eotgjwj3o
DR0=
`protect end_protected
