`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10400)
`protect data_block
hTX64IeLyHzfa3tJyS5DfnCGfI2VwUPJSF+Bc54ckFzfSJLvCkCAdE7r6nLip7WDnWUzhj3apIeC
Yx/OdOHI/DfHSXoewa1AmgCGKlyr6IPqfObhzKzs/us7+JCZpgDFsT1AgEnso0GTGAtXbjLQixu/
1BnMVgeOZumfjEq2p+RkfSbQfjyYo7u/uY6xDLROD7YfQ9hykk/miaVk19jI5tQMY6FCBcgbN6Pf
Hc5DtCsowgDbJ4wdzjz3y4/0PHztJ1JTfadXSmXSf6daFQQWkuJmJ5dpIOM4hJO2bOEGZKLioZ1x
+bBGhcP2ktvLv3jt5Yq5kSP67Y+O6ttg+mJlet9g4gsyd2EZhFPvhpaxpEhHPXyZSw7a6zYzTLPH
mOYHBj4FowJq3nmfCQ85mo6I47zXnUCcZH7S2rRgQj51qoocjAdLhH0MEpxw0el3eBlnjLcGxhQf
ctCb7tvsrcE92m2N0ZXaIzez1MxkbOP1UfjJIdtX7wmEKedV+vBv2k415QkG48/bn7I1T8tFFIqa
h2rYqJRIpy9aQGuK5fsg4QxIVLmIUKdLVs/SbGxa4Nqk1dfbxX4p0XPBdZD1ufAr2uJgyjiUyXSV
j4nXDkeSlH5Np7PsX3/6hap7jOPZYWNSlroaOqzOnP5vF/AP+5zDrkCwUOFeNE54V52a+FkvIryH
q5MXK6oSEhQZkVa7uw5hnobFGsSoNSbIo/hmQtkBfCuc7DS+efKNYoSKNSb+dIOjgIfoaPpIFJyD
BMXFmi1MdRShyW0BbL1lEM2oWhYog5IMfjMTzf3isYGQ6XfwTqCmPXmcahsDKlKn82JkJSLmYD/N
8O4QMI/66fe4qeIOxotK+e9blKZ2z8/JEtEXaMWIpLlvD8zvG1U4/Av7qejILlB3HVcQAs1vZuKN
hPB3zAl60bNSx7egsntG1Nrthmyx05QJbbXsnGoKXJU3iqTxBlxUxSNX+L5sMf9pySRj3FeXT536
IfYz0tHX73tMacfEor04gxF5LiR6DDGeBwLNfsabFksYXv4GOWUV9LUjnaqEp85ItgYrWmM2A7Ha
aXRo/Ul6P2nB5pzwTCWZC+1qjlLGVgabY2I1uLwajmWizIrIFAFCQTwBWEPaSPT6OFLC1pJ79p4p
30Ikp2exsJ02dT2XBpAqfNqARhVyJaITvlinJAB0yRo1Q9ivvT/0KLfLHYG30hyfnrQ+qUyZ40CH
qT/0yrXwt+XVo9KzpHuvxsLohrl9T6wuO/+IjUJpf3L4CvIr96c1i2IFHbCmt8BS270YaNHRBS5b
oM71LO84VsGjgLguqeCCsY1S5XQZJs5np8PiR8j7hodJIwvCbWxuRfvlkZgiG5jupsZnni1lKGh8
xPr/Bv0+mm1GHymWt+4KaaWQSWa8OLCtdGNetK2JAajMD7KKjtH41NAMMQLq/5EU/ehIYoscodNC
ITGH/Ir/KZwaKzqocU27S+HH/9bEi6vkZ1ni2wC+lxEpNzlkfrF3mnxTvcldDWCHiXEF5V+xGvxj
hUsDPBxhS2C9DbKmjJ3ik/Mdvwzz6od/rqaYt2gytTB9DVrBSqCEGuitp7LrweJBQ62GMBviWGNg
XizV/ctYjfwGLZepBN9TWWHqT+drfqDWp3+nd3OflyCYMgJBX7RYGeuZ5EwGRBOmv+CprFufTc0E
BtpzbdamK6WxrgCBLabZ/t5hDRfENPrHlSz6wG9qvmjyDpa5GfLvIHFGcRTmrmVmh0kCcN7nBQRh
lhOCX2CRmdJQucJ4BCjGdEWDHJHu9XQUuGbaAREbhmseA2ngHAUzVWY5MP5ucY/yZ9S+ZLZvBoUC
u+rkyQ+LjcnKLUyl7rKrNxckFvGa/ca/Wre2YsjAIbOkvwodwdU90YueuKjEz7sfCBMvWPZljwkU
Qjc2JHvTUkDrOy899XcWWrlviK7yhgmsYS6YxJhdi2gECM9P3S3C3b6azAm3NSw7SRO6OxT7wnNe
CDMTbQTKXYS3jBeU3Cbo58gjus/G3NaBLJRsJRHdVjsE7JFkwjcE+TOuSnPHoPFG/WUoTEam5+R6
KKNAwyK7DvIT6qhPgZX7F7z7SH/930eUpXFrDdHErt8TOxuMY8Nik/l1MUqR/6g2XnhORb8jSHvX
v1t5sO7uoz1phBRheuVR9T0aAv0KyFIN2Lvf+F6aDJgSWX0AUB4QqKpSIynZ0aFyJSAwf/+YRZ2J
Z9gfhuKt9mLBeES0Febv5Ty8Nkx9g2nPQlWUdWJTxKVUpMyecz59WNmL6HXuynuiff99ujMUizkb
iTCksqLE+aK3aE6DQgd39ZDRE+7YwgGOWyVOE/M+B7STZYkXIZziXxgIT1KCGjsVpVhCWmOjh7Vc
m0hFRDzE/eGYOBWDuHbq3+Hq5cyIsUtVv7TY8UPO+brOtzMo8lgMSXkpZhlQ/zRUtjNPKjmU6rYr
GajBvQhv0G83/pPVDttX5/QjPjCNbcCg/j5niwyu0oJvYAEbx1am+tWHos1tqvixH3QE3iXNwf28
dFsFGFwJlb6kclwg+zD0Nm8yFNMpLEE+6X4QBhExVxlH2mQOW9RLAx0bz0wAk4jTkfmhnbErC1PO
Y0Rn0eFdIqDXsvHscuopMRiSmUGTAuDzGIxlLQGSaUmrCBSibswX7T09E/TSm/9PfWPG/Bpashw7
iYq1C3q29l+auJbiQW6t9CoBVuqLdiIaxZ7+lXDkM5DAcqVYUt69puyxPB+MlcEyLdT8mz1kgyu2
Jy0bG0t+rl3sHMYphMJCbrbDyybBeEYwTlkf0oN1qQSZ97VpuwfQhsw8WInsCU2CbjOaxIqixiZH
RkK/dKfncHewmvM/dqhxKdRLi3nhpi80W5Ne9t4C99458q+HonkbVtSs4w43sNNAvQsrJw/sea7X
6NbF8Hv8kHrEgVxXqg4Ucyw82mGHuVeM4HuvujzskJFF4KWV2YsnjixRp3WcW4YC7XIRWuoErujD
02yPPgI3NWMAhcCtGBBJSTRxbI9K9w+x5jaS2m9FAqkyYZpY6O/MpMce3iL85ikYbSMX/BVnjofD
n3LnxQSaUe2d/IqQxPnx2jk0VkqNiHX3hB4vVpIXrCbwObqWnUQT0+72ASVaYiDVYcCQq0bN8tWV
AR01eHIw8ZWPhc3Tbq2sO7jGSK7eLn3GyhJshYHeXTl/CVdI02bQOOE4IE9zOGqqgoF4JFurwDhZ
cN2nk/gH92lTMTpcz9+Dh94JVr+SPByIOimPaS8fkFV6jPLlfqd5BMzAJWy0TSnML4yKf6ZJkzTZ
nRwwlCDoM3JQWOocVt0LfoYZ3aiTBe0PhBQq/Yb+inyrF8nBs705EcMbRp0AYK6q+5TjaXo3vx87
l/gIA+J+D9RaLxeR6hP6sjw3KcfFTw3DBEeYxMAkuh4hFQtlddYUQNlqmjBjBxGHcQceeBWPCBZZ
CSTy45AGNZcg39XRAQdSaMFd5pn4MCtvthtFj3pWlBLciudsm7bm+rl1Rg99FKsllTiNxBls34mW
ipPzhtYrkSo0Pp9YAm1/1tY5GS9MpDnL+SxvxnVnVBpUPqbGaEm7N/TiuH4HbTnQGL2fp1y0Qtzc
OOY8gJTkA4OThgjAVBdIM1O8EWVGtwlwkq7121Oihz1vHl1n7/5rbpfcOnBTg7UVGQW8oosUhMam
Ww7bl5hNM6bVtDLjQzqmpEAGKzf+aqMeSf2voNlKg7nMQrVqdvL+YfEKLoDgKzA44+KEIybJyfjF
VOkHQ1iwZtaKcnYeN0S8mE8TGVYAQ3SXYU3yNX7yoHDIGK0wXbFAOnJiMmp+mwhxQ1U52oek5N+b
Tq/yA7DOGhGzjafHb4ifbMUueRm0mS6CBsFmlMSzfnKtBdrtLd1KyUqgjiBEDXGUxKPzhkUTBYds
teg9bc6H0Kip+vT2cfg11AMI5RD7LTz4Z4JDWMC8ZC1ev+HKeU/UCmf0wSFno9MR206dNXkU/XWe
mIfhUY5ReisVvf8UnYOMDfT8khCG3BgIjv9LTCTwIMlhUlfbK6kPjUMYIDgR8a3eCVwboFgFqJSp
QTqKPoxk3bU531srY/Gtj6VwWDIakmI7TbOw+0VxzK/qaavlzD2yZhDK1FBH+PTIQJwXJC7haht/
KUefXTndMxn486lfabTJw76dC7NUpX4Kaug22TxTS9/vfWBcKrftvy7nu1HZA91weK3DByIq5/oU
NxxECwmFrmO6ZZph48hx2JRPCqLjGyVZgO7pQ0+LAeHOreqqMTeOn5/V0d61SWRjRLkB9S5hueC6
fWTEOJugqG/DmWm8rl8LNvmo9/NoQ2du1xw+GIiCuU61z+59a6DkwZulesZaclO2Hzg8+ocjtIPO
CQAQoQXP/kRALlQEFNMlTYxtRZwrESeF+35m/3HJCFIKiaVz5/UnN3Mv5QyYuBl97+XDygMR0HPp
k/r/CNPR46hww2El/cwdPtgd+B3qY/tC1d4mfCH9dvhxXOhFaNDMvbpWOTyORUhZLLtBz2N263XY
I6HDtE4BFbXgPcIILtpHXbKnwoMRaqie511ZwgvOE6O9b2N0XvnZZx3IeHISmQ81G6sGlBfYBWNv
SLCEdwgURrqGYt2aSzg/7JfKUK66aE7RjkmJiEzexDcoPsdLEPaAEpqstWcAsnty4agrkBXmY7Vp
t3WZHtJqRlE7asOx9hB7LLkw6+xA0Pl58bpNd2w57k2cyKK7878mU06zVdlglWx3eTyswtClXWUR
GC8fCagBkWcWwGdTJtaJSFkxZGXjjiOqCvY6rFKmnarz0jHRO36jI8yhE4f/T2sF+PRrUE9oPQ5J
pLwP7P9TGxwdXvLIvLoDMhS0ufb9+M7SzawXy/601ten6lfkYZ8wNkauGSvr9Yg4TE/vmu4tFKVB
i4r3TgZ1WrCJvWWjZSlwfV3/FDtVb84Jcy8AoAqixOz5hpZfYDANxI5stviEq33AXmoJkP49wHIQ
GKeY57QYrJlkDNJTt7tZg39RXHx2PGWniWgJGld4f7n1tCjzL7Recs1+hrq/MImgnoKHvg8oGYTy
TYELb9Z14funjkvSgAl2yc4/VMVv6n/se+7ofx6sSTeBrcxy8ffYjJfZMNQsWtTP02KooCuK/6cS
JW2XMjFDmDn6I95yhe5AZRW6w/TFkRMHLb/6JRaJMLA4UR9dfyLmtXITZFmedfahYHBYi3vjzeO2
AqwuMlDXoWdiqMvwurJGKIrJsrSbI29mQ8P0GbnYMGiBUX5RJqn8ABr09yoU31u4dQzlV2VBaqut
frqiuPr4VGRjBImk36hGcLdEsOTjq3tGGcFoom7N/wyz4ZXKr4txloxOH/uCJOKdAt6mYKaskWl/
Y5KQE4voRohfy1gmzDjam90LKRkyebPSKSugzY0DokLDuXHCQsOBU0RoPfpMfrcJz5NTZj/mW1WY
7qLNQVDauEGYAdUmS/eGkvHBBblSo1399A6tgVhTBfhS3T04xHE/oOIiIwzd6Q/okpP5feFMf3+4
4etrvCQMNvWOu2vJy66T6W/JP5Y/1l6PLBoXOCMuD9lmq2LRivvBPxOsFnQqKZMj/0C1k8TfmNh/
QHK0l/kVyIyutscAlYEJRYSmoBh8I/zQIvj6Ru+mB/a18bENPCt8znwzdbwPuAan4trB3uqSfOLV
5M4m/z4oRLi4hru3G7YXl8MX+qeeyx4eZKB3bzpinW/p6TLy/mwiCtbGMFDitoGIzwL1xsBDLe0B
8agCA++2B25zfWQOF7z9XpQg8RW5FF102TffFEEUrNuNI2LUyxUviWzMLzEMa4tUA2J3rnIdy8FP
y9E84A7N6k+o30sbEznYP7kMviHJf5v1hqIMGPeOUt6bcjA2HARC6sUWZFZ2BYmz7v1JnxFoC6dn
GoBNzxSt9O1QBir7aJVo8zDQc8g3gUo4Cx+d+89WC3khajcnlBHKC2GY2Msl9CtsnG2+FfUhUWmt
xx1KsfSWcOREq3UCXTlDNROm+oEk7icSwsXF3SEjV1oq1CV8LsidXuH/MoAJzWavshvjDyGWKQmS
rv/xQJtdrZlIDX74Q0rqgHY/otucQrr7hTOOnp6XEu+6zqwH/gpUDeaE7Ya9GVNO7IkRAtlnR91g
tPPdiHPzREhYoZ3cw6HnlUREO7N3Aw/ipOrW/MvGSk5m6QuX2H5HGE1c5vdJs4NbNesl+DlHhzPy
SZuKL08IssSq1xXh6w8b/F/HI/hFS3hiUaE7+jSfHggDkOQ1s11t9uumjaogZicOogP/0PNpg1fe
I8TnS4r8l++cSeh3B+rHIbZtT98rownyv9wZ6DV/as/DhXtaZ+4MxiHB9GmOthqS3p60sJCcDzh1
CbbG58PirOGN9JeOGV3+z3LH95pbkDtc3c/h3PF7ClAlhPhdwQyQlMlmQKxfbZENqNj/JpH/r3io
6xlJ3dbhPMHuhjiCSoabhWv3xVEICHbO5Xodjpt3KYEfBIK91jIPJ0jV2j8mubQoWcK5x29dW9xe
6X6ec4LTT8Ks52pmTPdLlFzhejYG4HLfKhkSCjj3yb2c5lLbjdQ+mkM1+cCSvpfM518gKuneiM51
gI762wfIieNS/FtO0mgi8L6YkdQMZYW/TYniPviSSwnNaxJuCQ8NafwYMQCvBkedaHPRyfnYV+/w
p+rT4pfYn+13wbDm2Sg/bUUhHwg5snN2d///UkkzVUcbXXP/vuK+s6MuMhXb9aoS8YGhMmzGqDpB
I8ZbggkHPhH325dky9SPOXIrZI+6lL56e7P89umeBR/Eru5hGBeGZ9zkanGanV/HpwgB23KQ9oNk
/0YBSUjeRpya3w3ancgbN5bO6lvWhN/GVaQQ2eRmWplwfTO94FB0KQC2Q+dM3I8EijlMw+JPx1zg
aMDiqNDD1EYDvavrHC4wtZfoebDcqOTgG7qJvP7tSk5A058thrWu3VUvQNvGFyNJBpM51OrEzkws
V3kKAY3O0SQyXh+D/T6MyhWF0klSUDvHP2kQ3BTjQO4i8oYjipljqugrRlm3ZPQWnoZnosBorZgu
7KX/WcOGGfq/YDbagwhqJH9Zy/TmzIvPVqEs+ohw6ziF71nazLyG/tBuS7e54TAOEH3OOzRs06q7
CgdSNziNApfp+rM6j/DHjdzcZRz09Cket6ST7Imb4pJUP7Ck6OL++AoSjZEyi+dvrrUyaE++tfYS
A6f7Llr0/Zj4h4G1Y8U1Kqs70Xkl9r5mHsZ15LT7u/xjgOIaorXFr0bYjOh1u8CQqTdHDbMsgZ7Q
FR+Ups/j12Zdw4JbCJX5HAdf+pmikYTLnLP9EG1byabhtrOeGFotHiDvmb5oCte+KFB0xHlWAVli
TgCpjcS6XJT4kIiFF3FxqudDcXBg7WWe4udCb8uQZO+sxzZQAWZYURVHAkq7DwH8zsT+dNf69oow
Z96LPgMShfbqgvT+tIOSDXZ1c5q38aHi7Z4nIo7quspm2Mf6XeuM2S/eCa/R8o1K3tTYvKZ3Rqmg
YuUSbzAeYVGL7zCAMeGSCz/CVRh0tbnxpPm1mtM9MgTb/lJB5jWSW46VoFv8I3Ybduv7u8IJrIuo
5aNSssfDa7UmEaIuvDLLHMckXiSYrjmtgoKjAFX5SqlXJ6PeKM8K8DcnRZQsMr5KNqVWI7HwpNK5
iOLktoReZeCKGe7KQ4W4BvenP7GAgrjERU9mj4Kur7RM/lXq7XmJpnHsaigowdeCrnb9FEGwVQbg
IN+kvk27mYI2RxZhfLzFXFzVv8diir19pNDGIn5HCnz4h22gPGZDD/seSATMXRm2anWR8Z41vl+7
fHnaT8Xm4AB5UWTifKrx/8+OfQZvwvahxSzJpcY+Grabc1K09rIEhW11IWmMKDZOtx271ZapCtMu
QFPXccVj0xUlEwNah3nuNW5iyw7T650po0IhNtb17tEfctLirAc5hg5gr0CfXQY84p8kHmqsxPrx
K4fPqeukk9D/57Vr31CnoQGNEeFtDbcZD5tPBFN3AMiZJcicn1xd/S4okxCf5QRtf7Ob046vy24o
h7TMCDzc2B1lJQo6aUFTOm/mMwfgTDRu3pYI19Uh/+9avCzxPd3a5+gZZ189jWvYH+gzBKLkrMz0
CVpPekfRMOxv1ro9XHndPse65wgdr5olHy82VrqD2k249Jn+LTla6PhLAyXRJv1BHXRMJ5cNKEuG
WLqh+1V25+5kazV5Zg8s+Uos3F3wbnB5eJQdDv51p7yJBKrH14La30G1Aj5pB4F9w5FkK08fj0R6
vySqIQOTgVEwqD90PHlMK3qlAzrWBEb9wz2rywrFCjgV1vHwlho10UWlkYKq+pKaYdRnh2LqACap
xBJx2FwuivEQYB8Oe4L0pTJxuUrXMTnkgfbZJRNaxqqxmLPFm6H1lz+koteItodoE7UQHv0Akxt2
oviYYIWFhN9p5LMVlT+qrN/AxktggwHpu3O73ZwSVpvbu1DJ8qShPWc1qgLb77ChinNzUJ9Lfdvt
g62mIVunbWHGiEDV00DRLBE5HU/TZlNRYrK+SIdSYdCAGvzPl8fM1ISInnY+roRYemjf9AtpPNQE
Zs+fx3uSfmClrxCAwD5t7AA8jppR8RgfEwdqkN5OG+3NNu5orxONWaYiQk3DbAuYzp0cR7ovmcGi
1PiPzpO5JidqADthrJ+55OO7iySR0AXB+rfxPB7wg1785nvViu6agoi+oY+LZT9YD6tqwzyVwRhI
o1Ih/ICSimFPQJnD1qxKZzHi/2MpDbNS2iVR33syutTczRFAPkxH+r46tFZpL4qutjFnyJdir9f/
8KGwqPdN4yge4hsJJZRmpJWK33siTHkR4rJyeBAhn23R4W0vjdHFh9rJjBqvt7Oqwqi4/wuYqd6s
gCwQZijC9RK+cFPm7aRLJaoIzPKqXfhtnM2weQF1ohNsdUnoJ2jFFUaTfqq6FBxQX9eomPBYFKUc
3GecktVRzLakKUkDxLqmXkMWlZuqYWp+13SuT8WpHKyrjd0Mh71FDxVQ4yxVYcj7YV+7V228XSU4
+YNDMB0htJxOC4e6pHo569G6RBlCI6D1crkS+IswOdij1/YetbubOyzKf5NKQxUwFNajT1a4rEyq
8448RDOxD20y8f3XwdUPcuPdMpdfwl+wfubvcDzAxfIYYrs421ep/eZ+/oQBd7I7ypVdfqDFye82
UI864+7rmJCIkvzR7Y0b2zKFzCVhze4bVGkDCWCPmMoyxr2th0RTSeYEJszEfiX1fz+iVZZeoGAw
DqFyp2lzqr7XNl8+78OgOZlLt9EZC/nBbJQA+1zyTs8dq+SiAesujxEUo4rEOwpL+I1kv590pFAE
82w58+gH1IsWT1/FIJ1tq/xFgqNgAPW6XqBEmF7PmJtZ+M4tV8q2csjkli7qe6no057QVALk2l60
PWBJjNlQeUkLRQGeMWCvJ6jS/RVp3mlL8tZdKCvd7UZiod95pb+TWvdEvgkPZIB2niWJk+ldgcBP
gR0i/xvTeYwfcguk+vx5e8zRT7b1ujlZ8TNzGvcJdhbg0Uf6KCEOReacxeIUI4KZeDuGSTu5XBTQ
EyCdn+r4P0zGqQKnXM74XiU40IvSkjFU3xqq1FU9AgfeU5c1Bfs0dTaxFZFhlJW1eTezB9vek8qm
cXSxYQ/xNRl9ee++ObNaXQWrc5sNo16NXuiRKgTL7/xq6dQ9w3cMKIjh6zgIBl3gd3XctV7xFnoE
V9Kj2Dbu4D3tmiRRcRkRjMOosPQUHiinbjJEjUxlW+S77ZjvBv3jq1mP63w+k+vUGx760zthjKxJ
SaGsWJlb06lmC5rhE8ArjB3MLQNAmplSBSZ18Cwx2VSIoAUc1PwQDm/gLsOqmresyCKT/YreI2hP
tKmQfG2O/bnJK9XwYzO/hxG+h/mnwZiaUYSqEdzMd27pALR5PPx4x+Ix95GF7p5YMnjbc+VS+ZwY
KtQXCHA+635r2EabuXAUZ+K1nM/KCabkQsduRz4oglACmdPCaVBOttwSbaWIwq1url7s+AP9O9DJ
jgYBGa7USfAWXTmsryA+j4rhX3/BK0Fn4nbQ29XxuuSka7EFesDW74kGOuvA69z734Bxod4M6I9u
uKwO4pVdppcn7eer3SW37hkKpVscPVO94WByLQXugsSqhPCSFZrJxWXIm8pFG5CgzfGzinn010A2
tmOc60gCWE9uTush3v2pTx+i79zB+EwBoo/MYEIB50b9kgriXtNk8WONOuj9ihc2WgS2jg06GEgE
eiV4Z+97eSx0vMBYpnZj1uo8caOBzM0O+dVRrWmgOgaOF9KhmU11rH0UgVx6C0cOAHTriJBJ1QsX
jBF+Z2iaoMWnzAb2rW41yCMEdRmvyOIk3UQwYwN6G5s5xR9E74Q8iUuAtoxTpPY2PG3eSo9wCYcr
tuGmWy/9dGe6swOYLLToNMKybB5wjTmOxpE4u+pNjntzcoi6WRb78JxZ8cyhoGIdKdrbQL4fzq8q
rkBmrk9y3a2XmrG6w9Wr5dztpKMHt3wICPdHJSQhRbr0iwr9pdF+Wy3VtJ8ZiwZfKULIm6M70GaM
g36QotBYnK5AyIrg6HDR2FrYscq6PlIwAQkhhfCDHvEASRW7d6VNDeM2QiVnqkorDQtbQhRImYIZ
ahZCvAJKrPZ/41eP53bIjp93qepuQ04yGJ4jgOtnC8P+c4c/nz0/1oxe2UGpOJl24e2RbxxDJCt2
cSa4qOgnNlQadEJUCU/wGWmvQxqv6sJE74zdefwR4FtRFouAc3TLrQ244GNaGC+hsKEz0MCCsnsh
MnFQlLyZ7hWcISnpMyXrjhYTD8gZI6DjhLIb9pSs+skS9DSvdQY7M5s4pIYW6uK5vl6kBxPRdGH8
ys11EIa9Ib/81WYjoa0+SqbavlILxkwtTLNUg1nEWn1cxuDDWyt8ywZv/InD6PUmAHqMgF2VWsHD
IGUS+YN9gZAPXP5I5mVP5N29Ad6CQeQmBqIUNbfG4HX71M8CwbPEvFlJuy6MuULL/yOJ1AnPtugm
rrgkk78AmlMSi2RIU6T/hX/fj5TirJqbGSdUHymO7p1Gt8znPEBLJLFSSpcjGGhzSMDdqUXqPcTi
RpfV7mnrKvUAyZoP0Sxqsq4X964Rn3ZlE5TQIMqptkK74fx8Du+PXJKekNi+Msc6NQlC8bfrCcud
cHgrq4BRY0Ga5NyXX4y2wy55ZYiyxnPAibRhT9liEvtkZAHyJ2EDIzhtcgcfK2X32XeGCT9LRFPG
hwE05/31+QYyGpuNUNPbBV73w1SX9Gx8RUt82GkwcnUQ4FbQnHJEpCa8anFKivfRdgJPokalKKcy
NwumKrJsyGIIOib+Kl3b6UozEmqdwpevOEBlBq5VxlAbTHnyosCqz8uhblAN4Dvob/Q+2g0BTEEF
pN8i3sjDMNrP4BMqUxRvBUlymXJf9MmEItHNw6L5N0fW8mAqM4W0vIwysujxzUtiQWzlNurZ96O/
sAmMKoBfc8cJIFF9u6BzEnE2RNd5GPQ2txKLIxJkFrX6cmGNsqqJLjVftKQwlfHJ8UWKtfnxrB+2
wuJvBGHBkwF7CjorNnMh4Mf7njlJwasXrPPH1scFJBhBwvPLyqvY7DfKynEplx6nqBPi0kU5dn7W
eJhoTlZ88YZTlBAsXLA7s/+u8CO+nG3JcqzO+8Y16RC+lPpcde2E9neTGnj48oGKOUf9GtGRaVa9
HUIWcjZotTocJLjogflb8336LDfKl8rlpiZUOu2h/9xMzf5ZKvLVlDVY3kQakVKrh8T/u+Oyub1E
0yFcFZQF5fYkDiGYVYURY8P7YZYT7q6KJz856OQ9YdKnUAvncN/X9HnvcyExrMJvRQYG1QjjBZc6
Lg2shZEg7UQx9hPFQp5H8jkfzGytxHnj/+4+2jDo1s9nz9LCaItfQ3MPgX9N0ASoM7LGQM2CX2J8
USUc0omYaoeao27pxOC0QJzUHXb1jtecPSiIFX8mYYlX26BuxZwe0haBAa17YjgQIXSIuoc56cUk
Dn0AfEWFuGp5jm+FZFnVhUoNE92w9/cDOeQmAVxZh3TtWVa5eA3iZ0HxhhGmswuaFlgqSfQWm2X9
GofhfSwV9A5LRnTA9dSRvzLuYdB8MYjJgo2ayqPjmad7bhrAD8wAGLWG1BtQwAxqW9UXRGuKIckX
e0Ot8jlHU/JGWi2GLOuGlsCfkD2Gu7lTnHZ74UPbITg3Jp9ph+LyImGqsffGwryq6TmkXNDaARhA
Y4BbuR9BOkeuBhZJmqZvYo6GFTQY9y/RYgmTFfTc/V+kDHC7fhq8r7Px9MMnpWeQRIumrH4Bfx5j
JhpU9e8crs3CngoRO7m/+bImtMMuCcI7zaJbL8MFQOpLHZ31+XMVPfDw8qcKQDpLKGBf+fG5kT/A
d0FYltlOiSuAXpyjfeiAdbSukHBcshqL4PEGC9+P/cg/7s9Dbrp6JSCtY+P+oIzosWFjs/nMV31d
90ilCTYAZELVMtocd+EZcQSUMJKCTW5gHecMU5LV8uIs8bJHCQAiOrC6HRusWc5Z0IC5Jk56lbdE
uUG/hbkW8TaJ3GKZ2rP+qdU8+3a3Bq9Qfs7imjl2OFGUsvVK7ezSAbFzreNL0dYWoUEVyupvcxOB
45H/QMMlqnpiLn5WMoFFicr4EYc57R+FZw7U5UuuewEw1R9mfVa2A230jOWab0paIKGWt+cCmE4A
KcQhx5ri8lWKl4rza5I9ZuviRonctDEyq+efysamwu0SBQyDKPI0Ni222CFiJbkKbuZEgu50QC2f
K55disVfBiwOd0wfsl7alWxR19O1ibbkdFCmF558qsnSdaCP1pY3kzg1rn5eypmWpAh0glUkF2k1
lEhU6ISPQrBF2M3BCpP+dP2HSFgoHytLf3ohPJcoIem2xuAt7porXX4kteuyAwf3ewj7XY58kUUn
DWyCcbduExkrZcln0dJpngMpAmSKlpnFWy1Ti8ywMCV/ip4BiPNmnq8TvQxw25eZPuX3EvHIf1Xo
NJhEiPdUsHP9zTgJcCV8Km548ONaReDVjBDo1Xe6+PbCrlpJ/HHQx3Gr1rl5v4wWbKtyokxScy+a
MJdnYMCAyAfGUP5D58U4W3a5vjVQelxl+Z7hVOvRPIbe+HEntwQYHM9YewitwtPqTgERewQL6OP+
5sogFxATL9shnnWIkjeSLQvjPWJ20UCBoOrlKeX37pI+5XIHJu5NMqZS9xQqs+TxrYXQgrU5l/S+
kk04Atd/s4JoyZ94ku34DhGj5mYVSRC4XAqbNdr8m5OcKzfKrqi5gBdsX2KtB6hblf+s7WDwxraZ
Wdh5/4xgEocGHg2Pb/seZ8j6Tn9A+As4GLiwD4nGB1PjS2zCqxlnQuXQX8edjEVbKvRabpmKS1Wp
IWe3BQTXylmo3eHKJ38LrZ1o3JftbPJjCwx9NM4dQIuc8La+dccUoyST9+bPv2OCph6BRzPehmhO
JFvMs0rHaUrxRKVzJ+aEuojZHV7djwXz0lUs8gHus3XMORKsjEEZJdtu+JLhsX9gVKspHqjTR/yu
+xMZuOqkpGnwSZb49317uFWV0sboPeKISMYd0Ot3R52oiWAfJnJl+l1AWIIrrbyBpjGd+TgYkC/J
JHupOWRm1CenRGX/PSVDMWLqukMFuoLEjkGFywSwuxO+v68y+z2s7lTh3B9eGAIBP2UgOdIbGt7d
+MbHgQIDfbhaB1vr1edC5WJPv2Y5DyMa9nW1KGs+/6FFb/pi0LNZKm4pBx8kCaI+GLCS2Epmg9ev
fIWzXEI4fTg12wbx7WeRLRoMXd8HDC7xAeX8u5DCjjYLeJCmlt96ksLsMBgZFXRWa04eholXUpGz
TcgiIGeSt/1ni+46zlQc724Xj3uBRLihLba3onTsZBh0QIGs1JLOP8I24ZwrDTHnopJMAeC+HUfp
+TbwimKxLxGs0udHKJ92lHagGyhBLqPNslA=
`protect end_protected
