`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l9rLb8eyF3AgALThasPiNG8/4BBm1wwJaB24bneaCtyp/I0xi7SHB/t0Ctv1xqonweX1MzV/pVKs
tQdRNspPIw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X5KWlL148JabgR5weT9wBUkHFWddJA7h4OZFLd8bdBf8Kop7kg1WdkOhUDgmpNTHeXS4I+xH4Y4Q
HjFAExnYrGUC1wm7p5WVL3DFzD5WTILYoEImzLFNcK9/mSAIwCGj+Wtr+9xrMpQDaly5jC8Sj+rc
Nr34z/YYnZpZdFjSjFA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XOX+x3GXJVQTrGGT75+NpApkQTW6W42cmWaYkzqsNsDYv4er+FitAoIemlb3od3AsSf9WRWhCQnT
6iXQilkemT2DzV4Xsw5A/7I/FZ1E441abMpjv/w5Z3kwpJvNtJvcGvjcX812mAAPcXsPvrB5LXuC
3JiNsCaNzfl0IQulHvHCqzDHmgFxZRkHPXNoL3EbdAxxa3qQNIHMXziT6TfG6V4ioLwZkfmj+nFw
X+PAA+oZbdjyO4IF/qvCl2mnZ/REv5vdMZsnEZ7xmZVfOO9rMWwJcGnuuXesJxcZqnyEOewdy0X4
g5x7ACzMTBvW4JyAsNl6ipSaUUNJcxvmP1Z95w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
umhSCUCmm4WZMMJVCjLiDlzFgH/9KhaxQqdvYM2gFaFK/BSZmXwKtVD0oGzsfgEnaEnfAZpnMH9p
W4FaTz2HfMA8FyEQD6bKpLwcrFDP6FLYTus4W9auRkdWk6MByslYcfESnbPd9BplDCjnq5X9FeJm
J+EfUISXG1WULY3BqQc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NcJ7q/waCn8/m5wYTzYlcTzCH0J7XhsrCXDcbP801wBgwPzwk6W1YaeEGpz6w5sg9/BVkYMZPdHy
s116tGvxEU4yIAoLSq1V4khC1G0CICk3cYOL6Am8EnS97sHVRnu2owQQ8/o01YRhaorvw4ApXGQo
FWXh1RTAkyoxms7xpWs910xGCq+5ztWRsH4I8eissSMkhuy7owGmA0f/OPnBvz/16ynnHSqeTcgH
5zrPaJOgTZH9aMea2bstTOpguVDKDnDoAXUHV93yikhxVZbDx6GaPXUh5fshHVEaMG3kP839Gx+j
prw3SfsWydM2YztaOjt4rwHOeUOZ19sYd2Gsaw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9808)
`protect data_block
GMQYRLdIBu3cBPESIImpy+xilfncLnKrvhSWmMznyv2uQpYKLA6mV3Y5FYPc2Vqnu/SBmj0f1XTc
+Z5bSo3nCRg9U07rEnuN7EcMhxVbeP1KBOwJhcaMwFEinh1kZa0ojPo+tfSt3fjUy0PpUm/iTAcw
8aBtZ+J89lZtHPC/vDIHl2CZpMhZEhEJCFm5CvLLhCOZxUH4nn2KqGGAfW/xDAVHYeyJtfvKnkTx
BeJThs6rE/1o0dRI57M8PeE15Th1+YX8AKqQBaNmhXmhoPI6ewDti9e3qhwkmo/l+co7hTT0FyCW
NdHouM5q3a5KK+nqtndPEJv+yGAutba9ZkafY20tQknFU4lcEmn3SbDnUj+np2I3qsEKtBzEvFj3
lZnGInbqlQANyQ6ymgSYiu5IIcXFjzuXHJ9Z5hOjgY46t5ErpGChRp/b4uz/3Y2G03VjsQDESrL9
7CW8ZsTJu9Ma4GFi92mnTFB7WdbR/iFnoyLMXVPzDwzFR8oQb7r4qdIaP9/VuhsPnI+mqV7aMMbU
aSwms7SAKhVpyx+zfAsRczIxplngvdT3NItqqHjS7NU0GqRIpbW9d42iqarYwoeTOH7RmMUtO7FG
KhMDE9Iwd1JN+XKCnWP3/InnxLqUP4Tn8GRI+6ZHP8b4RrwHySE5tfh0fsibWU1CzKfU+LEweSe/
aKU9yHYxQaqDuPp7x8KVZQJdMj9Jv87+w/YHEXWXjb1IeWoAhzmEGL6jK4/v6aA8CkvGoElULrA4
GagazIEMoMeHjWiigLqZqrvNGjEkbHp2CLq23NlgvGS8AmI/IbD7+xM3znUrCzDExB6rd+HYXfLI
A3JjjfK7eSXubW8CO1P5Jj9WotshgdTIZQT9OkdSsJxxxno7LHPxxSHrtAJ+ZDG/MYJUvB8EFyTr
0ueRtmcDI8nnMEKHGaY7ziF9E6TlLeBP3gangjMtHobLVNlVJq73gZ7NVH6reup8tRHbem46Fm9T
CDvqXChJYUQyyAXPRRWSmNl/7RyEf5bqLIg/IxBGIU5Gi5zJ6JQy2ii2WQt/TXPlm/G6WdbIoqgp
64DBd3ZXZlJ/hnfl/NTx7wph8sabX7PvOIRJNMfQD9CYzCkQ50j3RIUp9lQXbKEuYniUMrUKRfOm
9Yw/N7CzPJANHLajiNr8o8SaM1OMVxRzL6ZJC2SuH/6zf1YicGrBfuTnE47clktiYVo7KeQUauGO
A/DVqKoc0Hcs3844nbc8/TgO5oUjJ8YlYErdjQddwa7WLWeewjxCLphgHMMZtbXBf2mZZ2or+60n
z1ZKSNXsJfFZs7ff1KSjX6RB3W2W7crU52gJAiW1faMSb4eEeQMNgGSEWpKgN2c3r0qyAVi/vJoS
vXuCTs+K6fCMfiTBZVKgG9uRpkTS5sDuZpVXp0cMW9jBGyMdy7XhziXoesc0856JeAYzjGrHzBXm
m3ciGdeuuqh0ZAp9safVQQnkBmB1AMZ98qkFUoNztMsVHd52p7hG2h7OGdiOptl99NQerYeLQyHC
jt4JNg2UI/2yPWBVIwCQKKlQJ7pUQWV+Ua2PLR//EQF0xMy1UBIgUL5bLp9eu0n3CGe2OEb+NyE4
y10NWI8egMO+mqaP4NVm7xZ2EPBRh98wA4fueFEBNEr9btyjaI8hjR5+0ulyEXMiCCTFggTpbQq8
vZ/SxU7y43xilQEzjJI4Jj3tVb3hxlQa1AZTXofymHmTT17ETHxv8Kc8rQkUtEm4Gz0qrXTxFarr
FtuY6pugXDb7hiTGaorRYxjXOtzqWds9nDptOEooq+yvlcEQeeK/4iHUppB7czQ8jVr2DgqrxPx4
gFioKSyrpgtA5mymvvzIJOY7u0rWoHkIreHH2XZYYNYcBCR5zHxT4T7ce65DFXx57L9Arh0leWSL
m++3dKhq9zVplO4Jn/Y5FtY8xcMBm6Qhw3yAbjObqyfY4wLLOCpcgiR1siccEQFbuV+knrkl9lwO
nI2KUYaWTmgI9Vs6yjlAX7qy2Gq4+9myco2LRBg3XLLAVoMTdclh5JwWM/Mi0Lcm4GNqsOCGABzz
F+RQG3QNmFCRpI7QYLBI9UQ8OB3GkSKup/xqhaZETcFO+SOpv5+OXpshP3ZooNj+8oWMXmj6Lul0
I2SL97QheXBN6EarVwveFFX0lluL5LSE16qJDNaFufVR/ZC3Q01D92YDTBONJDJ5rXPlj+5MMlbk
ug6/X/VCiGhMgaJvpIESlDsP3UPkaKF4ZPgKZP6N9Qfyl0SwRVXaWHIJISnvzPxYhlPN6T2ERoLv
sQta2TvKcoESqiL537f29sUmj5KwiXnH2v9s5kpN+iP88YsInMSwGSjE1jsEEprVY8QFJLTePz0t
UEJxX5cKpYxELXRHU5io4M3xfR7n7H6WqDeRwdfxcII8tnsiQ6nr7ckvujvyDcSELVQyGrcHvrCu
T5nik1vYOyBMjT3JSZCoVw0ri0oHtOxrn/jgQg6BpuxQI0z728IcSmxRXIli7tr/oUkK/+m29bXh
XNjA4E1x+cTPvlFkt5QgKTBXp7Ok/l7vTBidphZyGck6nW1R9QU9mOC817Y1aDpVj6oqyg6ZU1fz
zbp6HgxuTRqeYRHlTtwW93RV9nJCdFvvlJLTJBovTO88hBx/TFGQnd2V/XEGMkmKwvO/dzzj0Y7s
V9qEH2Rm2BH+9Slld6DyWcORTpb0qxnYXposK5oCuM3TwqhiL3u0Xmc3EVgICTSUAgNDdydrof3e
y8OYDgSM6NG2A5pstVzQkXgFGfpb/gXinGq/QoNqg692zkWrcIy9EAatKvs+Iavzp9hqwNM8EHRh
3Ilz6vTT0V6TTMo4VTfOw+KAJh7wAlRE6PZF+YUWbXxjGaJcuXyJmch2kWvROycAptxmW0oSRhGJ
1zlyOQk5vpTyoMEnwyqYfQn3XCzLXkmvxoAj19ZMDODb/k8N0OQjk/SZoLFWoMF9rczeJ8laV2vZ
HHXUYPIi8k//XIsewwaLt9TuI+gwnjLxhdHBB2cbbfkYs3JSEyg02O8Jjufgo4EChaaULfpDRg1+
tqupOVElGzfEN+rklei/yTVvkG8tDyiGeYIL/h9UstFTo4AgAj32sHIySfJ3RqL9wRpLlWDa7A9X
UA0blXF7cM333uALWqWa7duIFN1jS7TNtVXYOJxhh/hMvoJ9ZNn5x5VQmii2BlYRAa3+RsSUnvj6
cJU3jdnfj/cdsKN6E3npue/BoqUN17Edk35g4uDted4058zpQCccPwJt00TzBVcwIaUIxMTf4Cyz
B0ajL5M1c/clDhl9aqhIuOwy9nFnAAFsX+nRABhWqSa9MdpfO+R9xdwXFZezTQt+HXAnNCpmumMr
aWChiKgQm73rGtROiC+G7HEXNbmZp+eUjPRpQvWHrpBoQ1dbgxfqslH92EGVr7IVS9lM1TgKXFMe
OAotktdwPKLe0C9rSlPf3zgDdICANzIX39B+DQHhpzieHSjUVsmlRIYoz+hrvkTuN6Ey9bdqxv8n
1IkyKoO/kPQgXPC5I4eTAzPTK8Q+gDS7tzpkOPTZ4+kIiEehgg3A4MPnH08S9diGQePW1ALlyeZ9
LSoPgtIvSH/b21vE6hrCCIyx4PE4t4vWp6qqbdf/Te1InEWsbrLJfJJrWLdzeE4yHyxqWmEQmRXe
6uwUQYxf2WznBghlEyyBZssxhuXPzs6WnDwMZHglq8wSFy2+lH9mBfokG6lnYPzUceDdCod8fmAD
TZBa+4+4eToemW+N5sYh6kGS2se+p3QjDq2jF1pvZlZb5oWzZpARBDj2IB4AU4QvvUuGWnwCiEkv
B/AevDwcdNu+l0vUPG01f51988j5qrIjNOO7b6sNa8CvTnpds3v/nKrXxofdtGrI6fRpp+TpmOlO
bAKyTsqxU5PuzQu9oc4slvTHeBpyFgtHOmAOiwu+P3F1JVg3VqxpUxKq615KxwFlDq4YMORA0nlF
xL0AH0TXRJ939uMkjnYkrMI+LA8Q/6fE1In8xezRRizZQKG1JEAEphMenIYdYUXladShC4yorgdG
fxsfyp8wUVrIDbrbHjKu4gvKpistjwRDBUnAZwSpsDjf6ZyJOna13LVvUfI3i+DixnfFNlE05hbd
K6SfNEe/RzEHsqXv4LNyd2ad6kJ2cj+elmZIo2xX3HWd1qiNWqmBNidJmbkHvOD+UGz4Ab/uhXj6
l+6uIr/lhL/n+seePp8o+yCylJE0pE1P2ka4E04ma5ot0tMZlvDl8ulLJySMgpq3QdBBW+Nvcdld
DA0OSiPWfjLUSK5XnsJwmq7HVNylcuzsCZM+p/yT30uO+YHYa4uC0/EXCfL3RxH3v7sf2Obh1Jed
c4uiVELTvz0hglR8Og/fSWE+uMTQgdbimGkuL8+c9LnHgfAWhL4mAp+vSS9Z8FHmGM6rn+93KJZv
os5+ArNgX7A/cT33cZfAlAeLKL/ZZ9Give3Cs+LEKWyKsPZ8xKt8L6j8fxAikXoRJiJt+4B+x2Fb
5l7OsiF8hPFGVSPtTvrsadHV0w+WvPJj8ro+OJtUbv8eZKZDHS82rRbfZ6IQBGZ9/jvIdKNSTuxe
qWscpdswWF6utO3yP/v6rtMt16jw+gqC6Ei8yUDri8CHD1und95Ta8AYl4mOBg9R989WPEklI7p5
FpA7jUEdd3Eifz7S6iUJ8vMs+OlgGn2ssF/ceJwiA3hRgV3b52IHg2xvOyPy9wbG1XvZTn+1O6Bo
LjCEc1ug+ej7MWloPetyAJGrLwUsxAxf7elnNgX9nMar0CHBZkEsLEWuHAeePaVy0xOmUPR92LWg
2OS78j/QlEpgaWxbB+9TxcQ8OyIR0OJlsMPfdj/MazCdsBlrFPN1z9HWzFQRbnK/2aM/9/uMm61G
3JAJuqSe8qZ7vyf0FgXcv9Py0iYcoH4zRf4zMyS5H48DkORzF/RBailjrVsNEGmmHP7ChDn2IWNB
iNr87/9khNqYuiUchhU2oY2v2twv39uRNCoZcbNU+4vt94VNtiZR53oaKKJOjXrBh+u+7Wqjthiv
fY7iTJYGugbNL6vyBpa8cg/MuF3xrZis22jjSirE9xi8jIA9dpiVMMRUzjkfWzafOJN9v2HgxoTs
jHJKCWo7/+2lMxi8DCb9aVdZqnYYqV2K7jQSNlRI2nZycf+WH+s7F9gwQ565ov+fZ4LzsEH0KpZh
g8w23vTE3pLSVXf6Qnfr+3aDnBsOvy4/R4UU1WiDtvs0dosQfcvEPXc/xI7FOcmXsPK2dSJ6R2jk
dqSNfA3e3MaR0Uh979x75UT0Repc05mRxqPFSjiv1cSnYsEuTpjE4X62VYKG3+rVV6Kvl6GYXKeT
Zdg7QTFMQW4EaiwIVLgvFw3j7131YhjN4ENRaNO/JUjnNz/kYIM7pLilw0YNAG3qOZHrLwvHhD5W
4m8AngKRiFqkquWswm5KHjFjGIFz/Zdk4yP1HwuQTSTpQtGTvhWZFP/yUv4XW67gmnQhoitDwYa2
l0Qb+OzJpErDBIV3pMnG7hiF3eJl47P6WKgzOcnlZrxmYVh8w8/I0ODnhNJS2cEk1QWgrwGzyH22
Ulqiw0N0+CK1a7SF6TOpRyb/hcT9JpVMfx01mH0ikyTXommIfjYaC3k9i9UGRmfigaEiVGbt1Uds
C4yVOLWoaZiDs5MdcqL24Qy4EjhR6chdrpmISLPOivm279j1PNAnjhSu0T5rlKU89++SZ6Vd9Jtn
r39acO2cRR8eaLj40Wfh47Ps0pSQfifZxrsBIJDkbdiXz+3jJIFgODbOMV/PCK2g6rDAZ6Y9RvuM
nRTEYxdhvbHMv5UHgS6D1WMrdPHlzH9+moMGNPlE7KofWiLNOMl85+NJsdiQ8aHaLg0jwGVMMtn+
L4rlHB/VdwpW33GBAJ7Jc4dttyXFpWRk5028Eiqsxvi4iOtGvSuy2CYC7AO+4OoqaqUd69Hz4pJo
licP206yrmGIFociGrWPjewXqvFO3u8wmqLYyQI9c1i/9qT/w8KVTy6bqUjHOfgnw67J8YckcBDa
9pUPjo1ONzG+pZ6HSNPE3SgPWnkKLHQMXF2YIaV+zlMlpul0mwN4w4Kd+7bd/iUh1KtH23fpikrj
hx4u3BrbO86EuExmBPjOTLo72p0rrWZ5BhnnxjTEQuWAFtD0nu3paWCIyDgzBFPaJZjSpB4Pc4QY
pe/ps/X/sfVX2cuvjYGb5hW4rU2wtas+vLkb4W7vScQLxiyuZCugQvPAn6znewnS51h7OpF9rAZr
Rb9kKVMOE8+kxyT2JtxisLU0jb8Zg2PZYuyaAXrQL8hvquhjtu9vNpGmEY8khPgRZcpaqxUswuYr
fQpiAxhZ2P71poJ+YGLO//SBVeYV0kC+ZWypWMhqduZkzt6zO1MJtU2RlpX4FguR5pNUT/qtvawT
R3TgvRx7vgClyOvkKQR/jPsqTytP/l+5g3BXlItfvOt9pKFxombuU+6FfCk6/+qSM04Zz+hP4dMM
sqXcB2hmwV3WSkjl2xur5C0iefvmzCSGU2LheN5FSRJwvqMfIEUpEaschK78y/UGGTf/q7LrYy03
eMd2iVhu3QQW+9j4SG1YFUcAe6PpGauvTD+e2sl9SdeiXrIgaQny3P2pRCI7qITmVdDyIKjxpde0
S1l5JOCyyW8Paj7A63yqVls4XKpU1qLmotMqMDb3lfe1UflvSPfWOcwKfDDG+gzCf8FLsm8mKPuo
ywUQ3/pep1xo0exMjpGMcrfG1q4XoClPEKjc7RVwRnRhIB4Fs60gzEV8cD/ZeHdFUWgTz3LlWmCE
KHiOKDsL5K0COjn2Wg8S4jm2n+5vNFAtUzyZKFJIPCyd93u47o/8JdQ+L/6lhfe1S7fOb30swnKu
jajMPVjvUqz97Qct47TSyTFCxuRyEqxvEydsRkhrJ+4Zf/BFzy2N/J9wbm6CEcGbwt4mwb3WAPX2
K95j30Q+YGCrsRYiNfwSKSf9oVIAJBFTfQd+B2/NlELQl9i76Lh+rbgck8OvIE/ytZeGrxnhXz5R
oXDCYzCPb9AZ3XQFEa7FRS5c4XUt17j5ji/KkHvZFebJEbzbjxUfBKLHpF2p7BvLbXUiQcAQCeDY
KnF6tzOU4vzz6PfOGEm+r/GgFV8IHZZnLNhjjhGtlwRI48zhHHH8r6BD6Dd10e7tsPrRSwHQyIt9
b/jOzdbHXxeeawhGNPgKG5rcnsRqQSlqWrCUNL0Zcp+5VI5SH4ETWzRd6zUiJnzZhbFdlZtpuUAp
+p3z8uLG+LnLudTTtPWRGU+/Q1gWuY13hhiHm/xQzBCn4yCu51ixVKr/glieZPzjOQcpFD813+N8
acSZ764zQ8edFIvfEadxZ0TrfBRbGrkoywcbdCuHRUwOvcBmgeLTqFndMpmvP8l9ML0TkgLdud4x
iO9R+4c/1honk79zsA5fMUHh0hWpU9UdaGW3Q52EN2QGe7+NKudmIi/kCCbIBq0sMp5k2+duBktq
QMRaRpWIh21B66zszqt3ravaM96el1CL+XF9hUv+YzEPpmdmHaybzK1kVcb8P2lVUszvGPAuz9Gx
EOy+mxnJ/bj3BACkhfqo7f8UBDBUkRUNVQl5VBAr0s5wVO9ju8o20XKvJHG8LnCLXzP3xxfbBOxV
ec67lO89VXXF3C8lOXwa3chWMfcbd2SLzAUhRzsc/RWAXKFa28INXzvveLTAa4HdAnXQtU4w5Mvw
sO0ITM4qRV7NuwXSUp2zfB8yr3hcnOLiA18ONsIFezWm2cqVfDqUodFXr/clBsCsuc0obg+eT37+
MHccTmwSTM9B3/N5VBlWaymLihedebImgafhWN07aASSVzBKMrn4F6Vrn4aTF5MhgGIYqZMWa2wl
VuI1VH5ay1ZAZXsfO1jOgNHS1/ywI91BudyjHSdoIzNcsjSuDD4DhFMrkrllnVrZR5M13k8ZycWI
9SJ//DuhhieTrY5mLhGx85bSD4tiNhJ5vWg4wIpEhRDD3Rx4wy+PwtoXRKNiqehnZ87O/4HaBQ8g
3gahNm5UoryuLvRkkDbRGp5ek4v3zPJZ1GvcGpg/sDiunkd7xB1eyfkLmYClpDikn45oLkc5j1Ou
BOrBkIlXwB9igEo5ior7xu24LXqYbOpwPKecvoSepl0s+2Ykcyl1AUEBmZmGiu8Zpp11MMP3QLjD
+L3tFD/d0Bld3xPd6MJzG8WX80MgBxFKhNI6iTUHRwKotnrtwQe7X2Q0U1vzPDPVf6G3UYJyAjzJ
lWlVjBh+knJ0ZYtQev1gU0iCiybQc+ArB4DmCG0zzeMAN9MFVo5OkBUHnEeTODrxrLlZAzOyOJmt
isAvDVu1AbCKJoNLErbXnwYKkPc6ohErv2g+rkAkqfFP+qYAx3A1rq+vvAGoaY6h5b97JCBib8uO
rokJ1pQcU3thM/ayNppro7VK54vwNucI6hyOfVmrr4FnLddvdZrx/TAKmHRJ34FZvDm0EwcE5Bwf
4x7om+iSefFU+xIUSflsX7dMZtsGUlSKYLLk/yMTZQ13xTxMJRQN5vJ64RwC9zn1MUzzcSbG7xz4
oGgs6Q///P+IEQ1tAfMVTzsMd6Ls+TsjSKxM1v4pfSElHgvpF+z6jz/aYqSTb6h9xK7CRzgt/6me
DcSKzUQCashLQKqwT+P3jiQWjTwxOdwQ79qmPuyf5qVnHiub+eQkBXh57rqQgAEePtAs83GfSXRr
y+VWecRvhzyJbC7rtfWvkDgXxgw8dfPWBEgE+YzPBj74yRt9FDIdTVj/H0rH8wFRMySD70ybgD66
+3jKsvO5Y18WtODezCtHGOrll/+V2aCat8b6Wpxv1UzkCb4gQceIhLTg8IYF3fGsAyhHZERIrm/9
IB4ij8crarHddnEFS6x0H3eJUfy9zj2bvExDSKBO5xAf+TMVcowezAdF3PnrqI7n4ZacTeFSNyMk
ZYy0EOxtOISlgUuMPQhAlHl9nkQVZZ6QgZI/sC2ePq2TuFhVahZ1uQY9dNcOf0ToSNv25M2c5W6n
dDa9CqzSTabKWEaCGlXhnCSkWEeELtmICyKS9j7+aru4X5UVcaMCGU4OY+1UQWjbKfNHb/Fkt1s7
5NVTsYDciESooVq/zBW0b71YqazOfA2YZzH3ZEi3hezTYpz31yrmTj/qQSoslKvcXkUQoEN4tK8H
mRnwlsuAxKey7TqjptZdy8HMLzwceAnpUZEA8H/NAhq3SEkJ/5s6sZl3lKwSYZkl8A+pfrooag/7
vUw2n9c3QY7XmtOBxpvFrLCz50GymGI1MWVv2ttIQGIV2vfZgNoVpvPnxUTOPqzVPt6Bb+Bcb852
HR/yuhoy49oGwkrY7tTwNUUUWdn6sFfVkbCfROxStrPLLaCe97zV8JofugrgDzYZCnWO7XGApkID
0SZAuXwq5O2iK6/6EIJoFyxVo1EciUTjls9gQEuhtdCHHD7UU19/Hybdilol3kvEuHqfTA4JV/sF
zaC53nzmtOVsHoDpzC2ugUhFXgmcWJCmNvmrHULiHuJFd9BzE7xxiAPprmaTW8tckwUpUFM+GObH
x2XMJtq70ej+axgP7zyv446T0h1B5JnuJ5FElGRQtX0poKb8hRyLa5YCISPiukcKHNVGzHSixgDa
XHPCWAzsJUGkT0GfhlyBPEDUL4aHgEJ6ZFNsaAZmUBuP+FHULUkKXdjWbhc2M+TAenNq8EJAUgws
vPww3LhfYhKEx3hFAgwG2XJG9HCcyH5KugRn3H4dKVOSEUkiNJaCrRVsmlH76ORr5XjF1Ajz/JLC
7k1XG3ly0qBwImizl0BG1y/z3QvEDe2thLGCs+sJ4pwRVwkOi0JIiFcQsdi7yfZx6jZqUfSkxlpy
+NBnNwp53qzOcwLRdnf/NQrr6tHM/SH5i4o4rwDc4afPMT8/csPVfipz+jWxOsNATKpId1yM598A
E61+Pj/MnHY4DcSSQQ+BVWO1nOhHfOrgtaY09kBhQPMCCGIrgIBLWwkNok1eylogQ8q1wveJRg82
kFa4sIuC6RlfxftzdCfel7fX6sdXn1Jkv8XwpbhJzDKsqqZnD/DJyCjky3zMxh/pUy4mkwLwfWPR
QKFkzoPnrlmLtCKrQ7gXCIopMknXplHMSnIS1pitV0j5xSBK2XqHVxjkkU1yVZKW7rXT7P+vluAI
GjEwDNYWYXXMx+t84FoKE5ek379MfK1aX9FBIvlIPT67uZO6Vjb2g4hH/qgXeIwOfPQbSLOvemBq
kpKy90fo4AqL0/UNtDiIk4Ek4tsQ5bptPKJz682/1cAdySlzojJlz7mfbqSK9cobYGuPLcxlYGYa
pinrUYjygzb7K9AJJ0kAD7PZ9X/jEpLgZI30JznUnw8NhObmcoK0Pu6ZXUFDceU6XXAZkwG6b8Wk
j9w8k92xJlhHt/NJAxfXF1kFkPqfZK04JM77KzNmmsufTPu/nqLdGxpG5QqLMZSfYiAqq9k2145D
NnQd/EMFLS/dvttRET+lGqmwstcVTGazkJReN8SrLUbfi3RE2Re+fdY1nPG61D3JVNFX6YYXJyGR
1ItT4fSDsUrSlNdM2hdf1C4Z8RRM46Bgo7PjxCJkFoHgWkCc3aLYEyNGLv46rvoX5MrIgt+ZUa+D
isSIL3EhxmL1Bva5dN2Q0AtZD/AQmgfIa+ZG2lrr6aMdJSobZywbGoX2uxI5eBlPVXg6kUQb6avX
MDcKhYU5WeYELU7P7PuYOX9Lb203nm3cLJgZbbJIpbPZxOS0dtKVIQJp+PFQ2sZKH6BFfoTtp55N
zqR4fxDEfz7XRR/rv9WbOhykKVdOATWs+g71mmYtwWo83ExLir9kkVsB1RrbNlmSPpnib6cnQgOv
baM9sGB+vVPgSeUsjjKLZ739DN8k/acjlLhRypllXO/uBB1Z8+RRmn9iCwWvN12ZRw0W/rFA6kfo
fUgr+3Dx2J5BNHPbQGYmBWGovOVcVKKozDZBJpJhLXYfvR+DtaJdFiD+/8wSsTpJ54FvKJaHe9GG
GW18gmaWXgVCiWTc8UNxvkeKVep5FdwQIoteOoSChZLCGdvcVcGnGT6mWKLNgHb43eimOT4xDxQd
qWC1ZAJnrEDWIEJz/hp2KwQiHGlVW6zj7YiXt8lLnlHriyZG8gFbWflf7WETih0anJ9o+2hdWDrM
A+UNyzI2PgFOa9LJdcXMu580CECUyXgWqxaW8JgUYVJXySI0T8VAE/Sn6MdR7YUYOJC0VucFnTbh
NdL0KmRIoj+LxM2Rxe/x4OdUifxYH1JkYHnlSwRVKoUuFAA0Z2wb8xvtI4ciI9lxOaZEHW3kz8mx
umxPgv2dkz7ZeXLZo7dajYwUs8fw55AAh2LRs1MlcQ4mhMg0gzb1JsOKCjwDEdYu48AT6pQXZCE4
oIMncBQA39HhrOMv9PWtlCTQOYZDC0h+WLnvOS9adqv00LjeArgGT2r5W2v5smlm3iQUTveVyPFx
LCsZR2W9bR197cK5ace/lhm1CzP/fuz/18v64Dy2ElTn5FjAfq1/ObE94fbCCCjFFDHFnC7Psq4z
9DCF2Iar6kbXpzgRY+7cI69oSNnI/TmVB3zqZ0Ou05cyNP15TRUZQeE8+QjapoIaSBEyaPrQFEdY
4VoW2LBpwytKiFS1I5cSxWTVx+SacTCTzecQLrvVclhHfIc/QeFM3nqIAeSsZc3x5vFgEoLATErW
UMraYh2GJBVgBWsHG/2cThfmn5IVmh+TAjUQvMmMHPtPbvU/xVLlboyVx8f5jVY5OhADdEkUjLr9
2QYdjosY+bDcp7H3clvLkF8h+jaEev/Kif84egCvDIrVmY7GxYBda99nlOjocKj+FsIh3KSW1pPF
VpENR6AbX/Ax5g8du2j/XQHDNvjua0zqVUOwuhP5/42LqM4tw1LnlL8Ce3KfxVIIWdXzsZcD9ge9
hwTPA6YO+ysuhBI/y348BM5c9ws2/SXQ0sUkz4Ff3Bf2C4NR0JxUXBA7kh0zkIHWxNYH2jCMuu9R
3HeT2CPhQmWEV1/22dek5kaek/msMM0FxhhtoSHDOb0XoHjTaD4Rt9QSKH4uyUfnos0Cn40Gk7AH
MON0e8a3EUBQ4oClKfFP6vSH4dm2zQMLjjUI21uDCjVEXUEmQbdKAFIds6W9X8aN+n7viYEEWjrF
oaBicoKKaCCBWK1vQXsp45ZdZUPUSKamxyuvaiMg9f1av/tWuWO82KwXe6MXkF0AQY28FxK5wSPf
+zRgXTcueEd3FuEjEcMFrNnjxrCYVimmlaJJsNRGJ82JdE3BQD/ODJV8W/JF31fYAH8tBtVF9Boo
RgjYURMlLsuVjFRRdARETl79N335QCaTn8jaU/0IetVJf9lYeC51mEWdo2lwcrB8Ea2jw3aECnUx
YyyOPb0QgbqLfWzi8GjfkYGwz1AoLZxwjzMp4yiqOGRjlZ6yonE2+cc3Li9Tq3QwcNpfGQ/i377c
uIC6aWWDMJotOwqZrVqX6/sR8fIFhTlq90ygQMo3iMCHikZe7W8YDauZh0wpOO+wnNlLplGsdSpF
fbDnpQ0zzzM+j4y83nzj1OJwW+xQknCxAi4riUhhIZNZMxj58nlv74TBeheRslTdvo/FHZCWWZ3y
Y8MNF7YvcbD9/ysAUAq46qy2lT4wAqszeA7IIvHAqTJuYsJW3Q8D5Yw1AShZ2iNrdhyARq1Z0AbD
dVof/wL+TwHCMikb+1geCMWHjv7pw8uviIB+y/JukrcKzuHPWsqZR3LwrtxJuXwHisR4RvMm+uZ8
Rd8Xqo03/NltZnp6usPjaQyaOqo3Lv4lcxzFAm997Dml8r6HpSQ90bjs958t4lRLXapQLEHrR6Oz
qVwRpj8+UfYsqbevtPHeA2w2Bg/N/TcEPgVHfCy961GQ1iQqEn9xmlbEQRYOe74v6sC+yVR9gM0S
6IPrP4XNvXI3cNzmar93jaNimdSvpGjGVR1oRy0vt0C5EjJNHKdyH2Hi4ZVxeZPZszZDgnpnrLAt
XBU8NINB6XvxyLZgZeKuScll+FORJBNNJfnXViTbhDS423+tXRkyYu11uiyDFAC8AW79n5QbwVok
4AL1T5gFBVI8lJXw5YJxKeushJF0G2Vbmk4Penwq2IXeQz0iwX6UpkrxaPpOgDfcgI91uXxM3/HU
rPFMOA==
`protect end_protected
