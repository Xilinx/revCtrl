`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35824)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbkV3TO4Ee1mp364NJ3ApJ1FbWY3IB
02vUs3YLSDgyj9eUBKSlf5PAlIHujQwvWVgSVDz+iJJGj5Wzr5M9Se9oxXmJiqBPOARnpsHODap7
BzJFERYKqccAykO4goJ7Iszqq4uwwoj5pwlPqKSo8bCySpVEOnuvsH4pbUi5Xr18wcTwqLpANcKn
kbvOkSWGCCDHU1W7lIEMhqsj5W2cYCrUxKyGLMHc8KOC4XPIl0+SwFK5AvYU0el8tZNrcsyAZT/F
fXyqxnf9gt8m3ylM/tlEiT4wrmIvUCkQIzc75P7MGX7vrJEufnIC/ycHAmwBfTi3P9H+1nD5f943
vRMlPl9Twl+g/v5g2ccyLSVr58MYqooPCgmsSpk12iwg4PBRsItnoWXvGQlcanEa39C0UxH2U1zl
UfF+ad+0uV466VJLx6JroClaiM4qg9cHrR0CsXRlmD3QZoBACpidTXN9nRn18UAkCt16AvQVLTj4
hZZAJ+xwfxCDrjklXU7OXT4IHlXjVMDCwho28ohUO9Vk8BEq29XcFmKXIUyio7iUsmuJO+iLXzmd
Cei1GGjHvct19WuMgWxjFtCBJTwj4Wr8Eg79b/az9hKAHeOt6B5KnbXqJozXotnJpqCMrAM7/Eqx
C5grDfJg3ZWs4lIsKQaEgIrkxd7mkZg37keppx5lXGmZ4YlLS8uHzdO3vQAbUb4N7PLDUzSySydB
kOT40u+NUjt+B7IpxItpUQ87AvOPyS4r57Ps1zedSJ5VTi9Nf2HChge0h05jKZHM/t7JNEN9sVrL
y49qp3vbZgPD52fDYZN6GoFqCuAMTxuW5q884lGHgZKydF2OsZcqB98kfeBIyCZLsfEnO6r5VaiL
akeQC7BXSqdSBR4EakxM3ZHRLnEpbFewedcn8xaYpRIQx9J9b+l26u4h8KcsZ8UeBZ7hH1sakrlD
Jd8VhOTpRV1JSOGfIVODnV9OMS8NwEXp47aUDY7EOf+6s8O37cZnbZHwix/Vd5KRXlfv7b5wo6V9
If5Sym2lCv2n2OegIUIuhAOqLiB/79zRxaVkQ+/EIFkDP7pN9ureuWQ4OKIvkRG3JhBhhzAkrhgq
A5ptG617zYYKdzCHt/GpCVcqlSDd5432HqMgyDfdIG4Y2ZkWgFqxlFbaTqJ0aUR6V8/fSxly3aFN
1q0J6R8eP1PdInEIZTfFATzva+VcRCg8eyCM2fG8M56aeoijFzPuYi1/QFI8sdqCzYOYUEjKyYQZ
cqtJHT0JqAjUpLvejDQxoL4OexOPNFlcThFn8Xt7gjV6brVzh2z6uXL1BJClT7oWJ6jeQh/Gh19c
6Sx0QfMESVN3ZP16FCgT1GrUahM6Bq9iKfqNz6yXr3lxaUyIYYwHqU3Tp1aWLy5CfC8MApTcYXjL
rN4nWaJYBy0mLU3PSSjvFKzduJnD6v0fOFYO5c46344Kq/JKkNJ/KQAdp9Gy6ZwPLbf3MqICr/Mh
pErX5/H3xwszzyDFc3GQoOAsM+4f0KlGCber9/PX72NFWdsZOVZfhqEHXIdKVcfxSGBQfCKq+hO7
ZBB3DoNo2dWxQ7FoYKsgiY+dg6hoI8DIS+1MJ34KP1sS2YkkIWPmaH6AuNtNVTvD6AHnIuZR8Ktu
YjQ/jexz+X1UNrN/YrUvN2CCPTQoN8+sTtdm2kaYZ6cGE8AnFpKADIrlotW+aYDS1Xyl6bp44dbn
IexOg65GnEJiCo7QvB87CLKl9gHakBd4DSwN4G7XAfgyuiCZAfo/rPWVLUfEoDGs1mNTrgQCm1oQ
czXTG8P/Ai6mKJLnP3u5Ah7D01QkxGxM9J5G57cq6O3W4vnUZQAY8a1OTfE59XiJlFRwqjWpGFdy
JMb6YMYa92TKRYfU5msHrme/cpCqPdv5hT0zJHWXknI5qZWC/Vtvu2M1iQzX4IAuk8Qj4/N/6KrG
eR8FPYMKM2vH/aeKSGwjhtzPz2vgWHTVWcjousZD70vtvURYyutVDAnEpi1z/XYEVCQNvt8kBpnZ
lrOk8SnrAdJXnBRvegV8C5EAyytEyzXPh6gbWWji8qSf3syHL0zlAVkz8/VGZC9oR589Ae3t4JXX
4uM+DGnXecPMg7CeFubYytutjKxTgCWWbl+A/PFRWBg1iljPfAXsIbcb09chXmXwkd+0YUYEv3Ir
bWBtJB/D2X3ElYMzzIzGCM8FTc7idlHVnjhYaOa9IA6i2+9RXpatnSZU/XDvLwk4g+1zmfKaGOPj
1ln7ZmKZ1aepF0kPSFMIUJYzRt5cH/2epLWw5UXyGD/gS2wiM4nhz0vIYRlZUMFHbYk6GTfR3nAN
dTrTG6pVch+52waxzke9SIy3yB5QAvXLj02TaH5+5/Fh2llMVffsf6ACF7G8EG8chWlr6yWDZhPh
zGWNWtFa7lpDXSXF1wEFm0j9ci9U/XDBoVZ6TB4BiMNVTQ+kcVlKh5zK02kPQLFWGjjAq5J/ZKZ5
06Jieu39Esi80W6trlhxWOvsHNBRxH4FUCfzw9F0FOo8XCd5SugiCWhw3FcKdKvTgWJdIpYqBEAU
hE4Ea4cLsrVj32fhFzwk89VMzsQ/Kuz4BpHfIlbT/eLrBhLTQ7sFEVyGT9KtbZwnKtEWJZ02y0pw
uHh6FRo8DqXPiNdA5TfT/Fw2GV1r4iWVDjNkJ1IEenFlnWuBHjFldFA0rKFEWNoOCQnFf66tb6MR
FQkD3vEAdizuCp/9feK7ImXcGtrvo4h2n+X+G5x+ZiJi/YeRVMgWKxTYkFFM8Xsdncrk08glRWyH
0+vHFtuYPGlaSqgGcaNmuqtP/sg8qfZeWkw616sJvv3hX5VPIDZILJH3Ye8nuYshY9WM76IzAC2g
aTiyIPRSCtenpn19GcnRgoFbUYJjQ4VFDK9jea2t/greOkBnfm7UQQ22CclwH45GJ5ZYmPYZKJ/5
LYML5OqjdFsYiYUtT5cl0YU9nU8xyjWKj7ROvvId/yQEl/T34YFHNYqr5IvW40eiTh6fQn0qYl3P
YiVJAhFcuZjr6XXGRnr2fmCcXYb0VZEiiOwjwDUn4G0A0er2DhR6HHvLZe0DR5fBGg5eGSY0LY/h
eeGvRKHpGE2M5iPgAF/KxmII8WFuasr+VA+kYgQOiJ3PTasoore67f45KsOuA3Zt7/OJdui99Xbm
mcquS9unIudIY6a4G/j2kAPV/FTbGuNwR9PWifH/aWrJZd6vB6KWwkFQcR5kMe/VJIy9/d2vxUkN
6YfIsb8RdhR6FcRr/bSFA9njlgLrrM8LjXuesUW0trbc3k91Zmfr8FVuusCJqNNOIW3rPZYQnfIH
u9cgiCNfl8mUltV4WbYvjkxYCoyRH2HhUq/P484Jh/LXUgBggpI/LnofmjPba/SIHvv6VpVZbyRp
nXdgyVdePfsC3IU2OHkA5Y9T5lh2hKGKnLyLCdp9mdNdAj+KrUEJ9CAyFEW4lxbgZBWQZIwqCXFN
EIYTd/mZDHHEcUl6nAAsrQKeKkfU56cIMkvRSb0u81HpdYmbkL18pijpo5NrD6Likby8xNW4bs7V
rcnVZYZ/2dgGaok9wZcSnFVBJp/JYGce+IOphn56F4SQ0Ii2Y/SxB2YiaygXkolE1qrUwbFKNaxf
7cpGqfAIwPG1eouK57NIcj/13whKoT341HCWdPuoRmxoONXHVGiFJzao0IGGnUVg8onjzHq2YeIz
QFcUe1nREPcv5TUYKfHv+9e1YWF8Ni0yYk0k5IBVzMZDOKJOYU7mSwAmjwczOuo5ue6kyvHhD1H5
4PSzRF3OnRIaVhXy8Ob7PAhLBT6jX+FthiDDmFNXZ9EpKe228/k8qC3i0fFkNuRnnTxaElMutPtQ
kqxoCBtdn7WjXrvikRSoExkSxsB80DGNft9Vy05vINycPY6RZg+/mF+lLdIiInEycJO9DoJ+EAUB
/QSvGrA/ZvSEYy/rMshvG2f37Ma4w6tHXHZYq/NUf8bml6kNAQK4E4jRpttltUSCacyuURO/Mu6K
pqbX6N4hllrBdq9aE2aGHISTWljHxAiat9gR/oJkJO4i+gOKcQfDY57v1CNYrfCcPzgihSYmwhmw
BHcdrnc98KJdoL/mymEFxIsIzciS/LXlpuAOeLykYCSb1aPifVyzdLwEvF01tFFsrTMzPdo8JdO2
0IZXrUrPSoTaebZVY4FYK3k2+loTmibVPCK4WaKrq/5iNCtAsxxbGthxkl3RX9WnR+OB8+6J+OtQ
o0IIu3yIPe5OnrCOkHZvtCgwJtdM59jf3lUCUZd6CZ+0yJklnU191n7IJr1lyHBFGGxW583IciAc
oZzfF8OsqyNbhEjN3+sJ7GHGryi5ZOBxfiamNmx7weFyXE+lDiHd1aCYZ8dJJwWB1omFwnZ+JBZs
5proqAYe5cvh3cPirZiMmsuLeva+Ld6/EY7mZb0mjk3KMIJp+G3USir5zlpfkMoZMf8knP5I+qtg
ONj0crfCVEKF0ciiE7N4dIzkzQ8fcwMyOo+dP6/4ymw20jn8mDUdwBwa93wjxkz8TMLxc4mNTyGZ
NN12A42nSuKzNicoSBcEfMAhJNoxKhE6hmGzslFIKm23kdUSlc4oGV196fOZWiqRb6I9HX5uC9oy
BrJtlVoLZjnsnzNlGl6LVOFoapOOfBEBao+d5ncUhfJDf1DuEwKa76IfB0SHl20jlhQN0aALK87v
V1nvRcwRi1AxMznHZlkkcr0DVMPE561c8AuKUUjQ2XhElwBXZgzEllFCciMeQuR3TwAiJSsgdmln
JSx0K7qEmTHAe4v2/mvKYq2kQVmBqisJ7pw6pJKaEtSYFQZeJYwqCXfinBdm4j4YGsHP4RtZXFWU
i1E7y+yZuzSuSxzCDNGrONjvwGfoe+r3yZ+lMo2ar/tl9lRxnkCvpG7Hchim3VzNiF5TaQNvAHzC
51H2mw18Fdsba3jX5SHbKejb3toFLflh/yeNGacyT9lrrKkqe9s+o+3p+IIO4H3OnMgllgo+zwP1
l3WEViNB71TIslNF1nsD/GYkWIP3n2agNUUt+ppMdovSgXDR4e62OXGnOywrtR3LHsgYypSa4O25
vxdJUl7F4Y2h8WGrZBV2/D6iONmS3gII4tJ404SCxkVndeCFF8+14B7CDcT6YYNTg8AU3rLawkMI
fooQa0RfvH4R55T/PJ9pFKDWJDJsaVXAtRHp6ASUzsq1gNKeucz/3TdoV43yv8C1FgphYWeuotYs
CiR5XWKxqZmuaGsyFlzEtoyoRSWXbsxeQuujRhPESbwWWEGl15cku49kRNZrhRyYUhaFJ7pjjIMq
qjXpWuAQWOgSgNvGpVUeKdl+RPRErsa6AxTo6WZEHNjHeU0I+7MhTwpX5WsHcNwSEGHqwJE84kgG
vxn6yemtOKAJzo63Eo7WdsnhEVsfwOQBY9BHCeTr6osqP1oNMwLU6q0FomItClv7AX6fioohirNX
X4HWyAAfqp/9rJ1fRyk8/dwMDlZAm2NhxiEU6rP6G/oBPUYxuHB4jfZBurF0pUsnQHMCU4BSs+Ig
5BuDNWPq+Y5r4B/Fz35TaLOFej+azKgtBmHPuYCmtCeoVWUlJcqil0D42Wn3KHbT14udUbHmVzfW
+K7YbGnhyYbtHptj3mFIZ4+mBuzC5JhaxvUZv8rDnpmGgUN05oqur5A4aSYQCU19oz5rOL8+wRPO
RRZ6K271DbD65Qs8CXo0bvR6hib5mhLAE62rvcG2Kc7IQu46N+YfkiqnxPD0n6owb4GyNjXkou00
C6h4j6z4q7wMyHnDnK10843NzmrhLo+Drw40XYGsLY+e4kU0j8ggt5lifkGpInvgBJoYwZys8UvQ
zWuvY5mIA6gkQS6V4d9+gtSStfc+KOtnS93g5dS09+uyhXjJ0PEP2lw6lO9dZW0kXIgFVpK6QoFX
gQOH9ZhRH/DA28jHcpAS8z4fIArgXoj5B3ieQzOOuZVe3gSF1gWP7LrSN+JrwbYDbCkTby+iQ3CS
FxA3Y57NTW/dRCix/IM0cY6vtMxix4oO/yolkGBM5j+M8wTU5ahTiBCZCSonTZ7eBczd/c6gogmU
Yg1CyEFLe7e3MGS19x/4asFmdPcOpl8Q//W9hBScJfWYGZS8TEA338uceMfTu8OmUO22xdeH/F+Y
3Sw3cf4HpxUeTKczmXXt2mID8CJU7/8UfTbZoWZ3CR3YogWbBMIMeFUsv2srrAIqb6zJ3TlyU+qf
cZbT7s+UHPSanyhlv905yym6QimEbpC9Bq8gFTJvbeDjpKNAc+ps65QOducFPl52u6ufqdWsmHRP
U2rJTysJsfCYl2oGM9c+ovckgl7sVIkxwODXEITgb/nqlzVIMtmXWFAsTcHXNTJnvshqns+G3yZ7
CQFhzZgW+jpvtjwu/JLDirLQFGg+No6XnDwag6EX26Fpm3ifIfA/mMpqZKI25WCnkv01pfR8BD09
rDqzBdb6xE4xBoZPg3+bg2s5/eSvpuyueHFz2wRejAR+QzrOk43GTjN89WHXERNQuokZu0wGZ+hQ
BwYKnAAKwgpNQVmkwI0DxrBb9Te5U5RaI2a14XjLQlDodXGLaubK67AXmm9mOWKGF0Cv9woIMSTO
AZu91pbkRoRYoJP/hAAHLfmqcB0qFKUpkxZR5MFnQBeDkuy8KzgkidEu9XjratRnBJFCix7aaGSx
AxJDX3ObocsUZog2vp7H1fxxrAPR1o0zUDq7AFMQ9O+VtyatgFiA30Jx7sPhQiVEhsWS2dugHC/b
v4ORAcGMWJjvVdg2bi5VdkWSFbhEwnTU8fOMbpwsSma65GKAJKuoG64Bc+TNqHOa+wbgQ0MYO6Fl
hd42mlY12NJzXhKfZcZW/KREF1gJU1k3A1jq8PIwLcfq3hfjJwM5P7f+zVLKgBIGW3NivD8UjuOl
BQZj2p1e4LFOe22u8rdX9xaonET8S1tDxMx6cLFfa7e3TQXSNmRi7wlIdefnp8HmPE9rlPNBiNK0
bi7Hxl1rCjK3hTuTILxSwGG1y2tzCYjR0N6Q8nEGJOd8mSpF85TvCXHWJUDPbcsKNEApNtrKFPt4
JaKrFpqd327rRxK07Qy/F89iAycM9OdTpam5n+YZenflPIcJGVUPC8MZnE85wiyET438ueFVb5Cy
xSbUsRLtkPjQkKX5x+rgoppI5+fXURvxOUZMlfj4AVLb0m8SD1SziI2NxoxXOTrRDEDpcmKAE3mr
ltZ5/I6BK5ZxD04vVIS+bfnX8hPOve5VL0YuaZkG0ZrleU3Q3lLtJoc33i/uBvd1XKvBFL44ApfR
j2DEDWPMB7uxZ8JJ5SOyIAX1ogDXVtSegb0TPihGbjVcB+hdxqtOhQ1Ee1NwtcTpY4ylUkdCVyI2
3nssPMvLp3Glqrf9ofC9lIyIJe24iKahGsIR9eTFiT96UrkqR6kWEjL0ESdCR/Dh9Nwj1NHK1TKD
DLhoELvi8QBtf4I34FpPGUuqtkmlfBMYR75qHJUjno+xLWV0PDhnXBj7q3uYwNyjZgjkmInv7vHx
igPdbLXSCWXhIc/AQEH/jYpGmtYKagF1LrPvRpD+GO5OVNycdZ85dbEcoBKX9HphH+tiukyf0qwV
lnPnd8+U+F/01VD8kdhqQuHVMz8Azd8tzHxSZpjXLR3c9Inhg2LCGdvMcuDwkbKKuMUQhLUY9lv2
QGs++oyi9B7oW0Li8GHaG6GcHVCFaG0DNLKg5MoprJqB+n0ps7G72iAtUR8NapYdMArqWMRkUUUS
XJSiFJ2cEfA+8e/5zVHPUc6YPrT05RVASwAe51Lq9Ap9pS3RlFreaSIXcSHOzJtVpwBZfE90qlo4
+PIWfLkPGV17F1Y4HSLulbbIx6fZocrWp+SUXw+fuepNZJppFmwdfMeF3solwCnKuQwwpw4VUExJ
dLPs9qKvRB1/JpxsPIGrF4cQ3/9e/z9z9XkyGGNZBZHRJf2Sx8tz0va8CySBW+gryvXZqehdBZsi
CngW0whICaVXEmJ9ZLmEYhc++0FS06/iUdOGxVfEOqNBWprgMjrG/Wgow38OHNfrVYrRnVwB3MU/
rPMX9A0YiH7iw4/YlhCjoxBD8Y/7JJ2krmlHlQBXGonTiCNOeuHgrjY+e497XupvEcXE0EqTjdFj
qphqBk//SFk66q3yWMkJAo2PGbijpddEwEnNA+odgGoaQr50x8DgB4BYYtH1CyJ/8R74b3J+OePZ
SJerUvzsCMmSYkSJ4J69tgetmJawZsktpPb8BgiJUcs7UcY/3zCN9mfvkgDMsPK3z4vYD2rDUTMg
2fCc5vzUECWVRs6tbO6py4qrjjuJENN8Jh+Mf2DvlpxdpUnfgKwzk6dtZT+qMX3wFf9E3cKjdamq
6Ob4XclIPpmrlxuyRo8fgiCowA9Qxl/FdQUshfNhi9LwgXgwhpBv2OUmmasTe/Bb9UL1OPP08sT1
FWxGFvbz/FhrqRLrF53DQ2CCdVb/OQxRygxmlPsiWdfnqkILPpK2CYKcrQPsBpCw+OvE0N0IUWxU
pmSv+f8Mv73TT66i+BqgihgNEraWSOLxsP53sjMGb6h6+kPSSN4EU1AVrGtC6w2Vlmj+DTaiBSke
hkIq5mi0vh5ec+wmnfwNFMl9U0Vnbe9p6NM5nzAWPX8qNFFdufOu7gDJntP1e+6w24Uy4UEIDHuu
stUKnx61oIZRqStnEUGf7umAd0qpx2hwhE4Lzy6tJaPPvvLC0YVJKPagNl/WI1a7Audpd/rQM1mS
cjQzwf+8CByLyIHnyshiHJjhZXeibMeWdon3EDpNZeHRt5Eab7g/0CLSAY2DUsdH+QoM6oj0Axok
v6qIHtoXHiJjrXaeFzu6NVQMYW9+1SThIqgCA1x69Q7A8CHh2HYwjlYdY6akzRa5E4yqhtF/N91O
cbaq2iZ5MlROb2XaMdSd4gJrgye59ZVGig3uZ9nsa77m1w5Y/eYh2mBx2EfE8OtkvcNJjjebZVFN
fOYS0KdvtF39byB/UwNhNjlJrK0c3wipcVdDPMvRe2BNIWQpJhNdU6NBf6TGDl8VKHC1cqtA3liD
kHYt/TK/WhyV4lW2znBFdjIX5HeO+XYeEdgKDZlzxNq6lIt0+ZKSBF0z6dC6vpVi3flBrNR48pDK
fHw71218hZETTQrfV/R1IIrKhyNvMC33AGon0EogrK/fIEYgWWKxW6boEIiBlgTVchu6a47Yt1zO
aaOckx9m+PS4ByczFeiGmh4UOmSCNby06FIDK+P6LqFeeHSp2SDmhPScpjzAd34GF7USdtY9hoEf
XUB7xo/SamtQSbQtnMXKcnwzmREExl8YXzi1YTC37kBSwJ0ssNo9fo5z2ot8LcIU6LrqhPNpgZkC
D8f7Ro1emv7ZVK63o0RIpncbB5NyaHHPMcb905KQX3y/c/GYthQxZed2BGoQ08HOwPyDw+gw0rLp
IJnNSn1nD2ghAoTfuFWZVGhlhjsjjzkL9RmZJ+6qYWk6CL2zWNoEr/pBSvRW+9J2okZ/vW3S1s6y
wdd/rgCw0Jec8lQsjFWEB7cPQx547x1wvigMmomJSCcfCtii8l6pZQYvJ9M3KQoC8S6NayfMSoDU
asp4Q1/xgxA8EHTImN+NoZnZVESAtnQptisxL+xsWjXQmlPy5z3Mv3XEveC1sfMyvNFKHwrIs5JU
/zSHvjJ8keuFRcB74KzEDAsSqwI868TFrMJ0wjCO5hIp3EROgvGhn8b0owNljFzXcl4WdfndF4oN
bCaZbF8cu6nefFxnLq2IxzW8OMvYq6I/D1sMRgvEXE4R+PFXCjXtcpP2o2qFclbOF/BeOSmE2hbi
Wh7ue87jqPZfpQnjJPRH8EVGVgU4ZfcOid5ZMiD0QcapW2CNG3OoO9VlmkZpoYQBvONjmtRJCRob
JaudTGrOzt90RHFVODLZX1QPR+taieuVfQxXHnbvZhQSC487ZWtgOGtkHmRIa6qfHbhDF7H/ZYEb
l0CM/5y0VCP+WNffkS0sEXmdrYbg9XQMlhVwISSSpnaSpyqmNvY7xKHTpGSrFyxn2Cp8IOaEX7Z0
zUyRTFjeIn5n2ewLun2WPraGvtzcnUoen6ClEkNWw2VjbGm4YI3GbEkMcWl/40qXjVFxRBIlptfl
qVg+bQnwSJ2e7DIklrqHAWMzJek4xxjXDseLwkETUulxxikPtxlBSSMLuSnL6xUSV+PqtW5u4JG2
NLexPIx22/svLAdUhepQklpBkC2lZLOuiiDVRGFioFRQwtBI6LdVZoMCyWckNqci2a7JSBHxckaj
fgE5h7ZxD3K+fAa6H36mMOchyplyanfdzzAgmGG00rU44l0qoU/Pxm3cjjuec1FpE3xS1RbHCgOR
ki3EXIeehNAL2PRhgPxdlACJQLR8rzvQnxcsWX/94VRKYebKg+7vpr7GV+fap9TXDcDSZEHA9ry7
2OPSl0d8WB8impc22xJJpl7DWiVyXtv/ha5OdswHVi3QBoEjEdJFMY3Lz7SY6IqkLMZMXX1F1OIB
qCZzzMcKZd3tOrm8BDK9Nko7ptLaQbPcAafTF2Q1JcFCgGGJkWnnCo9gH3r98F1jV3Hhx0agR7te
+n1F8qxbqR4NK7HmghLT7Z2uP4PEB2Ut6hPbrtJH+PylP8KHnQEeUiZwsKeYC2s3Zpl5l/h0WVgy
hKRYRXBzqVbE0evPgmJF2FUFtHhkPP5tdf0X/kb440cC8z3C2G5Rx1h3NUE53dujRJQVpUMVS3e/
1Vw4bz/XNhCnhgJ9JrppAEfWu/AViSpD8qGqDboIxI13urE9v/fFWwvNVwLXZhw7j9MaoZhPuuZw
cwPMQYo+7Wl2QxEtmcXn0P/T0faSvkRYBNhnODtkdWlhjXf2YfZO7pjRNy4ZJjcqHWjRV8P3CSiT
+qwbsCHKMrGrt7mSOG5J//1IGWkA5ylO3X9RdGpYV+/oX47GWfMLfmfC/o9FnCuhbvPfDw9HW5LJ
RTkBeTmeyOzCyr1PV/iTB/u84CiAZgLra+3+kknLCRiZySc8Nu/gm027H47tyfC4/JnQ1FSdybqy
1Af93GbmwkIN1k1PxwFzCkRFmLt4aYfBn+58XwgltVhf6iWurWQoOw1vkQb1Pbj56xq0wkk14Pti
oPbuXsjlTlDRM7i1LaspC2eAQ7FKiXanoV7dl8m6AIVORp0R9H76mR8jjp9vYntMSxUkYp3A/DHh
0+X6GmX7bpyTkCA9VPzUcIcd53swzlSGaS+9W+u0/Ah+iYyM8gVzO4sQubh1E6ughY1y88RlEJHd
W7x7fmbTvuu4C+NxsYHA/18+rExiAIORXGPh8us/ihu8nuxtT0lyGTnIJyljaeRILx5JcSLTumig
7/pz1igeZTBy17L92M81Rbs8G7gu+pKij+Czkj3qrXBPmSJ8zWBGJw4gkgkqsi8IcIUZPdJ6EFzt
2pJ+BG1l0Ha+TCDN61Jm+x+KTr3BKHMf6aPkwQmfXVIiaaZBgXedZiAftpXz3GmMpRdpxCd0VD0L
f22Wlheg/O2jKvEEwLDHVHzI4B2gmHQNHs6rdfb8BgxTGIoNv6P9zEM59mXc0uJnoPveA6i3n22f
NTk6Rggk4Mgp8gp/XwGSBuGMkDKZIKYJSGYQN4QihQprQCu40OQ1Vz5eVy922Cfwu6MT0XjKefJd
Lg/Tp/f7vycvTmx+QqA3+x6zlnVSYY8z+i4o6tFK0oY0FdhrxqjvgcVeYIKfVysxsytmPb7HgsgQ
043kR92f/9yMESf6NxWqEJmvc3dXc19ik6PcXaJknqKZFUiYadp9IIJkoRbdBtg1E5IddPzSRqYJ
d2HAdmW/xWZPU+rz52zahhm4nZ67M3wYsYdfVV/NTda4p/KN25XzTOuPZuo6Hy1FZEFL5UMT+mX5
lgCtepl/qKFdUnSogAA9tA75M7CoKxazW4CSyN3lJec5skapRTZINMyOcXbkGvaw40GAPKYNpqf3
uZlxvATDXmk82RD47Fx51NLwXsjwhTcyR1EQE70SgAX4Q4IwRWLYsoue7IXwl5g5SI09sMfcNh10
PjzttASyQa8bCQaPnCL+WTwvmYZYyH3sk3PN5twqnB+RUiCix0kvM1UATvNb2uVYXsoM5ROnCUBp
Z8rTDHY3UiHvxONVy9tZpa6knq6MiSoHcZHEGyW9UigXLgrQUZ26fGlYuaKdEljTrr4jZQgiWQEZ
L2tP1iQBIY6sMfhQ0WAQTN85K+ZhLLYzHFQTKbCxfAipaEtACfb4+2/8K/pbIJqjgGAgMgWGtF1O
B64txNm3t1DgkvEPe0BSuAHRdDuA/h1osLTqlxplxZLpAOwApUjyl1DLU0K/6saj/jkCF8ypW+CN
dwtIKvgWRcz8LZgdHgGMWWvy9R8eL2GRq2t5goLAWpHYwLk9uYrO4UVdNmucRC6LeW7u1llSyiES
/ywcNdZ2haDJOFDDreFJvKkFV6tq0hAxpl24stoAxj80iUcLChw1bjEhOXda5p5v+POXMkPlbKmk
TB1jNETWLoyPXuxPd17CiVvH5RwKrwViYE8XYfJB3PLTyJL7DyHwiwpcxQxVCa3a54Gt8Hs67jCn
SFHxq/kiOQ3VYH45ktWpJnn4mKCD+4LEcN5wObLuimQ+cFEgRNDrgwqcyS2KXtdXGOVVDbEhqnsD
1YJyODLQIuvVMOTc33vcX1oIIwA+c3M72YashI3tmtPQCIcMtXZk74Y0RQ6jjbT+DtN1OvWclo3z
s2pdb2/7AgPvj1brRDKFJc3BnPy7Ke0uScTSvdP6O4yumtLJDhWhCHQqueUtuTLiHKielWT9faPF
uBzWBPpCSmK44lqvkz04FbsEptULK+qjMbo53KWKzoP+dxgTZTmla8mCDcj/ENnb9r1LQjhZscn8
84DAZpiB723ltG7wsOxEnmHU8sE8NB32s820a12mYZGiQXzdXAwP6ddFDBlh5TE14ENK9xg3CRDF
ShnF/Cx+ezG9WAsByuSNdURsWpZpTGD9LdWVwiU7SYJwO6VUUbDTRA5zvZ1G9nfpSKX2o0w8WUQf
ei4Np9mHEfDR2sqWx0wTyHMBCRCb+c9QCfKd1UotUeN3AY8kyhc1c1RYInXJUkSD/qbDRa93wMtv
lmEGDDftfrXjgCEFHFmTrkGUZ1JcZg4vUHVDqj6e0xLa0r7tbWwz1bwdoHUwmZ+6nQl4UeX3+fbv
E/+8Q8SOvysPVyVKW2P2kcRkE+xyDfF2lrD4I8HCIK3/9HrfYYoZ+0JgSW6jpsCV7UpsWR96Qv9r
haqmKvhS/bl59m8OPJPKenHLPH7kqDbqE+AQXuRBqijSjr8wqu41B5pIZRy3MkNf1j/MElnSY6S3
lKAiK/FDAaRV3Ya9GD1JTWwKp8TLkpMZ1nacK311ITjBp45GyR9L/vnAlWaUSKA5CXGJnXbIfFZB
pNLpgO1JfIQqXCqxPlAkfrTX3L4tM/X1XK4qhT0sxgw3tnG5PemrnwlClF9foeVq9O3WmDWV1a7z
Nu4VKYJaK7M+K9GjCpcnTOqxq6ixKXL6vfCPwd3sxdj2kzQTScisxD2xDFMlq2Jh7rYtpXHbPt9T
Yvn8VxyhO2GkFCL1zJn/Q96n2GNNfUtwherI92rT5zMgQq/9mFGMKjvnInk++MkxAr37ELStl2xP
xtDuFirkoRb0iJi9eQr5kC9BJ/2INbvakCvHV2IUAoZcxYQaDBArv66Fr6B8bwfBcbfmK2DQAVnZ
z0TKmtHm9IqtL2Tjv6Byj+II6RI5FyMkHgUPcvCi5npteCL1WmIq59oIz0ViIrY/nTu+QX6/upOb
B5aaZctaMIA3/I2ZYhkzQpUOeOD8i2HwPiEV94k/+cHg/EEXd23nyvivzqU615+861kkbCiOZ8e/
eTYGbLI8i2zyYFQ4c5f8KinG96L5aYEl/zdyyikrhLmo/wXoIzy4+dIiKCsi8nXVWjebQpQ76+AQ
LpTQ7/Jku5lmp2qylsdZUppWzyIcp7UsFv/fsDucyfCPP8LtmkpJiX/OsmM1dnGKjtMOn/ffz2WO
WS14QMR1RkV7ymU00PzovbejOmjCAG0qEmrunv9W4m6O6S/u1D/agf3gK0GrtGV+tkLF87s7vRfa
oauqrmr9EBpyacL2XdKBy5Abw+dywE8DdPLo2zHyFd3rXrUccBsFlqKo6wQc5BJBOcutFSIubTlG
HFShy9QX5SZJk8JqVV9VM70442VqJ3PyMA5OWdIzqr0SB5NMyX9ZjIZCdY0UL+naXgLBCzOGl/hj
f9Mr8Dcdct/p53AZXbnEkQpo2rF3mtvr/pX7r7pkP6MUxJRoOPF3b93szF3m2nyH8uHfifsehjJM
o3C0WcerY7VzHwayUNEdSCtGiM9CjivCoD2WyqsDmZUAgSbAU27DlXP8OJ8NC0s0JLpb0z0rSxv1
HrkO1ov51EVCTckcwvVJ2r52xGzl5sQI3AFsA3UBr69mxqQuEe2zPPFp4ysUADKoxDGWvPfBq758
85Cu4WapmP7JxVo15RsQev0UbRXeFPqAOZR2XVbiKrnBxjhS1/RxrbrPXFo8HPtVzsR3dDBln8HD
oa51CjEEuELGqdJHjpi5IO5FzNri3OSoXsksWgzIdmiiTx/8PPrhnRBAS/XGCvK/ydBmWo9Qkmt8
nHrL/50g49fJHZa4pmoUesJmK9odn4/Ub1DP29Mlv206JwQVvEBuVPMVkGD0CkSu9NNqRwOxV3Xt
Mi3OkDyF6kCoXm7mq09tiGgJXjW9RrLpVAxr6VZFz21MJZHEviQ6pf/3FIhZ5Vxui+o2vl7S7KMc
5SLSgxiDs+FcpTzmLRV0OecpNgkRyHg3XAlj7/wJABrzwRg5inbsA1R67130xWaqD8AxGrUSfB3J
rvKit4qiI5KKIAfofdREAgq6e/fcBmjs5KJCbdEWtxFZme9pUJ9B1LpFZfJuFd84K+YE2m+PjS1+
unNLzzAQ/0phigeS595W6VhyM3odSB85KPDn1Jy1nlXMW8g3TnwRh3ACvCuEr+BJrTMUFgic3Wze
q8LUcl5BulNsB+QNjdHzJm7bHWil2cqqMi71o2cXVzWetvPUztPdGepcr30l3ccMb6EMrnlS9Jxn
xpYYOrFN8NruylSHd89zvGoDAQEGAaD/WQqqo5BSVFwCtzTdSdm5KPpGe7lbYzfAKmUfIiwixgAV
+uB6dSrAOflthDc4vNuwldkFci4311r31ColSH74Vm9BeybVLFztcvXwQ5F/Grr9xKjYedsz/TcR
GwkL4VgxAW2XjYttQAYBy7/fiSxI0DVE+d0/zo6LRVx87ffv6HxCIDNQbBLat9LulNGlhDZN5KrM
QT7M6KzQ+t29hDq62D1gtP1TyRqFRoqzmLWsHGWz6slnCFofN///jObQZDYf8VP2N59SNUu8jzwo
27om/aQc9ni4UE0bkI+eOb4gZ1jQ2CXwe0o0VycEtyjBBu3kgZE2A3hbNZHV/vbdafbgcSKfPIEA
GiQZzL8G9j3CpgA7gV9y9zuUFcierrtPlipOlsckggyjXiVQDJOvZYeAd11/V47o1vKiovo9jXNa
pLhNzaG/Av1ypm/5VYZ6sWVwfOqg91dNEoNrr3h5bRe/F7eLjAG9kkcDcWqdb0DrmlSb4MrOyBay
YDG1A6KVoDxiMPw+WB0Ewri27k0JVHor1UXhLOwGtap29c2YwzOvRv5Z3fb6BetWZGcRKG3PCrx/
EbCYaZDWPLlFS4AZG4bAZxmSfVTPuBPWlB7SQSHL9DsesYpw7fC9Ly1i5e1sIyND5FXT8Vgb5Wts
xCnsFimE8f2Ot6xm4rzUP21IP8erIS0gR+0CLIyz37ZjyIZn//m/IGd4qdsyhEJmiCOdc48jGDL+
wEojpaCvc1lDeIwNakC2nguiGVN/3hpiNXH449AwzcO+RKudhHfsNwVOBNBxm1p54xTW44VqgVHm
7DwYsQBbLVtBa5SXlH3vtDdjzhIDu9D+91MyO5BbduRcc/yxS2u/1k1sT+xG/Jx9guCzsfcNwOWW
iAGRx/RDWrlrJfyQMXFy07LQ2JAMCZNYc5aNy0qivZkUIzPt4PsZqmsz7fMTBMGBlTlQYBHT5gvJ
rr9KD/7eVVQg+pfq2gC5JdItZWFl3a4GILZTggQeAmX1UwsKPgXzdNYq7iuKoNZTXvNaceRSy+0L
pqw9SdZwHfFvOU2MxTJRi1cES2oEBt+nakBG2O0jaZbapYwubSHpzwCFInCvSJaFgbd3z67tma7k
Tot99Dmi4zLoXpGyOMdfqFiIXUk86IxlsdNKmkrJkkbpM5etzo5tTUFp9mw2Mq2/YfTTdskJEcVL
RtbkLk1/eVMz/L6pg2P+YTcyd7u8P/qvrX/Xz/uKyDDoN4BI0dTlUOwTh2ABkHQ5gLx7zO7PvwAV
Xhn74NSwdrSxSzsFRqFDzBCUyQVsoKxxXZB87sN/oVu8cjANYZPMc0Qr0APHWWytV/Us382OKODz
jYXkWxRLT4SLk+9yP05cblYPKU7sG3wgnG+wHXKG7IZnxT83d2cQWX18jdquKcfgBYIYqGTbHWn5
/WL7untdGIm3dIFal7c0vkKhxnhaamCDvL2lXvdO/hQHagnnUcaNMcIeP70qTQnyE6mVJzQAjJw8
1RJhyXv7kZfv643LC+wSA9qw9rmpc8beawXzBoSpKrqHT09/IjJngDBwb31GSa6o/aVjoYhl35SX
Rr5VQF9NxNJgB5Uadmija+EL/6jhZqa5icquIQIjOC4Fad0zd/WZh9uNKzpWG46/pN2/XFYb/R62
NXO5jlgDj2zmUGqzxtLzPTARnlKvUeWjCpwRVCSnE1cK2hFWBi7ZNmCjSnrsUTxu/D2bDe8VC7qf
lFJglIrPrAK38mKF3ge1xDo5nnlzUzjxjKP+98k0dZuAU/vHCZ+J5GtLhyuoccz6V1Kfp+RmbL9T
kbsWiMH3k/cuIY09s9rRvoP/nB3X7rlG9TxWkjUnIWqBUUyGXS5LZcHx341+olg0WC8UA2hVGBcV
WpescI2ibXrOcVCfftwpPkVICPgWsY5kkjyNfJ84T18zhHR5mqcAR5WqSaMrj8hpC6IAmq06H2jR
NVGJt3jq4XS+puXNNoMa6Uv65SrVXZ7mURVSvDoDQlO5iYOlH1KHAi/YR91i9nE1Lum+pWGqU9BZ
qLPiiyTkRbhphUxN+JLAuYPjayyCbQCLdzan10UQyjGW2H/IYqEP6DyzVCOqa8YOhDknUSxNx5LP
iSkTIhlcX5c3xkoShK6Z1UgHC8z7DiJRCLX8hHfS2srI0hyyE3VOoaQW5E3zxT+wiBPjGsLeDBz6
j/6Nbr5+R2DBmttWWGwoEkamwDqbQBUbkGChhmntnhhtFCDtlD+UcNeX9SJ/bW4vEkBObC65qvk3
cQtV+mCtvLOXrRQAgT9rk/mq1RRw0GfKvuJPK75/A8+/4hDX4YtxFQh0Tm2YpWlggM8pL21TP//u
MqFmhNzeqaGpxUhq7+2CMrmX4x4iDyNq8AzSSHfiLfdqjcoG2AebbQMaFnxlInk9hv6mL2F457Vt
bMnN3KFBjbnAmpKrkrYqCgCtJV1E4nB2asEqISA0PrF5O39sYl5h1rsi5YRztxMX7QkG2LBG3X5L
AqrNCUSw1feb+mGAHtvkYo1WJ8O0trsMKJeAkeTIBZuMsbVkX52IaXX4ecYL9Mjbys8U/dYRxiU9
iLDlKUsf7k4Di5597L5q7OJYzVs2fXWjGFzJjW8v+X69MGr8R4e8ucUKhxXCMtdYGFUhc3l0IZpr
4RAtE9tMH+CqXeukvXmm38BAKe9oxHKlFrBIUovvtx11zkW5ax7vkzvRMsfEtWyYFfJIX0//IlOY
Ga6XI1N+Ip4z4pgUEU88It2yYTW+hRYcoMS+YN/cQo7omDEZdbl/Qv/FHDU4VbYyX7SGIl6KsD7T
dBGCf6+03580Pa5f2jmnVJZulR11UYX0jyi7bVRjolimyb8BcueexBLRlwlGDbY5Xsep4l5ZS6BW
+JQvYR1gohqCUdtmY1n+1Lfjw4Ooov5/XUnN06qIvLJPYqRTq2rDLmJN/J7nETKBLlIp7sNjwt5i
HeK3+6FoAPi7qEDJvWs1mZpRY1Ki+g5Ux17WQhrQeBBIIP5wsE3faZKyswwJ8QhwFYQHi1TAp4RF
4Rty0KN79hfL71l8zF6k/EWE8J0kPj/8lc9U+s9JF8FTNBcBgCEkavprK0iZV8goZvtW8EDpiLWQ
8JkgpwmHvhk54MvxNFbFMUd7mZOhvrFYXLqJpoI1R73CBOp/TzBMpIqTxYo+uqXcQpuiTLTywoXv
vN7fMN4pbJQ+9sOrmiS9XM9RkZdXN6ffCKk6KlKPY17d8OhGMphoensRFUtcOwRx2uNaWUNq8cd1
1CDk202o4meAC/9lNXoGDENISk+kppTPPKksKbSu9PMcT+qXfFO7F4HTy5coPH8XFsbhoH0009Gs
iGSESIzglBoz7BwGkCyPggJr+P4Z2cPCbj+uttlreeE/p5646nQkWYeKV5IyH19GW00p9NXIBlYp
dhiB+JMJgiy7Y3PNrk/XPXCOFQuLxFuqOtAtyVoRKnE+FWUrSdeU8eDtQdLYj7jz0eJtbB/REEPd
EApzEd/hReiShrLgc3au/xwvIoM8VbW5h0zWrl1HIPM18q+ojN71Z3ppLBYFEyNewVh867u6aZSp
u1YLdHitqgaMIoby8I5nz0xQ3dUoDVktCU6oX7DTEXOXA0Y6UuHhSfIRGfrRwz6HPi2r+Ja64wHL
rWSC0dzCboOlszTFVxdOlqL5DwppJ504IYsEOCby28sdhxpyPKVDN8KsEF/aIK766tvBODkWqzw/
TygmSqYBoLQ/I5oXjS8tpDaqsF9pcanmSLHsJFhWh+NtNprAJJx1/IIM+5VS3ybe3yr6/UpxBauZ
zphhRjkFenw8JzVkG2+sjSk8I+o2F4g+V7wlUTIbubMZtA9t3V4zs4IqnCh0vpf37cPRup9HaGoa
hZ8GbHyXwR1LlhvwKP2GXPDJsi9P+FjauijC/fsLjWdmfgzAIDKeoHzJYwqH1TOvxUf3JwlhCrFT
nLGzUBDjZPckaufL0CMz5uFoL9zaTe32MWheZRc3BAPOYV13tPMljC5+Ufq4pBhsyKvoKQ/zg0er
2WBQEDr4dHYvyrx3yb8lqudv6n3IhWPZcsPVGyGnCPDrRseP+riD3hUGiVBfgVeSpSTouAfoO8bg
eZ5w4JGACGWJLtVRIa75Hi+3NEGBQqohcNRJSXEz8/7nz+hzR/HzA/YTtekjr7je/rZKFjM/BVxq
jjyEIRhn23Ht9ezycb35nqUMgIlRz1foRwooed6c/81tgLfQR+5+Hux5xmVZc8ysPUY9VnJ9tUGi
rmSm2SIZXIaU6w0nrDQvMkcacGGgflQe+Nq7ac8LS/ICbllrNQ7PmcNPfrcjKNQ7kLF5csavt2aL
QPy4XXMs+8YZzGLMJIawYHr9bcL9gEF+BjPIrWTBAH/LlWXZbJl+D2W949I1lmHWMFQElgP4IjRr
rs+T4qMna69+fuyZG3QlDvDZKqdTdj5WuMShyK5l9FuDqUtlU6pD3dpOlYywx/DmVprthMugVqGV
mkkZGVbj6FPn31C6l7xuz48aAgfRwJswMiEEMC8lCK7rxRe+dGqH7qExSPdOhl86fadtCibPDLgb
kVF2JSClvyGgWhqgNnfyTKKo579+gqw7xiYhA2Hr6ojYGabOG1MGFAS93zAsbrQ7fjWxCLTfiOX+
1o0rtzWn9K/RJi1Kh7AE9b29iREc4Ms+aEheneUvmh6GmMPbTSBPg+f2ul9Hs92bhD33YQzYmOml
9HYJaHvNhfl4zzjFHmvC8eDEFg3mLrCoiP0d5AJE+nM1BIuPv5d6yeKEZkm9wmfpOT5wRk6e0kun
FSybyoolcujT70SPGXvJfJ5eLikQ/emXOb89dZhPZLWOCTzXC4qBLEKKSnVL5q/EzO+ek7IOBop9
jY79pyxuWo5nsnisrUjohPZvH4vzvrvyCRxfTibJYXt+B6pY66uQpaVB5jlA2bTgJK1pkYJWqeHA
EP48afODevY5mhf1tyvRwOrn9fEFJ+VrXpREupY2X8KCDtcZqcT9X5uolp4K1XclWhkw1vIsgp3a
7Igsz97XQ+6RKTKeCwV6+1GTNn2VK7lUxchHXMlyZsxqvVhCjk32+hU2aaKq1Y1RIrnNCsttzGsL
ude7o6yGb61HUG/vd8LX6/yNRDJOFIOccYSZ35scqUmhODwakoDlTvVD8UbDEH06q32stgoWLlna
hiF2V5g8Kmf1PQn2Mem6xVcP1u3S+Ma3rYXfGXAvF5PCAbYZY+jULn4LtPQNFjDBUAhw5X95eqGl
Pjx2ygbqNfNwghCA4vjv/p5ByyKF8tKmTmd4AvvyTu1gjO/8JPjC3VBvkpFE7YxViv0siSOA2OS6
deUe7Y8a6DIvmu/IgciM1WGOtJq/DJWcRHlSkPwn09JeVerdm9E17p7JNIX/arsBQCVSY2+AJkUN
wc4qixOb9+ZswT8q9/Y7BLp3Pz2pXoo1Hro5CJ+Zb14q6lgBOdNVKliAjf6f/WY+pi0RfUyzUuzC
CuZSVckjr1nElBmy1AH/tWvF0DOsgFJz8kWiW+71UYiloT2gIq1mgaToQN2et2kcK/aERE3Tzr7O
0oYWpfZkv4XnmGczy0XEAliuSWlXIilChanbbAq//q5wThivtEgq630XlgBLZl9r23yGd/T9ZFUX
q4lB0RzI76EXWrQZErIIscp+X/UgC+ksq0jPx3Al85yvQwiWNa4S4Muw82daGQld2jMBR1enCDat
V7/N8lToJDSM3rLs5Kd5Ci6dw7+B+iLZIcAT32olLwHP+gi/GBQi0fzlMGbZXKKZIj7TYv007ORN
tHj5mbBjdnOmFQ79YNYaYFqZTjR0L9OrE2X3wpBGJ3ljwZ8ojmNV6BqTh17EJZJZWFHzrh5+zURr
a0eSKUC9oz7cdLudsCCCHnEiDFEt5QvOcGwTgqUtcFG7etJ1Lj2FE+iaaMdhLkgNYg4xsaci2Dml
BCuZfJG6RF9O8DFFmPlJXlwaEKtgWjjvEtFSsM44E4T/+qoebzC5cCOdRrZd3Yle+hW1gdK2Ew5B
SUG6767UVSBL0ZCXIoHh1/+LatuqoV68hPAjNtf/sbuSE/Mft5wiIaapi5OyugpMbDW06JG4KwcO
dSyglQlixFWDTCvUqjDj+UvA9OxyMrSoxKez3vQ/XHExyorTFGNZaAcFq0q5ixW9Wfs2sy347gqU
FbkgSfaY0WyymG5IGiFxYBMVPZQLeaFhpabhJDCVoLFsmF5N/OCbzM4MF+gpeL4xvyTvxglNbtrF
rhC013Gz/vEPDYWbEtMtKpvuRo0vXqrmvQ9ftmb3SBfuGkCi34GYk1Dp2tsPD+UJfqvE0EZ2o1Z4
jWSLQw4nl6kNiHa3vfeNQ/qw5V0/VuRagHoz/VXdwXJGBpUKOrNsvx3d4mHlFU3iqHIR5mIyfEeR
E0rWB6mbi3qBbbmu8dgvfAwBKemsQ/Ofy00dETVzBU0uTlzRZQU6BQIrqjGa8gHWZb8XwAvwqlSW
qZPXzFNW2C+KMrKIhAVdM+k9UV/oYOOBgDDASpSK4t68t7CqA9QyfaPiTjlyApQvsIRF6kz8HI6S
QHt3RFZMg4KXkOBOX/2jByUkryb5Q+yQwT6Py4EtltEbgE2H7JAIA/Q6/vMenwbPzjvg1FQSvTzF
9TqCTCXjc7cBzy12SGs6BHZWTnlEYiMz886vr8YaE8WUaviXSLeUqHzdPInYEUHxIp6ajwbnD3Vz
tZQWQTInp1FRx+KDudEXgkOhltlcR4BGauhTzxdUSqfhbGkdNsU8QCi/gG0j/PO6o7FDv1fHo9/1
eyUV6Q7Fka2NH2vyJ7RpF4Ti8hIXuuunvg7YsNNPh7FYhJKEvtIgfrOJQu06BF6UsGJKzND/IQOk
FS9JHLL52nasag2RIASUDmZ61ORcFH8f1Q9M5joKhHscPfI76YQiJJMHMW8mrFK/sNL3j2pq2Z1G
6rK1SmhsXQZCIYAyUfy5UZDORJKQMRIVrZfIo1TgTDJvyXm4a9ra1NMNNUSTMmWDcxODiPWFj3zr
mcZLxRK//FdR9/Nu48jRljxTNu11Uiy68gAWKXgzkhVge1Z2GVKwnMBGu4oLp60Ts7U+tNhEZssH
kkza81w4lJ09N8NdNhFKfuiyvhzCP/qGOtjuYDGs9Bfe4ADeJEg8JPrKusDLhhW3iXhwcQV5YfU9
/27Mzo5sjYyIHr9SzqO4pSlJEihdGqSSLGaoUOxDXtdQOjw/8e1DPn/y+6yX+V3rZ72qa/L49K4J
WfBaueUqE2f2m1MLr0cJIWIUgnd2j/z9amEGxXl6GIa674LE4TfGH8tnAEylEYyLhxB8V5mQCt7r
Sfrj9KlnVLMIZn2yhsfRWdcSQRULXBRr7fJt8THtF1sBieDX3bBzrHpTzpzmrHQxidRL0hT1VAJe
FlBBedQnQK5BCI5vjZDTx44yqLTo6r5XabtKX7tRVBnKXRlYYIAzaqLkNfRWy5jJ8NVROpPmQBap
f1k0MGLFeBt8XZz1eUJJ+Kq/NMws0jbey3y8Nn8UvxU8hl6PWyt3mtrNra62bDxOgHibLjd4a5ir
DhuG0KpQbvMcH9dknbeIEerhk9NCC0wHGPbz0/W3vBeTLSGVvwABYHAatXRshxtCMI9U0vhRmVOv
ffBj9BfXQU82tJtVhkJMFgg263+wbm+w1ecq9WBa52iOzlkNgFvVNMB1q593tVHMowhXi9yerHn7
1VZwP79+g7EB08FHHYOoqCb54Fc5noaJxZWgXexfKP2p+0SF1gaBYmXd1w5dC44WmGHZzNXxsOKO
RmCZSJeER1+1w6KlvLcclUcvVsq1psTynckJsJh0qJ+iJEfAY22emI6H3O2XylwU34qwWhbo3M0r
Hn7+7LI6OCme8E2vLV0OKhtw8dnVjno7YNc1MRQ+tTv5jtso7y43ais8/bfrHhOcDI8ssYYmPlyp
CBPcboMclVhuokch8pbVQl/+LIGV74JvNgTQeo+Yfe72erjZIT1LYqHmeY6ksXnEdKXN5Ir0HIBB
N7bnFavRijLrrMjLJrpRsw7uTYN9JCSU21wQzwg/cUY4sl6wbNrBvVnZbOLkM33L2DLmdP74vxY2
RBuCsF8jHV+0FNAVUUuFDDDKJeGWhcIWJB4UeDRSjvr4fczu7Rs9aYs1HbiY1E8q4SEwsCI7XEbp
Hb0ZtMtfbznCP2DuwFqLAYwQv2775ye0+XqI3o9HV1svA2hpXtBT5M/lfNWDsV2jna9amUbvNSm0
u8MsjwUm2DOTi+dPN1h6N8yqdI3LEjz7I4/dmgr5CP+8bmr9WMZPZXuo07Ci2tVLHwPUeY+LSMzN
+yxMnNQl7HN/UOit3TUbI7X6F1VmAE6imqzrM9EOfnz/I+TWYYZjjGoMVgm/JCKkb6vV7Pq5AWOz
sqiCmKYLyYMuZdwUvsvFB3xyzgPRobbKQXrEid9EFbVO1NSBKZlLKd+1otm4joEGo7M1KHnn/H+h
y+yjI4OyOAbeHmFfyDIjPfdApFoKWElVil7WFoim3WIUniIKFIGBV1C+UhS8D41A4qBWievPdnc4
ldr1MiCvBVMZokvkIWoEIOCX0T+u59qQdraN1FZz4UbdIgQPOMZnTI9BXZBnVV4jOXZANcPhCFun
ycv7QTOilbx/0L/Ca1hhzxh2trtX0mX8H985MMAfAsNTNjxIHmXICztxVu9FmyQazoFPPp9ATthE
gGG5/O1MoGeiGffCVYHdGaNMEy3OOyZnE09AB8XRws4KjaG33RPgXkFZrov5VEAFuhSnIYOndAls
rhZAcuS3K52XVI7h0PIvbavy+1Muhjm9SsSOWsX04xoH/w/pn8jbDKDWwcNMw/7fCHuagBZSMFan
rZgN0C+QKFtlFX7Ejo69K0KZC5YpUAQEbJQfosgkmUWPoPnZk5ca3+0NuEijBmiEk0FYNgwy5HDf
2x3Zc9xgQ3tBBvp4TO7w04pInVIQjxbYl6YLV9Kln0tWwwAaF7H2Wb8OFq0GNDwP63z51qgyifVx
J9/DA7oSOu1X77IJh8ZvdzxsLcOcB1rOJZscR+platetWHOXFOhi70PPXC9sREDeNB7znLi80U07
OXI3GxMV3LfbIf9GKBe3Aus3wrA5CT7CM/VIHnE6AwoeOFNQdkjV+yq+qRD6bluZWqXfcphuKU9Y
Yh78SWW1I8dnQ/mY9NOkQZRYZQqUibiIVkWZFf1tzpmG//BP/tP9d6nSv4UyS0hc7U3ZZ1W9Dj6k
ER3scXdYWLKC67zykhKO08Gf5jJYhSsk0jehTosJtYduciyR/MpDBIZRVI1NSxgCc+R4XvE3Ih4i
TLc5RNCTuVRlHtuKpmkFR8VjHNXxkrG42E8PRUgAZxyS6d6LMRVg0Y+wzH1rb8/LnSnvgs1jKAop
kNg8X+nKGZeuYSa+1qf8trjoOOrzwVue0+DrSfLeXKszQHNOQ/S+/Ggb2fADVYyKdhfyoIpWuT3P
YbcCOqb9wsVLK6a695H85CWnOWVDXsEvS80eN6yDMhdV3+d1PVGbcWKD3CKjP7305kje+4jjaWeQ
S5nfNt3SJuCa4hQZLLnTAqM8gQjP5WamLdH202mbBeBoVRXhbZGF1iYc9LUanGMZeWvIxnHj39yt
k+jhhaNYyKWbAK6vdC6bHZ/a4VLlb0eT48YmERzfu8VmC4MeS+ThoRA/W9lYPe0F7rG/w0l8yx8H
HAuvQrbbZZzQ48mPK0Rvmh1QUnSDaHHMS53iYWbAPODCmPWfofIJEUus59CgvNJ0MEbJifZZjmSY
XKw28BN8YA977ex3IUrqPP4ZBCSDhdLIJqYKjOeJuaQTKDIk8hU/BBxFZ7bFBrohbJvghiwsnseJ
z23+5pReEOHGMukwn2GMh7roE7AqlE9LoSn/GNDus/bsC03+zx8m/4FGSshC5VPMDor8pgW7NNK/
Ps1ur+VkNgzoztwEfzPD1mkIgkWnbnXG9rWSD88HDHOqZmAdZuTzpVtQCretjdF/0Klk5yHkP3pH
Z5p13J41e8kjeY8zYdceChHkn9tMWSjsGqbU2jFHfij/4iMul86RTCcc2WEJN84m5zT5i6Q9AuuA
J0/0nPmeXMNC18BseNhLt8TWbUCtwa0sHSMXwgXcxh4G22zRWQg4uQDamAUEQueD6tuvuJgj5gc6
e9oOwclEVBEMe93+hgb0GE4dFic4XHMe5/h4ihAUA/5zyZjd+zFuLa48IcwBXEIQqiTqef8cMnnw
S7YbKJ8m0vWZPLKR7mcGbQpWGDS30fikLcTm+2r5txV4clgQ0OqNHCyFpar3sUVRuG5VEeg+IWE/
SAy3ifAzvmN1vKg7NACa97TnzRHjWG2Adr/TJ4w/BnI8n7LGUpR12DVg8zD39hn8LyUV3wCi9Ano
6RPDBK5zfYKy8GKKLro/ZdwA+t4ElOTs+x/GZJaP/dWKWMNyDKDUCXnKbCibVa8BRyKs6aNp0cWo
9NMy+8DvuLBryo4b7NhUKAfVVbstDRgddA7OUq+fdUNXKOMh+NLibJAeyhkYCEdNlzebCeHUHn8R
kzyO56y8s8lZKy47c8rijcbmCvZlTbrGcoqT0p8JB7b6TIGQ5Q7Ibz1WKnRnXn87qPy03oeS8qhZ
6Bx21hr+acDxb6PpbcxXM1BI15o4XNd5g06gljXrknppSooSqxyP84EeyTSbrZNrlvuSdeVMTxBz
9V9PxwYH2rzFCn7OoAQcTcWJb1w8SyD/QoH0FeBidDLoaIj41v/h236ajxtfDyV4o3wRO5W9sLFo
yVFtlpl7RqppWTqtfNUoiKEfp4EolhhrLqMHkz0jWtAimWzFDW/UszvYtkexXMDLrVFcF+QMpAWL
NZJxF+hjcKXWfPEMu8vSefSmGANGiVsPSqAy16zvsggJlos8QkSJaUu8Q6inMY8GRkEiI0oFxGdY
04u3qHiJTEEfkkbF8HPvWAG12uHb7q24Xa+/HKrnoT3PWpYMNzn+uFVlTaOjzBQzDILWscuLwQLS
2Qw5TtvUPejnYCbYB41VA/f9ixwMfWkc8j/eCeMCMbJVKQ6j1A4NFrrtJ+1vtaqjsr39C+VlhWvq
048BM8vkTyczXgnpQ/CgkUV1cGFXxiYLh/5wUMxHjMR8UsPCzp0cs9vnIEvYvTcDjeKkXBMV3uqH
fRsSy0ABywWqeVcvzZWPyeCHwCERjFkJSMKJAPyWyoFNBwrUJuSPQGXB1QQjb75m9b1wH8t9MGa/
W09X+zNtv2pE3FmV1rJej4PQQDO52ElMarea4xo5RBGFNpdeppkL0mhWSXVN2D/aCh3pN0b+eAxO
OyF28l4z9AK8UYPf6v52+nCJknLdHVqm3Led3VAWnW46+Hk/xkx83Y0vtKwWlKsLvQgicPRziyqI
CqrpDqydV7aJUD0AxBqdHvlNPyif8l6rinKbXsGprBUeAZpHN+xmoR93vpYTE2M+fUvvKgzCfBiF
MHUwfHF2DCURMy1I54L83c9cOFg/FYMB3tGDja9eKr5Nv95QFuKSl0nw0duJDzTBN7RRbd+B6IVF
OoaW4mIWzGMUY+p6NkLJXmTS2qCl4t+8lZOeXQbYwaoohjxd6Cq9VPuryck08ey+UQ4fxy8l0M9j
dy7ZhoS7SoB0tdGSrYISbvs0Itor9/nLVUrYpe/03SXroB3MH6YoGvaz0RbUs2geWZTWYKB0H3oi
xgyisOw7ugZBRfTApRitu2DtXGJN2zoSxsZ71JHsAYmHs6lODG9fOrlZ6fYclPi98EeLrMcX+17Z
t80ehvgH5mbPTEOhRzUNnyToXvTL64/OIujPtHny/wZsv3IHc+mx8AuxHNyR15cIV2JOe3FJ0An4
L5l+SiNlTIl740dkGA/XFIKzfa9gtq/TQNAbPhnvlRax5NoDOmb8hvNhHnSGnPfiIpQ8F00NlAAl
WBOquz3rPCMfuXAp331Lz8SLA40kA7+TG64KDHE80IxSLzor0kduCwk6wowoX1QCNFLT7nQtFPls
PCU6SGnoqQxdqGOmFsCClJOKBixqug1lCxd43XKpfgWkf0heHZsyotPJfOCY2Qajul/SvRfMIGsk
NawOKP7zWag+u0Nkupjz8oZNq2/uWfXKl1IlrRNzgVkyuHm8WRWRmYTfOkb2gH96BnOrKeZ9Lzhf
/xBdpFf2cgamFz1PpfIYgJzaap3sUr896OKTN9hLeQun+qaQVc1Hsl/+EVpDhWC1NtUMFdPIph++
bnRZd91pzMQAgbpvU0fXw/xVYWQvNYfomUfEHZ/d23/Dl+HCkkDhXN5tler22TTyC9W2Yw/49ZKb
5wUFH5X0DHUMD2o3tFhwQ/ISNvRIfTeImaurB/8SxTpZe+8Y/UjvLjRc4Cy3YkV33AgzLGfxO6DM
WOawL7MiQa+WcAloiuFzFvhFWtwVbRIXhTEsjUHiHhknkSrZoeY3yW2iLbmhTMPyYQC4dReqWGU6
3mlvXPQDL9s+iuEwPxfCA9bQ6ZMZoitMOwiHGYxIxfrhLwsE4JJNk1RuhlfS8SKb9r0nwLiQhKNc
AqlCekEZ63LCs2IgkcLKdyIlcZatR6c3JEcmcG6jnBGHOgJDuiPAQE4UolfjL1Tb7D1BboiWhF7n
WCcVG/IQ1nBvqQjaMTxQTNUvSwcSbpQ9AtTktG2B4LqCA77/cEVJ09hAot2tnieiRahIgcreC7pv
XC9P80XxGLAIfmAiRN/trqIUvq5FUNjy44CtHF6Q7R1UFMoeLU358oK/1NpW21d2t67S1lE8e/DE
D/lCtQMc7xpH9cYX0Mxv4DUdbhmakbQYFdWZzdBQld6WXt38TmwKxdNOy1yaG4vAMnljIUjmq1z2
wywV/st4LJnw3Mkp3LLj+e3bz5tZX+Gum8X0T4cZywA7+YG7LCdq4BYtbFs9Y98xKlgcaclFtFGI
rKIX621NWRwdUwwskaeNwIMPrxoIiVUeSQaa2+mohtaGElT9OQKsTY8uQkcCDF6Hss4Iv8enlQbq
DM0gkjQ34fz6oQTGUOsVW3pT8q8tWgarLmyKBGZmYTrwYqU3rJRh9JysHzSG6I5Nwo8L2UIBSO4p
D06TlbXLS9HSf4DBGe/hqbfeBEkeEkVXj9wSKnDQ9frMAH0bRiVJS/IUA7JpbDDCvblGwN8ogyvZ
6ZmHTFehNBmLITDEuZWWLeooiTZf+NTO/veY6ziNYXNKB16oFmZPZ02Xbe0PGzeOUtHcXNpRf+sD
nesuS6t1TP9EG4+iakZoD/w+amBXC87JRhFS9GpfEkuWjjJhbZTHqnRACl3zwiDrN3LbhmmQYxwK
FlamRuE8K6JJz0JddFbP2mLaFC9PXjcqmOy82BCeC4ji8mxyaKk6H8UinVEwtdsMjcdWjQCKG5x0
0zejrTRJbocjIjYyAO8Z9uRbdbNQpvEopSCE8XYauUH76DTMTLmEkBEu4FHhVYRed7jjpDpUITuQ
1N/EnIDgssRZz0mmwESH/E7fF1GMGGshbD/K0okmuk88wlFqjNUdWwWPyBQIqoh+MYCrPLrFwM37
PYO8EYnFCFDemvw4nP+oO23OyXVTjd/kiOHpPahpI0GBBLC4Z3Lm28Fv7kbvpcu75/4bxKqTbLvu
sWjY/7gP1NO+pfJrSljxpZCZEu/xtCo/Nt8/IjTA3CsCmjAChEMY9uN3bDhFe6pbcbn2BC/rqxl4
ig6/oVv8C8RTRZohCFc/yM6JqFFkBc7pNAXJfyslDB4d1ynPIFQWzBeS6L8jOPaZbHTIjqQwZnQp
BWIxyRVXdl/JfcFQzhCh6XZszPRG/o53nh2h900ZXsfqkWC9wxhnUXJAGk3VGsS0nINrt384Qdw7
ZiobKfhjJuCYeza5OYw9n809Wn+NgVRGlsc4DMwWdCLj1X12lqcPlWcPMFENCZEo4G/eWjQMCED3
6PpfJO+PJhpeNcMwkEOOjYg0wdIfzl1d9jndoHRU1BP/R2mtlnqltBxGqLsdv5TRKRI40twl5AWQ
1jEz/lG6J7H8v35T8+pJd7lRiaUJUpigwQ3FCelIcvLyLl8P+x2TLtGWrzlOJyGQFObC0RnhbGoG
Gkg7G74crThUU3TZ9Sn9hjGmSn1ZbzNpT9xrHs85p4XQRry/JlahcK0s9zNl1JFJyHY0//YtVIhc
WOscoF2+oHkJaH5MqDmhaCI5/8OPN6F8iSZk65/a3gy1XV3feWgHHy/ZXVkXS5+pUbeNDuU9sffa
b5oKaaYNWY3ftTGmOSOYltdH5bOqb9zWHO0L/LBSwn9CJvAcP1iwqKQ6Q2d/RxBpy+dhTr0yk42S
FEXMgJp9SiV0Q1986yuLQrRPVoNOpojY5+cR4j+w/AKIX5gBAKAY12XSsW/zc9bdqNKAzjzG8aTT
+kAr5nFtcsZAukA9F7bQBJyiX+HRzC/jXQGX+TAF8axEqgUJb2fk5Ohcxm1WIdmnqd6JugyeNbbE
ZAAORStQkw7WlwuZeyPnNemi5TrlhwD5dl49KOsHEdDR7tVmkM5jz4xvpMkpmwPaBIjuBO9qMQoU
eEqIYvzwCciknnxsBt9lOn/GAyLuTn1n0Q36qxflGrVOlbp+CE8mhsvfVfoMySCfRn/iU4gdt7Rt
rxJLvmyED8ucD2W5Tg1w+DMe8s6u7ggf9L54Vpxmvy+2+9nTFY6cR2sfCJGejlBqwGtJlMLXr2P8
JXE6w8u9aKXAAclYxrQhauOTql0jMcQ26lUazd8Node8kvVElSs08N91KIKMKqsnFkUUzfgcjV8q
CDDvsLV6qkaznMSDbRlXuXzXFuYAzUSTi+cjsrKTEHukvW+HV5yi14/SbXlhmtevUDYYeICSZe6U
4OwHcAtd6xn9pg5FAznDENWOs+NJwV5N2owxEtu6uNJYKOViypJNPOYEBlyeyEJTuwLzgCIk1t/A
caL4dCUttghokFhlu7NKvUtFVMLmgZF2h0CDIIANCRM/pb6fUZds7lYoBXvEaK0nS6uK1dN5hwYk
YvxftwL3aZf/NhmBpnczw2FpRWGrWTkTi7wWlDbmZDFzf4zM5VU8Ely7y6qmGfsTHrzoBNIAxecE
nWUXtIFXgMVRTHQxOHt3Se55Zlahw/66Eu8UaCzljMXGSsvrI7vRGZeAmOdsr7uurYgjb9yqR0w0
8YX2ONk1gP28y7CQKcVwWKw40OttT6YOjs61MDk3l5ac1u39ej7iOHGMnHV2K5iI/bd8TPJoERJr
4wyjrS21bKdYcFrt9YJdOzIFi0pqKwc7aDPbwwu3JE6Imzd4Gs2DQduRB4W8LWDzVxQWwy7EqZ1l
OzXYLOSF45NkvDY14JT2WyJ7vnSx2HW5rfLjB7ye37wPtcqXy0nVYrkgRIWF+1qiX0KdKmajrpv4
poLC1ctvl8D5574SckeR7jWQg1XQQOKxanOf6wH54SQIUfFI1JxnTsxLNhGT7E6tkAnjwoJ/1/4U
ij+UCkMIIkFihP5+N8RvPji7dZHOUYrKXWFbXssdv2NGpEtBWZlYbg5CepxqPLgAbyVNRmNa/miP
I3oMwKzWQqiMs8JLkh3n38Id86sir2yaPQ2JucmYcQ5iWoS124JiKnGtKG9vKoP4UvTr1C/hqtKo
ViLvfXb9n2QZM4yZBoSvQOIt5HefGveSbS+MhwklYgH4g82MKDBgdZjgK4+DJQW+KTak/sVQX7nO
R5/BRhVDHL6OVOHPgUNFBfV+LxXm8/tPP5AtbsDdZCUBRzDra6yneE7m4mG9IfRWa+SeRUabGf7X
X6PBlHTKR5ms7kbXQFj/E6GaI6nTHS+8iCPwtdesxNm0c4+5vm/49sGpt3KrQvvkZF7hlKcOIWJf
OVQZrDrX+hhkINJjpxve6nu/HGqU5DH63k2uy4rX5iO412M4e7L5sEDoG9nFsio42wwtl9tS81PQ
H32tOAZxGep549UIHm+iLtJRvAWiPD78zrFn+VIYUszZSqEWlghPNjamtKzkFIb6iGoDqiH1lJAC
ihYP7jIFCvPckNZlfK2IhmgYmuCnrcw3NtBKubffulzSIthv5YIKpZPOdlSRwZF3ncVfUDSVaepT
J0oSGeHM8It6a48CxRqkwdnsqADsgCXBL7uw9lmABwqrWt6Vxc60pYYTOor2cFdG5VkuiuMrkFU8
+VtUdtEpwgCiDyzkLlLBCG3B9HUYORQKVq8NK1wkPfOMItAZdWte/mJTSELESXB3eFhJ+NURLzzR
7+0cAasw5O4eEZdpaJDM+2fjF9H7UAgkGzGE6fxNcIHZLf36BrxdFyMgqwX8AwlhByKHoef8QzaR
5Lkw6GYHk5/bGnV0PeYrbu/HIPXbf+vcxtlmVTLfCbRgyv53B5aGphSk9jpyGtS9o85sPWfI/gV8
Y1pxyrfe3xkP45NI6FDnKaStm4m6j9va6DYfc+sqLeblPyUKsDpuNngjHcRr6AHyWJywK4LorKD2
N9tZnebKPpph51rED372nZAKvsog1s9jMjiBpRIEJMQxBy1fFznwuN9eiEjzXLnvND990tmFYbgp
mtzNshCskPu9o6EacyaDk8MzKXoHlGpGSb1yKP9vkMN04gPJcO4hQGIWatWt9aN5sWrlS87q4AqJ
rTIL7anKy/87kCLT6z7B2Lul3JUoSh3OxAXzcrSntv6IKHeQBVCIG25DUFGtQotRNtlY2Uq1KWUr
voxLMf7oSGh3RI9c6Wl75WetsiVxAV0AM75mbovzDAiHSPmqwU5lBAo6tsdvAgR7eZ3xJ0oCixRV
FCljoY1Skrkph6NISEy2F+QqwB1+4hbbApyoaKiwVVZ1MdLb/t5abSHpzOikKwMVKeDFKLYs7a1J
+Ty9RmOwrZ9siQj/D2klC8Uv2VAslt7udcQjcIOMZ8n4yV7uCqoPyjg6Uji8tbHWpn/L6lEsmQ1E
W6G041xiG/KTsnk8rD/13mlZnJi1aJDYNYG9IfiDK9uUMjaO24PIlyE9UpDV9jqNGY3evY0cxviV
QX76ZSQBCEQNfdJ6R0l0EtaxfIT4l4ijy7jGts5n2K94ywW2t7y5+3jF2aOuSnxpH6VDd4q+VcgC
Dqm57zh1M3AllvxItt6APktX1nzsQTSxGRpWMLhY0EXq/SN2Zfjfj7rHhvtjZ3wdRFiQnqIK7JhF
Z98sjbMK9iylB9exR4TuSCtMElWDbw2s126B/lZqrcMHETUIi6kZptvnFpbAsP8PRnh+tIaTKAK0
Pyiel8M/dE9Pe1HrHqNMtcZyeS9V/8Lhyw9bmT6xGqxTrqeTym6ZILJ2aETQ/rmmF4VtBQQzW0gY
D1w7AYMjfAvFwT/X9ziyOLecaQ3CgfYIqYovZ8PE6LAzAlXv4zf7SsKHPwgvKbwoFV/35s9NGGWm
Hxv6nh/JzDzphk6/+ENpgMk3/2VxdYheVwwh2hM9TCcPOMSQNvpuHLfWtZkulk9DK/sbPQh1vwSP
6+jZN16wvD9J5VGP9l1LWBJC5JDY4KBKhhYs8ZJg36u7ehvAn9SEGlb3jE6lvRHt2KJ9f3iQE/k2
BvV+TM5DWIBVJk/3bIsXJr8Dp6+j2lOEHXDuQbSd84opor1d9cPd+4RJW3AtTR4pFTOtWTXJlBK5
13z5V5ZmUHlcXXZ8Q82khxMv92MEB8g/pUXJN9i1aWttby8TeYSq3mkMOLIcCPsKR9+c7nA6vCfN
Tnao+E+vvYCoIaLwKsZMrfL6qrZsKdKzKKq+4cvy+YdZN0fzCXocQwHhlzgSGYjmLXkbI6bLExqE
NGmlQdyNQV4W0WJj5MeCFNcWi/6IrC690W51tP7f9JKCYgpUIItXaJRaT3AebFAbiI22/t6CjZb/
aaWSWN4QpJ0FqMn08KkDvsvsA6R7cUNHzGiVwZgLSGi5+HtipMyRUWUvNbysaa6/As9oQH2VYEaY
/THusgNgXUN6P07nz90qwQCpaJIt5f5V003XnNDpanNa+BZw5cQj7vUe1ufOz3FsrzHcT05HUGxy
A8cIafYJ/pPUvuK4g2iUETLutW9Qjbrvy04BKx2xrMgL/Wp6po81WA/Fbwy1UyBPqqfQt1PWDrWf
IUIaCkc0AvYXYDouc2uMMxz97VM89JrOvu9gR/sDu2gKK4kPSREHBpkQy648qYN0+bx3XPwrb32U
8LQUrgI3+mx9MDSBXvaPN5nbYc0UzhIeC34WbUks3zSiT2ucNALhfSQ6wbn9YvJOAgXxSQhCJ5FN
eNczQ1OcbRKrd3+RetlDugj3xfpoDw52VjsHNezGKc8HxQpt32lu9EZk6CgseztpE0v73W1jYyPF
BsWkMj2lqWoVC5KhZtGLeCw9tVVWaDLsUHWJ73NaCrCGmOHbiUyjWT6Fs0bggU3AnUCwk52WVPTQ
vAhHwno+fHvsnOUSaNtmVX9NW8TedDXlDO91HRWvdooCx4zEIRXN1JeGGfrz+rcL+Xb5rheW16Ea
GhDcFH6PYdGyHj5FUAci6pg091+wIaG7LiEFdPIX2R0EXxi4hFdAGCJ/KXjov0Q8RvkjL7b/wn9X
SbtTgq043+YGaSXZBOiwJXAcrEwZoCCOvPkjiHGZ7hV0ZZaGVJ7EBZg4xvYy7j/cEILayeDIvzOc
P5E/h9zlvrWr8GtNnuuMnPjefwmZgXGBVI3Jw8BwHvW9sGaQSi6c2shuLSsUypcoAO21UZo9FPIr
QpK2dpqkykdH1MXceF2/IK7MS06kodzmJHHpXubJVqi+JacVRiknfEatPVOrcmXz8gdwcPYRLemg
nweXsHDJ8NX6gpx3+S0V92ahXW7R4d561aTXWZ+vX9g0lME/EEZULHIIXdciRDvTSPH8Cdw5WYxU
+PjXyl/5u7ABwV+uPyAHTy34YEzVcdevY1pclpiEulo26x74gNIL5ECywJAvkKDh3NVPLYxSaVzB
l/kVdFtontBfdDuXtOYTRcTS9yFVcA/lMX+dOuzymHB/FEZzYxyQtsmNSiFWB1L9mIa2ndz3FZPC
dAI4BJ9oTXHJy4QQ0L30rNG0nUjquaRbjJUUFo6pTI1Sw1Z0MpnLwePtzN+mKvc/tBIb5fgT8pUp
wveEQnN9gPcAQwVg7IaIxFf0lk1qOY8wx6zqaOn6c/fqoSoBwCXZvUpkZEye/7kZRDLgd/cA6u86
g/5MPce/tgikkQwhOUbuQ2UHNsBgz2VQWpQihk2Fa8GDota+MxXZRx/INX/Bt8R6h9ugZh/a6Fnr
2LhJKDLqCPdT4PxNkOwKUR36+PcTKGoyzmFASSKpKRo8UBYz4Q0iKhNKEvOb3ZvvTp8MWaiDRwvs
AoKTCU/CbbqT7XHdXazvMNeTT1VxPJ1m+qdehAAO0HvSSvm+nOWoZtkLYqZlXvSwJBx3fvjik0cH
cVxzbxItItO4LAW/h1zkzeshWQl0lpNsyb4NXPTh0PSQAAj3g+e+hxAmbD0+PDSXTWo1p/wb5jfe
GLf9pw7aObCj2laJCQUl2eYrvXcoCiGiwbReUKmbSan69q6BLhmrnkDpfbFyZgcAq4MlC5M79D0a
5EDsmEkj5GTJrJz24avq6OrACgSlTJ7A1gFHoXhQfi7SwXd+AONqMcRE6MrCz2HT9WPsOB4rCp6b
l2sKbc0KPSaPtsveLT94L4RWp574e1uv4hyDYtqZ6hfCre/4Jgj6v9fWOwKVloQyBk7LAAaj/3C4
XPysflPOf0eMmKFGf7gzkAvtoYfaXKZ+ulL0x7Mn5zslawxZH91IHCTMvvOdQTCx0VaLsJcG7gNo
S5qhGhfQ4U4Ug0bPj4DdvkIOG3CJgbHF/waB9lVgH3d/5H1IkWFg3eerz+gQCS6zsFwnwgLKh1fl
hV+7R+is2XnbzceJJeh9+d0EV0qh4oUDKvU0yugIhmwRKjwd80gplxW6J2zOMFxSn/1Djfa4lBNE
pU20Rn5wI6XXTu3t2irK4DQzUiiUCXSe/iV0jUCQxvBM1yQkXqSB18hiHtJlRy+oeuKRg/4miCW/
O0oXO7x/rQsPKOTwxh40KAvVXxkTK3/T7p3JPxq3wDAMBvx8+KNY8eUOBQGTdznMKbW+cZ4BYlqt
+zZbzMVOqPsrPdewcxwPQ/zScBAUrbRnPYfAdNlmqiw9LGFA3tERRzFOMMaTLQTTZp/0AdemYCMK
o3pkxGaCxZuqgiHH3FWc7MbmWu3O4lqP1VU7+kroboelImbpZvoxSLqSDkV4ZzVsBgGYVWjS0mXx
olDPrE+jUYm7wnGi1GDyoZ1FDILwwHlcmXZ1y0SxjVQ4rhtvPQgMxGnKVDhGjb2KyGmrWgu5uxHq
UXGLCQGJ6aLBpzS5bm/cvKcbsCeClSixBH4MTCmjGvaahle0+V+0DdoyL8FgnEKf9U+mcftm/5hU
lahnqspnnUBX1qwALCTs00cEPLW/oDTSs5ImMr/IjLDAwlxqimc/rkl/U+VnuKaHS4gnDyGqqXQZ
RxT6LNiYDdk/RG4St5Lywr0iBFWWKrkLRv+VUTLaf9zt8g60WV3KEQOiwedWrcPT6eOovE7ctT02
BGBCYmzQA15xcC34BM4nj9b4k3fm3Q+8Q6VhuTYVE7/Fg2bQxniTd7wsNemjMKtYhuMMMc7kNGCy
ByqUgYr4ZPiMmn0fM8/6Xy9gYLk5/+1kLf7kDncg73prDHCjG1VkyaUv2gtiSI92tMVDMpzibYK7
xwHsNzTBuppxCzba1Q/FInvfbg3BzSEGN5+JV+tl9sCL4VuuEJAQ7gmxE6a4cVypUd5iEpMQ8Tfu
Je214nYM/5mFGhUcuyNsiAaXdkAuEG6mh5M7KZkKV7jWGRSZg2PjiXWhTSxwEN94zA1PqnSyAOFW
XksynxqnpJyFm/ZnFrAqUkd9lvWQMHuC12lqgDDYfOFsuSENwztIyGsvCFmr9DPClWsXoBN59xre
EvQkKbfm9tW+7bn+vLwJJp7fcNT232qHzDzO4MZzXdItJBSs0YKWet8ql4RZOzeefVZaIUcKihkY
flT9TIbGLci1/E5ZzViauVkHUdjFswnbDNeMc9HOVhdJVq84IT28ifL9dpDuT6KyolQFUbT/DL8s
7bSSyF97RARZLrRfNKEzyOrHoHyilGjbbKkfNZdsMhttFeadx7p84lhMX2sM2p0JcYGn+187qvxO
lu8xB+jirWzjlF1QNTQ4/iMjofdhFfNvDDmpajFwTfQNFFATshRthMS4vYtv9JfK61mKqnAj/lNB
cdiWYtu7eCknteGB08TXkny0ZixgPM7z0V/zatiIpEW5+Qp6lURUTIcW8oV7x7G3mP1D8Y36NJvB
LuRnX0iym1+omRD9BWHwRpjJCrq6Ozwd7BUZ7Zk5GtC/i/IIoqZ0Xir2SOHD3nwsW6+wAXWoJK5G
kvFzZecLYAbD96KBXUs2ULEtLwEH0xYl+GIE95T0vnj1aA+KMsN8DfCda7QHgyGlbZwuezL532wp
BQK1KLDfw/mX34f7wrqdUSbmLojT6tzIH5bOVyKUt97LSm46BpWwEa5L++HvFFm7AnuKidXI0DDA
UGNq4cDmPFjIP048f2VvLoaghX+LzcdYGsA4vUKy/R5ESOsTtF3vlbq7C2pkIIhruV8RepW221NK
PIPYrab1lvM4vpU3VwraBGy79lverWcDfiYfs/FuaLTmyK02QmbnCsDEnWt/l8sPokemWaEL+kBi
l2x0wBlMtV0hnEDebSuXOqQDp1Rq/Sv4KC7LRV73Gm7UkL8TxR0Fhy1vgRVmiPIJ+hvMRq5Jo+fv
FanvQarelRGyGnwbchwlXzT1NB5+4onP1FX6YGktaSIIxcy3MyEUH3zv+VIltcvSMik2wax7BqJo
DLpP99MZuNS1uU6EbwDPLrmlPbxISm4c3GULEj9fAJm2JUj2POI/k9buE7jgdn4z91V8jO4K+raw
Ae8GxvOKBrqa28lQksF3/lhh0riR76qHOVw7O12dBtRVM0G1mqTa4dNaqMTbxeZXFyOWOrMBWEEV
rG2f/ZWQyZ8ec8p+exVL9hmGMJACgaAO75Sb7/vk/E6z9YTwlWxGpSIKowO+PXqLXw4XE2sjIUnP
hBv9pLRfw6iHbeVHRiJjtzjLxD8v2Xt8cPsRdzTnbBkEq2DsIXWNv9zhWKpVA0vfNeLYP/FanuHV
+B7oMWCU61eBgZfI4LwyrX+P/zaW24+NTArM56xLDkrQjlntKo85i7dtgfrKVB42l/FN0g2JTLaW
VSugDH5hgVwt/b4xhGVdCA9KweJoawz1mDdtlghX2MkK9Ej/9CrYBVWJavnqB2YSGjYUwMuxcEyC
8VYl5S3QyfZUhPM2UDaFLxiq0Z27g1tSac5I4URD5BVrAzy+ydNUJSBsVfb6iQxgc+c7Rl/Dn9hX
R9AC07akKb+fWqx4+DbgX4EkMdCQ63sydG92jMc5FcdNBiVM10M49OeUjV9BrUks9ngkAsjx3D62
xZ34vLEqxGvYwBS6x0SlzMnLNDjaX9AMfgDb1Doz9tUpES9rLHTvLTRcoQaQG+yJQ8J3N7jl0iLy
Dx8vW0y28HkyMUR9FtyyWmihHVncxiX72QwcBRXTb22VYZX+bN2+md7xq3cnaU8wji1Bmt7sxI8c
PA8beV0CEPZQfU6+5K/ZM01EJ9PZC7wIBU4V7UT4b/aH3IHO4JWwx2KAPv1S1b18E3O4ZmqoG+kD
QTlXzYnO3b3YT4LeJtQLINGauZEHPCckgfMncqDuUdDBytO+AluBlcRWQjVdTJI0gFRS//Kxhky+
lwEohYegqk3Air+Pa0McXfxQobIsKduvVHjFwqdecm1zsZkX+J9cuYBOabS/i3FdUgzoSSTZnrAM
NxoOfC0sYKceQ72Mjdzx5qWb/4/gafwCoBtpeyu94C98UEEhBJbcbG2LTlJTd+FJw8OIYpeoznKe
wdksxw/AZNIite+9IfjSn889Lmksy0TSXhWQfhaps84bsKGOAOHXaTjkrAjHyAV2LUCioRcarQEp
jXyKkJg8Z1xqNnKcI1kJDyAYlQeq1HKLhyyCQvCAtIUc1ukpWFA7Ej4fMWfQ+u36Z0sg+zalh5BA
UqQ3GpWIl/iTVfRTe50QIkTnKFch6O6Cdkz0ZntMvFhhhZjrNgsKytP2kUBMETHht3PRRCe5y/33
Nhsk6gkOngYlEpluuWA2AOnaf6MKSrYomSFr+T1kgxzx7XO4jdXqGfzmrGXQZpS0brLKmvTGP0Ge
WN0iCvi7QVJFybdlUvmDLDCnnERU3thnA7FgwUlUMayMxxSKhvWhJ+aQ6UWkovdGV0Be7pNSjoV6
o922f+rBRdSnCIIJO6dpTTChh8dMnwNNp7laeDOhNnQ8LTBNIijesDyAomfEPfEkYsuVvcJ13gLo
PaBA2xV6RzmfmIBr8zcJihlvLPluNiFnU07YEcA5OTD2YBKDQYammv/MbttXQMp9WaHHiGECo6Xi
6/rU6HRgpekVvIQjYu7sFLo4MmXBz9xf48kLi8ocWYrvRxcgdwvS9YnrQO3VBA84OnfgrC7L64MB
5jQkAXhlWi93IOxBv4Fg0+tjx+kGc9LF50M9XM7DY94NVGDF5HAxMMJAbxJmgp4cqd+7TPpmpOaN
U/HKo5ElW0mm24x+ViAqi5k2gWJDB4gzPkqjWBiPakVvXpUfbgivQ8LWdBxhS6W9jQ4MC9HhDAFe
s36zOWmSzPZkbLF5mmbewXZW5DWzbzj9VU+R0hqyc+q5g+6o19G0sKxhQZfRtFqKIUY/n20RBwZi
7D5wUB92cCy3RM09Ju+YRQljwLLlmWIud7NkqtIZss6pv4Z7H3lAck5lnpksvmf6N70Lql0viTL+
367lNTFBvOkpJd8pGotLCLOQyaFazQShoNEPiRPXD3pTo9v0aUjLEdu/odzcq12zWlVCD1DNBp9E
G8x4Vxgjev1Uz8HhdfTM723ipgXKvgLxKI+jXP3ubMkYYYL76jf5c1YLiC2YTzk+xQUC0uQpPEQU
Z8m6GudLEIxl86htzRUwdiGT5Kq2sDLGULfcKyBFAhH4RV6VyJRYvBmvEzBcTvuADmi4+bzUmni9
VPJq7BFpD+6f2u5MgjUQvscYRAIABmyS25mN5xIyK1lM7VxvQnCkqer+6VOM8jafJuKBMW/9sP82
wsEYJF+Qu9M2lI/Z/IseGQJiQ2RNWqXIxmjG+sg8Unw99wP72gBXz5Az6RNr9IWacS7bZTTPatzq
qEDisW5+LWX6pVApuXjyzSvgMl3FUF35RZ4e0q61zZC5PbC4Nyxk5MlBIkXcO/rKmIcPzWkbFc2x
FW2geansswBk3iNOUGcYKfakP5VZcMZFW+BxoSCOu9Cg99Z68XhPmJjl4gWGm2nB7o8/H1+6zC5w
osqQKQojq2vCiOzIDi0OcOnM6x06v2YxMPOb3xwq58UcoesBTNY3vfjTI20fVflsIHv4SjUJH91D
byLEOAtzdMatJWKAkFwOAUr55Ac455I0m7S4w7wkQ78FKAbXlk2C7xOx+Fb22Ul6lsokc4ye32y6
RfnfaJGne2cSiHyeLE0eZ9oKtbPoX6Pm/hynVlH04yoG3HpMIZiSrFQ6Oe/7R9Z7EhyDymfPZMd8
P6N7MK78s2ijLOeY9lY4PWz/Vmvl6id7BYARy4jEyFyIPNn6tiMzcpDDSLFt/lDb4eknuud2itcn
ckUbRtjVls1Z13ubn1vXa0UMjFDSSaHot7xay1D1cbblOf+kVwe/b+VCxH401bwI9wHhuS11izP8
mq7ln5Kk+NNXimx6OsaoQWQtX114Bvxe9+N6PYNaiv0VJPEuEeipu6aCbBF8XuwPjGtiGU3b+1ZY
mBnV2/jdYKqhCwh22zz/VRwz8aGG3E5xFyahOPPDGwfY+/HkQ+WEhzmvkPnTnhGyXDF2m5RhDVtD
sDdw+hGAUqYZSHe5ywfBZZ5EhTIg6nTU6vq7wNw3iGSj8agyPCJ7vEI2LEJEGZHc1anO/7vrN+AY
fN8z0pWD14yUF3Bj4QZJ+DyzELmVmcnAT0C7THA0Oi2/byhId+Nug8wikFy7z1oen6elDPQke8ap
NLTD6togC+DVDLyWYHSOLFlaBJS6hkIYqggiYKcdb9cxUWw/Zq8JxTKaMpzuguouRrtqdOEnAk3o
t+5MwLQYsq4kDsarlb2cm4KyiCRyfvX8ALmCbYbhZF9lFVoecqf7XyvuzruYHD0mx3GD6D5beTdF
5lGK89Em+jjqwFX75VEF0S0vKZkxdmvr+z7WsuT7QgAvSPkRCt1RUPTImzLwFaenDGHH6zM2tXGx
VU8ZJucCCVBC1VDhEDNBx/EfkjtpVYFU/OGkfWPYFzEJVdpK5V4a2UDtcFiOdyhhUVphR6FN6VBs
xX/M3vl985i/jHMfX4nO+tdL7yt3TyDF0buE3SD3FaIwoU96SwoKdUmrTFCqnJ+JEaPgdXpEDPd5
IHpV/7ovTrdEvVlY28J1gpl3lweahCFhtGG7773Qe5crVq8aPwcO79r7LW/wyvIcRbwRQ0P0HsWj
fotSFKt0IwBBFvJYYjGBfrupoE86mKPl2y10NnuRmijSF/4v5N20Q4DVVldBVcpu7QBrIFAQ4r20
1ypXfkSxChYTcqyg0qon/NedYirM7DEvhB03oyFKQ3BQkZ7TgcFz6NvSRRt69qlv82x2mia4fmca
w1SggF5jAOrOif2lePLcgX6+82MFvj4/FPoYPhhp8CG8HS0o/Lv8VydX7RlqLenphCZcqVqq2jlR
ZfyX05tJ//07LoiLkAp0o9IPumWhDiW0QQ+JcPoObz8/I9grJ3QvvhqopoSd2DyQ8nrOH11Mcgac
yj62ql6a2/bNXcB/9KCYKpq0xPXygGSHx5xGhsB+d8eaXXZG6CQkXyUTp6nqX7FsNPRP2ZM8ciiw
2jBkInrNnzn4AY1tkqsZY9bCNjRblLs3BTDVdNsb18DGbxvp6tmf4sZ9EkYOip9EwU3V0qniZ0Gz
o752VwkH49h63A/EnbUVSiGNCyQc/ZM629sWqnC//LwWR78iD0M2FLpfzZKvWI4bzi5mp6qZpyQR
zompxiirjVcGoG3fdO1nmwoWr2pH4lTV4umm75A3g+gIXMxn8CHD9gzbdGQNqzbWgkZkyK6b1Sz1
MDfYqpPDIS8iFC4XpLwkJz4rVb02xRm82uLrfPj3tdPmSZOxDzZt1uX2GRBRTg8zPBC/nmtbBSVX
X07Q2K7BNdPuUnSRRUyn+tmEZwhjDez5JvQYooeriVtf8i3gq0f2Qu941x48hqohXzg37KBXLehh
IeYeNlzQkH+q8rSliDbQRVm4tOhS64ae0ozSI76T6gZyxOVSE28zI3gLV5ZWF6mgt7fP4FfmQwmW
eQyMpccx7QCCKzMuQsyFIllIlRuA+dl9L9vil2EJfL5ljaV2sblUFtGYxkAPlfJoHMzkbqXq1BZn
urdiXNbfvmGnfYiz17frmMEL8817vtGvz/gA0NigOMpWADPAalWeQodE+ToVVA6LErKKTFoePzSh
r3GUpcogMaDaD2J+LTMQXuEBdnnrDRSEkfCYkPYliQa0znxh1uyGjkoa25D4OKE7WovpT/PzhzSR
lJVppBCRZE2s29ZQEejQ0MBgilDCxPWf8prPQOOVDqUaaQx5fybZmXBp3gobxcfpxNHE7h1/Ko5g
mBnPbMlRGjDttJU2e0RDS4Lv/2+p168qf6Jj+aUHDFOOMlx1B0mxoM1q9l+FSn8iRuJbiJ+Q2W4J
ooeUL577lIK/lBRuX9QDp3I5sW2pcjBTmq9x+msrIbeE/seKwm4e6fQo9jjaHFGaGR1WNjOHv+gd
08EnM41OyIbpP7LLCJHR5vtC1nYbvgkD7nZw1Qspuld6w6e8Ism0DIMilW2Pk3j6/9ekvtXll4Nf
ju1xrLYYpF2StUegjyqJxD97kuU64Fi3fa2iu1I9TZaK2N+8V/2bxgZPjmP4NRPm9kVo47aBLNkU
IgOJc4csOQIcyrb9aFFQ83gjtpY/eks8H1vwI68kb0xkfg3P7NthF/0cdSWAB0Tel72SHzEO0Hw5
8H8qD7x1zx7CRblm+roet8DH3emtci5Bc+fdIYtHZYTXHx3gVmTDhWYLOEOfI+oyrZHzO9Gzn23T
ILtghY/GI0jpy7Gj6V67n0rlllPX0Rp69lb+mi5nGXdNLHcFjG57Au+5GnHPDml34AtEs5NjT0Zm
GbC1797dRtF88d8w7IYM5Z985fgaRNAyvLHAJ8VnaqQe6wIHpHtdNS0a/6Fr79kZWbDgy7MMzQ6G
ZWjCGzlH4q5A5f0dvlG5UMbkRl/kWs9tFOQp9JgLr4HH8VAgUbwNz53pXUcMgd14WaLsdLqv7ynv
6eKDhTaYRbAS4vXBqJnuMB68rCpH1qy6AgBNv41C2HeHaXzTfsjcQlu72QSZKC2bk0i5Isstphn0
GRGv0FLUIiB0VMaUMSYLMhqwtDBpEZhBGOGe8F4pEsVPoaMVyE+yb6QsdvnugH6Z6qVu1TEiHMUd
fsL3XDBTRtWpvIF+MUE5p94/KiKN/mYEYVuQ7ERsyWzg6FAlxhTrum0PVP9mgIYYqkFWEkdkbP8j
lXG4hAFy0u3mnncaKOI0ic+TJm+01i8sqWkaaA9q7Blk0yusrvcuvlJJtQ9laQ9H+5RVKsFCVvKP
eB9iKPDicau8Y+kXIprRi1EqRo24kw4wFiwjCd1LtDVpuK6zW2py2ooTQABdeWOH6PeqAaaxMxVI
xUmLrni2OWWVYaX5sQ0IbOTRlmZqu6i3V9nOikeCMIkGZwfCCHZ4T3xqS9d8YDSYgWk+KKa/DKa6
psLF7IbXBg+PbM1GdQX3AUA5P+iWTzeeTnpUnoUG0enl1zuz1/J4vTFsbAjizTxnVQraFpF61vD6
iOacKLiI9o8JTr1p8B+3qJLaO2SunICl2OJY+vuvIQW/v5GJNZIiPwF3CePWOPBK3dBxvMinoq0i
15WgeWHlagtjznRzNCr2UwkEKtrXuNaV1Mn8LkTVli1jVMFkB2d+ToOLJsS8QtrlTIcFzZNWW/ls
IkyCvCPfvIWdsX+mov6PGovC37TpMJoI9xHl2vw3KWY5FY1asu4kCERUx/DMKA5ttlKolXkE8H2Z
fCzuLH7JA1bOEDVoZnASp4aIx8rnWf0S2VaEh3/j+r/Z1w37qHkXoZFpGwZ35iluKdIZEz9AgsAw
GGqBYn1lX+z5/fOudS+5xYkJNW3JawSIFwRCx879BDGJxezozptjC7/5pdPNk/w7PVCh6X99zBCY
q5beIP/ZSVqh1qeD2n9SAomWlbDcBTyciXNkBQD7hxPBnRmkL4oFUH1JjKq3bjk71kQXfAquBN+X
N24C/yqSVO9ndKOA6shW9t89d3zxkIJbFWTcuCMtnspVpOtKqYWnCtRotZbn4SlNFYmebPSO77/Y
TNYcLw/KoP44ueiqiaD2EMtPovw2EryQ1n/oNi1ifGmgkqd7p8rISQQSdSlHVCMVJ60nakvt+E4W
EQHwDI55Nnv0UUJuQ5PvNuNESOa+QlhR9GkPwlCmcA75UmK4p478KyQvdBupqjClIEWmkrWtT4lp
2a3ibvTlOH9nLakyzKGAjutQYqIUJ5/akQggRv/5wWQ3bhLb25z6eOsptxj+xrNxjDjAL5zzPQa2
a5dpJviLozQJ0ix7xtBlBZnW0GD67oAT2iTOm1+dS2sLhJqaQVmfdbyW+w1LXVewPRb/cyaKrxhv
wsyp6fExJct407spFCXWayA/Or3bEciCXi64Ke6sNA0LtixIJ05iGT6L6PVkiKJxIj7YyFXzotpt
17BEGCWXIaP2K04f+5n4aym9OYli9MtnvdOq86NmACB4g8Sd2/wB8qa4K0ZfQC2vTcK9iPPjst4c
7BYZhaul2NEsn9CkbfVfpi4lkK8R4XZ4BwCaicbnx6RKuFk8KvogmJYj1IS1ZjvolDc5jE8Q7GRN
zBDrAFVFTDYgYWX+Bw4pLp+aqNl7/Z1VQJoJUQWI9mt0nr9TiiLSmla4AGQB54UKXe0u3AXupuY0
b2H+8tj2I6QKoqWP8HgOPoKaO/C3kCeInDIfXtHaG7m9wjAFLRe1iS1ss1uLQLyCj70iBC8hq56J
ZRUaV6X4XP0oOvIr+daU3jTByMO8q+piWk3EpRg1AwiuM/pBIToH0FshRymRgOGkGCOEcQnbn7lx
Ev1inKjbVi8guM6lKiUPTaoKbmfZDVKXl77r3xh7Htw3fgFFf7W5frO5Daa2HiZfqznM7+IG9rrE
tpiJqs5qAs8qZmGr+HHeuyVswNzEhVR/Hds44o2NCaF+92MYRemUm0y7exbLRPeMzeK86gnLYzNh
w7NPjZYnfOO8M8BYSrhHoo7XqWnnxCmZH3WH8B+Nn58GHOxs0DI0ZHMwkPg8HBleGAxjVVib+3GH
9kEgawkCGw4wY/joh/VJ47p+BUNPLg3RI4R4yCxcmByW+H2geHEVmtGmcRndlY2o0XYhV6rc/p3x
N4KFtNABupotgcAeuHjrn0AQOfJJGdLpnQqAVd6m4eJX7yID1zpvlOcP6kL+uJaJljf2r2QcXD5G
DGP6iyH8/ipm6iP6FEO1S4tlZ9ItqUj1jRw7hw==
`protect end_protected
