`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17760)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAA32yaPLPJq32rSxDZfHSvXguEU9onMYEfLvq7I6GL9swYlsgmBp33oV
pjYp9Zp+ti5rq0Zc0FzOMs+UaRvLQH/7X/rfEmt/MRixoG5Uj12LDiKUJKbkwB6hhbWLHNnoxyva
1Rqw4rVYoQbQ9HxHjwT+gnqNXZg5+8HuEx8IarDMBMUqvVaW8t1SaCjQrqtm0OZDbQ855fZwc2+l
QKYyYMM55IYrP8rhhaiJi33t4w8Fk6lEMUbA/IPewty7+OReILeRrQK272IYBPG5oCjTD4QrTdov
tiM8zb+PRAD8Ztdlzru17zYHBgn7fC0RNQdbGWZgIltjgjmmWXKKesa/cHMVbS+mPW2hH4t2N9eE
+qVQI7Udt4F9DeXRAP5Q1UYUNqtZMHBEtcKr+O5ALYNXypBc6Ftr3MZE8VPB3pFgGWMKa0LOK2Vp
jYr44JUWfc9e87Zzoj38oq66pgA62xRmMQXDnmtZsEMITmEsuuZq7U7TOBPQ7B+T+Rh+fhlPoyvJ
P/7P7xM3RJrxtK2UWzyy80+n8hbaOuZwPLmeCQl00ZT4hXQ7c+zLATwc9ltOcONyH5BxLd9+LzJE
ukrO4e6LLthuJsNACs4BcCdn8iT1nwzb3r7VCilSoY8/eE2CgEb3x34xOVzW/gA8FQzicjjVN4Cu
baiq5ouy3NfH4ZT+WhWA037QZycqQPcjkyZ5qxCyQPTmJY1ARIIFLtVoOyQAJIsUfz8O5jd/ncmI
Z64pu4p/FK3+COIePHc78x4K7ckGBaam7u76cuVGJfpl2r10N3Cczekx8k1Mxt0uxv8+VKBvVHSm
jqNLXxkc+mD5xs6s1/9FG9R7Ywvj7kJ3UYP5GVNvC3/bveEjMVUMZIWGnht54dxSMCWuFtQTEsco
XRtfPNSxKEaGoD4o9e15MDSyQNkIgiRTUo4gHbTdnrkmXRrvzQHgj53Qt69OvEqDJdfxdcf56HiB
ywizG0D2hBBDxCKWBy4QTv/2eeDszAaGiZ+m4Lfk3M5JS7SUZzTdYTfxSvjGxkfoZ8hMX/iOj0K/
uP4kbdoZzkYqPg40pDG8w7l0MfwFkTVXVbwLtlrsLrOIfuRK32sqYRzVzg+fCkSTdxiC2679tZeA
iQtAH4cSPOLdul6QaLRgYC2KmJ9YhMAeugag4GuViLtyPUY8D3MQNFIkk+x5JlyxuNmWQ7YHddwz
ZJFDUL5tPIZGTionfimQPoVU1cisAe/jV3igLi2UOvQEzrFiv5vAzxc+aqHJHSZnvf7asrsavrPg
Z8qSr47Z8hRD1oNjxV1lFR7yGPUE/d0pICXBBghGkxOOVrbRRfr9qdn+kCbsdmUxV/BJA4Six/oR
6vSOihrhM1I+/o2wzRdwXpJaCUY/r5+5d3nkJ6s7iBn/WqQM6iC3Ba4XHr0PQyCXdxrs1CQ2hU3W
e6azEnZqSRNJ5Mzggu153XJT1yAoiiI/b04NYfMHnpFc+SOqmdDTkRCZC10eKuhVH6WMAXH4SCmx
2dYSTPmRodNGYltVSCO25JnhD9RYDlpmUsxGcOXOD87idLqlqTibWRTDSA01dlozByG4r1GA2yvy
rbddvP6ZaOLNN8953L4uRRC8LymFGS1QWeqyg1jbJPcH6qMhzTe7hkOUbuaeVt2xNQwjXBSN8fpL
2eJBNkK55jYFdhhHUFvEnKzkJoUVfjF8Z97nKGGzKWpL53CgWjIZBJsn08MEE70pfFqLD801oMjB
hpKUMK5QA/tX3ZYouL+bbvyH2mi9yodMcYZH+p9ZXeFsYjx59kckRu1B5Ri+/tISSVWhA+WiaSDZ
xl7kFQ2BjO8qkInw6SUIVvvaxsWVd7KWnTyOJAimyRB/P8BlFgc82pMTpLLvqSKNLB6rYDEFvCRP
XTgAnW6HXbtnbabDuF+3nGlkIaSfiFLslmq8XpWQ9OlaCRKB06qWkjNLdm1p1bA6l61rRtUq3eIc
YkEcuAZtF2H2zmA4HhTeJ+tyiEnwBFDv4IwDCzn6/It5reXq9DT0GQdNm5BWTvf+By85qB4xXRzV
CYibzmql0DyKXOHf+5GP1LW/zPQ5+3bcvTssks5pmAgaVNUTLVt2QxH5uaqzaBfbGSM0m9jjma/v
iCAnMRtBWNYeEH9a/sGeESRgv9INEsmU7pjuSAQPxBzanP2vERq8ouqyLjA4eq8+2VCoIX5XOSyT
ILsz/fX7zACXFXwxhqbCqfu194DlXUaL+uumtRFMZ7JfA6UOx3e4bMf0em1a81dbA5WJweCa3EEm
twZk0PiiQ2QBN8qjpQrw2PcAD0P2QHuYou3bNVO9wfihv6AYngiA6M3UHeVK8pn5ZOeb15V67GKf
LXKGcqxZtqYDanE74S7kE4ztCpGSpz0p1WHVMqIQ6/zJCGmKSkPl+DNbc7q1Zt7Zr6IOgzqDSIAH
nd674xZ3fxdbam+3LiwxUY/S+Dy3F4pQlH7SR8ST8+xLFdZwmvKb5i02W/XBxQSq6+wFuNXHabLq
WVeRL4fvo4K07tXOy7fMTVsS43OPv2P0CZHdOKNmgMCRJHcM/hw8jMIX8duO4d7fRe7TO8ILJiSJ
2Nzo3eLzcglabNahhWf+LWm4bDVy6yP+piuzhKrtasykonuMFrz4wU2EalVNKfwrwRLJOzyECdnB
7RCBkmIh6i2Ai6PvU8JHPdkkT66sIp6er5ht4yOAaU2bBlUVrnB3Q1zOe8GTS69JUCsDEjk2InCn
evF+zH/ExwIisn7WJHjg5JWj6VFQeh4T3kpl1fJTK07VuKvRT77T1QuYntVas4cRhPVO9qXBfPOF
SU5pK0lKnEbGPQu4TOUAfNhkivFVd9ca7r6cYcvNUvaoelszyCJppn6odimWHxrgMeZGqfqRiW5r
VTbYRZ/BnvY6Q3kx8brZnm+10qWAZVIoDjiT3NwJyPf02rTyHC0t2WZJh2d1NGG5Sp8L3G8UWdbp
uXGhfkIhigCFSQ4Wg48DszawOKDh444JTnezrCNfZE/WQaHwd3QX5vorejAknqx0Zny2G1+VNsyM
Si/zkRvPeXPtkFe8ALiPNBOkUlm44lx7sbqJ3dL3QJRFssAqenAzcTZje/lHVQ2FGRRGD96+0vr2
nCbGMBnNqTrzwUtRbPUFg/jn68MCr9kvxHMnjNX6mpJXMwm+CPWqS0/g3pGUvQEFoZYbKlK5YCNP
zvcgx+sPxxn47le0A/ooQEAn1XJ1QeFO1oPOWE7Np+48zmp4q8++i4n4gRu8LQAy0B25+Kx0g9op
kzZr6bm5cZc429PjzQao5HMPiqAQoRrx0Rtdz1UfWcxtGdu3mQ8nYHMUEzGoXOPdbmH5Ue1wU9p0
9abDS5FW8XA/fKy0ae/17uWN+naaQmKtbJ8coHYdzKJXezgyNNosTyUw+yCBv2eUDEWWPsWQ8/zr
FZSsl4M6WdKNEIPylWe73ZxYYJptMUp7KMlodACfv/G9CVqrDFXG2tIXkOQr4GAIPxEuc7NBc+Dy
u5qml/51VkDS00F12KzCAy9BJ1kYwaiOVfFvxu37Cp0NvNkCh0Dda1eGkH6LUP7WKtJoaZbOU9kW
zcLnlfV7vpkIrU/UmvOqG9vkztWQzMTun5caPehqmjziVgU1qnUGiVjA47q0vZPbEFfSnp+WS4YG
BqYc+a5o1tZEBqP/VCxcge40w5r/9Z4zxIkmH3abNj4eKEVTQ89kwiiwS/wsZWmKrTH5Wv+qEtML
f32Z2vmxc5lUBMkQBw3JSxGKxvIfsyMtYuxaMn2v6gaikdFBAWoDleL/jg+6eTA9xgmkzaazPWsw
xxBRDVKv2QLhuW8YG+vfGUQW7WrYstdcazsEFNdz5zGumVzyRqOAsXAFemUnkpKHRuT9gOFpHeU2
JQknwE/VXlwKmB1fSEH5/LlESR2OaPFILf1aYOmHftWZ8AyEKznDYItaBD0x1BShhxfyD49KrM09
heKrCr1gvdxg9xbwpm4q3Msrqr7uqHEG3JxycEknr8YdoYwxlMBhWlsVBvHiazXwVwWzyNio2p8L
NgVaaiKuwDbJrIOESHiwNXQTW1RRAT49A6IS8cH1L/7XkaeGgNQzEHCTGJK9lkaudB9wDrZd+CSq
LA37WQDoSxSCMsCiky5axEUiNAY3pd3PlzR9Q9QKZxaD9z9Dq2TTwv+LlNQ6xgwXZ0m7hdG6VG71
CqGwnGXRD+CBWcTGE6HropVGw1+8VQtAm+a8XfaC/azYxbbLancNhR+QNePVLG/VVnWa8V9WVkWZ
OlCPUE6/05N65ylnVjk/HZi/aru8l0AU2S3eR8ICSqVkTSX3HK+y0db8+nq7cKj5X/7XX+C6pzf2
ehpjDC3SaAgRySHMjpPU7GDraZPvEDBhBb/hoFvZM/bAFXyrrOW8j0cX+d8lCVS73/zwVZC2lk/1
Y7oUq4uZRUul1TbxUxSTE2ZpYjl2JvKJzjxtO0ADQdeXX0vVsGo5qmOLNdKqHTWhXEP70m6Zwm2m
hrXb1gElj6rldLqPEwcOo9Ljw0/P0pArqU/J/JUMBFoUYy0jgqHTaPbtZxIIYIIOFDToDyfHwF0x
TeqBZnR03e/a9sa0EyE3t1qhpZ4yFHiOmYVxcp5i0leIafU0qKLZlqFHpHqFL7mEyT2v34kXxibH
scQYjq//MiIvBGUZFqNrTgiESq2FJ3lOd6ERauXEW8nkq97ZULsHndKfFkHbxX9f88wJuiPErUHZ
OrxKKpAO45CPAEwV+KRvfUzHWnJk0vReAKUwbzKUSLI53s9UhM1CTCv8h8Im6bmahQYOuqtYC5my
u9/gSelVm8xydtGbdD1XZBVRnVhHCVYeKBkowCS2Ayb1CiHAqpiPHv1nhAcSzjICY3+NgSo533cP
VVdgGJT+Q8SOMV0itB8H5tiVSEhuOkeqsbxvT265SG9xdKyHgnXnGdjzkrJYyQ4kNM45rQlCmwJM
HtVO17uVWss3IthhKm3Q6ZzQ3MfuUbBqWMOF62oWN2oeybGvwU3p0bdXd4TwccxeNlCD8UT2TCno
PDkty2jF/WeNQaLaQLdVj/YzCVQl85UrRoKNtEZ9Hiw2bgVPNhJ7N08RAfqqtjysU6qUYZQEvD8j
ohGTTyWdKSqqvS3KP1al7PvAfkaCiHlGeHLfKwJw818NkB8ghMFsM0PScvcQpP43bOxbjMfcr1St
uWtlXsbcvkqJyKGhiVIrtN+NM9DnL8ypkEqVTr9ZfcYg+MhDRYI4m8MD3iNQ5U3h+rf0/3e/8zYu
PcDYxyBSXYdgARvHb4H+Ui7XZSBo0Bye5A3mpCSVyaQbDOU4ldjZh25XZNDlucqELsYPe1JsZ7UW
/BxXEOSSTcanya/POQ98ftk4yyfSEkdLfHlZ5Xx/Jjm6cWpUoVAP5TTBc2n5TB1genvBmTUv40Et
mlR2kA7RPWkYM7CKcSFQlSy33xMEtxwe+zGVeChCLer9VrIV4uTSGOKVDmc3XoXqo/JEEv/zTjy1
OhwVO0aJ6jpL1Wr9BqMkET1J3bE4peupCXe1mLKzDxftZ6h8fLeeVUKx1lDiiHZFO2W6IFs2Yf5S
FuQOvooeneinaTCLQeW97iBvqw1AxOhOISu6DmeBp1ETwMam/V+TNeuTRcx6YLS7hbwGWojuguCS
Xgub9zzrv2krGmRBkDD9vZtRvvEOzFKV+FhtBjQ1zSe60yzmBPy8hGYYch30EvJfd3X/4xIwLCAL
a27VPGx/tExkr4KeRR9l9GV7zZ4QhvV3dH+EUEtkDmiNk0YUejwvTocl2pl3MGH7N9oQ1vwsYU4W
B5MPSvhL7g5uDxX5sgrKZbpQXyfzYlKnH+8j/t2+FWPKqg4clZd5rLA9hW5YV/Q/MhpWM/Li88vJ
CeR1W5ErTSuBFZH1HsmIlJVgV7KOQYb2DUn78BMnHam27LMGxnOHxbRKWdd/Eo3auw6mPe5CLUc6
MAuG8yIBPBoWiC/yG42ya+U7C9X10a5p2v6Ep17JmgS5+Gfzbg6VL5NDo0XBQfHURhq1OVOGCSQs
ygZNNmcohgS8QWyR/H+tSwBsqahdoUzfLlW47K2iPWmqxpr8bRPYXTi/OI0vlC2qA2TsCAtuqe0u
gpdlakd5wdWh2YpOn1vXcdgELCwiyY5mjhTmeOCeqEkokvl/EHu+2YwDVBtkRAeEAoN1vAsJEpjm
JxjKsDX7kHYIVK67tnGbP1iQG0cBD+n4sKlDKOsF7Lk1Ol6DhiD1GbIuWzSJKWtlnPJJGeB14tgZ
sqXVwgSBSB9/z8AoJ3ndvQxTU+7aPjqdDkYBTkhTMYRo2EVT+ViIaHmHr27X1a6ijJYpyaX+k74o
jqUycR1UBC7nJZLKPxw4uGYCTneGTNb3ok3/xnrQUeTRExQsV+N57gjJVriZjAdyuiK4BbOoBXU4
d5YTfRsXXwzfUCjfWdaAL5b3toRzOfXqNOyhtQfzMuMQOqjQABmhMcjWGKYUShrwLLAI328k/GIR
jzQ7ipdkqqrRtjZQat6JpOklQlyn2uAPQ3cWnbm/1bkMFPa2yTOkJlz0qBPY9j/GI3ifQ9KB6y7i
gXiZ3ya7Tt1QI6WYeHeVNiRJacOwLQdEMjpAc+11nL+O+Vom3Bo0kOX1C4uR0yLAe0iaGJdj7Q4O
1TW3Dr2KnErPaWfAdZHR3GArqVNSbECn6mhP1l8xPpUIJRi7NfFFxc15Nj7xAStIVsJMJLLOrEia
WervwvzKAtpZx+s/d4lUnbxrkhQDHS8LeEQecat3xmjPWgsEnltL3/ggEaHUhVbySVXfeTEOYIN+
PTJI5fpra8ihLelKcSTtzT5P6c1zJiUoxIMLFFOySLNkGUM6q8ckwxwmetrLwuV0YA09LzPXigrs
DUNj+DzwCfPvudaiUnWVjmCMOepYR/VBWfbzOWzcodWxt1HobZkRGo7zVQl2CKwA813+hlEiCvVk
hf8cr71fL1GUrTcW8ORZdiV/O6/cRlS5BaVOZfSGfaFl+rf2xl7nCSgBT1p2X5t/GWkC0nq63pk9
F76vaAF70GxbAOFNI5q6NBnHihcmmX0QvNrnoYlSZYEUigfQPcGTNBkSO4WDxByGHWzBSuaB9mbh
eTENjwt9n57Q9wHByly4uoljErF2ibeDyfMlI3kXEkZCLTyNuCnJt2taiBnxeuThmO0Oh6JUFv8e
4vpg6IWVfjWsOxxK863xyUWJPdTo6/47ZFE0LtRS2WjKO9oNbG6BJ4nSA9E7u5FUKY9K6dHy0zsI
twHGHV5LJaiS3eynzlSjGg9hLgT1PHdpzyfI2VVZ1YyvobbY1Uvi8YiFpRXrolBUAwSVh45MgFM4
UnnRXOALkQDN1BchhDVB7porTVURQtyph089qCeRaKt181VvJEBQLao7FuipwQk/w4s3s6/jYV89
/1nHH5tSZKVGh9GyOrMpHFjQgbAl6dCpVh2PYlGGHC0+E2k/xHakKy8vLMJmhYQoEro/q7HCpaAf
yIyDgGAbww93RnjiGvSxGhTBs91bkIUUURCa5XWetWuBXyK9Nf5lC2MBgi19bnJB8yAULs+ixvBp
EZSI4sPgIIO5HYJO6PmtgPGewrgBGAuZIM95aWtwPmJIuuro+VSiGx0UV+bVid0Gnn0HJT9/xvqn
7pzCmGH60m46z9F1deOh91Gyw6h8PePCxTwF6WIU4SxfiHih+dyg6LZQH2Rwdx0lFZEjbZx/ae74
VE05ukAmBMo80hOYmc+Zg+X6K3HThW61lh3IM2ZakS5//NjRJqRvNI9uEqRcP7VenInhtLJ3PCw4
9OGGoZnV5/OR+s9dW3LQghAzP3GfYSr2Dar0waD7OvXu0VoIYO2hg7gP1WkOS8RGt+zSlT94mkmH
5ivHpxuBpngclUN9g1/7SLUrD/aIlZXpdt7Jxli6G+LejQuI3zEnedV81Q76519wtMm6XFhZko7D
D/lzFA/VXR1vcIxsfpTbkqNWud89P+GL9zBdfvkIlBq0TRICW3HO5w08gnIulKzaP+ueCGGrouzd
TK4vj3tdvqVkdTusHCiRpSG0Y0aXvnjFt4kVFsTZFdHdst5u2HUCVBP5jyKFYY2wFyF9wv/V0c8Y
+rwIkNF7zSlTgnS5Moh1dy2+T3C7qC75qdwKTOZ7gBWn8l1KYF6yTfX0Nvr7emtgqjSxG/SAbtiL
HJTWOe1kqs6AuOGmhdpfb3Nv9YZWJyXkYHZZH7+gxAMI1dtDOoVxI882pQsemY025trg4idM2kLv
Tt9dqrdUZMu77h1BCTzSv1dQE6K10nds0PMtw0c7CjUW4ZlpYYNjnp5YP02V0J5I/FmRb0QbejvB
hdBKkFpEzL5TPy/XXHk82u60SzG4f3iCLtmztbh4B7CVOIgpyTklHUk7MrjL3Bb6Ztids4ZQtx4k
eYTD3a3M8Slx9PnwZqFBWpuvQAoR7KEUI559BRAGi4SFqgwoRLJ9wHx4KEkYp5KOg0PZcwNmDlMc
aaIU/TUXpGUXeqnjWGeA3LesG5Mn8Zs6jvlojPkvimYxRpd+/T/F24eDmOEc8OOkl6hQoXmK/l+m
sGqe/f1xYLWOnqNBqlGTURoVjmrnsH+SFS/k6obBeywzznjj2OpMMHwBd8Hpi1OZNu7UAyyPIRK4
wTCypWMOMTYP3NFLKn2VT+mR80kEUUzeSIInfeHA9rM2TIyQFoYSgnVZ81+4Z/YSsDQxY0aFudHz
GuzLLjFOGA3C2A8Hk3Tvv4comoA1lzAoGYXxnHqhGi4WbfWbkRoezprCelN0L5h0wSydjp66XuPV
g9nAAAcjsR/kviBSizpdEZrqTRnYNKeiHoaeeqYM4WdYRpWOUOQPD0m9XHNJY01Tc/HZIZQQu7oq
7SuidyDwpW15NHtMdtxkDwVIxe/c1p3UlZ+3YVCPna4YLANK6CvaMKJu7U8uVxRWZwA6VyGeBt7e
KziwPZQlG+nsZx0nQzdF+F658HCtEy7hMPtwRg8gM00zLmQYTOU5AjEsOEQLv/KSo288qq07vgzS
6X6SyKXmbZaiPcYJ8u3vWg7v4EMWyh7JQwv1c8Tyi5h1bzgfgGtAGuFuyqBj3C2gyCZo+ml1H3oD
WbmJl3ezFICr8lnvVtMDjTTBv5o8I9fdWvTCj16FkR/PTkkzdIPqaazrm2ilU8TKneWH6nJrlctH
ZRs2FKXBloRPR1mCbj5KZwhq3s2MRKiRVPotYQ3Dn7h5xQgw/V7WcLA++7jpQ6zuwZDcMp4fuTrS
yfL60nel073nys55vR/CfEwH7rJGg+Map0hSmVolHuvY0QeBCN1WfN3SEGlsL5DHukWWJY+wmlNn
kCuunTisFxj+f0GkPmHTtt/ZLc7xDiUbT/m60ysIfowXFZ0ODUk4OEuh4j8aiybCw/geoHima9vJ
jfXcbVaSLJhD/v0e3xW1EO3MZhQWiUFnJfu6PRAlW8JKqfBRrkdfWv2Hriy+i+Gkc4kK4UeUdFqy
q88DQkR6VdU3a9MXVoEjx6NO7KYKgbGsYQgQWsFGXO691EqpSrIygM2lDcYnDjBGhDjhGjQHVlVY
jsGyL7lMkWTIehDb9OvhvXZLaEFpDIZAPkqaT5Rtda4OwJu8IlUaMP3veh26JbC9lWaWlr/Pfwl7
nKEFrZlTEZi7nyvEVL08AIao0qkwcnvCoRApTNjagi4Qj4z/hRG7wfUgdKlbch3rL6miAOtM9p7f
K7GopyG1u0Bmb8pgZQ1eqFNNYBkjD6MxndmzUnoacYBrJaxOychjAv5rxUNhoElIKxu3/jNR9fYf
qepgPECXbWUS3k5aI9/sK3q9yskC12+//KBagVOJcpE4EYvvWQrwWaF9Tbo1ZZvGA4STu0Yd4s/7
uyrK/zAMr27LVb6tqSW0pdNRN3OAvnVNhBiPrDj1ywHzlSwQt8+y5IjNXARwARnT+syy6NZEaYjH
umfks/SxbEiR8sD6m+H3mPGR4acYKOWIwkL87N7MCnfEaMYNMnya0FvLLoeol1D1as/5MTSATETf
9X0sDq6oDEQQPNsfPNKE9ZuS8Tjt6ACh/smuVhDQqxSv17orIs0lmhFTjIO4gxksoJLuvXMi4GRG
BJO1ai3bxU5CPprmG59pi32gsA3OSdHxgCYATO9XYqRAArm4gq1leoCUQxDE9qOvl0oRCPoSMOA5
ZeLm5nY+tIDz1wkmcxDombjGySh++YMT3Jvar+PzOSIewoTXJq4Zw0OCyJHTbVtxnsuntz4zmcJs
UswIKNzK1PtT97hDrTMq/wa5/Amd209bSEPpgsWswRX4OjNnm1S38ScXTJEnxD0FGPKXogOW4rYY
QcAp7YyvgUkqE4cv0vt5tPyQA0ve4iE2Yl74oxmdeXL4WuYwDCJYxQNJkkOEwWSIryv4G3zxITCb
kF5cyQZtbXobHBcS2xi3Gmdca893C4sdn4OVTAn9A1uqLgDkyrvOhJ8LvCDMvLsj4L5Cj0QYEp2e
sSz3J/POvZy7rF9reJC4IHbCKuLpF5cgR2u16kDn8TganyIFhI31m98i+2rHu+McIeZB4k1FbN84
d1YKWX6YJBp0+s9kYUD5GRicivjbdLShbGr7GTB3AjP1HcHpkaOwi/KuRGJeR+GlvhrNAlYsi8lx
NL6QTJEmj6KYf5BZT2PwoB8+Pg48jzkyXtqExICwoSUtuQs03Coah73HUanskQy4jK0yHc0JoaBB
u3XOtdh8TBSSOnKSMLIFPJnI6lwGGoaYEvhooecVLGEOxjH73RRsEt7A4ToC/M9xMBNXtBgzRKeb
2sJ8a8L6+W8Qs79I/L13tYidvmIZ4KzpSubahjHoOydBe2GWs9KHp+MmMTaRNpQuvFxuatKexzvr
UDSVSRq6hXTv7tLkEZ5zRGrcL/IomwfWYM7tyl7umU7liStC9U3uVp3KGqmkEyngqvOdAcBsEaY/
cA0sjwCOjSvEWs4jC0EaDb5A5OkvwAMxFjJqc7kOxTdZIF6WQ4qHnwdk0dDjfXc61fbgLorzpsIT
1fC64ziU3QFZasrO6ySiOnqHsn1bwQ8KDUMlk0+jOIhD+15yqvJ1lGVX0AKshl2qQXNyAq7hRW2c
aWJGh6uhZo7mxIhtlXqKGHGqVF3GX6F5+ad7nHls98oOLQYi7STfyL1mz0SrXXZk8ThAvMufdH9L
990RicTPj5szetvJXmyLhyhZ0AlPnfQerHZyQZFCo8IwDtcx4cJJt+VbGYATgPuUeJ6s//ULWS37
WHRsoe+96rxjGHgnhzrI97K9oUy/QnlbJC4fyJSVsmZ1ekpTY8zEPO+pDRmsDHIAMAw1hVTv9LMp
hHImA9xp5MrihS+eq8S5BNe/U4KTVnUtKPgW6KsmAUXea3kSnMU7EbcFu001dTBd5BtxTLUc+2Be
tJGmYdTjcl00PmQhHHbl5w2SUVP7lmvzBrnSXaUfRMvSLd9YTnKhO3UVMCLlnaoCP/XkV1Hi23AI
0FItyWl+iMypRyCqO8IF7l0N1IPiiWlSQA61IIqGlIXtWIO7XV9CK82L+TiCfg8tPjLlNqrTv2Gq
Zrh7ru3kQvnW6UB+F/o6lh+eT+pC5qF3Hpf2c0JwnyDccSG+qu6/2rPi+FYunmdGyCg/a782TYHU
XFvCBYRVJTHUBYUOYH2K32tf8MoUK6zQ6EDMBLfg59FLHCcCnWQHTOoDqrG5uw3UG8xVXpU+D5Xj
/tKIPiREFuFr5hH21bzrQbkqkWhUaEAX+CdXgShvVA4Gewg7q82C7oc261RcYrppODtNgsD/PjwW
yUS8CJrQR9VHj7KgsCsnb8hm7/r9TL/Snou6yieRRZ+KmMw9zJ6+47+v/NnuBZXdW4b0Zs6NoUzF
Wa/mXA5tV8aNOXFqDsdAP6GNRp7vs32rbOI9GFQJNMom7NogkBnrW+mE1yujxUNLJtjiQHUGGp8/
raJ36UimMGC8AMOck1LV9ZEqhoytYoIaIjEPlXX/zTuTCJ58rSqeiQ5pORDOvPwvPV3Ci/RFVjwT
nSjTilmpUCNEPErhzi3ZjjSCOWVSWQy0PDpN57SlW02AB8qfxSpR0tWiI8Z8ngrRZU+ywVRCLO4B
N+ruaszxeKkk1Z2ExmT+pSq4GpCi/E1tlnMgxm172DWZMpmvwc1cDNxjzhWgDgtql4+QtlbGuv8R
+93mNRGsUqw6H3KU5MTIOVjnPLyb04J3/GfJfoBJUVqHY/uB1C2mvQf2jIPe4G1rkgzWzbqz0uNP
iePbGvyJQRlcfwKqP7ZCdU+sPjGjMu7fiWSprOJIgG2m+UhjcCYbmb1GXr1jDnCSETZ4Rt/IPAr4
pT2LkezriXiq0mDI7B6BX+N1KbENFB93msbBfwAnwo1lCyHbH75ZB/5Awb883VSh+LcHt6jEbO+n
EuONjbTZwk6b7JmKtAWogJofhas2tn3iih6of9Gcu2JiFqKemn1nnx+bRVaYxHpwsuvwzAgvBISv
3hvq3nkiS6MIwoxv48qF8ix8kLZDrgodOKZpj50c1R3RqIdnWTmeqBUfI/Tb3eWbh0nFr4yqJ5Zl
U9ryWKmR7sWzyqlUeFPkg/8exnszlzHWGLicAIz0UhZmRrFNxP9CIS0dIXzmkWZLDJwHg4NCH57b
lCVhGCBOsMCPCxS4l343bvvpiCtrc3MCNazbk+KUO+Lk9ScymomqCaV4UJQiLyXXxMdQtdd/Ajgm
dJSN+DlRpm216fVE0fOW0WWH9NRwS8r2JR8OIKGlP8+CCwtNuIjw/cuXYWaAuNPEAFm5xC3RqazE
FMj+iOjIdhTRAl33NZKDAHIaJZXrmS/G+zBpVS7D50bCbof4Bad8ZA1LK1caDEgoO+Lj9nlxHrbI
VmjfW71OTH144s72K6sxSwSXq+drv12nx++ZTpvkkK+IQHTr4nT0HxiTvMU1N3WRUcLnIkLYyH6i
bFJAyvELt7v+iyuXo8Pdj818nCx46kZjYvRY/iclurlRTjrLsKUn/fJ1iWn9SfI9YVj7p8pepEr5
7EDRrWcw1k6UO3nJiyxSsxSGfz0MCorbU1cMecQmHhj6x0hjlaS39/GGmcbT3eLAgAe0McjeEwaq
CrUsTICQZd3Qq+6sXYXbtqc/4bwc/MlPydKH1A0g8cRnTVU1OR5b2Qfhvy8LkCObxv6wGbS7Qiw0
NNwkbKZ3XK0QEpApWeKHWiUBFWfuM7ovY4i6rni1C17JUN2CqgtobP5QaR6F1eR5xXe+JXu58Ag4
pgNrXGieYL5fT7+FDvTeNNCCFENv5zkWfUrbjp7DiROIFsZUGQOUXe8FNFw1HTReY7zIFJ1ujFBo
2FWYsNNGlCdv/6ePlqB4JBMuZCN3sh+o87+0q3jiWspp5ml/fzgliduPNy+SmqF35BJr225wBS+Q
uR4LQH7oNrn7brb9+mh6s7J25MNZem7eU4KzidhFUjU/x9QCwat8S1O76JMr4+pGtYFjzgz+rDs3
e96pTg84V01/4btd/ASlGLu8jsGXo1qUWR/E1ncWfPfLaf6H05OHteJ9OujVUMbUQcwD5LvQeE3l
eAyG03uzLS07fs83aR/bk2sbMXd2mrae2KHu/DwIgkvGOB6YhAzSgxU9V6weZ2UoiiEonalu/jwa
djnq36YEvl4xPWYAe19iNJR5pL+RUt0JCE4gg6prFzGSTaf54UyiQ+9jBzIU2wn2S4pJ9jUTJnCz
oV5pkUoAPRGZ6gagYTuAJkplR3zfv1SKYHCX4ibijGgMbE382bbjdt/gB4JBrf4hfSKqi2U5P/Xi
HF0Q8VbwmeCs/O6ltQT+inUwpkhioreWHzoYFGTrPMsE1jLH28pYsPl6xBs9b53v22yLfGfVbKSz
Ag9L4rwmhe+ILCVmztn49nT/T9Cpg4Wo0D9CHJSbkCwg/h978VDaWBIthdmCJBpnTXw3sKwoCFub
jlqGd7slbh/hb3Cubj6ZMoLruLwOiG3RZdd+zyTTKwQEZl8Uce/yBwLHDynyguWgp6prUbqLXIcg
FTJp1GC52Teyn7tKhG4m5Ld9j+r04bYUzeIn0RjBgy0QjRZR4GZAqWRxe8qBI920flk24s6VU4HC
TgsSXRdJHEkCR/vlZLSPHeLZrEELlnoNBanI4xr+DjufIPQfZWa3Axm9K5/e6swtWrt2NsyJZGSq
vYj8HvhnhSp1qUzLDi5O3qyh9c1tE0mcgg21uFxMV6R7Ax2T5Mm/Ajep6mzvABB8wZ5myz2ZGlMj
qW6luG3rvEArsCYZuZ4/W5bjCuDbpDFUL3/BU8HpOvaHImb4yoWbDT3dRNgiWZb7qHiAr96bymyq
ZNarfHa4TroZsrA3Ra+zVJGoZ1Kq8RuT1O0sl/zLVatvlZ63I10zD3QztxbwAlLE9+H3l0sgDGPN
o2CARuKJQhd+1sHsOLyEL3hUkGDa1q1RjL1R5mi3gqapHghsoT1jx+iE7llD5ZuojbB1KMYVRaaZ
pAyHFduy5T7dCglr/4FWWsuKK21ltnGoIWtMMpNC0CYj7C4ZvaPC/IOenyiiqohGMfX41/tzL7Vo
3RqCvUHyh50pNrrX2Loyt6v1/Kb25Ws+OfwzfpO46hV+aHUqkqnW1z437LZ68Z3LrjnUWeqdzNQe
hHMi0xuqKjBh/VgAXJuw6TxGBHkSjDB/dcx6eQ3Zx1JxS4LBjAeBKNvXiSzJAC51HLZ9WVyBjWIi
eX0tLXFruxsoM710O7rltVKPdLsixa2A6ov9CaiT/9shb/5AJzWi6BKoUnSvEA6yfzUElr6BCORi
7JGpArbG3GlOlpy2v8wh9DSCg/TxVt3BFCNev6sCjWmt48wEcd6yoEq3KkTUB5NYajrui/mLMEar
3XkRfmZMc+FwYkWT1r6WDqR4QnSo5sClPcb8elnxxhj2eDulCySA5R4XAaeD5cBpf1nQ4BaynmD+
w6UXxhH8fL8uw3h10NlT479exUxH+8HvmuMbkfUPn/0TOi9cl5KWsnA+wDM5Ky+Y8JGr663MzBwa
YhH2cosVpZPSVqBVgVq+Onnbn2Gdm5IajTm58szb8qPlyD9ccW84r15XVo9GQt3O4bjSod0PV3C8
MJnwfUAIhUkRSgOneuIpt4fXtmjVpWzSvycTVn0lrpN5rEVBcvvkH3dPiJBJYz0A4cDvCAQwMOvr
DQjEqYpd8bEsNSHz4H87t7XHvcySs8Xy+DyWSae17c/puZsEN8LX2uPIHOTA4wWEi/02OFzBGDKP
zbcGnTOZF3aGtMLMyd2Wh0v/uD+yJej4/QxPvKLPnk97f9JvV98iJjPNmOeD21m8tYk8LXi2J9DF
pwEtxhxylgKfcR5LusD/vCarJ4FY1Z5a5lgZOk/pH5NZ5zhJ56uA6cKohmAulDqQICeXgxpftNIf
6Bw3f4nuEPUAqiFgxEBBvYiVdwCmJZ6YUrZiya9RZYeXwTS6AM8qkfkB21UiITDwjdwHiD9ih/EQ
Ht0WHeGO4ZF++dtmK9sK8hkTXBN0YyTzKgMNZNtpu4RQsMXiHwZEQsZ3RjAPnZ/jGjWHl+h8n2Tn
WKpeVbAwCT83fpY7QHaq3QLrZHptJX2x5WzoMgc/dpCBl3aXm3wqdMl+i1eBQx/mH3P60EszvTTI
1stOtSmBAOVXaIbE4/r0mwoZOQzbMdIQKyN5Uv3IbUL7gqV0K5F4b70TfV9dESSWuAtPuvncFwcj
aPlJhcvR0LFp7iQuAZ40g29Qutcj8gnGGu0r1/Cy7kTICAcXwmYIXEXM2vCLs51eAz4cZAvVj+cX
OQ0ok6MYUXmQQeO1R1VfpNuYbmqod/FWaGNPmVR/kELczuIv/l8WpqBZPfmpdJ6MzTtnva5uIwOg
xiRrTfeoH+4K6Hei7nZp+jn4Ej6LXgk0z3488BLfDBAMz0OvjWfAgQQmGQ3RMX4tQT2RWypvi515
iH7Ocvo/lyQ/8HNB4ri5w4o97vnK8CrEOiUCiU53QS+CbIXePAWySEunTcRJvuML0iD5TgteVcD8
Rr+iPcdLR3ufH3Dx8I1yjL1Ge45xEVep5Y3IwYRqUlGJyjsXozmN+61naDUNvcaCBbjtyfuzflOy
OSMVleWfBlqXwSzDiYru+n6zri53ydIiEHT1KgT4JVNIZVmoZyPLmZI3HKGibMYAbtci23I8bK9Y
5I4uTjPXUB9Xmu/mbxcpT1sFHns9PVSfPf012F8AS0b1+DXvYFq0o+MpFzJp8laCyqlSPk8sA8So
vfbRKf2x1W9ALij1fH0/G2DFdesUeMKWu440ePJ+jB8NQmUb6/Kkw2wrIhFplSmOXUEC00yygNzH
E7T3f2U5MmwqQCsU2jSCHheg37Cd4YO8o+czDdNExKYCbLFICMxT8I/cboTtu4NcLIcD8zd4951v
sdJLC6n1aZOAuhCqbb5vH/wZoX9CJBArmauSduXX3r4NGiz4WMH25HotURXm3mqB2J1UB141ct0Z
qDCHgBsEdJQqkxPjm0ZUMPZnjyRK1Ji0cGHYCNRfpL5AqeGR10NJ4HtGC+srMGinolbokNiTsySG
L3AZmlAA6T3NXlD0iIOozmipY4B0mIemeNWVWEdnDecMFdynnHzs3ggsBBK/VGZnrf6nEgvmImRd
wEisK6UveH5IiAvk92VaX1dUGc2VNbT50U1ub4ijvm5ydNeWlWFlKip64I/u5JKqs8DxPx8NjC5i
3QmoyoqLz1+C6gtvJIvqzeimKrcPHQrwuRxyb7d0Al65q36GjeLdIYWrYDyiYZG3Ppu6llwjz62x
CycrLLu/l+uuGiEm0vuuYieSkvuViU3xgGhp1E6sGgoCjRQBnpsaILXuBbzCxWSuB5EVWEmkRFKB
HF4Q8i2GZ8E95msUE/JMfPqDelC2YKR2MQ+3jXGY2KtiaCu99jjZetL5sHjW6cqliTP3sR+Od7Ut
uwV2jMA+vRp4vU2hBeKuGBNEZSnKPDpzdEY4lrbFmKpEEaRsAu3VS6wxLZ2Q/yW4VpSCSA/ElTuI
f78yW46mjDG3OlgRpR04lYP2Pr8Q2Mk2m1lpyLMSQAt3EFevBT2X8LwhiYqfIWdT2vzq5l/vjZVx
ZrUwBvaFP8aYbiwzLS0wIysS8uuHfMgbuEFovWrpUoM8l6wPyVwkE/gLc3B4oa8S5HMJJPe9C+B7
n4UbwJWC20/SxUD0/FZbtrimDeaHOfU1gSpzGYA/+hao9uIisMDhssIS4/XTF52VWSWkX1Z8kef0
liAmdKhF7Dv5NlNIC0pNmLwZzDQBnY6e+X8qiUcYhKmJ1t3fzvmnXUt+kbJ146zsHHDqoG2DxJGM
oBYnWGEQ/zEtnHyTdB5qiZ3+X7ALB8GPOyWVozv1tx/bzH7rHsFnBKT9jTvd4Dqms2vJhUIr143j
WUECWr7W3kYEujeHFLO4ty0q7ZPVP8qactSui977ZrePMiYmYydWl+Jekb/Bt7wFYCV2UZ2ojNEg
miDrlE96zZcg+PhDhGjNfaOw2Cr/AnbfEE9AWt1FALba3ef19rMPTIxAYzdFFG9sZnRYDmZPQ/v6
v0K0oE6GvjoUieNTlCSRXGxZIObp51zh6gd0hkHtxTe/a5ZzYdlPSawlV9pD9qR4ES5rcgCWR951
OAqPuHH1KUnHDpMobY0CfWCU5kS0TT5F0Ppo3yzw0OT+NcCnGJK/TqHVnplbStHhnpG0bqqCtrK2
0o9L6Uz+QJ0MQEwqQ/XqyEhnv05BNX+sfLK3vb8xbp0UaKZd0dF/BUadNRMbP1b+gCzH3dI/h0VP
Mmh3UT5FCqeiMbeG9jTb3XRhz1isdUJCsPbfcwdi8W6Q3DJZ00a0R6L4CPwE14h8Q872OfqqF5XI
aLMfkZeMOqwofAJz6cX0xWLXiumaZwSiD0Qzv5CGxZ7yVV1qiLHxNaiMwietAH7xAnDsK4loD4Ci
e5YhPZ4SNVpnxSeSlnA0S29czhyzan78ugRDvQoBTaViYtCovpuf1ywJzRjNsdujbl79n+GKSy9a
tfHrnApWnVIveBE2dRuIoEKsxu3WoMeJtkhGMH8IYmaakvPrviKJzFtVdICiMsmDK2WNZxa4u3hJ
1tykT94q4DXQBexHUVo4PJPNy4+K0K8l7cLr8DwXhzUo0HoZw9SVXfHNkSjOK86unXXuXINI/XXh
FRW5PvqJ37Sj23F0ZuuNv+6i56nWfYAYZxD4/vjY18c7ffFkVybxg3EgkBA6HChj5d4xp4BQjxDY
pAo4+3c0ETTOLkgSpuSFU9C/vsklc4L9ZpIV61FEEYJDHQm4sa8YbfsL4lbzsqRVeuRe7XAGmLDJ
e6ZKmbXHlLqolGIyXMKu5lBZgDl1ymHCoMe3TQBSihNqrGydQigj8p8PonkzfGVrv68DruS5kPf9
tnm9XO9IyWYciA/elostyF+lIOj8vFeCsYkOXB+eM6AnFZ5PZSVplp6vBpWjz07Tlajp25uBMTvK
TTYDa4XU9/lBQpcFSrfMnprkACLqo/EJATsRVrfRKCxahek7lTJbUZtHLzEt2Bcx8OsNJ+L2hOxU
LZksnBYrLRYrxgfD8KEyk8F02SMVxEvVEGLufDAwum0LFrmfkATx4PBSKLVNgZwW0BNv/bxvE9q0
/Bi8eAHs4DY1lADelK3REYH+cEKvzB+uVPPnHZFBy3MpboInOhU7K5K6NAezYnuy+dzWwgdxm8HU
kHMRc4SFKujbXM8mD8ilm8sMoCqPgFpSrKBq3SKMDf6wtt6WpJWlZHIkjt86XKs9/bSTx7glnPf8
rgFK5hWUIIUFKJSZ2x3S/85GGe0In/RlynBuPOXG5J3znAY4V6jyXqae0KK8pHtg4bq3yZmfrGov
pg+zkNVPDOuzJcCvSyGMg5XSq6xSwHHlE7bXWOE3ifVJSnM7K+a4AZ1byozUOnf+rUpNO1usJwaE
cdHsuLpkQUCDAkfMY0jKPSG5TWUsldapKZFmIp5rp66bjM4miQgdC37ckMJ17o6kHmTbB69x05BE
ZtJEwNv0+5bvCEcsy71ucjVJAuoZJydoq9APlrWVohwZ0Qgx96ypcUPNvQDMCjX1/VP6k2hYbiiB
5gpb0Z4lG6Ll4UI3BPspLhpH17bSAnny2x1+51/TK8PCtiyKgLsuZjRX9Im5n7xVM+caz8AlyJG8
DRtUITxayQ5zd7GV8IEA9ZNGk+WKcGlWsciVnck8H8wYQLA7n8oGuf+2YTBR8rRA30gHdX+Otupq
d7ItLtVYYpNy7kyhzg3n1PVwJIivRNv/93Fibv1AYTqKrdePQuNeEf4UY51GlSVpOeyp8FaXZZ5X
ivpYmChTeELn7T2D3MFcQs8PRjD6t6mR6c05nBAxKcmdzufVO5d6Ss7XLaJemcu2V+2LOHfapb8H
Vr/6PVK+aSRbqps4ZFCjsx+oX2ERDfop+rK9lcBi3w21/I/M7b+mRDI30jgec+EFF4R7WXznFq26
QXGw33tD7M8zPhHH18Aua8IJQngSbOZFurgozdb0kArw3AODugOkPY+Z6lzedqBwGbbOFq4g8iV6
7gORSWD+gDZhU7x3RTd8nxN/mbbpyjW+g1v6F04bFZutaXaJ27u84tCNG/KJL2pfHflNEl5E+jgL
nHMUK5EWXtQQbOb0jsTuuNSxr+Wr/17t5yaqGLWNbn6FG5sAJhWZHNVupfPuDOs+jbVp6OnB9jYc
VBW27+CRGYas7r0++3AVcjXcuU79v5XV/dtwptkVnZmVQHWStSe96msSq1QBX/3/PR1ucRmhprWi
BYItjkCSQKNaZlMjVJV7Vd6HVsVvUP1KY1nnUgbHZauv5Y1Edu7XROfpSPQGERXqvvH2W5VDbKQ/
dUKYB+ePmnuX2emb1gmJd1o54tyJ2qfJJL+tIB52JqgTwrREY5HuZUbP4LofHa1NxSeQ4SQ2u9Ug
XGHFnuRxXKShLHBvtT83oDJD7nBu11E2GnHNayaygkZEfXOd/aynLkXrnkJGAfZFdlAedkpH33AI
+may6R9XEbT1I61JvqMlt3xri22zyZPgPbMEHgFfpo9YtaL7caHX/axsCyle5x/Kaq/oypr1kN7h
23FOJFDXZuwkPrz50U3vGfE3s7tIaOvkMrwr6OKCRcSPHgFPUqY/9Ouo+Abu9RtIfdzWGCEIVBeZ
qc6cDmj2oLHIQ2KWJXU99RYZjZvrudH4jcA9y4DztLtxRI3Ns762rlSZbJtt49U1w3ZmWwiBeRQE
mE8W8JegJRS4PThUsMKhx3vjhQYtzv9GLUmyMYnkXUp68vgWChQYhOQE59tYULungTAjc9dNit4z
wsgwTZXRT/fk6C+95v4RpaJLrDYx7D9TPSMRQ3TA7hELatpjswiEkwaBYNjp7FFdXN7Jvo5nDccA
y+6phPKOVyLsXLcuGvouWmwK4P//u6yDw7F76Ehs+QTU/1JezcjhzpQ6JdkdEc2wN+RP+1Xu4bHi
wg+09MoMmw45khsPa0EbevUBxFwBKurzfHUN85gZ0gY8r2zNwVeLQY/sILiH8qg81YU6IlMylLW4
M7bhaA+WRq4soWmgD6+5yZHQXhNzazKgYu+rHEStCKDNWdG0kXJwl9VGluEOZ4rLJnDRJV2Tyz/c
mQrLdezXko+uYlS6vrVWF3+/iiVoeUE/cCUx9S9xzncpTH6BNMslA3qN0o0faWl1Ckuhi4W7upuS
GKSglgJruh01DWzCAZiK+V0rGRULHIg39/wzAw63+Z0VuSLYVROTiQ8fqnXZGcNK5hq/yAItZQMs
OphfPK/G0E01UE+6STXAnqgagaN8pAkCKuJgbqyIGNajSCgZWPg3CpzfdVPrLd7NVAQKpi0DqAng
DskfozO3oUBM2IMpWma4IifOa3xNQUYRvv7sgbTVSx9uOXlZlSsKrPg2cI/E5pF5swz0jL7/OuIq
Bh2ZAoQYBMlx28hFheeeXSLv+f0hum2H1Yr+yV0b3/i3cHmPQ8d+T4bUjyPrvK9xdGJXyU1VD9xL
14Lp8VIVvVfXnJGqWNsHNwBlYqw+yVOd3cTBfaRB85RAZSxS5HFXze/sY4KxWbJ2Tqd1OV6l6jfH
rGHUPk4jLlvPOXEeqrIMi6VflURXgTwSa7vN1o4cEL3k+omdycHGyi0BExautARMdgNaUoXdNDDz
q8DWckIp9+Qsrf/ibUGrN07eGl2ZzwLq8AGYcXTdruNBN8BDcmtp16vIq9kldOuSz4TvVhT/tkpp
z4tbGq5tuWJ2yi0+Dq5DNOsR3CWuhk7gv+6r3uZ9J+1BXoHYr1UQeAciWur313RAcmTVzeIVtlmR
5um+lyCe/K/4na+5bSW7KnV1ebPLrs57VQAHzI5VOCj3KAnuMiQwoi8z1nmQQ5LGOcxLmqA7kYI3
JSVG4lsZeQCngmM3qQ0mnvAVKblqO1AH0gtY3sdGdHp+SDcMHXAEGEKJb+F5BOPvASSxeksTcBI0
41dnl8anA3GdYsGdrQAABntp+SfqVTlvg8yUHXCalik6C+ea6IKAGKChMn8/G4mgwzpiob2Pb8iz
bBkWSM1XVePSumzvLH4pEGFh1U09OaTjIcm5yxbEtW+uOCafY8uRlTbPlehGi7VTjdAE/pTf2D8B
X5yE8CoFvIErM4Y3S78gC1rDSfuM5QMZ+OdjpbfcDSB4XlF2xboqHpshACA8t0AA5PdufiK1DsAa
5Sp0vVY6eBP0UpARFAJtwwyREvqUM5zXr/5J0P3fmQ8UmtC7zKB+0BD0gwR5R1BoEBdlgiZ7lXud
q5M2MJesD1tibXoQscggkvd+kUtVEK4BBn1CgcPvA9dJYRC2IKoM/cV6HAWh4rRI/0VM+0UVc9z9
URmUqVf1a02bMzJJe89F72hp2oGfrtXeKkaC8kGetG2bS3eEGwxz/alzhMFhwggEwWZfawoTIlKT
uLbiDZpGAO5hBpUdJaV3dp918iVQzrmLJrznquLcGBPQQH3ilJM5ob1Ye0zm0MZoGrjuBLOgMuoy
scOnNm0gKpAbVzAw6iReofIBv0jDMExAMJOGy7E8ckx8WY+kCQXPS3IjBv6HhJbj3bv/+4kJV7oz
0QOcf+uvkI+J8Q0u3o7vfft/yefiPKTEJRYAgo8vZ6jwtVbfM88dX26qxbDWg0H+EeyIdliR0yqO
iWG27j5CU0/o1w194AGPhFdand8DdLJ9HdHT1s4LwywNp1wMWxKmARtKynpZUWrO58sev1A/lES+
RYDvo7dmE1WHm1P9WwkNIjxlHmiHpI8kDOzNpO14bvahCKLyrgK2eBDSe95I6A2rxeOONSpB9EGi
PBcuWAM9G40ZVHfVKb7bCTRUl7KsH3A+1fFXwVHYs7MCGossPsajdgqrFOvSK3Q49ECu2J+663CR
8lLlSIZONvkDat8ecjcYpTQkJ9qjOkxCsGvujpjwxWDUZz1kftbAQfYz7qOzQp+zaDoR3ioJYBsb
ws4xypJ9dANtqnomqK+PO76LMQ3XnmnogVLmIPd2EJGKh3l1vfcctC7VlPnAuM8udvE2QDytnD4a
3QU7qYnpzYgEQyDNhZ+yIrs+Ru4Tg/UxH45KpBhg74UaK2kncZwg6OPx5de9xfeWknbzSew+wnDa
4XEmvuojel+aWALwG4rDwBByuUJLhKxSa/PG1cQQEwK3hHGujmyamnjX9SfIrmT+mG04DbUtztON
O5PyY5F9HnIXfkAGCrNZajyztKxmQ4nXe5BGFVxFARZ1LuTWbzt1hkkOU9zvOOG0Q4zzPVnTHbOL
/a2dfIQO0kExFsJBB9k2ORb1n2UUwAddT6sTGQEN2f8aDpZi/8vkNIi4ZbgwnoO+7oIBS64L7RwF
UaUb7uk8BxFkcMt8hUuNpggnclDdC3KO3zWi7iDgTvJrFEjg86pylHkf2lYUC2ffPNCarAdxRDZR
BqrwaLCTAQjKmyVRpitvKQzQ/ox0L0d5JC4kd48d1Nd6DME+Oz4aGtbfKSIF2HvvmEqjmfksnDJD
LCSfdwI1GvxcWEYKYBBWWvgU9kU8qu8hzHvDyBKVcrJBVJYjDPXMY07r8Kr2OZOcVRAvjvUm/Pt8
6c9bB2PFD3c+JEWmKJUgU8xQ2W2uMEjH1EVeU9jY1WjQX9n9F8uM0JKXSpS74NDcr45HPd636M2Q
NLUmAQ8h8W1Bf6vWWMx8S4PmOcpEtBqdfuLl/XptfHNgRHe1FSgVIbMOZ1Rzinh4k7TU4w9K/6aA
92T2T3MCA9Yz3elMCaAQlvGpDRIrtkhHb88nCpUNDzBmYxCsCpO0S+UetHWsTaA7USC7hFxUio3t
pDybxX7TA6n+Pey79f4NYaowjf2+1dtpX40mcveCQVEjVdaiJ8m0/e5yrAUx8TT5dCneV+SR6bZM
hd+2KMigx4khUq25ws4NF64zXv6IRSskmNaIqWxvGLTmUKjeFdkPkcQR5Ct6jYNT5fmbP2XTSLZQ
k5vHpEddsReE/PN72dFXWyR1cogCmbXR3E4q+21vt/PIHJoJBjs4IXA8aonZMMMy2bfEDsBrGzoC
w8ammv1haSBIb04fBz5QnCqMzUse5Z3rvzUs03TjEosq2pihE5yGhZIdJtiA0fAZPchaD6/DvUXD
j1bFdhfPLHIoswYcQXl73RWWfFDprZh/omvuNwEqcMPtCTFmeqfXK944ETizcaaGvZYkYm3+ptYH
ITbqdHp2+kU2O/e1Lp0ePlHCw5G5yD3UADNm0FkmrYeTLuCkIZP7h/HwJeefTBtKkVyRBn+3IKeJ
4QKYPaAgVjiRU0Nhs8hf1X0pUtE8bTUFY9QvEXAnVRP7vla7FtCbty6lcJTk9dD2mtqda1ZVRyn6
csWOVunQK5LAT9/eqq7OPng8MeHjfUoIv7koix97ixG4
`protect end_protected
