`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ww1cFCaKpEaygJUT+P6Z2OD0uzJ4IJG8iyHDm5UNlVWbTWS9KXjZ9jEg11wJmlv8lA2AVebHxIas
7nZJsy/GjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gy0/aj7fr+HoqiF2MKC2DdMRffpsNgkz3LCA0LoXsy3oP+ExvEwYs55sO8KAxVdJaUPMOFr+w6Gi
VDRBmTTzMTTD1KvHQEhDppUtYnGyL/2qAWb6xHvmSHDtiAjlHews7qZ26fM0sYgNx48H6LSqgFd4
hai7P1C8/gEiLdaec30=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hi2M/LxF9qgAZzAUuc501Ws9I83yzxDz1ea90Q5QjM7jLsFrH4fLD2d0WWY2wDTdG0Ih+QNnE4S7
Oq9DybBH0zvBRUhAQoExlvdlIfU3Jr1YKpM3lLPQTLIhhCp1eQgIZljQtMN1p0u0HDYYsZO5DBeb
LZHGhmPHPWGqNQ/iLmQ+PQu0B5Cb+1VKyvK7Ipxjf6wKC/NZlztCmWzwV4WC+jY2wHB2IofyzZfo
xRBIRCIpTb+tTiKgZ9oAjPNYVjgXC51YW/c8ZhnzF0gIdh/tD6GDSX/DdrrBN7Oz/gtduYw5jR0b
WsJx7lVGCa/mgRPb2+p2mjuutW8gGGnh6+Yo4A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X16goI57idQ5Yk2jq4rj0BhsplRtdzoYr8oOU2lBTTonp1Nx4fK7AS7KgGuzY4UqvPTHmPTfD5ww
0YcXmh8hr2Hk6aIz+aWFV8C8XcReGDrBhi5Np0Vi5hozuTfEPpWuDV7kTmarku7FYKZbPt+lsAsd
f8+cIo7ySKaxPnzoHbw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RA9GWDJZOdw/NASVbYOgehelK35X4QCDpOGKLkbLHbvCU34C5eqCOlazH25KMTrAHxM2lx7+fAsw
HHb2ZWqK4pB4ww23gPcOsgxVCyXs7Dx/H6E84snPbj5EBFAp1p9GZJoguz0skOVQzCSeso4vwekP
kvLqf3Ypkz4/BbGmeIV5O3MvxWppwuIHCb+NDzDYU2x9uQ7mLUtu7pYCzPfN1FeLiv9ttZaXRuYJ
ADExpcAMpFzH3bwg6Tm6wL+J1DzA4jLGZxI9jxK+L6xNTv2NtONryX7sLla9heWPJCSHR4TT8ow3
t3QklA4V7oRFEhlMh0Nv7QVOAHjukKSZ99LumA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6000)
`protect data_block
2JEuFaTgqghMsv5lmjCzRKFTRu9v2Bd7cfnnEymmK1IpMPqqHVgKVztK8UcvkN/cLu6meLkuW+GH
jEF+IasLsTsQoEbARf7iGoWy/qxr/Wx8iI4qK11niwKvKRzj3E/VIfcoFWMI7lDjskoNrB5ON374
xdQdL472o5haNrGgEzQCs124gMoZrq6ZZftrvXJyyhHqGqmNNfQbG065CYcPsuRjXxzPltG3oMhc
7n7pQE9F5O4ObyVFgYrFINih1IyuB6ga3CPJSEZRwp7Gz0bxN4RD0DBaR3vYvY1rH6jZ2As9bin/
g6/KlClzLL3bvhOhJCW+iV79gXmGA1aOoqLtf1NI51QmIbHXkGVKhdf4Fu+qQAKs4EUswx7jWcaQ
i8Bnkz3wL35Rr3fFxj/dijlYjHEaTkmvtypTrR2ghzE1dHnqBbQgcD98qnR9ylCwFQZ0za6JJmY3
yJm/xdmOi+bcWMjXAIDxRp9aUo1rnJaow8zk/AkSPz1tDwJ1uqsh/4nhBQTnLz3UcOvmWCQ5+JO6
eMqgBwdrpDHGFxipPk+h1Vv5WGJRIJlkwrImcNrYDApl2ukdjFm9EHQHC6R9Ca+fobaGIVX65bYd
65V8ZgyZHJvXbk5HBop6v6RnwdIgyGCKyMT7Y68XMS3l9qWfOAXagtQxookF4J8prZ/x9uWxOb8F
dyLrAX4C9BisA1kyVpR8mwTLiBTnuwY3NxLpCss40iU7i8YU8NxlpJyv3jCUwy0Ppzs+GR0aAeLW
AmXpMMdQbekBmftpD4P2FSrLx7I4Vplht+sBGuS58Kk8UlYUh0IuNNxmJqj58H/bWkaAIWr4ef1P
/ETERYjzzLIf5Qww+S+AXmzZNQHUNnJ+lEY0Be9gGA6bVwoCazRHFrLI6AlG/x0EhJzWmw6WAIcQ
XYN4dGjWt+JAwDDoLhqkU994TP0wzMQtBA5vDX2nYwOr1eH+7lV8MmFKFNsA5tBuKxtq3OAFYoJn
JCnrKNFkegcUFKiXNz52yMuAWF6YC0eWRw2vtYVj6jfykEsMpAsoyUqLyR8f0/A/KlCkGyuA2V5M
2ktcdUVnNs5nGCr/4wXQC6076Gr4XOH5yrzOIwwWMtCJyTLQQET2vDMHt156eWZsAkf7JERp34bp
Ga29TJzx7NtLLL2AXhEqxgXiUHvryyadcZhrM60N9InAWVIJoHjSD7LwHJ/XQpVHK8WAiCdWs5T6
mYuS2DZyOaS+xH0dAUl+jfSdrNiC2QKQxnhDDoMfjh4+BWe/wVZza5yJVdmxN5FwdPicTDKgcanu
wsEdSBh5haSHct2eECerR39sv5g8j65VRXndSyTkbDCWTfbDaNpYrCDBn7NlLea0KyDTml8DiSDT
2TaKan/VlwXAN/62TE0KczqPW0tICaRaJ7aeWtVbhxXMBplZMk+4qzeBFFhp0RUoOoBjz8BejXyc
R0XReElWOymUmNoFU79L/s9wNGU1S6N4WXK1OT++ZZ7rNs71VKPFus6jK6TFBPFkaDDYKRmmV5rr
0kFUvjC8TgSaqJj6Wios9dLdCfjIltoKlC+4EqtXPfcL5DMt72pxaVT+HHE1M3cBmb03wRuZQUFs
U7YoQWh394CFopW0j9qfoRm9n8bLSAU6VydfVLxQPAeUhAas7MS9JTZ4va50ljVNLAv19WpU7OHi
H2ipvAqdfEC9fG583MPABwc5pJbrPuA15VDGRHwtwIAX/fDMFR5K1tgB2qukLWVOuLAYF7gJRm9P
EzTzaNbzjmrVzjL7aNETS9obGLjkNMPUA/H4i3zTffA5y9/22HvDPx51h3z91xHkvGl3NjkbqobD
37r5hvgvKCId894n2Ycef0UGDGjh2QyA6aVaoNIzbWJ3v3csl5XzDxWo58OL/HuqPtdS+4FP9STB
Z77VoKAkSozxdusECXFq02033B8TeIZFbiuTxcmDyTpUqCEV5EOcvNNcoHe936OsHkjGt2MmZ6X0
DaifvNDa20r6oY7HYhN/oSvuFHsgFvlqlBYvpR7VwQMcX4Xk4qghfj84sIxyX7Liu+N+m+aOmn3E
rEs6cXowm2XWsOVLUVWAaEtD7iXD5c36f/Xpj3IIE6p3UuLdiczNoXeyr7BZ18gvfxOTavmDT6CE
PwK20cwFSh9/AucsyOPj7BRCnaWQvhGIWzIth6WzA4SKvjtF5c/YMhSOq2ESMyd00w/ULlrTxXpl
Tavj++iTHbCExHJlPguMkVH50qYZv/ix5EdDNqfqSBa2jsWucQm+K+XyMbq6BR5hBd1Xhb0oQUDT
xb9pOcEb/fXT9tZRSsC2aoDa9nyk19jSMDD8e6e3iLcdIwrZTmWzZ1Q5VBLUUbmtzgGDmH67QJFw
EHaKF7uH6bLcJTxHlXpPNmEwRRE9uWa+sc0LiDEw3B3A3TIHcySKM1lqChuo7Snrs1MNnFgfYplN
fWJLAHjGL3ycfAjU+aJ9wY0mC2e1RL6hkGv4jfEHiBx4LURIkvbHSJbHJD9t8DYZsNAMWYWQQl07
vLJ58pmkIdTEOl5wPdakl0O3iYYB2dUW22ZOcoHbU8JyP2NQlMPXhjwcjSlpP9RtQZgSvOedqPRS
q+3WhNNtwSLnyHu/oY68bGLv1+fudD9lq9+lkQPJSv12D6zaP9ww73zlxodGBiKVyrxHCpopSAZ6
efUDe9fV5lMqe652qWs8ZM7sTYnkHjpbD34/CcpyE5bCBWVZkoaUbKXSpDkFnFQ8idFQAdNb/Op0
xbZpo/XBzusupiijalqqYGlAKzrPZbREEQMLDA2G/2hGHZCsga3XTh6+5aH/YU7uZmA4yOpKrQe3
Ub5Hmr5Fu9jk8aNNSmA+PmgvTGIf5/WonPvfLEMxL8X9dYKAFDOC/P1ZZWPfhEw19F4eNv9FEth3
xEXbRwY0OpGmoHQQnnDYe0Od4CuGj5HesOaoequrgEQ1/paYKORMxI/yhDmXqCLCBlL9AQk6kUI+
/4XahdosiOavbQumk6kCde5jPtvEcPMPU+LCECgWRImekOYIt49ekZWi+fSrf+SEL+T/SCqQYQAZ
pl0I9rNfKM8vDkt06Tkyi5SYj0jvNN18zUy/X3MdZChmFJowRtucOj5Qo3NSxA6/IA0CbrhZwX5+
VaVgVXZChU5XdxunagFWVoOuNW0XuTPzWJ6fTrpxXsEFxHRj+qis8SxGcCdB0TU8SZ0IbpaZ4MDG
IFHiU03uocFtaNKY1LKgZaTSvJZGgDD4+ESeyz0klK261Y3e7cyRA3LFEVpgF3rjifY7/jQr4/O/
z1Bvd7LknqUIbq81Sn/ZJIhjI34qZEDQDr90s/7FxTt232PuFhfk2BilnSPDziNgTjhFf0798fk1
GzKdoJBbjQzjGuyJRpRaCi0JdbfyQq9jnRQmvZZaPmkQYxbzUjMX79FTrIsTaMniUKReXlArKErM
5XmwBv9m8OfTS6UCehvlPv+CwH10S8yBp9suWuGDb5BrqWZ4fVaj2dihwRxnHYuHdbVFwQB69ExB
+MDpErKefYEyIjziw1MNQ4hJmPXtym9yGMGicsm5ufWhKMPIPjOxPM0E1XsIbrb8KH/otnXaInfz
BAeRdWktPvOYLitKs7Y7zoXU77kApN3v6x6F4gw5MwcooEhwPfRS2D2V1ySDbujrQjis6KiUqm7y
zj0ZWdUywhROSLKf6CP+D7MDjRprfwTjiRDLvdtyL06zyGbgTrQMJiZO5+VQ8NNLkVWcrkzG1H4J
sbZpMsFGBw6m3pUcq2zWnFfEzlhbRTgDfLDRC7RNtT3WabKlbRKKLoqwTj6YjaCfLec5QZ0xpRU2
8KkAvO9L5iQezWySvPeJDU+I7ubJfL9edvOpF4EydO8ag3q3ERRHtaJw0WN8Wx1YH8CNhyNsFHwg
PNzu7c9hcBzECfvhjCgJeuUYAuIiaVqWlCg9JgM7uC3RMWmzAWRfkpMQg94k4Dvs+sKvFskUural
wv38reXI5kSat6kDcWjWz09gA0H3cs63a53ndxhSeBF6PxC3u98U/a3jp+SS8waJcXVT1RnZkZlW
go9m7FHq+Yz4Md4gLG+ckL7F9XMRgdVzHFquz43o38z0nw7c9SMoaFTsyDY4Z6ZfYeUNfCy+9a11
uwgar64ZmU9z+iIPi78OVPNQqlL0Pc5a7xjh3NbuBg6KnIleQQ2R78qY2q4zXoxAIChap8sjWjit
YUBcg4HbQ9VfJPfbM/XDNmyz8mN51H579RJA03A8/6y9hHEXo+SZP9KNb90bIu1Vwy8NprbG61O9
Gu5275vk6/kkqUQCVntqu4fJl3NQqzan/OcRJtrUjMsILcRmkEKgBogXke29TQV5vtgwwfqshDjK
z5kyCW+EDJHMlCmczm/w7BQJudBPkIM73ewvfnIjFb641boavoFwY65Mgaga/4vOrNJ6kTP2o50C
I/k5O656g0DqHWc4/4pnP5BNQYlT9eq7OzjVOYFueJeDQYjXsmXhlkztHigFLl28Viq64xdz6YvV
z6YHLaNpcfOEtdnx7s8mc/HbCYlGEY4w0OPkEHoqQYSlmGljuf7522EJZV+XUeGfiut7PL3XEKVi
sbVJeLfxy53yyEx3smLRyLVxY+NPkfkcQYBP6r4eNSe+dsOxE7KxyBQQZ55TviWNQ3NIqPNkeo3U
jRrzKLfwE229vpm5TVyqgsKhtB+JEGsiHu5Ko0zxF8xlZ30bx55FQFl085ZS085Sq4K9mwe0Y4gW
oy3/Qkit+otjteBKKijJA0kDn0uvzDMj8L0v57KUhQa+jShQu5Dc63UBATr4dXnXz+tN+2U7W86Y
Us3YD3uoPRt/RSiGZMrazRLm67QVgeMD0sV+AqvT766anTQgPmqmHe2zBfrsNQFIxy17vutjgYWb
83okrMWiDrPNstvD60/nH0h26zmq12Ith9RbUfwE1xNl/TZr+GNzLtFLxAl1URhg9kf7EDD4JP/B
eJ3WE8cX8rj80D9L+CDnXuxBN5xiNRUdoli376p/H2dJVDnGcMmRjeWKjqdyr8YA32sU09GJm14H
InoahXpYLLzEu/Kzi16cQq0vX6diZjBLD/JzLyF0A6rRg2n9Hn9/YL/fJclCOztfinhS8oehLbNq
r/89fnY+hxjN65M6XK9G5UVhwntGW3Gmux0lAkvQqltAZQN/gv+43HnzgYpzATDX2OeAhAZh3XTO
N9NePGy61iFKf1zBs2L00KrdUcxhlQQC7OSTesJHGk++715Q/MwNvwntgIWZuz6b7JuMw9Jo6iOj
nd9hOBBI9WZhS4WUyH237XaYEvXgboh9FakhRHyYXimJvWZIzhBNiUp9i9qxCbg/KB2++R4quSm6
Vh/FnsvBd/lwWsYPhh/u0CGnvtEEY3JP4mG2C6qt/V9bwDDaqeOKqdT5gxCcxaJT1wyjEqpsmjxL
AzL8kOCkPvKLUze8/zeIusmH9XS55sQLzsIjgR94ckvTSCqwNc3xqulX5w1hpNhXUjqXIQ0/nni2
ep+nPiugNyJYdxv7131Lcz+f041vjhEm/GhWqNd8v9aA6cdcF8XJO45rJ8UafPQO89Ba8Zg27IV+
87KaBLDaS4VpysLXm6rZ7fZ6GgPYoGv+98o7SQBd6GANUFgt4uub34YycTTHdKGr70uOA6/qUoZv
yZsAAhlZ5rF1BD5QbjUBLEk2YevJhqEAf0gZM1NxIUM5R6v/wY5S2Yc5qWLvM5BeQqjtB/XTrT/o
eWbzOkFHhhMeIZdZkDgw9nUAZWUNkJcCzxkDByX2RJG432DfF9eJG1Ex+F/YXigbJoNnmnEaIjXd
y8AcXC/it9gmNnFgHryvNIviQSIoUk7zhIf8FOLBS/OKBZTlDRIpr9Mu6W/nyhdpwsgZC7WX7YmT
DL2leQhBcQqWWSrxl0ttQ6WY5WUD4ce4FZaybxn4U2KcENy0hVgBTMGe4cBAKUr+BnsieKQR7iHc
1Re2IO3MR3HVHj2IVqHb4sUIcQ1/mHgpkcwk7qtyCPHQVYmvae+YlGRZ+bDQ/OJ3wtYtqGcnqYwF
Uwh5hsjhLeuxelslIgt5xi1AGGtWGMq1p1nxZkALDtnd0rPsmdvmr9OZWC6fWeHCCLMbLr+uGdFk
Eusi41aC1C0tMKaI6KFwpc8Q4cwTKUF5IoKdEECcxzs6GpQpITDC/FizcqeuxyBLFAojkUY99QeM
Zh7n3BUckymhRsaMLR+7avSCR8bDjhWH0klWdRUQch7Rb0rantlvMhyvInjycxxZ3u1Fc+TohNc3
0q18jleTtAC3yR/y3BqcDK7vQasd+sbyl3H4WOx4KskjVD+wyEwMl2d+W/Z+81ZECwnnCaT5KXEE
XbwLQsKGQpS1PxCDUeycRmg0hbXvfjZvkJ5Q9PE/nyUKW5Th+Yo8hUnW/YqylA0TqPxfFxlh5jqk
9G0NAHxDYY3lN2OqaOj8zdRoWViHafWCn0BIqMOV2ndqTE7AaJiW5ZdIa/WTZHbM6qgpdaTAZAiU
eEYY0k1+KxmXjH0P40O4Njkyy9A0GRzqN3uRW7HQvSH8Z2pw328J+ARBuG7ow1qEyoA35nQXyQwU
UQJL5uFsz94DDeVpvEwFZRzKyMuc6b+wv5CmIv/a6CLIIPGWEn6a/Fhv1xAc92eYj5bf1jXH31o0
T7V3QGAJaUBDJuqaO1pc34DaFk6S6Nou2Xs3EKLpw7BdkuRVvPy4LMDvD+Db5KEj8oL4W4Gv16jM
eBWAjv3jdaJZpkOnBYTPI4HQ23To22HFVRqyqBxrioBmhKXFyzTrjQQdhjP8JsbAkC8Cb0ojZH8E
2w+xQAaKWGxFBZoNfUXoMLqo1O2dPT5HpfoyvVUa8dXA5E6hxonZBU7q7PJy4wCvc9rpBeR3XAFW
hidMAt2r7RdVryvtNHmp0kVYTsAYfbT+bAjoizB+4bvsvO7Zg/Oj5k/QZNkGgIPd8Lcn9LWzadY/
UqQtepNp3Wk5Fq4zmIxN2AV3sSDK8xPTcWBRs8yERYIJ576SvNhqGy6XeMoYRCq8/W4191u94Asy
9yw4jWQMG87dIjblCbXrfYx1/KtYBKeBcNCY8k9q2nIQvOVCIzErVL3zz66NYeCJz/Nx8+xawoM5
gBwhTvMDQhahbolqgP6Fi0utd6ZZt+5Bu3g+0SfmFf1DjGpKOzslp6Gu8exC0miMCe0iRp0ZVXE7
gDtNdc3wyIdLDqjJlx+Ss2BwW02dHPsZaxC0bmADESlZfIwFRcVnE5arsGNSybFtaR+xzJqIE2TE
b3oaDy9+pW6QDxfeQZl3REpmzEiMHZOBF2D/jygvxHOxv317Tbmb2i+1+4GLxpCGh/4FwUAqCdam
uSK4fuhOB+mFyzWnsnzOpbg9h4hMMggGY7G4Bt0Tmig4b9pld1k3loM8ukrdTkvjFzePFWrEsCUr
TvUrGksivt0ApzTbtRfQzH/8gQVpzTB0gP56feFRij9aowQvXx5fWyryAkN2w5eH6L5KXuZsOWmD
rPJeDa5QtrhWyrOHQyh3pNRMtOh+JiOONY0jBENJOy4986lECZ0ia1W4BLppf3c6DPhRg4dVxpfz
/8lV0T0mehty/uLM2zQP4GOKjqkyE/XNIxEUo9NPiCkAOrU+rYnM/JJKVcNbCZy27vWA0ZGqT6ib
UIejQz2L18GouIC2dtB+5P9ZdUB7yPVpFM/NqblNkJO8l8j1PJVy2x3FGcPnFSlDU4B/yXDmNphu
71rIaanMQACbbhMwt2WLK48MpYEvRy1Nm/GjJFFZWOf9OamII8F6HhPnV/V8pMWg9nbR/i51T/5B
INLxL/WD8e4lpFPcZjZc02m+12FPUreCj9ie6re7IQF49IZNY64/8vkhhG536LFa0noV86OV6yqs
SNAL1AS63keZSyQaLXbrK1gcWAl0ZO8r/B3CWEEdHhekrpw1PFQ9UOso/B2ab4BMGemy4oL/TYLO
HTs+u/PSwBl9rBLeBGetcOr5IXpNNhKjhN7/SUNQio/Hxm+Lsj3twhYD/QM5P+VsTnuVrsxnULF4
lz90xmMmhuVMvj74wE7I
`protect end_protected
