`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9920)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/Y3
LeD+qw2K3LM++tksXDWlRgF/znF+Jw9c2JQAPXKM9TKRvOl/czmCOhE3aNSoCh1FUwlKG7QK7XW5
1i+Y/6fuS/CW01hotPrez34/+2hYr87se6GBDorysLqVAXMsLY/YV9B7HhDUSw8jyNyknIEmI3U7
WudHo8vhLWlCkMQkDcMf+Ivoy8TEGZRjbwDtOXoE24Tpyh0y7Szqp8vQqEDariMqKoVn6oTmJYLq
2DpWhIEswln6tRI/+zBSleCqwfAdmXyYA/Icw782kOJqC1rm3rVrW/fPVK8K9QJVLjxlLtCOUsdW
MXHfW8zBcf+OJ6M5Ps5WfxcGaSo9F93JhZJwtp16qQc943Z5uL5S7F6uhx2/2/JNEiZKR4nwO6YF
9lApKneiqiV4lMknv2GfPf3Z0yt/epCJ1D6rwzHUxOS1WE+QGHCe4rtK8iJJPU8gdqWBAV0E38zX
DrRSC8OcTDpaHRsM4h45UtUZ7QHuncOnjyjfle45UXlGJHuJmqtQtKoBHlkWLaWs8IxPTRJdashu
kUk0S37b7qinz8QPzVNDizIo7tt1mrqBCLYTAlFjqwSpg+Q2GoQNpEbhhjJSmvYKPuGddRJZO7Wl
OSphxyLgZzVvmxDSH/t87kHgGHsFgjp9dviohojl/U/zWNmgRey6ALjcz02ZkQE6vzh/zBsU36oI
1XLzZdPOsmsFTW+hi0YtW4QXrws+XJn0lDvqAm7a/4zSUan/YXPqgWJAp0UJnu6AAEQbDjLTTbka
rmLtzTc+KBM7Qh/MrR0nLXOt+vB6+4vpyFW6VF57FxmXcsdwTMv34b7IGNAHXV19xTd61xcwO0FS
hYiDkPuuZYyI4HEIp4JXLUgW5zvyHVNvmOFASRRNUBRiTkDYHnHp7Z/O4tBKX1n17fF6v/fg3mwS
2JeiK4If3PXvktkxXJaPGyiZmPmt5A4Bthy7HLbet//JHNLV38xyJ74gKq7QU9oEASiPXGEAhbM/
x9I7SkQ7MIJFc8uqyxac3MnFNurIiDEeYdHyaMERPao3PN6xhb/2oFOdOfTFP1ukLGNEUsk0hPd1
LgkUtfW5A20Gbm2UqEhuCsZlhhN713pRuj/0GuH8RmIBQvAjd/LXyOWfuP01wImCTKOjz7332xEc
vYTB2ZLyx0dZNiESt3YthzquQ30BRv2JZ/yMS2L3RICN8EY6volLZIQ9J/ZWNZnto43SN9PZ1A4d
KcVhHcitoNxEjWlorIlUHZeWcgjrKzRKTms/5Qvq+XK9VFq4xnGh7Oac9iup4UOYCOq/mhqKA4j2
JlpoYNdiV2q/qk1GYiR9lF2o5Ecimhm4F6Qr/f/9tQ8wUUD6qfkiHSEpOGq0Z+43W/6hQ3pmdtRH
CP6CKYahbYpyAC5P664kR3KSyU3BSn/mcTnKBa/6NWGyfV/dwudwQZYVTSGWPphViyNhg4NXBZdW
VpNjfiNyjHV/WD/NL12VW2Cc1vUJznM7Ohc7WOPoxL3rTVqMbdkgPi1PL7rVXfy3t8gZU9LEOkRW
PzJtI3ekd0GtH6hpTLnCd4KmXpUwUPsqehrqFsbkKH7YNuki4EFBpsExEHrPqDWOzpH/kcA6Kdrc
YH3a3yqe7rPGOTbbq8kMXtkWN+YItZVlgy9BxRaEYkXkPwPE5k9IeceOrVP1c98Iv+echFZLGGt9
j0QBJm/V8zqFl/WSHqF+eE2suXsp689eqNMH9JYhg2llYDoxhhS7WHFNPfDyoEWMj1/FlOG8ECsl
8hbPn81Rxh9ZGPDmnWU1rLYxp70uYzLoDW9knjjlU7YCZd0swAJvYRhXsXf3VpO1kz3iv6W+nZMX
Brg1+/LfOSXBphl/YIzzMLzLBGrPVYuVX6U60QduJlfeyJj/jsupLa0YCq10Y7+A2WSQXESFHfnp
Oo1bNau5NhQE2DlB0tGBKT9+EPIslfIrUiX61m6Dkfx7lrqNHGsqror8LWJv4D6YsANdMsKop3y8
ywyUOABWxCDeC4c0Mvj7ZXbQ7mSXzmcBcrunwbWP74A7PloqWvI7iteJV7lKc7ctjR9u2w96DihV
W/DwvdUVHlOVlxCx01PJRop9W1LKbTZpY/0ZzTe7UocPsy/89bc9AcwM4aV8BP8oa3Tq0MJrZOMO
mP8yNtdJbBItrltMSYPKOFrGF8h5Z9v2p0WPw/sstYnkE2z48Rw+6hSemnVMd0wzek9T/E1AS1oE
ZrA3f8QL4jIonmJyBqQNSc2KVR9ezwV6djyk6MGEmqbDiHCADFai9EZ365ggEep82nSHyOwH7e7k
WAk5TUhv+Z/kHNdp52dLfVakxOtEHSbneCdm8hkeGJ7HytHDkfG0EsgZqwM5A1W/2scrmPjhfeMq
Z5gZil+FLHuqDgpnlqk6GwlHJoOLR6TnOa32UQ4VybJP9TMmBagp/su2C8/eaMBKHBuRVk39v7FX
8dhO0ZLg26Y43Dp/r3gPiA1p/bUv+HokNtQflnLHrnfgcNwAFuo4ChGQr1suF+/6MEZ39+YYcLQX
aZIHry63MB6k2POVKN1jUp6i5HvsZkxmE+SYqfeSDdTzqzoy3kdlF3NsS9UON2EiPWysa2Qu1opo
tMApEFghS37Yp1yaPg80jFeZRC2laiYChE9ZVjVUsteBxyUf277ypkGtcghPr72TPqQ1zQtbODEV
01nBZ4KzeBhaYwC0n8+Xh271Ug+NcvgaVLmitcZexDBHRfooei8SXKptlrX0Oj+5f74mAi29Jmga
Yl+J4Ze7y68N+bzIJgr5GmTFfbhcQWOQtM+BOeiDagj3eW0qeSPaLziyW5Otu/hbEIob2UQETk1p
onrFt1MwZK1hw3fcZGOjClWT219Jhfuyy3lsb9z/1Y0t7kkhyoXH0NKDKRuDurkJ0bKhY+0GCyGQ
H38L1GYASu7gN5ku/Zk7VkFeHIldz1l6oisOIKm7UGg0hicb5B93f2Pf12QemWqxMQgJ63mSrLMV
boU5NveNGoLsYDtDnaV2YNF+CNcyA/sJMBZrLAgN/9Y9uAUXs3U4HPLd5x0+voXUhAbX4JvYJBIt
lCVF1LiQZRVoZ0CoPFcTPy0oqZf5t/B0waoz6o3QOXzVHLjS+SJmInj4IqzXOmBxM6t77U7iDZIz
n9W3Sa7sPbZyUkMw3waxCzEA5FoNts2Qa8bPOznr0I2KUnvgB4Ks4TFz+sZXvm70ikvhmrkvcD+9
PIqsrhbfBFUMcppQi1BDycK8k8r7oyqFv+lu1E273cnxUMf1PdmyqY0tFJKKB/jfUqQcGsELlXXV
yzrsMKGF94UB4/QnS3rY/2JXj3fytLs1iF3gUrveswOcn5JRuk4jkfrwG+M8pxQWsZtGdzr0TT+1
uqrfVl0vXB9nRt1lhce7cuSXcGYznYPX3mJaANlLWK0B6dwQWGiWY/xuGAOiuXOaCv71+cvOYZdD
lJM+qFIn9YBJdwpvt2Hun2nkGsOSFdBwByRfNVvTI6jaypdQFI63IrcLWto2k15bYYO7K/iTUR3z
ngVJxLuJWl8b5nNHQ0dG/ioODLmf2kaI9xN1cML/3Anqgga6jZYCNbos7d+Wjqh4+db5a0ubk7Ro
xwU7SDAodPMySyOmYYlN9UcmAOlK5r1U14y+glvLgs1edeo+Xxhn0vxSmZmkIrp87ejZtfairDa1
xriSIc5ED1Cx3dWjBsKyIc7Ix7PX30AazNCAu7XXemheQiCfMwX1ntAE+9HBr+4Sab9vWIUMQQC9
dlo24dQu0w7V3nUV932Nsda8phb9htz2td61TaTuOJzfaTCrY/OT2HBt8HR+rp6FTk+48LL2aNT2
EDnWQZayhdCP0WyMUXKgnvWCeYeMDzw+oEjKWOVB0bhgKHiV+B+VIvab/nFNghGfzEZPegRWEOAs
ckW9pi0WLKtIrwdvpp8uDh31ZDOQo2MBGlNU07AS4pXA+737z2r1v/L9D7fY8rMKrjh9FVF8L/Cl
3eZn5lWjtajpEZoQl0UOXLJpa8TlxU1qLZYR9Ojlr0sJBckeviGYXxgXQohGzgwBOH+FxicQgubT
wZtx2xRb8X95GAh9M1U23B3KobRfVG/j/2exYCdBrcxe7KUoFSNrD+tS157g15d9xR079V4BIgqC
xZy7geMeD6mrBwo4PM3ehNG7L+6EIsk2o6jdxrmQfZzmHYBfu09fWiWuU8+xvYsIOF6rgI2cE6xc
BZXsbskAQFkq6xlQidmSPyqK2S9Vtx5mfsNYCjIw6ESaBsGr6MPEFoTMNWbuou8OBGqXE2VmDIde
Hk7G8wLlaFn3s4D6JIao6hBjw7/V/KDTbvu7LQ3YX2GD+tb+ZdpMTo0JClb3pvD5x32psO6hGbkj
TS047xqNKeeSuNg7JZ5LIr3hAeV1HEc1sjnougW/rjM4OM86jrhtDnzoHhJZemkDvHLCawsPM0G1
cjRUzZLFMdLxVSxqNfR7krmQAOifZLFEdKSXDjVfa6pIQhjkArOT8MzOeBci5uE95nQTaT+Cg2FF
Py99D7prUlOY4CoqYRvWT0Sm7Z7Hts0OFupTcZ/1XIVTR5FqtTSml9NXZfnD67FawArRMVZBKrAf
46PPapa9QLxoRLzsb98BbCe6QfTCWWEjHlEZ16L3mOYQxku8aM1Ya28K2VZ2lO5pykOghRkOgbyR
HdYbiZOrq8Pkx4Z96mafAplxTJeDjxtsZksBDl7VXb1MWqnPdJGY/7HhJgkkEEM3RbEQO/dHJrIo
0qdIx684gpJvWIPWO7ajLEqFj8bGvRz/v2Np9Ure5x+uN1bRUG72/8M539bF42d5xmaCX8VgKk26
EwhCKGOgMH+aeLCHn2l2XVpSdC+3zBTZUT0QZsXaWmterd9WrvjcvmKPMMOdtG3qzrfI5X+cYfZ9
iug6yj8Vfj3w3lOkUAhim5QYuyY7ZylHqPu7DTrgSkVZmstOsQaL3thEnef/R8oOW9kxItzRfqcr
BvOgicP4UIkPNtzYFA+vXwErYG6Utpd3gDMLuCUoVA2/UrI5XYgT4/SJ5F5ne6+kWxruzonvAe3a
ij4h2B3WJbYhj6z+EE/bCaTm/U+YuXtcd9q28okYqL6dRODH5IYP/aOZXhpcXDpUwu4TdEfce8hm
Gm9ydS1bWfoCJtmtpK8Sp6ADs2hpnzNCR8GL53tvxpdhKWR9NX3TenWFKfZsturfKwEFZV1LqGI1
v8WWAv5xQGv9YkjgnywGiUViu7mwR07y8dU2wHivJl2p6+nSuqD77IxP0ROz9Tc1m3kAvttNcR1F
cde4Acg+/1oPgeIFUwSYkpMFwHK/z0PdBr/z83hRaOw5jfXkfruOqg6hBUDaISyAvz4hamN/y/qE
6nu3x6hXWVuXCANA2iZk5mn3aMtmkI9xSo4ph+ir3rw7PDJ9JutePvmb1IFDyhjT5FhQfCAK7xHw
+8zmbPk654KnjAhCg3tYWkE/yhHp0VKxL84VQtqfSVdG6Xaf1jsdYhgD+nxfNgCA6yLabpebk9Kg
g0emdp4UbVgm/pMjfwHDorO3evtZlh+qcc9Fkah6o3X/EPDQfXUn9aWmXwteS6Z5stV8HERrs1pa
Dp+tPrMxNoS+oXw1DH5Ld8LFSAWsXU3fVhutbPwqDRmR3hN42sy7A1B6HzUSZE/P4tVSAfUGbcf2
1C/Y34+ZfcjVNtTMy/IW8oN1wWnXm6gyqfToMmeIFYEsap4xlcVF6pqLw9m7efLjUNrhQZJ/nwAA
5LQrmsCzNbbChG6pEgyF0kqYgDKXT8XfgLQ5Ot1vtbYcrFJDF6Z2S2c5ZlkEKy9cwUKW3AyivWza
5PopBEPq2epqpPikJDwv2CLY/pCR2PEeT4BaIBg1JVRZpiJzDGqs2yhVTS+ZopENlAsrKYPYgAqu
a8T4MNJt1p0sDLhUQR6Hr4yDrYRcKKEA0yNzss6cN8RA8BfhSSOOMjG+Pdz/u5EL9wlNFo9EauXJ
C63hoTOjobLLhbLulOrAAYSsmyfOpW47j2Uw06wuuGy3419RqWdTFckJWCYEBl+g5w9sIjngqp5O
dKPydRC0L2R8JQmdqBkr/Ti+OxJRyE4Gtfz9d65V/YZXqLpUSn3pET4gwXzabBpqEKXyYlNj1ABy
jT7SQzBuKyTGwu745cO6nkr6yy0zca5nvOZseS+EivcEs0Mapks9+HGO6vxwl5cHN2t88ga2pz6H
9SaEBleWNJ8uUSEt9LUvV3hp1qkTVpB/QjGkl+wPdCPfKeAg1Jo061pwdfntkcocDFin/ntEqc5V
/l8Q2T0M/xaF5f/AHw9fkKZeNew3C7ufLkFmkL4jBhQYKfZg7CM2K5SCUvpzboryiAejDrZi+WR2
1yE02XSG5n2NiEerrXbOXjsH9gbyRF8qQtMqWYq+L9lTgFLiLQE9Hefth/iv6DbOchoD3xp9w3v0
6LsCFM7bcKiGZdfXTBfuH4vmJyhWocRaIgdSo9pyhDOsyU3ZY7j4Oamed/T0wRIYlIQTeCgULIIF
bYtepZpxBbNyluZ0na3yGjGTyX9a2bCrPyUk4c++ZmQeJZbcUtnVi3B91k8FynHcINgTqaBJI4bz
bbakkGo0KdXBzBnOmlp4vqHded774VhBKWUv++Lo7r6VmRSdv+Jr5RITXNwD9dPBQPsHhRXl24H/
zJqyvvH5Kyv+149X/WdfmjGNMYJLeMGOPwqYakRqsZ2F9SSTUsVBAVHHouNSSqfG32NNFLp7S+1+
wkVIfuispfN5KiZs6FgW9KVE41M0Erky7icPs2EgSM8KfLDLmDGhsaMWVv9WMXe5+GlFJHXwPydd
GXSxTB/uM8XnZG9fLQIz2Wu6HESMH4GVTrI+ve9diaCPa90gkctM68fHPSaREAOkLCgpF4fCDiGb
EQICv9qnmZPyEsbzrEcz6r9mSW5AO9cz+gjgKBK9To13mIsrMEA1UZVeagRHLg5RcS8Ems7Mt1r1
ZiME6Y4KA7wn+//pZojTOSaCFXOFgb6Pyii+eE66lBY5gl7VfGuWfhfcvREOmDpD9Giz+twVqyqX
DtNx/4OeU4KcEYDcJf05kCAWoYYWcli3aNv9Uh0HKmlFLK0HIF1HKXViCSC1Ru/Pglw4MyxgmIDO
XXYZSUtD+WfTZ1pRXYqtI/NKrKAh52HDY9EWLXrZjmVD/U9aN/SCO23aZXJDRzpvVNDVnr8cVE6D
sov6vCT4PxW8jmjuSplXWmZhm5Bh35aL8lfHXCKRY07ototIohRXUPlS3wXiwoanyQFS7wijm7ph
7uNmhAOldUSsKPRSiJrW1paVJJUtm3WNDpnARBBpADLgJF3WfvPR63G9PJmeD3rGXz9rW9gg2ctN
y0GjOFll+2EgXLJ5GiNVGpRX+Evfqf5phLrPP/vatmJk44l7XW4XEbEVUTbRzbe20JA6o/cULMo6
JSTD9963BAPJZdx4CySRCvMNu7mJmHLlyIlVFqr9IijgiiiJeZweuWzciwLuJk6/PvpcCcow9j5g
eShrbljW0R6vEwrV9oI0BX/POPvZcBDg9IqCJZNdjbz7RZqFhBUEB9bBjrF06afH7yXoGSAxupiS
E7Ms5+JLh7BplWKjNGZ636Pcc0xTcWPUA6neVANxkdsxvOP0tRw8D29oO3qhAbY6IIY3P5+2Wort
P8h1QRI8OKU30yO0FGIJ0b/EYVxrLAp1QSpufK7MljE7tErLJPtrvYoGcM/XfVi+aGBCwNHiR0ND
3xie8kOGaQ7eDi1w6zvYz0W8XwzUrfhU9sDgR/9iZF/Fd6NjKNErEsksCIBgYDe8hqFeGce74aFr
2XyYAC0aVHDbeaedfETG7CZf2pCocneIo6jMXrvhlW4737oq8AuHyKkfDYLY4wrerGTSrWYAzUJB
J9RDawaQGqHwXntve4qTT/z2JPuIDHrARqIi9jOnN2JPkt34Iudjq9QN4/YbHofVnVPhpkc2/0/+
v5Nw0/M3SXDfcXhuok+0wQO28UvW/ekGRJBfhluGbLd+SX41oawYNqAA0YCFEb1yp2rfwRRDUun2
b6sNXzrQTbzWBShSjeq0wZZu/sgmDrB+FaLfEQDenbUoaZR45fbAO1Ws60n7kINxoNAQq73GSyTa
3vVPG/l1DeUjiEDiHskh5qWpOKELcG6xY5bF1uyEL7JaNpfHV8+PnFyj68MsCJPuXo4GpOBBAFl0
U287fvvyTFcXvnl+t5Jo7IfFA8QDLEIRA54n/3c0kCTNWX9fmfxtZOw9Wnt7ISnT1GSEpwCkh2K7
K+fuq/PXKvQf4Wqrd5Aq9gwLT1N9sf1KopmHyrGzqG8MFzKzO/ns5wEqfGqqTGv+jLSBfFGkcdV/
Hyockyz3uJbVPBF0qzGX62DnYDN1ukAVRmtXqcLL95xNvHRoxdHG89yEtZxo0BbZdGX/qAe44F3G
S4g+TRTWgTWNcOQly0M53u1B6+xIc0mFPOhPFPf/21GQOzBMKLCqwnAXvKwMfqSVF9hfvujaLUsW
86w8MhjFHYg4eMy8KqLM3Y8SNz3mPCHkpEoW44JjY2mMNdggKu3rOmksdcpCByyPwi9iObe2IHNy
LylpOad3XEg93QvuKtLFkQ5WcvkBFuGPMbPArEi0d7pnKGfvUyKDMzho9LJ8ixLnNhDEGteTPCYp
f64PKjSeEomIyZki4M+iMIKA2MQKa6vKmtci7HrVhKFPI/UZSVRdBDV6C2As/iy/MXbOJ2oWWtCq
ODI1U/zyUbeJR7rojAN3AUsgOozFwLF94L4IXVr7w4MP2B1bmcaqf+IqX0K8u9I7RbvqYsiTrqpy
HfGhC1ubMzescZZ+pT0qf0Q6YK75/8wK0etVBLmAADQdG63yKC42l/A6+BOIz6sJT+qR23LOl+lZ
svdZh7Zw94XDR1PCDdM6vKvPGn187IWTooq8fveH9ATA+7n4mnHxXrEEBHtkLGnurJTvmFM/Ubwy
V1g146Gx/w6LyOjrxRRPCOA2baENH4N7dlKwSf4cwQtz+EYphhrNNFmJyEPtgCU413I1FClOnwAt
ODBW7KzhDXwdzMGnS1tHXUby6tAjhltZFasl4gygyvP0ct//aYcDaVVbPSp40DWKJbmlaBSwfxsh
5+4/Dfj344poCQVgb3qXvD5r6jcCQUdQtJgR2YO6Fsb8OKdO4eR1a/fdBarjWJAp/e8xHIcC0uaU
waUiWocL1um8FAAD7gyN4RPIGSzlaha+GXKl4k8ccx99JPDPI4qQrtkzzzEkkwM74IJG7DqFrG72
+sYtsWKLb5Hz5I5TObuwetNT72xHWbWBJIrnMcaLhR6BU8ILlJ9ioRqiRPpx5r1Wy1wDu1/c+bf/
4bEgo4KY8nKek4o5JaFP8ehMrtCZfKSTLYNrUpM3ROZjLXBGL62Bdp5ZK4aJuqO9hH7v5ntasKou
mS9YSjjT3N/hbNo9vTZwDXeifiJ2woLws+Uki6GGa5FOhLU4/qWUPcySyyFyY9FaIV3gOOPLIQMH
Q+MCJQOkn072u0fO5eORQZcB36dOoAMaGcMxaYvvo4yiu7coqavbjqZNSihQ3kBTE6BMYY+E+r9t
OhXjutCRbJVoLbcm9n8Sf+v6QNvF9da5p8io/s7cM2BSeU19IDeO5f0ekyGJWJX4dqjK0OgYoBeg
n2TBw8Pvt3NW6enRDcb6QM4JAE1YzRmaTuyJBvyAf5/2XSH9NsG6TF2FbqFltQZ1KaM1gi3EbP1L
ueBHBJD7AkwA38WgxmwHsCR39AFESVwtPuK6pBetmMmDY+zf5rGrxa7h9KWokRCRlgoLVlBUOSZk
YEXr4nPbMNQ+IZDC/egwppakKgLMBDc27mrSLR20YQ7hwkmcwXyNFhkjBaJmKDpYQOmcS6UH6z4T
4TIQvP8ryS7I6G81TdxP0rf3imIsn9cR2oRoU1tEkDCRxtCn6el3DOMohYiWvzf1XKx26iJpOJ6n
/dPBTHgnbX7bDGOENrlv16clP/e2g/seVrjJWFdemNg0JBIcV9W3Ee+svt6+RPxIXLJpfQs1PaT2
/8FPvgsxLx374wtNT7eAdlT3WLibqcpUt3FNZ83t5H3sJEe7QwGkaZX1ltVtO2z1/PCZuD1+sBrf
HLbajd04ktqdHX6TyZyIer3IBQAv7TFoVuk2OdBSeR7kx2pzgJ88899LXGEiQqcKgIJgxr0CQKOj
ZY/iUVbKbUY34ni3PF3T58WtS4VcbYG6sOcGYGcvdToNbgXZbw4UzubERYA5XFS2N0Jl0RXtUO1B
2SDpXVJ6oalAKsm8O2cCgbo2E3ZtKAIGoxqQAj8YHThmL8ziSaJgEsC8Uc5bV8mBqktfChaErIDV
1Spoe4XCb5u6mVQQx1AGtnNzgsAuLviUjaYZ/KGGe7iwEGQFpde7hOnUNWSkXQ/JbCtOm2frJoan
twaDe+T0ynBW3JdgivCXjHeoU9+tEmyqhFzX4MQj9raJfsFWE3E9amZ93ZqFvLh1vTOLHqmZCyyb
7OzoYipSRSY7at3H9FHO6HYzEoXV+jAuC5XeTI2mtcjfa+7LcCOjR+eNPImd6bNd3DrC4EFpRAxR
n/qODKxYeh0RuzJw2s6RaooeTdCMHfNkMOCWZS1ETcjLTsZJhpyVkW+wJMRcFGuqpN8ppkO0CS/t
aGEma0EE5a1LhI2Ae9g6BhUEvg7k/HsK4sWdsw/NUj6l3B67fuyTXvOGMheIbruOP08iQyx8ICz5
C+pqVCJh/D8KSJECBQvmuAqQ/IPgD3E+UL9rd7cGLfD4x18yOSnsb+VwUPFqZPLjSSwILE/6Xy+f
lBOyL1LrrYxQKcXP+Ja4aCDGN35Dt+YgFjeyyf3Qh6Sobmns/qsoZfTjhHRmEeSj6sDDekQ4bHA1
z98/RXGFfyFO1R9tmBBnWxB7CXFUADGNtF5IquQHCUSdjSnzAXQjsN+gNpQy+O1xiI/XpkwH19oX
z4nAzDcc50U87OKF39+wrX79u9RdMpslRwZFLVk0a2CFg9axStlM1l5Gv7SBm3jYh75cJJGbd8qN
ouk8tDYz1TRmQjsIrX4WnJPTRkjklS1ZhRL/3BZ2hRx7HYGe9wXzrEgxg2ms0mOGY390IqJmaDd7
iGgdlCFaISmLvKs96dlJo5kkmxhQnIAuf3yLrQq40F1yNgk1zZNNFqkOYPLId7oaw0PFdAnAtFgu
R14XBxTi6RO5HJu2e1pbTRpLy3tQwD0kjEYe0Gg3Ywv5RyIgGkJYrKtN7aNUTUV09lwA/PcrcSFy
vaKPfP9NXk1lS0bWIT0WyhWahroQnja4w71ojKesgyeVVRDgKqUh3I+j2o+Zgubcn+qLpNTdg53q
ZJXm/fkwyuAEFAlx7a7/ip5Q7MNTVkfvDT1GT02ktOJJErOzWQkidP3PDJg+6zG4rZtyS02xvrjA
3jiF5G5/EzQzLhaDJ5tP7HlCyiBVoreGdNs4JPZaS4rdC286kE1sfBAzTBebXpbJGwsS/JHTdxYP
hkhLlSq2xeL7Y5tzpdtoqbLxZVIPxJK2LPFDL2q5aOovYBu/KJeO51OxiTj75aNhqxAmpJeYTbTE
SITyEDu8aOqYunKMFyte0WNDp1jdH9B3wbxGfAtDLnVfkN47wV326CwyP+8dQksSQ4Hw9Ae1lUDQ
p1LL2d88aXL4Hx2X3c4QqTPnZssAqkMeLEsloMecpsIzdYuc11qIGM9Dv0ZY/txZ098nYJHun9++
w1AxKCNnpzuVNphWw7Um5GF6ZPVBHdw5EJIlW7HdivEWwHD1Yo7lB/kGL+veM/2z3HJK7/rEmU1J
t1TwVAJDe6O6dYIoqMNICO5piqK0LpKf/jSRg56Evcq04Rj7s3m5xMoI43mo9t+ORDYN5jyAePy6
weuqJ4hKIV//Fmg6dE913MwO74wnupSwZYvlZmXHQHzQzGA7O1PxYjw45j1yIM0i4OHYTaMHGux4
peAeqchJESCFFfIIwzOEsFleRTWjdd7K5wwzOieWBIr3DKLRDmWtAbPIqRN+zqRsZzRj3powaW2H
Pf1pLgKiYN653BmEbVMITGyXRocoHA9tFyjay7DGj3vE9s7I7oE3QKxDUjGB4DYkJTVBlLvMGg4e
ZD1fsj1RtwOcmn9aUUJCkgCbvmEGlc5mWiC6+viWT0Fj8JTk74ax6BghjnksDH+ffk/jU7GTXmBF
EFJM9ZgMrrZaw/+/pANpzfA/ZEJdaPfjrNc3DpwIjBnXcWmliKlFl3bawKl6Ad8iVJU1DczqAG8x
bci9RSTdiifkNmN9ATgQKIldKoW0jvgQimv5dbkvn6dVjbaVo44tkdoEQeHsZkUfyzcRgIQKBB6Y
KFBIicPsCU2sNWFdYUStfNmsWG5wQ2ua0tP+jIGcvL7RjPblmMomaKB2o8xBnzx6gFMBc4sd4oQ1
kAR5wBdUeKxPqqT8lTg3nc8lP1CW6xroj8gXL362gGimrKWwwk47AzwN6BSMNa5OJo0DejSL+eJO
tRonIUs79ZOdOp5yiE4V1XumEpN+vT6hTpBF4WDCP8yl9GVS4HzDYhQ3OwtJkC+kuzEK+C8rAlyh
Bz6QD4XnNoW2dxHz6lvnvJwKmuSXk/t4/sW0VpZ8M/yVCYhuhVjSiEydT561S2JY0Cph3WMkp0j2
CQPr+P3D8AA3cKMA97ZdQUkK6nyagXTDh+Hnvj7W0TkcV8pPqsxb/LhIYZeoVepJrAuWddbtKe3Q
XArLANdYeQWCu7OiFwFtd1qwKvZim3QGq8b8Ob9yl8gsV68ng5Dtm5chEU7m5/9C1KvQ4JrPRAoR
k6csZ/j6ey17j8ruioLfibabRX2QOCXsDxfXdj2obw8Ey5RXVpX7rZPHM5GXC4ViZyXZ2FJY54ib
Jg708wkjvcqLsbIOEyDp78o4STiu2feOKM0n/3yPrwW0nwXMPhjnbBaCTQwrhvUP1oBAPh/m/6Nm
OSflSw7W+QlDl/zFLC6TTqYVSuNic6gcalEzqBiK2bjozWWDjAMNaX+7s20jyAqEPTT6LAcG+WCb
kZ3H0Tc+6fkitsup0VvBjiMusw9/cPmVkOH/crtm+UjLoQXAP5+b7+pR0/XNxEKfyvpWHEnqcOFN
UFTq1/sLXnVAKyuJrSnZNlIbLN+SEKCAxGFod8LSZ3P2/4LBcIajtzkGiZ4jrQG+mIJo/VtoupgM
DP4=
`protect end_protected
