`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ww1cFCaKpEaygJUT+P6Z2OD0uzJ4IJG8iyHDm5UNlVWbTWS9KXjZ9jEg11wJmlv8lA2AVebHxIas
7nZJsy/GjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gy0/aj7fr+HoqiF2MKC2DdMRffpsNgkz3LCA0LoXsy3oP+ExvEwYs55sO8KAxVdJaUPMOFr+w6Gi
VDRBmTTzMTTD1KvHQEhDppUtYnGyL/2qAWb6xHvmSHDtiAjlHews7qZ26fM0sYgNx48H6LSqgFd4
hai7P1C8/gEiLdaec30=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hi2M/LxF9qgAZzAUuc501Ws9I83yzxDz1ea90Q5QjM7jLsFrH4fLD2d0WWY2wDTdG0Ih+QNnE4S7
Oq9DybBH0zvBRUhAQoExlvdlIfU3Jr1YKpM3lLPQTLIhhCp1eQgIZljQtMN1p0u0HDYYsZO5DBeb
LZHGhmPHPWGqNQ/iLmQ+PQu0B5Cb+1VKyvK7Ipxjf6wKC/NZlztCmWzwV4WC+jY2wHB2IofyzZfo
xRBIRCIpTb+tTiKgZ9oAjPNYVjgXC51YW/c8ZhnzF0gIdh/tD6GDSX/DdrrBN7Oz/gtduYw5jR0b
WsJx7lVGCa/mgRPb2+p2mjuutW8gGGnh6+Yo4A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X16goI57idQ5Yk2jq4rj0BhsplRtdzoYr8oOU2lBTTonp1Nx4fK7AS7KgGuzY4UqvPTHmPTfD5ww
0YcXmh8hr2Hk6aIz+aWFV8C8XcReGDrBhi5Np0Vi5hozuTfEPpWuDV7kTmarku7FYKZbPt+lsAsd
f8+cIo7ySKaxPnzoHbw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RA9GWDJZOdw/NASVbYOgehelK35X4QCDpOGKLkbLHbvCU34C5eqCOlazH25KMTrAHxM2lx7+fAsw
HHb2ZWqK4pB4ww23gPcOsgxVCyXs7Dx/H6E84snPbj5EBFAp1p9GZJoguz0skOVQzCSeso4vwekP
kvLqf3Ypkz4/BbGmeIV5O3MvxWppwuIHCb+NDzDYU2x9uQ7mLUtu7pYCzPfN1FeLiv9ttZaXRuYJ
ADExpcAMpFzH3bwg6Tm6wL+J1DzA4jLGZxI9jxK+L6xNTv2NtONryX7sLla9heWPJCSHR4TT8ow3
t3QklA4V7oRFEhlMh0Nv7QVOAHjukKSZ99LumA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4768)
`protect data_block
2JEuFaTgqghMsv5lmjCzRK3A++11CP1BGktXmilnPF3kO3BNw3Sq9uSYJ2pBZAfEozFS3A53Ggxo
JqnL4GngMEQRrYbIm4bsZy+EZ8TdSX+tLWwcGLFK8xgP1MrCrEO2M8jgZgRKowlZiBLnnN9nbuB6
nxtcs3raYYmH9szuZ9WQ6dQn7mRPAN2iVXekzs94weVGc5a5RYSV8nmrAhSET/Xyof5NP+32b1Ib
jJZ4OSENKsVi2MBjmkcCOD4XcAT7+TN8lW5Kb8ffx0Hn160YgwlxiNqs+c7NthWrAV5D3f83dwEU
7Ev7vE8g9k1AppFzBmytUuyVygIPVudbukhu0s8BAsEN+2tgiyb7vuQz+RKiYhfTpSDmGsmH+Sor
k0gnchkv/3FsAQj0cdZhWAcvu+f0SPljWu7fUrNkYYZpR6LpiCrkpIgzK7RriE6Kl4uCp3xTMhIF
Ewwf9pQAJCf0/ljmqlqk29H5MFZzXE+6++NaDME55d/t+B9E27ilG6F7+9pOPpubjFsuU29AlSi8
LWZtdMNTTBP/J7+w6UzE8tOihNlxZu2CbU/SBk7hO3NJTm6n9JSUWp8N+ubkknxk4o5xS4MgF5eB
QvZk+4q6OqM+E7KwuEYA1lyRXdPJ5uizxCcrTP2YAhWUYdn6gxmU88XJAHHJJXDjYQ1B8Qq7Gjdx
XXHUuUkU/08WjP3X1rV+mZdY2QEFCCJ7Qtp3mmZcaWNyu+HnS6P6fg8L/2cyf0NtBpGUEAnYGyKv
PFXuIiSLU+XTByhn842Pfnex/KL9qa4mncxERDsbCBPXzbc7ica5wTXw3r4BMrJhs/o+4NSWgnco
6iU1iudJqYpUXEHbPzGBPYc2w7eJVVdtPmW/ljb7z+KwLI33DXLZ6rdDwbbiUc6ihRH92qv7vzgF
2EmbQoyXuqWypuKaodptcjakK425gx7s1x7lq/CWF/+evb31+ZOiQ7PUG3JF5ffTdNHaYs2+pTt+
lX4e3Nsp0QRfNa1RjIex+gcVn1B924cp+pWsnF0b/EuwQYlkqMdjkXpo8RptfsBdJJoGgFQv+WFf
hxXIpXY96KPtE+PUCFX0RUi7P9RCj4BJDZFDfidSnfZtKkEiUDSzWp+hN+a4f7qPytJgU/SXtGXh
hX7ha9Ntb3DhRXw2Rg4Rv1W1vX2V5Uy6uXzc2yNIqQ1FZ7rQyYk61BYQh70MaL+H02CGpTXGP4jt
Hlrb0I5D0/TxBVYLNWTUnSwnM7JfXE++VPYBHu/Tnngo4H3XoUWZf8y+Lb2IudxbjySbJMnmiYCh
XCxChX5pWU3nQBLjdU/YTmN9uIh/m/2uymfLkcvVok75JHb5HLdCsiVN8+0zVvDgoMf4gLcA2s/A
apbTs+CgMerjGkcM1YB8S5GuH8u1ADr4mEjiNIU6U2AsKV1Z6+11hE0En7n5J6BYEDGI/PpLz7Z6
YKelvFYeGf85HoMqNYTMXlc1Uoll1d3d4qbLN+spvmx28UwTDv9LSAeX2miQRmr3w2izB5HQxNqs
0T55MNXf36+/TpzW/GGTnvvmjEOV2Pqq9XmP9zZNEmHQq9CF0UapO3I9e+9AWW+HcfrGRxt9Cqo1
ZoNikvZe2VX0J0c+OiFtf4bzHHuyDwhloFMTFXHAAp8DLFLNA2RDilXXMJKRdFWmzDdSA8GV+6Bk
5XWnjwvMBTs4W198FDcgaExY9EdhXlze1mVibA+I/ILGphEdf/gxM2Yhp13GWwjS/LaMxguyEyHo
CcXcUmFcXbY2UN+urvCMearnDX72d1WHUzDtcW/idnakyTmfRfmW3g3UtpI4eXE9NJ+kqrMp9mSn
gtazjLdv04i5jDZlENlmOY/zIYl5OoiTs6ajhAbCd0pCm4nD11iazjykt9XwKWDWquqgyb7jeAVB
kIjiwqU2wTS1gJDm3YsXyBVF/covP7t5TcH8jhzDM7+q9I5SI/MPxOLWwC/eCgFetjchfDw513Hj
ZZxb/bBrMSk5b8+QqFyGIbsZEzdtsu1/hsNt7z6peLZHXZv426b33aO9RKClSaZ0CdHNKgu6KX3M
1qOFQ45sUXFjT/oMmo9CWHl5to4vIOUlwZqdEj7W/loP8LtzwB9Unuqm+lZD071kfoyTxLjFiylI
eKQYXglegrwZiDZQnrXHCOfkKcomodiuMnumbDLtKOjTtdIz6dmeK+sn8D458JBF+F0TU8s7dHZh
2gdKobnBkgaGGWdQ/dtaQNPR+0wBuHYYWkrwM6jDEL4PDapFQSR2A/fjTM7/B5UqMIuwAQq4mgLx
o7kR47TwUl2R/lbFOSFBeWt74cadTOi+2dqXlUC+tzinkztHHcw9e84G+DGC9nGz+SYeg7q0/iaR
Kh0ILeJZC9vj/9lOA5wCZuHP11boxPJOMwCZZ6UZUXFiYtakC5YjfoSi72A6rYwhS+4K/MZ7qRT8
47LP+/EkToc0/kOkmBfA6DbjEl7S7ZE02CWZ6gx/uBOhBGXAfHu4tXLT4eh29L18lmV2zPCQ97F8
V0r5BMbBj7zMGdUBUwx7a9S7RH2ome2r+BS8ewcXd/wnN9aqWNzmdNUB9T+1zaCp2NolTZDDL06A
fyRo4U8XvK+sO/9TtkNKANMPJtnjIKxjhd+da14wHYbLrLXac0+MhesOtgQ1u7NvnTHnLaz6OLVr
xn2vUal5vXbEZumWcQRgnXPkxeViWBEe9Df5yKEtYWUC0NuB4VVSOYxKgzf8J+DL0+oRdXtMRIJk
WBUIqOMHsFbDKslE+LiYlXZ4/0g8teBNRszLAZ14qVOKbX+SBFCAtiX2BP9MIM1VI1KcPG6yp9EQ
1oz5dt4wOhIuP8HkZLKgwWSslqc97DA/Rzh+DCg/v9pDV/3P3/BixmtpFPMsPN5+nJPBFrFKcG5m
+9vRkPesTsfR9O1ou9RzELyEkfaaauJ7cm8LhbI9EnuHdufpVFFs5nHC5h/Gyd1HwmsWYC2vbFGN
TY4aPTzSI69ua8N65lBXDr5zJrAm00sYuZ6OHpr2VAAGERHwtJNe9JM39oDezodxpgzHjwCjtLdG
wZnYc75r0rYuF3emAYJoZiE7MB7eYyKqBFkVXUwggKK8q8DFE7Cpf/XUzWOpo5c5mhfpo5PIkk/7
hdf2s1ViyGAKM7SBth+IsjZJM4p8vOBje6NFOcQojD+y7EGycMolUZLZsui0zLNhusOMatW4Getn
RD8Ii7JvQQsMxPOYSDOYQrTy6ew7YQtSfqGMjgI0Q9Vq5xxPR+FQ2hmUA2+lqJsDS44kXNk5HzPo
QioxeqqNFnWK7aSIFXUw7wjFxjldfEsHwaMGV/DGokOAIJZJD4XcSKfrj0dNU6ksVWQjxo3vwcg6
cgCRhZhPBdXmuInScOTiC2GhaTtWLAShbiDYWJxdHekYkwU1XYMG3F5oU0kIauISZR+Q8Tt79hkD
KgZlhEAUVNwTMZpjoulWTv7cwTz27baylHuffe+3Iu+eS383Dychfe0ZjccqM/OJU5jl0IRaYQ0j
pFERn2ea6RMbQgbSd5ollpKkxrX6rjzBenuo7R4CsuWc3mBlzMwTDBG4Elu95DMBrpIz4bg70S3E
flHRfOc4X7qU0wBg4PuS/dUDgCX/dPNpa6wtrS37lcmQa9RJ7/6gFW2otF28+EbeAkgQAAk/LbwZ
1LYgb7w0muc9VX+txxkphduhAR5lfp5bmLVuQ38sTtD7kyOANnmTwnz4kKUFnkVV7VEoJf/zf+LR
53id2wXBlhmpAjUxh1UnvkZGeGFYRFng1EkkOTVqxgwp66tPBHHLhRPmqzdfwg+PyaPvlhuv1KQv
nDPukaayg7aXI9xtdOeYFZncSh05Zh3d+rsuTBZ1OjQabQFNuqUbeOf1vsp9rwVjZtWydIIc4I5Y
0/f4vt02HsQFYaLk4h8rzZ0fSbyY/h6gB/xJbRRSnUH5mxRTiDAI/jOpu7DazfkDL3LyD/zwCbd/
Dd1bRqsafAyCVf/6bnQXlKBFVOiaooGBP9RNHMgEGwcSblQ25jVIXIv3bnKVXUosfsBjPoajqUCI
JT2iDl83e/xWIH2BhqV1Sc9urOvwpak6VmJ9XWVL4ZGXYbWaZCyZwYMzP0V6tj+4iNqmm30dHJ5d
ffoZPZOYVHmwWLa7xzc2faFtOsSISDbxgNhq6IbgzbVkFU2xeGZb2lt5zzDuBVEDs+Ec5EYKpUtW
cTZchazqISjbh29Md5nm0uWO5ShIP7AomNVpaw6ZNskFhAWeXj5l+rCVfME4B4Z/sxBai+Z3+VIy
qrJQZ6CT0apxKACH0/GalxpW4Tw5C8z3kE6DGBZPhZ98F5FEPz+nWnsKQX5p8eaZaFODKUUb+J0A
gVocn0CC++WtOC9zzkTdg16lAC+R7byA872ffuPaaPs81CpziSljU66UIDltF8GBbLVDq0dQbYeD
qontw6SBESpobjxvzN9CXOssSRQYnj3ZVi2bznQ31Oft6phNXR275UTn/KAWgpF+98IMXq5Z3wS6
rtq8HTTHwNv1dxEOt61s1mqIoiJPLmz+uHmZBFEUakgXlXiZ71FzqMsWvXvKpHr78+zaLrOcwyRZ
fG9QXhUYHdBAUbu0zl2Hbj6iBaAoCV3dQuaaQ5Vyb9SCjWHzJztfcC+sfoU6x/IwuMU5sUsmMVH7
+jwEaNH2FMN2ulNMWwncdm/dZtUIpmtWfQZI6K9IRQf6vvpoH02QwvYyqmsIa0I+88Yfgh88ZKKD
1n85imCJ7z6WpNs8ggvJcxkugJ6YVZTA78ddBNhVYcCVDFmd74pn35Ct2co6f2KuM3hY8uHyItpn
baJNpsAGcqfyikFMk4VXE8I874NGZ+4Okodx0DR4xUgFQ4/Cm1BWyzwVj4Y/8NugtP9MYKq0rYB+
NwSCW2J5jHZBFhY4wwHHDXrvivOx121eU2mE4kDE5IHOiAXLtPBxFt7wh61Yw0jIdUT17ZAinv3O
0j+zYJHSi2Hw6O/4+mv604jOaY30Sv+6NhUxC9PiHgaGjRuRnHuRBTvEdAYDcw7YFwDyO9a7szRl
kvngGlY8bBgM3I0XeQxNpdZneumRXggCSyEgoSSgjbTGK5AJjAlzTNlcmh99PMY7LfI64QEc1Bo5
y0DaD3pNth8Hf9z0l+N6zvro9T9gzLZOmPxvD5WQOaJGcIHOMvquhZRR3OWXV3FV6ckbrFi6x02N
iPqPl8LVDUGpn522bGAIKDO3sSI62sqCOES6ukUQ45RXL4BM04noozehWboeYORgYl74ViMF9U+F
QCygWMjE/q4SL9Jw9Rxc58CIy0a0p8mereHazfB/JRwQdrRnSdkLdMnpjx6x2BIlhqJ+pJf00grT
GTLdTTvsvDYyQng+dAVFOj2wiUHIwf3R1xkw4hRvydv/187vqGBtlbhKgfZ37E0ge1buunmrxh8X
U4ITI6UidVGV71pD868/hOQMKFUBuBchs68eqj2DuZEEVcr6Br+PhgUvm46jjRFD97IJyhy8OobI
kbI9NgFfX+DC4EYEGdp4ik+bk4OfCZVI9fYd9TfriYu463wkTEdmOF2PxYicOBBAZPLYl7uI4Cc8
J6I0sCQb3CqrasH2z5WM/uWhxZSMQrBl6KqaRc0jtNSa1AF473EReASaPKkuqxuJgbaqBL6ncIvn
LPo1v8yAHnxbuJ2Q9sbctT1Gq6E+xXQXWaOtQIHlLUidyv7VhIB57/C6b0sRO1fJ8D43oRATmlzN
f1b4JruaTF4QOEhpcV/hq3aN5G3PrBln8VBuc/n0KSDUXOj9roUJ4rupNEaKxCNor67jf9J5YyiG
gnPO/Z1gpQwudpHTkOTOxNNRCxn6BfdVJVxgJfkYSD3iliC0iQUIb/2ik3Oo8YVcK9m2PIYWQmG4
S4S1avG12/wksk3VCs+JlYMYJ3xR/kyaKTxXVvUaPR2R83IYbM2ajH4kxWN0Hc4vXP1F0XFW8B0i
ZuY51Lq/rjOkebXu9m2CM2hHPnb40E5Mr44FhfjpZszfkUBNUNCh+WtcCmjfI95YZB8zzCsd/ILM
35f2Hveigxx+eUaHh77SYxbJrtYcxfX/a//0D5902JVnSDowJpqnL6vaCSoVEkFx11+/2f69X7Mm
oo6nzSpXaQebPbOxCLUDI7dmj4E5AWuwwYU6nfjYD5/eiUPax3v5HRx+VkiVRb7B3wxzPwCNhQeu
AQylFweVze7hofRtn4DdzlAzrc7Ax2nuhk2Ti/DGkBFb8jCmtK/ryntUjpIiAGttFS3qNB70NBhT
OqEOQAlWpFvoLVUnfszmQpBCyyE8Bc5SW3BHLHMJ1wSCUx9mx8OB6Hoc5xoG163a65LmsbDzb543
NgJUNaJv4/mOlhu+dtyl+d2GWMm+svuq2N4vunwqWl+5BPgxzw==
`protect end_protected
