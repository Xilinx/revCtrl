`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
crsuNbGKr2+HGjsnrWAO3ApjaENLE5lmTkmDpqy6wXOqFQIJnrktoh4R9l/TVlY/BEwSOhFtvEbq
RKvf5np1ZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfoL36fNI5DjzIQX15YYPTK98uQI+Z0aMjl+hiAVWq0lzClrfpDjXWaPyQGiPvnYkkUnnCNmSyGP
qGrNm7GOsjezCGzMgQVr0792OKktWuV2kt0zVP1RUZuHk/37eznwh8N2o5rw+1YzW4dGzl1QbJom
tmB1UpBcp868gDBGaIo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nZKDyxkYA9uy2Xb3FwpEri9edMFM6SqsP4Aed0tRsVeeX445M1QANBu8GOl8sJ4QNxr6T3VU33/s
FK93SNbe96iXZq7rd0ZTftDGFn/wlb+m7r0WSjfp5pkNrLXaYMROFr5Y+cSF68dabG3s3COIhufS
z6LjxtxffkVZFl10/p5NYIyhVlCgj28/qTLowb5EYe1tZ0WPUAxBFuTyFKtX6X8Ha+x+nETiYK6i
PAhbV564AhzWOG1ohxDJJcn/sq1JfdeuDFdYSbNKycH1TqhYGY4rODz7EB10q4+UCVziUOr4Tv4R
NCotWnw5vu+fF2mIxu+vVyyYTSX+rhEfPs2iXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZ2XWhB75BM0Dt/9VMCHTjvBqUtECoyfIkFt8UyDN1IrerieLUkQavGMJnAyOgfgB2F9GkPnzVQV
7H9tsdZ87Y+A3ybRmsawN7gt2tqx/GGsvZlikuuSepi3sHN1vWxch8VpcI/SFn7CnlCh0jupM6VR
707+yLDj5AJkQVyH1LA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S4eCKuneguafnmn96ntdnponlGVTmyJu6zrxyF34ICbqsowM9Vhvgm6poU8XDQ/BrjS+RNPc37Fg
G4CZX64FNy0IB8M93ARmuOVvrGN2bYMf3jNRnVO/z1hOqr23u4iXXLcNjJcX+q+ntygTqDn+dkJa
tNf5JDJd7KcZbafDC5iOu1RcjafQnwlpqyaxuvNRdQkJM7f5tDyB/fmqWMaeSiYSf6cbwC2Jk6x0
7wUP2rAkEzcYQjkJqSGT74QQ9ZxpJuO1xNUbfsJDlmWbSmEyg55J46Q3XRBw9O4UV1TNB2XnSxvt
0rRnDIzS8sn75CDPR31VCmG8K+PwSCayofA3ZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17552)
`protect data_block
HGwVbJA7sypyD5yh/+WUmTRH1DY0aA5L7AQDUWr6ClOGIvnn0QaYa1eTlxZLj+z20JIGsk5V69k7
V5RrBwgRTd9AGKcOgqujCdZ69suN7QVFkvNqjJrKH6pxPXi6NySe7ntJGHeD572hTNMpjRFAAz5T
fAhKC5uUH0r4CSxkEohyQEzRBYc/ZEz/mP3uPxyx92znKJAgULOhIEHyQ/sPZOVCCDwFSGWLMWhp
a68zhjTNn9BJhESTB2e7JhCuxoNsVO+AF5Z4johBHW/zNR05aKNZI0jNXxzMIdB0udTnWuwgNqhj
6wEt/U9EP67TIIzq8RJ8CiEc2JT2lS/DW5n/pTyOVL80BUU7SELhSc+g9U0DFBLNJ9gpcoAKtQk8
Z5N90dEURqLZIZX4ue3dijStZrIlPpTR0LF8FS2mBrqCMqkVPEZJHAPlPhV7dN9M0gd5LjrAod3m
6asyOEZHT4ZPcUVyTD56l0ejyvMxy808erMlcpDRoknOq5WGrJIQZvtYvYR2tRBbf/I/6LI46h8x
hEW8/NZA/OUhyL2YB/LFuYK/fGBRieTNO3okXXQsx8i5Dj1waUFs4axYNdPUp9SKLhgZGv1h5biH
IeBUn6QRhv8SF4wrjEWSua+J/hqjZcoJLyGZrE/vcO7KRrDmx0T5C2TNhMDjhjxOZrvAgOt9wk5Y
CXmY6iby0slvT2F5jfb/RPS+zzugA5opdRjJhwWLmm2WXGWi+QKQzxXAnY/5a/151dvJ1EVf3QRX
UNFddVtxyYTnR/a1e/026gmkIkM86C08NFp/mUYKV87b1rKdbZHICCUEJdEAuJYlTW6ZyRWv4/5W
zvi/dHKu8q2rrmg10KhlJMuhaDAigEb/z2dYMJ0BfsplXgvcbfCOFyHgKdWwAww6dZ8i1tD400JE
4QI7gD5FKpIOGcx624Y7tWKpsU/dZCsMKHaHShzmp9KyfKCjhOQ9s0VMI6yFK66T6ldqeDbAU3Sj
nK3KOmQmWKdvbD7kOF3spedbECZUiCGp67xYvrFPg+lwlDUiYQUOVxDULYjr3O6iEB2i/Htv5/r4
yMxrHFCSf9uqcJXOmZaGYkDl0Ljk5Kel+Yu0M06TjLsYqtyqKSwHwIPHa9faFPx7+x33+5iTthIB
S4IQ+BxFLYfvDfSewE6IG5AKdzp9Jv9Uhfwt2LVUjsq/ReKR7eBa/2f4Q7TDnGwsS0dv5yGHHbBu
DGX3i0CxKKAiYUH5uWENHVYU/9N2ZoOUaYE80z3EZlwXeEOzs8f3pdHuJfKOrwWyx5UF01qDk5IH
4k+tsTm60a95foZcQrK2ORDWcWA1gJPgn/QxiJFcrjHeEYO4pvP0RKneFz8e46U2/k3gtbHoJ/8z
HdRTyaTfwXz8D95bPbfpkPkdcamGIilA11P3CEAnA4BjfCb4zCCtb1E9JMoNqPpuJ5YbMdQJy6cX
Sg7RZlAYgSoS60KtnrPwV9m9icNxqcus26GxohnHjYVjZoJaDzzbWjj7hnpChy4byuAiVQJDW1kB
8lNQd4RqcfrX/sQyDUDv/O9d8M/9BRHHPz90c9fcl9MDuQEgpY75ybYkWkdp1b8eezXw5BVWjFCV
uNOkBZBU5X5qq/11H3gbkzsYWkhWXkMYu0Qd5w2tewhqRGYGobFgw9oK1+ioBcUF41ehqJvMJJ3X
8MXHyuSYubNlSKHGLXkgA6x+OLmLg986eI+MqyyiATrk6rc06Opzy2x6TrrWx42ZiNlZ6J0deo3l
YeWpIBufHy/PGSUNDbwlRhXBYqcE81Qg3H20gg4zS2xvyjMSH4GFt/OREMLmqWmq4OVEjJYQ9bQf
IAq8U4chFm0PwQQRtP8yzilqYbmTQwIaNI2leo5U+SCo5ZF2/buVqg7R2C+bi8ceOl7EsXLvDD6U
rDTrQWbldBxIu2Lk8UGXswGTt/26BCKIcifHzgg1LgIeMA8MrHB2r71s+k+TiK4kFb6ePJLAF90k
JCuAtX/OytiJd2JLF6JdtDQVFnKVKAXCktGQR2ZGOuCCZnBTUzUSNCkyPkawne94kK5HLLQCosCY
iTwiZPIVLcg7xQdThtDxgaGMdnYjEPKWkuE3MpO1o17Fo/ZZ0BOcC+ZGVi7JCta7k2F4a0sh6ObD
3MRihPPAZCClz/yTXiF1OE7VaNRxYnO42TMgC1iHeFOb9amEMyYEeZDE6xVzZKD1KbDodMjp6ijT
txWva1OImH/OY+E2+e10n+vVIuBgbKvoR3ZL8fxZAazJqzYc3G4jtHjRBLsC/3K2vBh1DqYJiPrn
PWMpr2rQy3nOzVBPWqW1qXIEjHOw9md2AQ9Hfx1i7Mm4VB26DcnJ2pH3XRDOlKUrOmdyipqCaxog
bJKbYKSDL5KUXiAo97bum4+/rHIPgAcKA8p+oT5pGq69/7EiE3nGqri823Z1quFH42ZZfvZYau+G
0trgbZbgMbTPmh1TM+ux8FUFkUSM4F2iyf2gb+uNzN4b2pJASQQo23ftFP9XyW5Tn0M4B6fu+E/K
LQ/eeG9laZh4fDqtyr+Fhllmxq0SLi6BMMpnWLLMOwl5IyNBcHls23X2nu3EDATFA/8rghjNkbxv
jjepeVHqY5hFYrvPsEM3t2J08QqJqEXOyvnjoQhFvKeN7hFZ2LfbhGLpA6mpgyMYzh+GuqLE/d4+
mKX4J6zopRLjkjzaACPdDojnEZtiNKLcoD5a0xok/vza94Yh3bpP4JoSjDhHoHiEdl8LUPVTqBVI
b5+ZaJsB4bAkVkFtx9BNBE+1U7Ar28c5QBDtvTi4z/rI/SXRB+hiYW97at5eX0VoHEBDYf7tpiQ4
GgAXbAXI5fzuwicyc5zmC4Vih6uZNrE5GJpSuQ3d2VeCqkpkp0Kwm2OV/opHYgR8uAHOSDL4WmJJ
No0dsjauG7MrG0j6sGZmrTqCI6kkshhMCka8AiOs64OcImLGdNSPZIgChYHbDCL8aEKBetD1efoo
ViIxVNlPP3VFFifxRIk8+hihJUo6prSuVDJK4WXQ/o2cGVyGRseujVf4PEq1lbVjB1ioe7955FaF
toa4M/7YZ2LsdaR7BMWle1kvvWy3SGVUJ97f3N7Ox//H5RyubpyCSfhYOBee77Kx/EVE2/CNQiVm
VhrmTG5sK9KOTtWWfnfSSGZPls5n0JBXepVT7foBgEsmOQkaN2TZwx7/CGT4Ehh94ByVzJUP78jd
GP0rC0D2pMDV4x6v+daA134+qnrePzOxce2zCZDkIkpRw02MVmRRA8rXkOMMVw3HcpeDoOCR/Pqe
V7xf7XrtM4o9BtLE8l0pzNUw6EJNolkOwz/sv7J+jo8T6j4U9eXO9T4SkAxxccqrb/NdMdWZyhFR
vmt+DjtFjJN+CnUZe1JhcUiNoleTrkhMNk1XIkiHuC1aANprZqOvF2kZ2+1wfxZNPtfn06K7ie47
HvZH41LgcIQP7g84WWlX3su6htC7XM7inh7VwEpuYMMy8qNTh1WBDHkwbkUvB+klgqR42kgK/2dQ
KanzUuBbTYC5vNjp5zxYcgNBcjbfgF2pMmuXX/Pl4VBJ9GleWFKmxPenSsZZlRxo2Pq1Azq5Oghl
oFMeWHatYRehb1wmfUcor0DfEoesqUXlKXOnNQXraMU0W/GHBxDhHgTG6jOhXTljYPRAELhckp8E
12WRQKog2qD2TTEFP0EzT2GQtqKoFnoy/ih2+D3bhIVvxJyPJ9Sm3h1HjlVN4Oods8vf7CEcGQH5
pAMMtygQKuB8OdKHtTYtit4RrdR93Ac0nbQK6YseIWJftc1hU2PPE3Eit5Xr7AI+DtGs7l9ccr5s
hw7EeMW3G+37Msd2WcTOrtAVANAXsZscQc5BYig06iNkBiqExSP2XypFAmNktMp5n/7a1N3E8a5+
ztu0BLqcPVx14RApLI8CFeE5LRtr68aFB1uvg2xbDUk8mTgSbtyBLgNGhOeu7MvLV0WXVU0fUXVg
YuP0eGMg+oMzvqxtccRFib3jw6eboC5hAQt4z47pw/vEwZez1kel5eU1q8wlHd05ADzfZA0KFbv+
SorQpWBZRW7sy2dYu/uKSB17uNEgNRNfTzfZx7SCoJ/1vNdMhiSTrinIcN3lq5m4FJ4Wzn8souVa
QERaViIUQqIcbXU2MYbqEXPcm+9qWm1EyRyLIYO4/pKzAs2YjkZJo+5ytwRxoYLW/cMzuUNsKqbg
hPgtJip3zH0otUwpy5QfzHtl/TqWk0MKARH5Q/LgrRYyJarYucwF+pwkVwsLS+JZWtN0vW7Pl6tB
JFn92eHKZj1XFt+5/wpAm6cJZx+R89dXHxjxj9SO6ke5Rw5ImNMlQ7AE47uaHz85YA1Mu9+KAs/L
ps4UMnoy9UgZ+2Gd5Q3SA5QtnGSAQcLT20NVwXExVE1aiBDfVEbnzni8KtHSGBGKd0i3aYIMoKuN
nWOtjhuZvkpj/q0tx7WDsX9pOYW77y9SvIG48ZXsjqEJl/GLaXJ0Jem3xBEbbQpKglo+cVqXLIub
6Bd4fAyWWvUWjyoE/k36em4V8AwB5lNDV++7/n1TQ+GoBlNGOxOAB1cLuNS4H4SKdoo0jsl0Susp
TwZjq4lA36gcXh6Zrw3m5fCTk1d8twk5dg0NunX40zoL1NBC5zEUfjiLZcF6xauSwBrNoS0Xkb1p
/Kzl36UiAF8ThTkshhTShtsVqA606LOYZZfKpTKAAHdjgWUa3qp7Nhe4rEGBBDmIHPcQOYYiXjdv
hTM499t7y2HNvh4mJyHoO60ATUm/VDN8wXs+XuS50tNcIgFJ6cen2/YDeU8Kdwh2JDFu5qE/2/cD
y57P48Zb8NEh//mlEIjemsft8hw4oByjWAOlDaAwGvVkJxOcZc8Yy6OUREPGouskpMU3Vb+BxlrS
EwU+uG9K9naRzm/8SNCt1FR/0S0aFVMJf9QJNvma9xOcQyo1PD1ZdJzyi13OqTeVYxCanqlOEELV
jYg93i8HKRHllK2Utg82GLCbxpKnthu9Pzy3InB3E0hqVrJqOpvlO1qC+UjFyprL4fVDZFUSqLMO
v2icCuQVMEoSV7TXRyTlHAkL1abnLgTUJ64DLLoo493A8Tdy86xsgOUJ7/0F8kD5NYNQPAaLNx0E
2BfUQI7sPXPPPSbrLTIEqypTT9UiyaLBFzB7bYW26bOQvDdhCn6l3PHOP2mASz6zMcuzdKPQHsur
5AlPpLKPKEp16oYT156w/3ZQl76/NC+OIouirjei2Cv+Ci000xXVTHSR2d2Yu3LQQZGdgzEiwJbT
+LBgO/apkNe8D6ahY/UIsp3FbZCuoOP2gmgULdCA0QFHDi6TLxagSOkU1UcTho0wRdQJy8kk4NYV
DLx9J2PGI8pGpGDXEqIIi4beuVV4PMtyrB2KpgcXd3qgQUeVS0aQ8hv318WOPNIXUCWHyFb+7FZY
6b91GftN2ko+tyv4fr5wsX3lICqPd9xd/AbNUEnGVEvBMGi6InkGKrxeWzFUengAQdiZHBqQ2TiP
iIqxCGQsRv4IX7fGptVuvApARh7PgvbKm6O6ZfEEn6TKABBvx10QhmxRQQwSVv6NR2a7GNovJRFS
8qobgk5NUjYkgGlhoSb02CItalgEBm54XV8cLVs9Aq/sYvpK8ew7vm3LKjdnlsjEt4DnE9j5j+RD
ouFlqnv3L/fJFyg1wzB/zrgBXuUolG5rXOJ/HYuFyFn25VfaZN8jBuwOiHyXSkbCvkt2jtUQ0rkA
rwy6hdfRyf/zRDMjgCnC/YMrocNJ+yCvKyBQT9k7CuR6ofymuZcKq1o3vpLMCvaLgLRtoS79Lo44
wurs/z31WClKdvenKbqJNEoYBMW+ZwGGlU0hpZ/dhrBiGw4KjgT89HO1LWhjbXn9omCXvxz8Thci
mMd8RogBBs7pdBfOSFjugwn9/7rrF4PgsEY3xet28q3jVIVxAq830jBcd/Og+1w/BWyX3mRZuGhJ
MgN8BXIClM2ztuHk+6xMZ4sH0cePCJiTQCqWiWNOzmUx+C9i9tf7nL76aJlf9l1q/9peBYepFZoB
hPE7sharAL9+T0OilZLpIMdWvgYlr5p2VtP2hrTsYEb4EBfQwVTcRv0qu8biffmpioQ8CrUHP1JY
x0OqhNTF93HW9XtZU67TR7JbrPCsKReqCdV7GxErG+HGi9JPJJnmv3q2tt53D2LLMlYvJ5cJqvOB
OxXuo7acm0CJvB/8lRcQeJD35jouEx8mvMOPRaPLzPUsk6mWXa9m/8tAlgN4QLF7e8JJBP58nczb
KeMqn2CJ2W+aYuma+VVJrPaJEAqkjOdZl0uF9hCtZ0AZ7tEvUPuH1CUO0AM1Oqr9Qp6uEFPZ5ueT
L1DDcJdryCzMmn/NP2V9uyMg2ojUFzr6z6D77a1N2/j8YV0qzSpEsQQp/HVbpiPGuyIA/jV0PHqT
LfimVot4rB6p/cdxZMZhhMXfWmil8kLy8VlKA16ClCTHSuvmy1QjMV/Ur6RfptJDUHVKxoQUdnVn
7zXI7kgRq2RxiFfbwVzYYKN0sdtOT103qdySI2WPkvH5/7iBIJqS8YruAWeVqMsRIYAE932CVZyW
mAK1nEEasRUhf3RWusIUi/qMV0FcSE0cuocidFtD5dHY+OqaJm3UKUGsFIDBrn8xz/1UxPRBPK0L
NULKkMGLV1nrz8911GEF4d50lrGAo43eIPQvlEmfWhwH/kS2Xp1/7DTk4CX51RNf8NJZACky0yDZ
eEEdNWHVVkPMi5yl8ywOPxIsxstAuarmAVbvhGYjrm6JbbRkpZuJvkra2/srq9a18oKEKY/Er5aL
F06aKX623FEUnGL9MCb0azgghSRO42czqkpioE3lGp53HWJ8gK4qo6LQVwBbFqTu5DGfWYsPu4V4
xX5xvfoOv1B4xEI7bCmq26A8hkhFVYJ607OOfK195dQEfODIEhdqKH4+JypPiLXfOhfxJJbRxHl5
w8e17IGrK6S7Eq0MMT3/Ycnw/OkvHA7YrA2vWc6FRUhfBtCUzuD+yApi8UOJv66G9Ftppr5UZxb7
winaLt+MllQ35YboWCTpJlNotUZMqADWVqHCkVSPutyL9U8dyjHMDsbvcCT0smbbBaSjWF7vUgSd
4O9hzeGZQHxtY7tBcF9efLL2QnkIm0kfE1kUpv9B9Var+zV70AgSurU1PHIPxvG8pg4qTmAIm+lU
eJuS/F2L8UyrLxpwdrAkYIR+dq3TI7mrRPt4BroX8PC8ggwiX3eVOZj7ErpCuTDNawG2HVb9zfNN
QpWoiksj26OdlTdC0/nNWL5LjRev25LbUoCWc0Snj93FsoEp/DOnV8P5i6+1wpu5yjJmTJAMcHxR
/KU5ACLSH/TDzRgCdcpHypKPDuwnAQANhN7TdAQV8KShPLT12ixrugkuAyubATGwINqIZ85Hj/+B
u0ZtNwQvCE405Bgyyh6JYjfx2xO0W02sTc6lsEEzpGb9sU/eHajYk/cFF/pyJ3eM6JWTKw5NA8Od
5H5PPI5vjXDbJWAVXKZWDe68PWQLuX87J5O8JR5DaxbUMWKpRSE7owltZbaeTozlnLfufpr7XYCd
sPkCWgCyH3nV5OM2+Yfr85qKrmkdhH8Q1t8wBksWZL0FKW57EUvDorY4HYFI9L3wbJFqPfwHF5zR
HpR6K0vLsbdAq3eBbluUEic1nKROYm5JAnom0lV0Le6IlV1ZB4X7zOhvNcMuHeQYi2QdWq/tDjbm
ioPZ+/+S/MLKcxmx21uVFbUiwZ+aptlHqDrK4Ge+BOK5zqePoES4LAuDOo2SfsOLkPhjyzqhcAfp
OkCv+fsh7kaggd9uDiOPgkoTZMmFWmYbmLMUZfcdxR+eheQEh3rSqcKsMGBn/wOZyFm+AjRz1xqc
wQeqlPmqZF+CpLUSTRC481ND7MUJJPQBZn26VF7buDy0PuuGJh7bD4Oa5wFLLuSVrwPCkTTkBV0v
FiadDwV2wy7tFonOjJsVaUC83RgRQvjZiU6PDyY91hZdohXAaKfYmWToYcdLBoy6hQ5yatUDJGan
wQfqlFREyzmqIlVW9g98sB60a+IzB5j2iVV1h6/Cpe1LxjcVbOAVEXj0k27I9dojiltlTsXXtN5e
20s9lTW0ExuLKLyhvkCGOBw4Ek9IznhE6389BnJIdB4Ce+NDD36AeP4/qzdIsNs50ag6tv8HTeuO
J+tG8Nm678JURdP2MsRtH5kKIceMuKGTSqZwmsinyK4r1L/MqNf8+OzDEC6RQfjWbhRgYIa1Ep2X
imn7SbmhJjaN5iuohX+gyJPz6+7ZvZsXmrtnkED7/1wfQD/jLua3y2SO8WIdg4T3Vg8scBMidLo3
zuo18Hr0Tku6/HHjlWt+5nkqPo1+fy11+PCa11wg2wx0Gtzpqe94Aav/zQJy6ZC90RMKNkeuvtrG
UjW0sAy0egC1IADaPzxYaLuBeZ3vu7c1PBGJCVaoXs2jcAS9COAvWQyseFMmmxVp5We8h+Hz+1Ly
ed+04pj5+BBp4yFHF3tnHD3R8b5jIzra+g8jNpaELIPXuVJwDcO3yzEN0D4P87mCETfYeYymH8Ep
8NIaLGS+Qkffs1djaoWcfelAd6dT0Db9/nEonaS+g7horuFj59xbejQ8exq7rnhiWm73C5vhlXXr
0AQDWr07jFIgN9BCY/OQ2gDWHLzPmcrt9QfHX20L075ggEh6b1dOzJ5DwpNXYBuswPsXnXFZhI8u
NN7fiXF5tYY/CfpgDnroBCh8DxD7JhfxaM6syVabjx8AblWJGgNc6OSOZuTXVxiKj58P8AF1JGiy
4NTf+j/SmoF3YeWXPq+7me9kxkUW7rL4uGZa5yssk4GMlvbrWmhbQUqa3d8QomExlGRqu+ywnwSy
XQcnASrV7jKGpxka9I6v1HLuujP/t0IKkRl6E50ZQo2OH5fByybkuGy6Mn0ivM/Xfv26Y9wdNjIn
P/mfnj3VrKSGwT8SQxE9kR2LKW30ehoEbr4XCpf595p7fBQYmC40bKvuUxRz4SkWBPJ0DTbBFE+l
gMjCoTzNOi1xk+T0CNOWIYP6InthvEtdNXSXVVw+MTAhBTpcvBq+0/okjhCW+9+SpSJT00Se2ka6
JL09UYhf4vo5uqXFHEyR05VPFWefZ4CF+Tg3ocx5uyo2wA/DFvvOHJM6WEY8Jf+NVzgWpMHZQGhu
T8hTusbQUlvIXv6RF6jgk8pKZCVmCSMmTl0103tMOhxhZOlcJII78RRdhgRZchO/XXiZyrz7q4BB
/u5XuRzea3o5K5biXlGcAbqHOVUqZLRLowhNbeZzR4md9jOao5cv7lnNRm6Hf8yYFLA3bHQB5kf+
zBCe7Fl3NesXvlrfyDzJEiVGlz5MYOqI2JNw7PMID1ru+WtEZ2MNOSPGQbiUdxEe9dusREU+4SHi
AND21TUw1gj76mSizXI7zDlh+WdN7IyJdrSTrQnl6vpDmpAD/1sYsyFfrCl4BGLmXxuKZCRtDD5L
R5Ep+DoKydrm+AsyAsnIv5LBsP5jOYC83uvROsJr4H2/J30pY0oRLJ9k7e6x0i7U0ajPzCI8APiB
ADpQBZCMND+ffvIC0uROosYKaw1Wt3yHakdqRiq7nmOk/GKnpAueROkwonIcigojvWE6GiuNYzzm
wwndCUN8Mh50ms+aH+Ly6lVQbeTmZdd+nphdd9zwc7vC4jq24dXBEKE8n4afnzxlG42Hb1p9EOfc
vQyl3PpXWk/KKy/cyv3N+kxIJ6O++0BoJmhngYBCR0g/7OuBdAgH+i9fAYNS98KLcbJf+4i5MPWC
DjAW7oGSJ1wdzcR5aelI9bre/Yy0fP+sg5kNHz22IX0LQCfMP7+Rfm0RzO1lj48NR0NGNc9yoM6I
BRJ7MdKUYTUOW32BU899NdEx0oP+uFEDV2RZXR6MGBQeQekr9Jd9c3p1FngNT0c44aeAVTLziwfa
1ufmmYT98p6IQFDOGvYkBVynrg79mkm7P7fsp7UzeeWfcYWqysSM7f1q5xUvji99XF0DRgxBuFoT
OyKNYfyR+sjJu6mivI38zK5lASdzDErt0DXceNoyN2Y8YHEZm2cutwTbw7PhcZ12gMX2IM9ESMeA
NG2xgEKKHweYs2xnGWEDoyVNzmyn3sSeJcW+pTLso8jVeUnn3eSmu3mlY9OLCHeg6k6dqVbCVmqx
is+r1K90GjSuxUdjnsD9phMLZZeuocqCl3ymr2PXPp/wpcAzIHiWkYYz/d3AYtgLvUUv0JNlnrIU
qOL8kTWsX/8al7JpW9zGJojzulg7n4Syd8qU0FNzubWNWGw1gn/lJrsPq5FEm1GTdf8R3lDfVbI6
t7FISZLdQhndzpK5gg/5XZQuEXgxNniEafE7qpYuCf0qlATZHM2vwtZwbf+PdvfZV7CdETQ+wDWP
/EAir7IEysBa7MCNtyS8sJoRW5uW5xBJPpAFi01tBq8di+McDYmMLxPcmnJAZyJm9SqFO+KW0epd
oSe9VFj5uaZ1OErspVsKUo9v9aFnIp0c2QoETLM63jo1//HSs/oxqMbrYiAX+3adn5QEUdN5hevC
IkJRYBqIsQ6jkFJuMxGs9I41Z7tCec37nZeKqR2UEyjo3MqHPh0zMbjGCSYWXP+XfRg/rwZj8ttX
ysWAiQYB03ZGjOFO0mHKT1ZHFn6apKoHErH7qRTYx+WUG3edkDuKMXjSDRO5aeVxZRsux/Ewq6Po
+BLCsh0gYzzxjc9NYL5b38QyYwsbc9gM+h7iDKwrCCcXTYSQoYbcQ5Rez08ECGJHsDl94Qg3zgd6
Y73Opddikscc9XK3ldg24A8BlsROo5t7IxEBJHqoK8KMpuVFRdTmlBamjPyb8iQXlcYc3k2ckc3C
AdOHJAq8wwm30dFBifH2j4dwmZxZydJVXzrHGEPA8IFZVti5YmJO4hD4qFkrRWFBR6SLd7sZH2hn
NF6OA9bY1C7YGwl9BTa0jc8jx7MBk9xCyfcK1V0AGq1jrwFhvEtxKaZgfnmI8IN+ov9mtOmkN/dL
X8ZeW1Y8PuXF3NTsUdX1SEGpnzlWG4l+GWZAY0KGYm5Cw2BxIHQ/jB45hHCIoECr3sbwNuDBHpzB
Ex36hYAGQ520/x9uQBPpHhPKvxzEXkUbRzgPdIBQr+U8fiCT63rK2+aVmNOpOT7Mm7NrO3qBOBjo
diAKmmm0EKdPg9MX6c3wjD7m/IZPgp+oneY4CYBPP4GQ6G/ZgPNrs8IlFKnl7kGZmFxngSX5RJYM
npyIjO0dBUQzQxvRNLVaaF4y+SAWhnoZh3K47unYta/PxG3Dk3dPp2aV+Rs1DQBZD1cvOo0wYMKQ
KcBXDjYzPEIu6jw/fbQ/QDis8Bf2FBJp771XH4IoZejp0pRc1aEruCP9+dKtdtCz3+xEaytpmBoK
f2u85BHpEQEFX4cN73D7DF33zssxLfjkVI/7L5gt8wGuiRHGajgn21QZvVqOYoAYQhZ2h71oWqYP
qyQc1BiG/e1+qIx9YnzNByj6kyoSIvy2t1t8G3kLOrngXDgYBtuHJx+G9YtBF85e8oHa0dl0oz7J
xbYC1swbwXsxpwXu6hmIT3dtbRYAk8oW6ft6loOb90mzkbltqQsdowMRuIJ5o/VlGw48dWGO8v4u
8z3k9A4ge4TL8gcJHCxn5qqZy/jVi/c4L+XlecJcVePx43Y/SyqHGRoorNPOKpKGcFXz4pX2tFWa
wx1sKATfzCBZyyCxwh7qsR8D/tV6+0mC2Z3sXB0vf7w+isXz1oaHI5CKi1MbDJRHOreGt7raFaeC
yNlLw7eNt9+fcwhmU0iN4H6GuB3mXRGPYqQInUyR/sJMGNYJhEd8rywOfd5oeQM1wLRsxBTuoJZv
7T9SXWk5GIbMfrIaHucLRPKSg6IiyJiinGLUrjLtJatJqkWwEHQHBxGM8ty7kVnL1jRidEb6lx5u
rnvoX1y0PxXKdkU9+iTGFfYWRoPIGxWByubFC5PK7A7FeW+6uJoUhfNu09qRs2P0ZStZSqwnQ9tj
A4Q0wGuJUW8MWRvlPSL/2xg0WvDqDvueYMcPNqHQNdgDfZTSDX0U3uQ3uIylM3FBt2UUHX4DVWZC
UbdNPhhrxNxbsXJ0a+oF5avP0IfOyTdpFlOm0ykoSuDR1XnFxE+A8o1Fn+4VEC9DPRb9FL6PGw7F
/7cj471OhriAyNeelkI+dfHvgZpAFuRkiQ1a1qdXbQY0ZNfapp8GpaEQZzQWEwg1Hx0RNdlwkH2N
tiUHFhQqv4ZFnzRlNRKw0/DQm2xzfhbsxMTRvNkEHVzFy3cF+Xy7QJjkA1Z/7pxD2byBBvbt44b2
Iw35zo7VBfBUxZLtYqgBgqyWjAXl7SRQedQm8gvE4ruvuKi3MOp4JsJErckPZDH4Mod64txW+AzL
F+hzNAxBDCzIyDoL5Dl8SWvIiM7h0mY2J8rvbDpPe7/gNGIqClVqpH9Z7UHa2yjCpJJflMHyyI2L
+XbcsBcyG/JRmiEJaa++xI9DF9X6RtxRsbcteTBEw16pdZ944c4u9eiigEFxvycZwlT/5eL3FDdP
Nrpf1ECArg4ivSk/jk66o+gczLyqecUce4vyg/+SyT8Ni7gGJT2AbG0Z7JDsvMoPi1QWR1wIw7Sl
9+SkcC3SVQpBv6m3R94ZN/TPTDs6L/ZeY/gE5x02fHPKEMAuZiD6955uBfCgXKUtOHQZjHXnySud
2r+QNaYakRh2klLvHSli5+95LwRO9m+ZBhMzr9Y3CanZ4a5z1DBIVgjQDZmxmb9AKL2fDg2X37TY
fFsb497uN8dT8PUw55rCLTdGhr77wORLObPjdlkz9FVpNRzBaNb9Be+wxMFEKhCJecfBy4VsrT2G
SVdWxRR6N9ORZH43H8WaE0gTxlD8zy2YiQMyqoE40hLKuYy5YYACWqvlehzPU9ufJPFySWB9fIc5
OeK8dkK1e6N8UosPCIDXAnKCRp7ka1J4oO4DAbEngWFnlCaf9+Y9weD7JkazKQVYF8jqt5EEKksB
qiD0JoNZ3lJ5HdgpB9lP2vgXpsMRvwBdNSkXDKNBfJqA5C6mRfJvKImz3fDNbZBbn49btYePz69c
mMZROnyCIE8h+XwPrZzzPiw/yvp4MTUGorTLpLr14gsWTEfliT47PbSMdCtHdoTUwgbBOCIN/DXF
kkamKq+6VdKTfmC6s89JLD6kriVUptGL06RDLIBbEol3CCOGM+hLKipo/uF9qwCFsNwhx5LfFUnJ
B4VOBJ7HDL/cJzQhRkjIn8SQgM9w8ZqAkt4bflsavG9nyp/DRDzuOa9dKxs1+2rhy14RARE1wgM/
iSXrHjdiI9sxX95q7r+ioC93Nshff6buSc6Kh18e8GDZtq8OQF+UoAwmE06AR6CeWZQQzL6mHJKn
uNRLbkkVcZBrUmHtfUT+QHD+43nMeRSq17ne4ReJYNvwY/apNhvt8JI7vsFRRcJ6/H+i/nYkfLY8
G81SPEUPMh3ZAS8MsSWcNhKNDOEDcLTp9VVGGWa7UMGBYL7+q/zrC/WvmvhSg3ZZDwMvsMIulnzB
CqDRghvIkh0bUwrBTGskXVOnVLepJH/coLUPr6WoHwYFxaYolQEEuiBbppt7he+7wC0FVuvu9M0t
lV7dv/MpsL2+W+ZSuuZUKDyB4D9erGclEecN35o/q5aWprSREOhqa6RNq1HdOyuKfsyS5RohNaXT
TUP3mA4LcvF2NKCp6zMDrIdmbFY1jgK5lPK4CCCiusD2tbFQZ1Mn2Bk4Q2GZPk3fenrjOAUP7AqH
mEhUwfNk2r5NnU+nExeDLLjvs9uE8ZTURE+qx9FyvMLZNF5n7eY0HUYSalOou+OLKBjaL5DixWZt
c5VgrAJRka15F6YHiUohQ/R7Rn8GAUnH5SNfQPL8gP/yVaRgU6KnnwbsXepZkXokx0kl5ZAHuJWb
6hcal0jSf45/IvDkMps10EGxlDvNly2SwdQeMqe7FSiqRNGunF9npZjJxjR/UJIBi68uXCdnLZ1Y
c9mye5A2opNuzclsqjW1rDcMgMbqSr+JOoBvBDJ/xLDoV5cPb2L+Yh9CBVsaHsJtmwUetk8Rmkx8
lK5lTnS+m6q8KHiM51eLqyu8n/T0Y8g+aOhH+HVq3gNGTWQ3TFuNI/Mk/HOdi6y1IPyIIpNzxjsW
inbg5mhH0WutlP5BShx8eZ9OBgSYhftgOLo048UDM4OP5Ze/K1aJcHgjyPIXz3mWC1bIFj0/UUYV
j76T7aQU2CBGW5zYJwLNNdxMx1XA2af5ANs0ZONhDEuMJswhJuBByKnSTkEWJewi/9AOZ1WjI+gc
MG3qxty6co7SYoQRRaPA4d4p/tdyR5C+AWIn5jKDPmo9u9BnUK/TtBQlfFw/oIkXNC8SpXk6Yase
7Pb/2RzhOLrWp2xreI60RgeoGR5ET9oaL34hQ65rPDW1oa8m+8U0KBC/BBA+YIljz5F75RExlxq0
qNj1kdfD1Krw7OkZhVWba/J+y5+3ZR5SbkfHuOivwIlmuXE1Ve+LpUFV8CyXs9E3ogiQ16OsvW/N
KpxKzw8YXYtTDkiZlHbplKu0h2OrQttX4PjCQJIqMoenORz4ktWxj1oYwcK3dTziVr3e7K/Vkdjj
QZgrEGq8ph1mHzTja1mDjfGaK5nE4iyY7gipA7P7ZzfQLRf4Bj8X7LsVEfaP1QHg3JbcStqlxjcm
lOOwBQ9sAITlvu8Q9tekWMhWxD2HhXgGh/q9Tm0GjkX0y13x4XsZ0RqdQUSdhwdMx4MgQvibMtEs
UOuN598TgeVQPFeu116M6qDF/bu4ot2Hq5ZW9IcJugN0E9pWFJ9IPJvEAczZ3Gv1mXcowi7J1Mou
dlEzzHztTl5poqOg++Yau4YVC8CW6v7L7LoyKHcDiJiN3u3XVLgHrgptnC6NXlXxoypWwLMx55Jt
Xa7pP9iHm/+qMI8KXTCAtMjZ8Bh+cd9CK0Zpuas0+nejU263O0xbu6kRSN4pRYcyXs4+Ume41HPl
wfQHu0f2m3efOuylDS0jKEtoD7XKKN1kJhl1EWJRllmczkr9yd+csEjfC0AsVv5ymvPqANnBrM/z
jvZTZdqKWZkn9AeJJrDQzsE7HqeUj4RXWgyLdwhM49NOfc85Vj3+pI12VxuClXv/qHwpKOlbdsXG
oLCTxRN5bbnj97q/SQQsUkEv46oHXlre3BOLfOVo16PM5+rHrQs9iz4EoJOyVPRfwuYncbzm/l8W
BAM8Zj/6DAbi0iUWuYnTqfbfQvhgGSTlB+xlwqMoyFopsMAxgflqTn/FQOZvzb+vrm0pY9UO1mLt
38df77D++8UmuV5MwEKhFiad28vv7L642ythguN5WTPPsAd3CpNX4pdesZUiHLq+exL/26gsrzDc
gpCgoPd28dcvoTi77YYPoYOYFwoLzutsvTTUDnkam8HwLl8gmVa7OXGhXeAsrufSxPUTVxHwCly+
Fmch8PTkKHFMveCmFE4b2yTwnkWDIvNWUxdgvvzA32d1BPyy4ANg9/o8+nzEV7z14GtoRvPd6IuZ
WWm/Ut5IfR5o5l+6SnWTbs9W6eOza38Q31OT2JdWGAPZwWvlaOIIeQviAEVxs410jlz42z1LBMfR
ntAF/KrxGwiqvHfhkPlxGYivNdkTng6X8Ff4tPrETQ6OQmUyTHxc/B3xLcrS2GFGR9PDt3YZtbDD
gAjwy7FCl0K09vsn/egnlkneEbO3ta4zbRMuki0z6aM41fYd53XQbgCoBxJIWlIS97K4diOqNF6y
XPfp7ZmElA3xRuyAtfbLKdA8grg8PS+/KcT/f3xAgX4O7NHzxFLKrdLYr8PF7NljOLSQI55EIONf
DP7AOdrL5K0t+6ulehqFb87cvl9BY0e/llxc4OslWv1ZrPzRJbzWuJhIdnwujB59R1A1moDPLiXr
pyJvEnTSzUMTlT3p0lbLknct4wnlmyIl3DBqw63a6P9vfZNoCnCimLDgXetarAcC5ryFGO08SsNb
BXDYKO0dt1TKiV2Qt3WroXGEdDSIr6tg5E626rfyy51Y+ludX1hFmFrEK9tOkPfQo5PF6eCIUPs7
vI3OaoQTTsC0Y6WiEQm/8PcemdynhoWqZ/0Eo7RS/F8qXYW3mAnD0sTYeiuVSm0F2KueGNDoheh7
gzglwylHSZCnmpbHOSPwD2aeBSQ+KEbTWqLTWmfZAnIogoBb/t9iGkAlvsdCS+GPcsK/3BG0GPsi
w5JR8ulVzLODn84bvPlDwY2K4rnYDMUKCUMGMbPRaSBsb9vd1nZZ3Y6hqmLoQ3W2LrCIdhbzLw2j
bqkwG8qwMNWIq0Fy9uDdU/nTeKVxdzavSol9byisIUv/+NC14LR8erIcdMH0e4mbOd2Su3Tz8MFK
v5nhgnc0AQPalXi9BFiyTVtwohtIt73BO0ij5P+ZGxMgrJQkEtbhiptdBYCiF3MNlzmGcxZaf4JZ
M03REp/VvfBciNag6C3jQC78hVBUcJT7rnYPU1IrS9QK8ZZ9kQKohl/VFYk3QZambBE5avcVUUmN
4vN795O3FU+BtWa+g0xY1+peTgDnYlJe5doo7i1yZnRIEXjP5pmilHOFtqjyjmC0yw9d2aNehnjG
A+r/e7gaofPcARJj3FJa1BgKEFup8QdvZ6NZJTMhGZeJ0v2SbtZD5QD3fjAWxIidxZ8aCz0bVKeL
VWBwYnPW2QMDuSmSu66JadhWk1ZpRN5lPnGBt3jtJbED6BzlD4BLGsap7jvtbGa/t8oZnbWqcz18
B45yTSzvmB/1QKI3KVnTXXDmu/6XyKpov+m4Cnvjvhc0Gi1bSMg54NIIY03VUf5VInQWFcp+g7kC
XSxQjJmo/J0/SGoIOhiVyFB5wpdo64D0F7ad0qpan/HK0JhqHl1Ito3zndle0wP3OB12sYVMoChq
t7nT6VFRnOhr1y66w4qYRPBC2l+9HYaYwewxbQUltN5ahWYn6n8hLQGx+9raN2FRO5qx8TkMlxdE
cpz62Xxo2kXa2/VNihz48pDmOYYAfUIRI/GrzPq+m1+lUKTj+VXILDYPA/6a4+sUwgmBUg7vd3k8
bgMzw0/AZmP/dvBDYzk+nAGME1VbnW6VJK8U3wPF2WKndCaPJp1oTVUOTJMi+67vAEADNbMeMv48
5mpeSMAm8Jm/7XL06H9LZcNcHoO8CJpBlPMHKTO1pBWO5PsWrn/fqTq5Uw0tcuCscsNsQL75gT3A
Jd7cTBCrCwIcEMLg1OunyotaUD6xWQ+h3R5wNVryd9aLz79JibVxrRJIafO31MOkZ7AfSyGw8GAl
Jc1IdZc9KAoHVrnUde5JRfeQW03qfKCizd2o0yYTefSTizs0x/0ZWlAk+OsIMZMcu2sNhrZSBv6x
njwgVgSSFmKZ4LIFkK/21Nb5fiGltiWGexKk74zJZadS+S16a5nv/uxiA600oKAQworN505UAQWH
ZW8p+ZaGUCPK5ttlEDss6MMtUwzhGSgulCdZuVTqP/lm1gIZsRz7FUTWoBcG4u9EPqhLDnUr9ez4
YilB1sR2fpJnRMXbz+7iofqWULffowsbOQU3zjDMG5TfkkMft4r5OskihzNz8ruLFYUxrcoOHlz+
Bwzac+2fVseJiK3oX7zsaRZ3sC8XbafWhXMxoDFYmxRvnDcDh1JVX9Vzyssff6dkaEc5lVlKNvjY
9yyUJ6+lOr4hAiAnXtrgNEH9uBYR7TlgdrjzUcTjbzm+Zx+tXmIpP871m6rkhrtXjGd3R+dKqeqH
5X7NFU2YNsFcfKsB47Zc35751yAlbG6HI2qLDZvAAZJ9l0sJCs6b5RE6PVZyhlK3WXs/ZQSbQqHh
cdU/M4GzkM73vAqTvcG/PRmRX6vEqPF9sqR4o+sREX6hESdt2M1yN2rRqi6SyCsQ/o2ppLWqkCM6
yOsEjgFHM4HDI6BWrTyEF7gHMhyJUqf5gd1ks5TRh4m5ZmXR4gpNbXOfx1xJ3L2js7M1qeqeTM0H
Zm0o1BTp2uovNq4SXk+2jjmjsczsylk8W0lX5xOrecGEHpwtjxdRE6aE3/ktf3KduU3+ZmJ4wCo9
HGRO3FY7068lAsg/myJA1XrZWGTU8LDk+B8a0D3jGPYz5+qgTCXhFrSW1/jPKOEvoBXBPlPweQx/
nrGc9cbUvioUfRrB5PTruyZz0rW3Ke/varqD5lF+9LuhvxoJZtEq59BGXjmn8QhWjn0GOVBjTpuD
YguWE1u8W5v39nD2EcDobKbkdyOeu66pT/NnXSYQFjwZcmsDv4br25G0yqlbAgVvTb5BRWfnUo6i
YkBmCtGwtXKuzmKuZcEpny96I9nILhi6UmxZAHrb59mzkvZTy0P1z2gRNku+NQPESaR+Q7UbUYmx
H8+1YAcJhLLseXOD88umxUQXsPgXkgrld3lgp9C/N6zdyPBx97ogo7euHRbrSgFpg2XprpoMNxga
O74MlTWOgO89X0Gri9gync67pDIZFV4nRqs6Vj2Glth8c+gnl49v2Vpv/wXsrI3vY7vI+b4ao6Ed
Rp7Uy0/o/hMKaIs87plc65kua9/b0JI6mFSJMKahMRKz0OT0+JnSZq9kYMLeOYe2oI9HAEwbyR/F
2o4/CA25oCOD4bS43Gt52roOPgWt8IVbI2qUO5qmG6rgDSUKGTKqE6SPK1BIGGVXlpHgreKG92z5
3nqDPz+WGbjTYfQUukf/uH+X12HJ9rum+9HuYMh9DfBQObrG/daio+jKbfHC+S+DIAsk4m1MezD/
0QElKxtWN29LL2pZ3DShLVmz1bJoFLlfNBBZwRoP/hlM3J8q4iM8lS88dd2l+wwKje06rvfw9YuK
fIerLPL2oiu8mSbBtb5+k5fgHphfgCMyZvpQgZ7CZ85jUng0w/IKlPOzOedL1/DrKVJg/TzraiCS
u3OHDZ77t9VOBP++PnqAuXTDMlRbWl6vbijlUoO+RLt4VQAGuZh6NXHifcOFJnQbUexDAeyQ/C88
OKKIBXVOQoWOJxPW22Q6qCvl4Hmfnz0zfbOfgcZ2NdcWgnSWCzdZtHXOFgF2C6g7OhyvAY4erd58
lvsbgP6+lsqImzj+It/xO+q5dl492M17k0+hyLV5JSfif95w3ieesvMMVRpjdp6AazJTewBvokTF
nfnK/4T5Bk/duoQ1POjs2oCNH4h76EHbAiQgI38SBDve5MMU4juhetei2kjWDxjuAW13UP+d65JB
zvK6d4rv2ig8G50rXW0JIFDW0PbOIt4w9lJA5Nj6NBpQeNXoBQxmbgIpnBftg/Ej995mzysUToQw
fe2NlyxjIoYNHevGH7vfgejdwdHUuerQArClCMeDThILMfeQ0MRKC5SnrZLGgKEFmAnjhYYY64SI
pJV/6ABZ6io2Su0pMHDLo9lKgCbEMMvJ2aeoG1/NyUdNWV85WcHkU2ayEAkfgxA/TDv/UnLns9PV
ceRWSWYHVGUxnCD8bQr8vhF1BjLtF+sk92Kb1dy/I7RLgYAO39vaPnEQb2kCYYlpGeRYRo6e7NP6
gH8HboZ7pCqmE50FIbT6CoqNDm0oobXjVWHX5jQ3yZLhU1PgyPNi58FShydLWoU78l693jOoI9E9
uz6Ncnr8V7wiXDQ2w2GIKwcbBvKqqwzQClV0pt81oskqkYdavlaUA3HUvKChivtdr/6Pr88JMczw
psH1nj4Ozvsbey17grNZLq2y7YEQIe98vKktp0ApwQwQpufexYetjrJ+fKWJIysv4+Jjh++uC20g
vVELqjdV/kUnJyrZWwvyU5pT3j3wdO5AxZ41YUYnUH7s3javmupg3z5tKXAK5kIiOW1O9l23oR3c
7HnLnfFwh6+X61IEapv4Fk7LWUdQ9YauExRFIkD/hi4MTnNg/XqxF791AFdEnFBYS1x6il2OeYTv
Vw4iT4XmrxV0/t+aeIG2or4xxOUBLMYnMHAwFJTx+6GXyIhXAJt+hQJ0ogNW9ABh2MHwColDFbSx
mQhsfnHkLfxr2FvotFiTfgzynOC5vAMdMgkhEmtSO+5ktdCHAwDsTnS3K8s/xDqJ1jDVWaBXRWpa
kkqU4h3+Bbqt2fwzSESKF3rjedrmRxDS5RK2ARBjkNNhOo0ItCmLG+1wChtavRMritP+9FnXzo6c
Blp3wOMyBEhIdcoZJQoPDo0CRUiqyIrhuNma+oHtqzpghpDsmfRw9AhNMgykoll86C/3nAg7fHgd
GN4guqexCKf5Q3APeGLZ34uuAXL+efAGr7JhuLPCUH1vHFOBUvtIzGofgFXfjFDwRjotdTUuDZ+t
MsgWkWUeyOiESErbjg6IExdKkhB3XwUFWCJoJli5oZZOPQNYwVgb1rgSVoMD7IBHobCanl/9vXuO
BlfnXCLSTOrIO1DmcawJ89BpkXoIlQA0VQDcpnexbxp3K+rASYVEW+5tVoRUpAaAeN/rKeeGPnrA
eldDaI0DQHh8YwuWqVyRw4R6YNlMxWGzknL6obggmiVzf+j8hPm2sEgvrezr4ApiCovj069rS7ft
qGm7WIxmaxWOy5MHnaIK10ubLQHjAqkNCBcUMTtlcy8mQos40x9dCD9oxOWdW3izC7zffAUiIf/i
OaJBRO1CzorzFCY96gDHPJWFoTCuT7CgRr1VCAoH69GfQPtWRmwCLG30OwDesQrH3Td4WKcrW3Ep
PBJ7Ad9bR7goV+VMXDOmf7C42X/SoQNW+XxDQUcXK7cId58qSl+ebvPAeM9Me/oE2iOAvyG+H8NL
nuBc7PjLE3D2hENrpf9/9S9iHsFLueumxLCkdX5EAGJv9eqYFvJQ0UQPJzVX+Ez+NelunASK0pgd
wbnDGm00D4OtYIhNrqITCBVbOKOcEuMaW2lIPpx9vEA8GPPP3026moSlEha53EdFIIen2LPYUFY5
V7GdGeqFZfQpY3x+za9ES6ZJXbrR2vqOpD0kketRd6IDuJ53eu7gKdDzMnl78QUupPHRxn77tDLz
Y7LS8yjMYwAMGvaIlFup10j9SnMfKWmMa3w+8Hc8ONOjBHNTLPNy9Eo8BtoMBCo9no/vu1QQ3GH7
hXHJsSLeUCShQhOXPa5AYEgI6m9w+9MhrctN6vqOXMr6Kzeb5wtzdxW+ZecIXsROUas+lsf6Nxtn
wpRj8jsYDaU2pPjNewHTGzQVSwXXRubDS9nAhiW4a14JK7xLqndvvCBOCsGTzdQDxX107XUBSrk1
hRl4FHVJO6wlVPis77NaYZh04h1PMxWdfkd+uw0zjpms6doOgR6VmvbMMltivBRzR+1NExyDsMdW
eD305wJOuLJjfEQcIyq/O5b9isR8i+AeW6yagt5RaNQ6ZNfurKktWXy/8ciaUdUV5w/CDNm1wliC
Zcp/57TfrqTyz0go2fIH5m/ZcFvBkUBEv5rhn1SQhs2chTaqreMs1EPGxhPrZ+SntoJ9rfaQwX0O
xcU6cXmA5+zNVDLyK1Kn7YpGs5uwA+CcP7gTFBS5kzcd4Ri3zN0tSCGPzp8vkwOcteINT9ld6XSp
zO4SC3o7KMx1h6IeRSVBENX5nRXGZFSp1gkcCoXBezFi3kepSrV1xvpbgdmy9mO/cM6leEkGtw7m
9V8WuxU8kJbYYD3Tnd8aXbjCBfpkk1MQA+MkeiNZ1qsIWMZo9HSGfWcekj9gKk/yjnSIgLedZX/a
xjAO6b7C9ml3/VRpXI0EXHvhN4tk5H6tFUWeg+LfDdDLvqAitii5ZZrXuZbIAjCn1Ggivpl57gg6
FjP8Aap69YzYGEHNmyVE1k6pLC4R/Nhc4HPttEP46ySA9y2atV7EVcoy1P1N759yx9ZPi5xK++EM
FTRJk32sKqBoqa8WVYnDO/x5maFYAQaVzdpkPKQOQcxvA4GBlywI8UhScJWTgj5xp4I2zx/lsf4t
hBwESj78oznWkNTeEp/rvbr6scXsie9P+G3W7xAtR/p8pWrmWYp7ykUaXBAtf54iohhAeuysflU5
+kSyCZkWF8XMlFnkAVToGKx9R9FiZLwnGWjYSw2JzQZQL7oJ+eBP3qqDOn3Rv7TTLa3zndwKPRdD
sZn08vsxoy+zWtyqtEM7uhHJ8msbCXXFlJRmWULAYuZiT9eh6UwRmqGSUk6culYz0rFzBIgVSkec
dz8ZuPYwsv+2BXlPn5eQJG6Cp1l9ykqWXc8tXihirf51v2vtkfv6ViNAudVr5k9+d1RT1yrlsYYt
lWdeWmL+aZbwntoWiTerM0uH0dfE068qEdOuOz86hmEKPg5+EWImMJRaAikzVdoiEsaoQC/yFdSU
0CnuRmLYigY2N1uQEzAKEH8Z+MzRbzRHrOtcowxZpR2c2xNK8tgeZ87LhL6yKaVxpXJEPOqEvoqW
JZytzJ2v2Y39MdLr0WP7zUtHC7Cu+nbfDwaU4nSGW4REXYe1cbGJfOss4FK57ZX/lJ6j8GPlltLU
6hRL84VxEq+3HqP7g8BVuKzFAi6M9qeiXXPMzVDuFMKIq6H1xKr0cPSkUq7O2amsXp2B4ffQxYK5
YxgFEvXy6ii4we8vPBEH577n5L8Aaeihwt6505fV7TmXEIStmUOZuA+HxWWGGjmYHKLZrtf+a4s5
81rQtEfaczR+dQHbuM7Y1+Ug633ywEMvFZR70/PKv0E7ql9aTFoBELBDJk09KDKZLTU7X4A5C+b1
zsqlb0u0dLd9c73/dsThQ2BYoDbkgFYd/ehmTXSo3HpNfzXJxSQL6agCldho4GnWXiKnJvHKTp7p
UEltPRVzg0f6bnK9+AvDPGOh5V8Np2Pt7HycNHtfxwuxALXYU9ItWRAJPzKY+j4Eg2eYfQUxBoKg
Sp87CQ5bpMvk9Wh+nKm3lcEEUIQywB9/t5C/qDcSNtRAHQ1YYnkn6m9bxjN4vKokAzOO9QNPK8TA
UHPeFjLWooelWvVGDe0CTTwBSdaFfvQX1hWp/gcyynmU2iuC4cWq8BFGa8+ldWDqAhwOB2Lxihzt
APyrYL8rpFw+dbzAIAFPHRnAAS0zzUtIbJtH8rQF2OfbPTi/kPC6CMaT4hafeMBygMPKjrPvBzaU
FjecJvP4YmeZLuq90RA65AowTT/Y6JLkRu51uhCEMIviErpmuqpev64it8ZtAw/1+31BCTAJRIbE
2kt10zPghzqYoDJRJInf9qx8N4fqBycQzHfdMXxUed6YnJhAjtpwkpmcfjvcBgts+bP5dqLabZtR
o18oLTTL8lh+8nQXZ/tNgOLKgmyl1d+He+dgYzSczCJBxm4wqGAEQ/KQ5TYTKQV6Iwpgz2HrGzbX
p76+TBtTWCgzvUK++SkX07s74ZxneOJiFOXvfEEL0qj8y1rKTFJAesXrK5feIIfSvCnkBc1fXY6x
Iow1vPbok1mfMxfGvH67FyfPA2S3Q7guINSbJzKJiiuqDbxLBKykjbl9fdp830mn1lWsqXPqkWu8
FpY/uK6c3nl0zPpSI9Xnfd0V8KjpDOqXpvVoF8xLjI4jw19SCyjBpvJwt8Xn4ST9k7yJIlZk6rmP
iykMNhY9Lw2aypjxj99fy6hjxa8OC6KvMMzxF2SUfzgLAoPq6xsNuUYl2y/KStRuJFBXIxk=
`protect end_protected
