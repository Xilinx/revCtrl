`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 81728)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6u1
ohLKFYtbCVY2WZpIcrI5sGMANnIGUl00Lubk/uiRZWwylQPRofhtbxrmgqtKEl1I4qq7lyyg4t4/
vPl/2DyUjD+T6LY3cj8Vnccf1dfyNNmacsQmrpxTCTcm1rvC49XB6qq86h+BClvoCmag6E0KY3qV
Z+rzQwMMqpmiYaFQ6i8WJYHvAXjEHfLMd1U2kM3731g+48CUibsVfd79wuu8xSkJdsctcoyf0siN
LXoo0wsUO29b9q86ypFNW45Ld75LIfNAm81PAiDBmV3mtjfThjlQBWOWNDErATKCbZFIx7UoBqlB
NGpKMvx4n+MR8Kc0RiATAhDtFHwyH0dfOBR8VYtwLbg/9PbOiR7HlXKYQNW1VuMOdUOIXAaWAHTy
1IzUi5r3q4quLWdOzOLiLUYUZ++FWPvDMo4ORpuYtG3tvQsrdsBiFUopSCMvfEKnOm/fhzH4WFk6
NuZjyCs4llKPr2iGoPErqCqaIhi2Sm0YBOmHYuY3l6/vg6BHnPEUhtFTkKGsMWTvCM/u4K8cIGtC
BLxmMo1EJlTWDT23UudBkE1j656pteAE68UiJ0puFAWmqS6zRBBBh0DIBfBijadD6dwIUktdXTHd
eS75NR/URJ9e+TCu9hULKnqRYknkxSxJBMNcS3/wtyz8JTgiVd8z35GxaDLbobMbYgXZbQFdIpoG
acmO5WG9QPpfX68zAiEpgSE6lm7IMieAr62jF9Vo3PjNsEir3jVeoizZ5HfwyIncOxqR3SrrJiET
vs/VLcQGkb/HPHBRi3OeAo4m3uSDGpCGELxJqFi7gTwZv0HGNWT08t7xTRmR4MKVYmHB4ZWqHJbA
MG0ekFvjkJ4K67K8e8mQDzBj6Up9vn/t76oouUTZrOgqGKxOTnh7XzFeLWiy3lVVaDl5G7ZCLgvC
T9uUdVP+U6fehXsIr29RH8bmcZySo+Ovgc0Zj9Pp/xgpH+a0RDQrXHQ3gZ5kypJ0n4GTYt3sn8ls
sR90EpWgqy+0KIoYxF1TzbzhAkoYEajKMyOOCSNqgrFJvdFbySnWTDAbLYhnmf2yOJ1vOHsHQhJ3
wi+OVqPe7njtxuEN5PtsWIUdJS10QvHCd7gJ2O9DusdFG4wn9gur9SnIGCZ1D5EQWPbWGImYZ1CO
TMnJmG20YIXIfrbRHTLAZfDFCMbXQ6NvN1S7sOgfPfvjVEcuNh8R6txQdNVzETueo8AzzVYzCDjW
abT1O7lu126RVu+6v9QSHEO7MGG+2IK4Cjn6mDz4LikBUiWyACjzsvv8zaMV5EaDpOfT21af+fjj
NM9W7gNNj2n6DKGIlCufIbzMUgIVvAUXWlGZQRcrOsyvyA40onaYgIFnhNeH5wsdGUES+CG59pbU
QeqTalQafQtN81dsfBKLZ6z88p/829vRhqLLZnGUEuiCF9oaY5+aR5ovJy44JIIWEl0kz5fD4ZYV
V/3AxvHO+HagyrDD88pwSU84D69xoHf+CzOevaNSv9X+TjSgwH0sPOlMMGk8HJLdgC1y4WhKsRbs
NVYAdxuhfJTNpPyy3JV8p8hEs5krXg8ToBWaHE6TAnuPHjvuZWQqIJj7vNNI+1MH04q0Ud8arLdp
o0C3U4YVv93PMlv6zxbhnJdwU5naEP4Rxf0mMlqEHIUCIW2ihGbiFIi/OaVpvTWlbc5wiFGTcb46
Wna+1rn77rH6IX5Sgx5N+ob1vQIMei1vTdKJpJPklJwZqHWyCFevlTxF9AGYdn2NzFdbPkJ2TyOz
5SGZtBvavQx5zCj86fx8UY02v/yqBRYNs7YHuwAB0twVdel7rPyYSr5+6OkCvj7Z+4xBF4W4+ymD
jv5KK17r9hNJDGfzUdej6Z40hdeJDLMRNQQckkJ/1qPHcsfxXffT4pUOfXVXnBq3/yfThrXBsxNO
Msb/H0c6BWPDjc5HOXWKmffuvEka7Ig/rd73Fpzauk5GV3SchikdOpP3kt00/VNC7kOJIdoUsxnU
qiSLHpqnrFWjGy69Txm1Us9K0ncB18HNlNWJdE6mDoiG1pPgjpI8Vs/iVdJ4DN/kHnz7UwTPORdj
kB5v3g2fuKfeNab72mO6HrFF16jaMnWTYs2Pemgd1ObgChMu9bSFaPAlNWNm+POtugAStEsxHF+u
4FSCf4bYonWz+VAY92mPIKC9c9XzAmgY0cQqarzqCRThUdtbc7h8o7Mrq2JsxdOQAsKDz+eBguqx
U32Hys44TyrcsWmnoJDlpuY+7/yri6VVYhYhIMQ0IvjD/mm0HnUFiohy96a296F08+DHudpxLzGk
nrhbAS88MpRSIvHlEroWiMbtnFBZlIRaRqFtwM6xXmwXXQvmVMo/HJSD97MC3e5YKBXnqX5y70pR
vsIYGf0M2SAtuPv6Te8ZqTPilQ+9cZTIfxkgSzisaaoA1kE4wccZm6Lj1JlQvqtg4qR8WhOK/O7U
Ip1K/NWVfZZTinZPok799RJ5BZwy37OUiqFXc7VGKRVxOAwh32pOh0Xp9gzetyjPC9DMVwT7/D44
5y+UNrlGUPx99zCLNnnQqLDzX+qOSFAz1yJbgrd6Z7oyZJ5yb7PFz/Zpgj6nIXpV3LB9IrRr5YUo
52JCTqjsaudM24rnniPjYer08TE/9xZ0SL+0ZsdmGNqBZvZrw66e17vh+wryzQH8cbT85RiuvqRW
CJ0//1YTr43tJd1L8fZ6XFtFMPdqi08MFiAWDjOvrj7K6a2pIQvp+ob9wcMuDmCIKLTOwmovcs8y
DURuRyX8gHAHzCZoQdQ0x4dZYeH7b7bXjx6785FQ9dMXJG9P+U+jP8GWGxxlhyev4D/nICnrvcPy
awsp4jcdHXweDqb6Lvo87MKe2/SSyP5nUAg8zhe726ouKUTVPkhaHT31A+0MLClIX+ORjcIYNepd
S4yekhq/NbG1jJzyl9UeZZt69O9DiwabM4JJzcDGaLjep80z83KNyK/5NHIwpaTDlNFgot94HIxO
XJUjaU0kVx4LL5CxpwbZG5LPuei1enXo/7q2PYtj8q0U8m8sIhmdbzVurXQAKZvVgvyLJwqg7ICV
kH2g87KsYYZ10SySsNnP1Nr5X6/fHUvYda3Au5sIwPkMIqiNziL3K5LQzY+DcUIH+zX5Muzojc+m
YaID5sOX9sOzLWgZLcsbfhHzT3AW9KB27neJo5fvGPOZ+QMnxVxzzte9TK3TEo3DjFer80siT/E2
n3gIoBIMsvN7G4LA++DrChUZydDWbD5rUpxb4wf4eKqxmiqSyAqpGIT6Q67QrcASwaVnwErYmeVf
uNtxBsbl0Ps6LQivxzI8574VZPbTQqrjWolL6IfmgiKi/hv92EsL9nhveFH6GUhHkkhlUojoNedy
hoGFp9N20m/t9xd9N2LweGHmqJCTaUKBNFLtb1C2diAuiQPtsQUZ9IfA0WYLFMqCdtono6/5CGEy
Nyq+F9pPYFn+yKQgPorapRLfA3OQmGCUc1ibc6EZ68h82UNveBhzKFumwWabfEBQ18mqL6vun01J
cYT2Gcm3VNuJ7giiNDIv9j4vJSW37i9Dyo2RnqrS4NOGasv7Vt3O+X/NTyhplqJeR1dhyhoLasA9
3QvHBJh5fUied4UFBltpVW3KeNfwq7huzREUAdtTZoVtRJXspmcHij3VMDfeD0BGswF9o+eh0lrr
+2CRugaav66/WSh0zyfQ5lXS9NVCjm6c8WA4Ff/CX7/gKb2/8DH7rkhx6B5D6xIp+2nIl0YV1Ruo
IxKUXf1moxuaql1FO7llonUl06Ca24FN5+fdJAZOnMXQTYlV5kb/C54VhSa7Th7v8QZwgMjtMbXZ
KB9lAsNoeBXQuPQioP6Nxe0gDmXPAh1JA9Ks+UsOpEvgRUUxV6OMjymz6o6gbNN2kOrUQvA9TLAV
aCMxz9UE+mBSQxHO2dlsLWGO4yhIjkCOqSNgcKqLLMy5zrO9gf1iIKW35uBWco3FEidDcnXfuDF3
Qt9cPLfZpgyhM9jc3vpXVV5oskV+E4q4KoSyouHNBJga0VygCIEXtOgbEvbJDCooDXW6scJihfI6
/JmhPuwCulLjJTmAnApjCwloVPMdT1Wn71P8m/EFPHgk4qfDPWFNXjVv3PYr1wnBzsG6FLZxJ0kk
dZEUR7a/PpCWGT1qUV3hT3yyGDDsbxSkQSsCmhoaWtnJ1bt9fvh1tKaPShNPpXgNuDnPmF7U7Ewj
DnZUhGSs9Qh1HI15fHX4m89TRZElISOoL4Ynbt7Rg5/gBm8gjSwEwZdiE0rRm5hiUpopMpo+HFKE
tOHA9ppOP0xjFFK1Ud1ELP4CHNRsRznecOtISy+4VrAUZ5ORDedYfe19hy/4TpJAibZm7uP7lFgL
SusIfv0sb6goL5EE9v5nlGx94SMoGnjrgqN5FpucNWK5RE4MRqzkcmAlOIs1+IVNWqKxKwcvMIf1
CkVUJ8ivTf4yN1JHrBOaZityCgDrHuPfToHXfyIm9HckP3fWXwszWbm4LrS8BZ9kmFRJBuhRN1FI
uIGLyAdqQwWAFWtCVXleMFnGo8Im2arWqMKoBec1Dtg6lyUr2f3soq3whROWzTtEyQjcMwhCzqjh
jt2gSIcHrbG4qW9rMOdaeDAsQfDMKaAieMIV3VLEdLmkCziJe/lZLKAve5NQkM0uqJhnae00Essx
+nrBRcinCsgvKW57+yUWdRkOrslV005vjxpfArfp0TNhqxYrtI+2EfPNwMbvP+8iDqVKnTsmjGCd
qS6exT9mjk1uRz+P4TnqRKtsrJuI4Bfk2bbj+xeOUI8TOyPD+UgT4ErWvACDRrP1OJtchPI4H9jA
TPNix+xbRGLzve+CJQoVQF5CujVPAmAj2JFA+QBolG27jveO4L/jZuEygw1PK4RQr2QMBMquGHo4
S8knRM+4QL1Dec1Nv7FpBuErRM7OX/CEg7QeZqmSvkCv0X/uJgLIuQWtyc6o9fgYFjGL2v/+cWkI
nwTWrS4xTWJmx3WcpJcU1mONpf8R90aXn6Q7YedgstEdiXtlPbNhwRKdjZUj9h5A71DokKBHnAHQ
LB9yLdsIi53zvpUGMddbDFE4yVdZ7kfivbMGRXwBUPe1pxJRZeTKb3AvZlKxKkXdVPnxbkG12UDw
9Wk/cCga2iTx+Oy2FhPKQKXWPwPaifFMmq1jnHPPwCGr/jAo6MsbqrU6Jh5w0svXjUZgM/r2mCt0
zYYAqgBueigwPhdKHiVwkHZMpPBARKpDpDFLn0jylaSL59aWnks/2kWpBElvRzQBwhEHsQX48MEw
FwPlZrn/bHpi7m1aiGcX0ajBMg8u5p9EB6uV4WO1u01BcV8pNTOMWvk5K6qwbCOvvFCj4piy5mBw
vXVtxUrPpGVZ7dHgbCyXAsGVCnjMixdxt6z1UWyW0Xeg5U0VqcJlmd4RZPWqZS8LLpvJEazz2wce
ieroNbc53a0lryK7NAEUfxZNUmpC2QvVt3QQ00GCnqexXN0aPN57snXWufEksldvWgLULL0FgFEm
jpTauQZF9R5ZNLhIcGG8s1t10t/rQUz7fY+LhQdEKSD9pDLfN2IQAqZwxw7u2718v3kwdP5RtWhy
zj6JyIfXXKfqjYkUUmo4/dhBQ4C4RPoaVGrh03wp0WXqfbIcyCOviDLSZf35blKaA3VhX9MLmOdu
QwjQJ4mGTY67tvog89i6l0S7hUdBzgkKYzfzpguINFYzx3+HVVrepk5cohfDFPDWa4dOHhefFhRo
Q/4yFHUXIV4lJ8nYt7ChN9D28b46ty1zfHIcvLQqobsoazGWRyytQli90UrY1ZME01RrWeNb0Dab
B4ltvHSTPshTX8Pf8UvKXoUmUaz6y/k4gKcDDQtmnHkd79X4zlkKzlUhkxgjGNw5HuZ6tpgOeIyT
VFoG9JJDwgVG59QszQEHV/+SFxe+g4+kD+2TwBfa34Gd7ILZMmCVoxioI3Q5hf9w6OQ52QdTRO80
4Hw5Qb3umJBLO9GQ0skGsnW7Sa9WJ51LMsNCbfpGaMsW21za+1i86LP5DbUX4kc65qxfCWALkice
6/7KUPS2zTklaxMszQ42AipMpY8IiayyKWVGVkRcIK2kJMr9Xr5VEdkE5pYhgbPXo8PRoZeQy0S5
MgFndFJ3nttVisjk3rgvAV3F1AkBk70/HlaI1P09BY0V+F/98E5pnnUilMJ2dMu3MEIZRRFhgSZj
wmECtGcwKDBp7puhT+E6a0sV7nNgysphRi8o00nPyO94GsiFRa9oGtbwoIaIDMBYWD5JiiSV+Hsx
/G5CazhQc29hiAWkhZD8iDStlbamI5sitXIfcvAsS7fQ9MewLzeJDPkPasL2JxlavWP4Fl1Seu1h
R7DWRZjuT0FsZQ+Dr8hqaLEh+TpLGHqvqfVT6ZOOK0ceu3Uj+lbru1Xpz+lKis6yQRidiivI7g3b
/5bJbFROHZr8LC7T+DrDjrcqwbzJ5ezzuCL2e9lq5pfBiNOfJ29SAvD3YJVPoKhe9A+0ZY4uCvWD
p/1pJ8tShNUYQbV3DNwQ1/DZruq6OKSR9BpVmyMYnqonpviukUS2iEMMR2nQ2igvJ5T3QU+0WR2J
nEU8ABSrFkDNMll+lVGe2whyV7Tcl5l6TG4QPL9iEbuSN6VgEuZSyFccQd7HiTqBtrL6VjA/n4A/
pp50CNAlZKvREEXKp9Dzn0AfjoRx+dOukjcBg5a8OGRgtOHCDGnYlnIXlw+0Gmb19ZcP8UjMoVTl
quf5/5NtLU2gZyCHuL0+qdAwguYBBdWcxT6iZCEBy0MGVcmuUEvKlCbXY85D+13ceNauMLUw6QE9
GD1KSdjS/3HMZsljTOiEJXpL8a3UfVrmymhlOhZr+oTl+LNAVob6XB6n3uYs4FTP5Mio8VZS1D6Z
pq2xVKGKOCA9l2/YzOwMUEGUCk9BhowTk8PWwE/MR6kZF10dPsoK4xJ0PNuitMR0aCKGW0/XzHHO
RSj3t5AQNeJo059Q8hU//7albhRNbEaUstsPPC/6cJb3NpAdGokVMDmqCzHS8wWnTEa3mUUd7zjJ
hUgSSwxnEG5deEDCQJYRbtyeB1kpP5ny9I+0jPC3fNYUaWTRKjKT+0ciJo5VB8sheVQqyzZVG5sR
8CmqCv2CN8Li5u1kaz0Cf3BDfAgm171Tt4rJnefwfx7CJgSZqPy1Z+pD85JdPRQT8oEKqLCUM1Nz
vJwkHQnXC9+GzYmr/pLCzlz44At+x/fGMHt9eJTYqdqlzZsijqQSdMcztrhAOhFcCLLTv7dR7HlP
ufcx01Tf2r7d+vWZAA/EDiiwO72JRuw8J6pmOTy1QBi4AROwAmIIr1nQMIim0CXrqEeDEAeSuYKo
+DlJe+pTI1nhqmdnJpvBWp03WUCZ2uF+/YUVE+NypGDOUsyGOdzLT01xnMRswsXIVmVAA5C+tKX3
1OepIVTzr53PdUnZ5GxlheKbNypk52uwCllAIAg4Cm6My4c8Ul100gLtIDk6zS9sc0ur/lCvYI56
G0nQXXjMr6REqIfHlyqKiAq3vK0ot+x5RrJLhwpJH0WvOfxbcWSt73tsTTPMPz41H15eLjMtDtEI
KN8LCwuuB7sZvvsyTrw0pJr5XRp6qLQLmWIPpUzBWvLl6Ri1A0ghEbiHMtTpwJIw21CNZNVnANaV
xUKuaeSC6Q5hzyhpq4E1NeifLhSVci7/y77BPNvpmy7l0nWyihcmqno9NCIO97tDs3dSe+S9nNkU
ECCWfwH3sor2LV5OwuN5nOfvfLD/xjivoHW2EmZ9FwMaTprXwgWXE/dlB3HovTqRXwtu/iMQYtrR
n7sqWZEz8ftcPS95aXq4MzsCmX7ikXRjcYzqkcr9I6KgHX/7MqsT1V9fTPYYBtn3gYsJE8WpoQj+
OQcD+kYowejXj2K1hqgEl7mHLjnpDYH0c0DanmDBF6usXgZLG0+l/IQxMNiBbdfaoU+jounes+zf
XWUTW4Tp0tnibx4t/bhP/Bo0wQSnStEG10ejnpdepNzYrHJGIcRKUQgbbVYz6oi7IMFcRiX1NyqA
7vCWOIsfddYvCEVvZU/j9siScQrDX4da9GdhZRupPucCjzaC1yBqrgC4/zC6xouqSGVysSUhJhTL
Jj9vMcq37BmzUqDH8//6QIpDilhOKG4aVTKsD81DDwMSuAZAS2Kl5+0Q4DT0MeobgP4NxGKHq1lL
VkWsqdfOVbLRSJHjvIU0GC+xPjSCbIANcW6Jqna0Z/JyD5OQ/bXQm7JYFNxPssXCQKPTsRHYygBl
FYWv8+7SnMu7YGhhCLQ5VIFz8XGO6CG/T08uaSduQByjfmibj3pvIUTrJrMznRCjJZcNFxfU2UxL
zgqMav5yJBmfm2KDPJzzHg2yq484xwljGJGXdCGMQ4fTVe6ic/T+HgtLEQTU124gZIa1JOHYkAe7
4kt/fE1xbSqKuFDWSHAmNFSe91TsKXOEkijv9SaOhDFXu9zMBqvMqk/lIz7VnHQ0I2fQiYwfoxgS
ttCJj/Vpg/sber7S2zVY5CrELWhmW2SA0+cy9ElwEKeQ64gN2UZ1A9ai0AaKGF3Al8h+Bt4d/gIn
g55GkaOP1634bEX7E5imArsWafmdy/9Pc2NjNW6vRMhPOuYvN85vkh3ZFkXt1Tit/ySLp1URu583
zHizhizilV0ec//3gKdI6xsT4REVfAGgWuejjHF8/vl6o5P1MysCl1v8HOQWbPpxyhKg0tKk1p5k
/prEgyU53yIus0W72xne5kGaLtd8zeALX592TKZZ/naBzFzO0dm5UsayGG9VnENVHh4OjOXkPFQ0
ifS6pj/EXRGXT8K6hLzRvdlT3QsEgL8WgjqRJxBXWKQwX4gkhOxwXEYNuKRayVUElUXbdmqAwVto
GT0sD+xI2HMMqqUYRDsZG4dCvpeEhu05W26fusBrwq/sCwjMGNWRynwaZ/61h9cjap1Mhhopcbgo
MW1tQBAImDEG2HMalE8m7fK6A6eoGecQmz9cKAh43pG4rMrdvkJc6k2LWLnEI65RrB3DGdvbCMx9
RcawfwObP5zwh+uLIgF55tUw/lhsyWMkLSMbN06qFFTIrbaXrFK6pdqH621qJp4ia/uRWO5laH8I
HaD7u+Yv5KtHdtynlNQbCJVIccc3o3e+BH5UjlllcQMY9U73vLOwEh23lrcvLpWSH368zl8u5HSL
4I2SkAomvpou/EL0q5Fpg4VWtw2gGAYccs6q68mK6FW10tgcM8dLAe2fhZOD5X+mLv9JIXnaihtM
LO2iYXQjTB3iGCdzIi/BJ430oNZirbz3T57JC7h74gAraFk87u/Ap0BfK/YWHgaVIXwseHfaj60y
G8tZajPPbrSaYYYWfQcZZBjHxbvcz7XTdlKsYkUWeMtn4L9J7ROLeGDSmlbYJfY4WTDHWeyGZuJd
HHsIEfzG9WN3XspJgGZKrH/JXoHRS6HWpwAZDMyH8NiLII/tb9Ye5IpGFtNjyigtxn+Xrf1Rdfkj
rt++3HrOzmX84YL4riiZFsWDRmOJPWHtAFmYSgD9g6OTnKi+ZHd81Rw0vNER6f3d8uRjOHMv+5gX
LdIy+NfyS/A+GskUeTaBwB8d3klMD+m/HCBKYIu4LMzUwd031ePGbg3ntgycPQlqS4RHN4iYoGMX
sSFRb8NsUyBmf56rJizCRTJWc/x+1hZrFLxP+5yM1/TcwTQURg85kcN43txacjMVPZdxvR47mmEy
k2drxlepkHy3t/rZ/Rvz7lZE8MV+/dnL3lDBab09OojwxJQ7nEJa/e6v6cwkSRVXTMz46V+dmT29
NTlFlfQD1BpOLDgav9V+8dmol6dvs0DbGwqOhyY+/ECZdK5gv1eoipxWsIOy9HkGxnthdhvy8L2o
CXNxqATC6Gt1ZnCfW45jBtpmR3OR9Qs7JgpG1EIj3MoBq/pMpWYLk5uuOHZGEyuMTOAs2ry6TUXi
uHgyZZ0/ZbFLJF5u9/9WzaCU6dKpr6dpnXkHDij0YDE6PIYBMIur62RxKAB/J3cdWxTYwHjusMfY
LDrX/1Q6iyZ1WJx2DOpZE5A276fWJT5B3PCjpgSv9YNjTnYUZ/jZ1LMC5Pq5uP1ReVj5v34+TYCe
wyNqdnE8BHdO1yGc4emG4PrIrnC/+1vz8AJ5VnkByMw+iC5LlnVzQocnT1sknVn2Rns1w+lYi3P9
MiP46wyI7Seyt/ODvRK4yRaEMSUWDxfMHyyrKqiN1w/HITrCJ1gWvLJCeCgfvIH26wKP/cdAHfs+
rO/IicUOfTR+jxaqRYMvz32aKarw4kFxdfKHIJsa4jxySjntAeZ1iUSH7z3rYHejBskc+6iCObyr
9UmU/39LKQEZMmGRW9JM2GI7CKDwcTI84AU+byvnjESt9M5tUm5juP8K6DTf0lkUojTK0xFb6B9E
DRi+TWmyOhd1achUaJfb8iSboGdjS8mIXpTmMnL+6h1yFrqqiKWRM+fKNxc3HL2vH2B/z83yXkXl
bVVJcln3Q+yi3A4PkNO1lSkWZLCrYWxZhc+4cZ3H6AZ7pxARu2vhF5U6QjXC7sKcBxVMvroWZbtx
aZ5QgaVn9Cq89pqhtxWCDUe19GbEDHkuXz9u33+rou6+DlU0nyv12YCVC5EU1OPsjAiTSjeWlcUG
UaWAkfHU22ZH4chC74DgfQkAvLrJxouoez5lh68QATcQtz1wCyC5miT2ahPdyhR7s4hmG6qeJlZD
k4uTW4nZHc8B23DNOB2cBW1vrSbla6jbw3K8A4IuLkLD/whJYk+vJSmpyxsUlSFBYGMnYeH0NLl7
IPLcv+AioaEroo7yMMJQ8WZHlq7zrUc2s0IaqY/AmUhcQSvRnvrBagTM4xwHH2Va473k+ZVoei2w
VqieOciJ+1WXMBiiY2f4fcO1IATigbtRfANy784TSl71s404NOqFJwDjXhFRYOrfROjvud1m6MKy
+PwTGosxwfzoKeS8g6qz2oM6Fe0ZO7hrFaYAy4rpCAXPzAj8Qke9FdZbBZL3kt9Z2kQq6Z6kfeM2
dcPeFyb8XcHIBKGOXznG2KL4qaAMlF8+8NqAlB454OkPaPosMkJDD6eXEILybqgk/y1RAu07mU1C
SYyj4jOxqCSuBVKqL2zcI8R1OKNxX4Z2pqenE9E5d4IGMfSa09DbTkjhqA+faeYqRZHw/1lwSE4S
BRGo4m1kJpRMUIXfD11BrF92aiBO6qhn27lO9xH9m6im8QvMQzD6LaFnJFdpnrPbbwXmcy4BEQya
xYn3iSdRRbR5UCGVmautnQQO0sCWR7LCAqXw3TVbaDnffbT5mmjRn8fhQ1JnjHOs8INRuPKV+dhE
Srrjtk/qL6tdEq/kDEWqY0/93gAAxeSHDhdaNC78yjXhy7+n5XvXW25QHGrNcMCU+a5I3graBcqi
MZzrdfYG2ziErx92C6x121iT2lF6+LSX43cXH35GXBVfvYu87tvpLQZtm4S1HRsgNRrHNw9YujuO
vueKrq5X7p1LZeawlLuqWihyNUlDm84PQMYprH1ZvCAd3hL8gILyKLRJmBPSDfAfnw41SEQZyHLl
iM8MZiUFR5FYDwvs4++yud9wUq9wTV5LtE4gQ3rqVLQy09d5wuR1KyxtlG3HhUMZEyqOI3ieQwB8
oU60Db/+UG73c4K/JZbgfb3SWvM8kKkdACZMMp0nQxA+KkcL+bDBtp22M2Qc2hLYZ6EzLtQw4ZRP
6leqm2n7WpTHn4bZwLrDdoPUyl35+XK7feVAZ6taYBJtdBZ1tkrne02AG0HG176zX4f7sglMRJXb
eYMVyVPce6aMqRohmeOUgw/M6ciw/nwKBAX81GG2mQT9mOM1+DRCFv3pvO8TLekwCyNDgFaqlSNb
pCKEOdz4lOZXUXSX2s+JPupbmsodyhEal9HyY2wpT/w0ynmUU8FeFqNp/14ODcWGFEKdhmDR4RrX
hbu+kFpJPXVpLRBiYwgZcVorX95IZiREr8vnMwSP+DWwlnMr+sqHSSK/uneTZpQCmWqzeyHbpuTJ
bZyopwKaxj3LMQ5N+p1gF9BFea3ygGpcJnYaXslVNjExbsId8H+Y6lwq47m/3Mn4AenL+QdvFOlD
AD+43u8p4QveUtGwsA5I3f1jb0TqXwSQ/tHvviXVYNaswSylKEguwPq+5d1MpqFNg5+XuwnW8Dmo
1QGC1eUc1XSEGjVIyXqEYmiybGW2CdLvjnU6isPmRTzZSn9z/5ayMyM8iE/m87CeHZRWtwBVyfZl
R2UT5qUquI5uujI889KLe/bSfEsOhMdk84ixnOG+NxagCdx+/wbAR8Jm41z27Lyhh0JBC/CraFMx
1Q49UQVZlWfj89+Nn1w+7aAagKBVKrNy/l9eIR1aRA0qdtSgXduEJ5qbHZQYp9jLDO/W4q2OIC84
GRY3GRubc3eWTY+VfLKh2Cg3fjj54mVdGFDIyspQ7dOBnQ1piSSLjbHOWSQKX0a3vI7osvgnA0Fl
03o8dTgwlpAr6JZpLZeTYyozWxJEhOyRC3eG3PW6SzsvEqwfvAG5Zp1hGFA9VihO9W8VyWIj5Egk
bI0S3ihHVPTEoFvqVAvs5LGDAhqOBa9B9LKjMi7vpM2CFh85LJcYY2GFtLmL9ODU8q+Jf5D7yXSR
VCygIwaYH1QX3+VAqmYV985S8bqh6SUJDw+qqGCLjRNFhzCY+ClcdkDxdYmzj6ORrEnNbpIGivEV
cBaeK9bAozxl8weq8aEgX92vmFizn6UGXX96BSZcnn3eB1AcH4rV62kebzugCaSzAC/1nJOBf/0m
K/j3uJF/Kx2XmVP0SVUV50nFImdbDEQoYjr2wg0JhR7HE8yD2roe33TnNwv4Kz5woyw8tDDlF6JZ
1MIg5gCDn/LglCzFo4+pt4mmdohVrrw58EFfIvk4LHoXKC/nLk9TWrIb7q/pxb8vAVBujI7n6G86
jPKQf/NMpEU6JdxujGdOxd0Bk9KXSbhSzrKMVWMzaw0ReCMK2EHPPbUpsvwuTlxvcEtbJwTfiWux
ha6quhLUAPNTl0r+tjHSogMmiN2wl5fgQoZDEW4ZFiFh1iRytUeuhFSpZPyQCgpUhiVLLFDZJh8C
ZMbOTvNgT3ZnTR1txovUHKcgOrzL83GtOD7WJxNW+7RLn5ce2Z+6JcmB6wT73kfZI+rBvU1ANFco
yxs1yU1ykSebgORtkNFiLVzKWgD1X0+uQS5RoHQIC26LobbbUAsLfujRTfvg1iEluWJ+V9efYYXo
g5dR0fjiYogZaMHeYKiDiHmHMF0QeQb4f5on0zIMpPcdbMC/F1qaBnUXL6huDjeV/sXTUwltJ8ii
UQZEwjqghjbJkFmxfy49ndjuUcmexOSci28GZsKAHNeMR7SAc7PAU+ytr9RKBxTARnAkwk65CvxG
dKgOwieHlfm2Xq4YrE/SFajUjoJ+PqBh5URKuWdl7uB3OwjLHVVXO7fmbv7Lx64WrQHmkHrge9bR
JmaCNzls8UAprrdYNqI3U1ZHYR5AxKf9aBEygQwpDAQdNsBEv1CTEYr0npln0ov9GaenDrbBZH+O
fpoAy5P+Xx0y77ZpVwFwDcY7J+mXOk7xdomAL11Nudm68HPZjsPvarwIUSIt/zPNwKXQ0DW3w8fT
hh5pGBu19uOq+f1eR0BTgZvtQWhDyvcgaZXz05PXSgHxVxy7BbPW+jH+21HeO9tFbSpqV8VPALa4
tA0W9ZfQiBWHr9/3/WWBNWXExJGfLww3LIV2XjfKH9yC7q2SQ4gPKtlyEJqXakG4Ijkx4xBHXRAl
7IrN722SRxF86iKbMchNzNyWlBlN+jP5UaW4AOjQ223iMRv/MKw8iPRclZhaBScwMY3RMfErf2Hb
GlTpUjQDcOmbaBzbg8SP8a94yhGzLlFWezb7foABtw2oRuw9PDjjLpe4mXp3aXDknTGJyn5UvwbM
pH/LdGbRjcFWVjqPBNd9tI7apb1p9kJ91DPLvF6KbdU+kcyoCOmIjALT7wgy1h/sc5NG7vl6GOL2
2y0EVkaLrUPnSc+CFzbDSN1xum1JTxqT9J12wLVBCE3U9NNR6SZ9QvscWaMkuzHsJ4r95rorRP9k
2izP7pnJnfSYUpqo560I97P60rgKuk/vX22M58o2mjYX8NarcrOlvc9SnnDRklhxps2+2VMvm03F
hjEF1RnHtLC9toHPWcAOVnHlDX2tyGzYleP9ZyRF6zD9w48jbkZ/vj/LZI2RAJ0YSB+OYaGCnuEL
jYAcW16VmrbYT4wpz8IbKgcLXfEQfDBM/2XfpO7cYKFtGZDc3d+6SDdUybcjkZ5Uv1YL4BOxmZ/D
MuO9PTRYzpn0dgfapxIkPGRl072GCNNF7KYra72I9k8uRJzNY+mDrX1iS8MzDKcaZo8+G27dgKRX
KVxFpHZ62oFdOGDbh62c+gyjNva9uzXS0VwNuD8JHdwthkoD5XJjK3ZBiqZeMwrPkTxBqOxKJ77r
tlNBgyC3oKY/gfhxbCK6HD/mnnMkFRg6dGVUH7WQHfwW1das4KFvwKM13dnRKfOr/ImSUAt/NJt0
WwCR1zPlH2Yi7d6i0ezg9Pj1MCCSUkzg0WHlkrzpDsF/rkJfww5VEGDj/5nGEGcQ4tm+/NvltLii
VIe4akEZyo/ieyABwbbUi9ZbXZ5g8Bp8sgoj66cv+nKdZqKUk/PL2qSyonUXqbQ601RkIQ4J0Hxj
mn8vIei5QYrK0ZpOd6PX7E2vMQ4D94fcwsycTHNJKxRGpYaQ+TBcNS5DvqcrxhabbBbfYHyfx+yR
74ldaP5Na26tW6mePWqid6xosffh+hoFLfhGmSLctCXLLWuRD/8Yf4N8tArglZNvY74LRDsWl5AW
kSNzXCO2GNUL0HLJCFArspo5YIsv8uYLb9qgwcQ54FnRuWmGj6mdxUc2JAPhkq/ZU8Hn7k8E8lXS
eJdvlwkrIjyT1VSK+deWq8/qh8QxmvpjklFkLoX6uldJBrzqX//Snkn9O0JqphxlYX3DXC+nTJC6
TMC8pZ6/bASCE7luN7yM4ntwpG6Be8T2rsNHOQb+Hlus65qR6dny8pHuM+IHXmUO/4saUSUQSrGI
b9K1D0aLMti6ThMT4t5O5MooyfI/ad6giGqv42/4hhCeinqETalEpijt97P2EzUoPooUar7Jn11d
5jhuh08+KeIFnLwS1tSl7u20lUV7x4Aw3nhC2h9IEpSQrGiGSDJT6BKCzDtmihqD17nhoI2Xngs6
UqJAAZgrPHjPIvWWvi/uicQN8lte8tyVfF/FiR43vX4Nf+any41am0NF15iWulpSK+1E8SnBfP+B
IbUYGGQNWmevrOduVg54/DjzenTJOBG+SsOWvQoj0hzwcmwhU/s4GCAL6VILB3PZZ1tRUZudUgHE
aFpZnw4KhkafruhdxidbqPhA2eQakR9adkP2PwBJUpFNqK42RJYRWyYNbAoaj/K3mNMxBGE99gG4
gPXeu9ccy/Zfm5O45qcMWUPtLiiIz3CohxIcvIb/B32s2Ntf92EWdwtsqzMpZ2a51pJPchr4ypuZ
MmVsvcovN3WDlFuavvF0Qp7l91xGMWYA1vmzaN0TkEPBBKHyybi3CVqE3CsJybkMYsCmDlcgwo/t
BO4qrHQIgRaq1/TH+P3QiylYOE0sYqx6Be+1HZo8xUpw4EFmZ8kVKRM1ae83laQURGZS8QKp0WDk
dMaFZvAKuFJmYhI17RgCkN58L7j4hfIymEIVP2WxRaoUvDmrftRlE9XZFYCEN2tLT9JohUxBIrLq
epf/xh9Nwze9d22C/7T7FAsAGQsVPcfETTzbHJgPnPb+owLCmU8skVjah5NhUVfY3XptXVFw/1HK
GvTWufwn+TwO4bLR4aDYklrPx3EVMcJwLjDq4gk00lWdL3+JzvwhHYvx2sdIRvsjM5Toa/EY/h47
A99CBFxboSYguHENIZYog3z2F+EMS0ZoTMDmxhOiLIottz2ZR7DXojztS13FpAr58fIlx+QVIntd
m1lbJLNiINRhw6OHu2lwPBRT96J7R9aHQLPB/hk9O28kfpHJnzKMDapWkThRaCLa0VizVuNlNXGN
fk8n/D9GAd5ITVLPTGNO/dOgVLY+VD0M5uw6EKHhVKUeMqzaqRZmV/5xFcmy+JezLCjIiFl2EuyS
NFyOkKCP0/0Qq+HENrRDAC/pDfPS+CQ4lqlgc/pmxRlPgy2jMzIqUeslKtjqNe9PM+JydXw1CvJg
Vx4X/ARLur4nxrUJFjE0aSh366xF90nGSvpQOQGqVXayiR/KttczjpK0ba1wNQIfgitRiH+A2lTW
JnNTOCQ5XUUOunWMsMLDs2k8sl1nEWU09sA9OXdO5WSwlpZhzAp1sR4/Nyaz8QedRl2rKNiz/AX7
Bw3K1I62L5tWlvqdVYsyWN2jAlaS/AQkgmZwgItsXHZkMnuLke1n9/rrIRe/bNVHQXd6nWcG0OPZ
t+Ut12H9qDhNASEpN1nP8gA67jN0LOpiZoKuxnUTQCmn6f7ihLgR6F7LTo7Do7cwMLsHcdjl5ivO
t8z+4zoyhJukOP8k36UGL3gSnOp4Xzm5b1CZMZft0cPSTDWgQwjLgVkKX7yg3vDz4YzRR6OAnsnn
aMVfbp81qqI3lmv/7WPrUaYnOfZ9gYj/E2mkMGpsoOfI5Mn95Xqekx+HGR1L3luoZkdZprlK+HKo
ozjgEt7yTRXPrHro4pEwXhVauqGL3OCZf5jG2qz0ctPg9VvrjpAS7nh9IVGqbLfvkAVG6DQDEoMR
G7Zek0Vohtl9veJsy7JV/asTAzZw/8CED0ts+xJTYsEZFrjLoqQno3J3bP56qye+/E+0BR2ebn2c
As3Pj4YTc5qBkmBCh49wYPgQ2zVGaFPIVoLovAR4poWc6Lcx+CWq4/gie7Wr9bm3HwPejkfZJ4J0
V+3kKm2PJggwk5AbrcKE4MN/mdPBUwL96vampsfioaejKu0KU0ubGiKQsLCTu+RPhVCzCCNejB42
NxHYa1xlHb1C/Cm0l0UikNVONLsBG0zeUcXhYnkC3KHh/7qso7kOrAY6EeyeU1N8vRTMieMotWEs
RLRmWqAZl9kXR5dmZWq3HtnLFaD7iUxyxoIsoaCU1vGeS0u+CKB25OwhOWEN5eNjQ2DTMC90lCzF
vZ/R3cYmZofiW83Ou49exVdG9/jNh72TSV4dL+vsSvCjD8hNkjc+PyUYKvK+ZiNdipi0+BnHiTFX
/tC3Znt50I+TuLsSRUHomKXT9oYTKeItGIOyGIjcM7zDxZIZnqd458oPFgVWS+3rPQz+0oHxFjtc
mU0sLMxJv5jirHjW4wKUXnYQGZ+kqtvpdIXZPeKM81odOULypFjBAO1Pz65P23JVvs+d/nG2Q4UY
/68KaLbg5hJ7CXZtsG8tBp1tQnd9nyW0Y1cSKXeov1raryIfY3jGxZnAkgh1FRW2fe6bg15mym2J
dolRjcTR8prrrZQjrROyMU/kKt8MGfgfsyYEgHr2+jTdV+HAvgKaIEBPnQ8FVcjJdyZ5yFApF2Rg
OWkTKdMhmgPurFxrgH7LamVqYtjqHNeprjTkpo5wbq7kxPcAvn0n38Y/4tNVN6MA6mwunDb+At1G
AaLp27zszXGMgmSGM0nTwyINhxt1PtDKWmNtHhybx1FIk8uhVz+9apBO2DivToZf4LUXpwuc0nAZ
IVcLfS813QT9Xn4rw2e/VU6wfOMolMUPYOq9Loalagkw3pEZpW51Vtx259ovV/Z8VZb9XUsMjQBo
Wle0cyfQfL9sVKcW78NWeY3QtjpMIbFoyMCcXIzYMKkFqtDGey4G8/DF3GMTKKhAFDMOTZtAKpOP
mMmdG7Zal8JaSOd/SSJNE2eAvl1bKYgF88khydDV3BDwXC6XH6ras9iEkO0EFvgnIel1WPh4zkuV
QT2ibT5UxVVJLKsi9n6FqT8Qj8oxFlxSGe0u+agpJYPPYFF0Tg2e4m+IPB0xGs5IlOc0o9r92ciW
PFkG8tMsneoRzpE6sFdCZYHlAdtibATaaRyKNtl97Q0p/1VdHiKjl8WT/gbaI2FTt/wUpPhT4Ynr
sm/kidS8DG6/O9kO0jFlTObR5LcmXcK0XHwJ7rIFHvG1K1R//CjuLa9rmOErWWM7Ll7gFNv3soLg
nKR39DFsb63/5NwsMHIbag3i35/p3WQbhsjfd8fAeB1neHitFB0garYWMLYsdXQrSbmrm2ecxl2C
IN3iQpSsJUpj7ELELDZNzURVIMfITvB+dv+QvNsw6YPS/w4EYSpw6Vp+2yRUm6W7CdWTLKACjWH9
dpR/RtX+UeY0Q+4G6v3M2zJZHcl5K+SyCidVeg3vQxaLrkXQ/Vv3aEEqqmKAltA6pBYrW9E/Y0kc
uHxR6Rj5bLJNId4QO80Xldb0TqGbIRpaDaS9qNusYlRe6KaApciwYiaRqyWG+stZi5lsepr/8FZ3
BgGhRNM3tn7R5E6e0bb3aBybARHUsO4rp9n8i+xXMBhdOEg4b64rUBqzdjPEZVc2UdtgzMbGV9mJ
FeewLOZhVKDS1H59SzkghRD8pVPgutKwz7yiRubSacVX+a9KDsfKIbJQ549VkE/iUDAYljfrDGZe
ZYjOSkns2Vqiyh/gDJ/BwLoqudILu/1hmPbzjPWxa7xxy3XLmnjHi0GgoO8bKqCvwjbExkfYPBvG
p651sno07mKOK2+3KitFGJ8g33iO5w1pyTjLO6JdRBqtZpmSxb6G+GaSdWLOXHTULTN7zNfblaAl
fTGRg3u3DulfU0YB14bJA0+vfz6wXh7s9j1WEJzOTUyNDZgrWw9MN69C5DAbggKm567K0fwKhMF/
p4lPbHtRsjXrplHPhkDJ9ycIFTAaRP6qh74HRP7fospVVcB8mDUP2vqedOStZYFk3cLH4cIbLSRU
P+7OkW66O428EHbYDPr73NMqj9wPkDy8s5GHCtvPjJMTpzFgyxq46VES97nsQLv796kJNBFLLdCy
pLsTh2Kh1PEiywpnMdO8vGz4kSUaqRK7dPJSwfbpemdOXEmL5mXIG0Qn3WsC+Old2xeaXKLZZYjQ
CEukuD2hEomQPssjNRwFkNym2gXdmhMg85mA/FJcBqz0F6xw9Tnnnw2z8CWZpGXQYm18zHp6OKVX
3drCGz1oJSJ6TbOCrxF/P+UhOzt4k5UX2gEGZwTKS9KxJj2d0qui7KZpc6uB9F1vLyPnlddB1d3L
52YIC2VjUrg6VKmQBPOOjhmPiAoa0rjiZLc2v1Z27fB1pyS7NxUHEq73voEkuMO3nf7WyVj2xvak
vnmos7fN9iuOEZuwuo8xbIJNfmKxasrouVbWtTdJikQDbc8zTN7WxGFwSU83sGG32WqNvvEfH+ih
oo33Pcx1gncKVyFv8bGs7YLEf5sqCib73kuHBgH/ZCtwXMi0KKq6ZXkV77sUct8xsnw9eaLP4gu0
dm0p2LAG9mM2YkSlYslvUtNpbr4a4qhb7iepE+tEhA8sgBraw5Rr0uWl00UUsmw1dImbF5qcqu0x
q5Sfn49Rl1X/Dwm8udMTRkQNMR+/A8wUS5isBLgVBocGWOcL52TbKj/vOiCd2rdFsSSNZa4+LvGk
ZZAEBdA04XZ8CW3EWq3ew1qMTgBjXgCVN0v9qIgxuwcyyXSmpRXCLX+2jQ8N689dh3vCK87ahZoq
enqHrazUOf20mm67+QUJr+Wgo19C/xUMunOBqpqif8mE5a2HGENAX6tu+JF0YTMu5b6MpdgrpjKC
4hxWaJUmOgw05DF2ngsCH7KIH0p961vV5R+ebD6pAzIBxzxh6u8bsfgpRVS3gCa2IAZKJb/zdXgL
AmIS9zRGkYLZ9i5gEegqFB56YDIK9OGgFXfhIKQKt5mh0MfHY6YyVhJIqEKw+epwwvktfL/ssIWv
eFuq2LB352Lyp4ktuFLNY2LqYjYJzQSi+SiI7clnxlKRnMybZEIwVuqh1XT396NL3JNKZR1GJfLu
D9pwkxTNwCbpCwsSnIrjg/tfVMKU/buC2liCj4QZdz1tyu5Zx5oAZMYY7zJJHd/BWwoffxB8mUma
rHWt/1bQJRwFHy1h5LcC/dLYAsMFd+5Ci/JWLeUTyq7E935+Hnq+UmL0UsPMQDLzlOA2ZJ2YLKxP
Ql2i3VwkzLVzAnTHZ+M43pUNjctYyiJKwS1tgNIb1M7dtWLcPB+ItekPz9NAEAVWrp+v+n/VVQuG
FTs2/vpxwPToKT3o4AW3EYwHiFZ4dN16Q4sLeYWS9AhptH+NtQ/3yK5HZ+33/+EjjfT4ZF3vUnnU
HdK05w3bVBVdc363EFsjeYRV+IPoN6w8hO8YVEUhPxALAOJs3sR9FvCnSQxIy6ZbFbvOGQPKLgF1
oskqJZfm0THbJN6KGvQFnD+Gg6+guuDoRjWVnJnYotFdc8V20xSfkVXxVUH2YQlsvp6KeBsH42vY
w8YgJiQJ5sldZje52orq83q+3gqjWGdiKgDVc7YRCBOzj8kp4RVeSmki90bKxHO2GwnXFt22ANE9
SfQaVyarc0d/BB7yuq3nRl1XHNBo+qdmUu7WBN7oVpoO3oatdE14yJHmIbr1xi4E+TqB4p/nVXVG
+i2dx99xQzRSc6x9DzWJ+hN9BbQc8owTFv/+LhVj4K1+qmEm0ODERIITHvLxRSX1ltTaDzyO3rmv
9Dkh0e3mzvGBaWiGrwVj9E0slVMDRc+D5vx7qHydS6B+gSIYIEchGCqQQcJUR/2Ngdag58v2YKxv
JBZA77BfalT8hxCO35KyLpn4q8NfVAt3KpBDj3g8+wZ7JuzOahNA7DGU3DoYBr4Faq4dywL7FfVx
oG4y4a3PwR7khX/NiofgMzvLPRx65VCm7bBd4X5oeQq+tsBixB22LJ2LjUHXHVPZ43vbr9pDS+H9
QAWt7aMrMGhICMtrTB4zqoGkP4DdO6ddhrWPdnKRBxhsysgazTMNgSRL47/1NRvH+zPfr2yUcn1g
xNbKXbepIttVJgDvm4Z40svPYq8Q9mqiTEjLaTSV6S9F4OEpLRaByV1T3BVE7sZQ4Nvi82w6gPYZ
J7gFUDidRrusX7dfe15V+0F6txhAVgivzxPZhRHkx7xZ+gNJIf352hJ0GTbuwNko1WibXGcsjkyZ
mBM9CNzLvoAnCGdsg6u0UDlcYJjcAnwDcUjVR+8JSFTpIKZqlRA8NrwybAA9WIdZatIxvWBrzCBD
aOAvg0kZXwjLUIzxjgsmrVW2b5k2FRSsbKC5+y5byMgPN16CpQ8gGmbcIyO9b+fcvIVi/2Qbz/OB
UpOqU0qnxrTu/0C8glS7S3uHxuFalWZIMLQF+jLvceQKvwyfqYZQQTdMTEDFurnAaNcoJU8F9nxB
TPeCpZQj0TWTKbegNa5vWM0KsXeQIvEBZhd0WseYzEcJVWhbQajgcHvTf86cJR1pQ0TeMBbsWEmJ
QYa8SXVKQBvZxJwQ/cKSSl+/GIkSKui15td9wIiKM/0Wm66dd7NXPi1ZeShKdojwItK4BOsNiDLd
zG9crNC0BQDTFgnTMb/s7VjPWAWPAdRUol1A6BdOPLQdNzUKI++BSDL2nHbSTbIDbvHRs62Fttv3
pVUhG7jky3UliB58LFntW5cgmc5Z9dPuZiaEvju80Hzaoxh7bo1e3jU0iugxqT/5N3FIHfBxg27G
Y4vRewaSwEhqWM2zgVdvfwp/8usUMFqhT030SAKlNyi9VxOCZsvuZDGf6qo6qf9Xhh9yIYiazRcT
vR5rcE7IWfy7c/YSdLMQ8hF9jSVfwbUtir5XXkkeAzrefNAltgF37g8gJmASqpUSYKqCxCKOrin6
AHfiVsddmBXVGHvpr7c5bRBSNKTUvwwxe5Yv4kqXdvYvVBl774Ck0tP16v3MLn1CJqYe46eDZ73K
WOdRh3XQc2uZ2JCnIPHqR/eFxVtV3HgayczVTE/RHFvgRxb8YhHTYwpgWPeHfK3Y9Yfb/t7uIyWX
wSyfgMJFZojeCEx2Mteagak54YfgEh7i/fNfD4jULbMzPIgdXOdDB9TDLd3GqLmIivjhnS5Mgro5
QtBW4oJWiqVLtTNAPHi9z2MG6/P2BE0N62d+rZWzT1GkfUhdbBEW8dwxM2Cgj8K7QuLBQDECenNp
V9QEEmba+KKrkl7OKkRnOdTKF8IohX+JLemhffkK+/miZfaQ9+tXRZtdfWr4rw598lL8flB+M2ML
cTaShVbzAO5aIc3b91tOuJTGnBB9fQYbnsQ1/YrxvzWtAVLcSINfNK9jpO0Eh+4uAsanniWsjTYb
IWU65dg/tQOtWZsozNCBKp9ohGC81mI99Jd0IuMxfQiLiOy4PTekAcaF71ptiXGb3bE68ss1Lon4
Z6QpnL1EUYaOtXPG6yltKRCwrsgEQ6a9/rFXXnYA+5lCvJB/if2VCMlyaf625azfA9DTKpRaFJ2j
29Vbkv+WPi/0flv36FMz3mRVc64taCVxs1D+aloEmb2wjvqudSwSp17mFMRvmjFCcXcGijQEA3rt
+q790kN6vRaF2LbYNKvh3KE/IKaWIBljLxW6/zjb8Tg8tTalWtI/SNz2/StDM91vDHgXRweDn/VW
gnGzUDTFz7OyvmQCrEG1m5LjuuU8tkoB/6nprE7DK6aHRiAWcFRysllfCNVJLURLHXtyrcM6AveF
ycYsnPRowZdA1/S3+PvZwmoIFmB7/aeXl7j/DbFj4wDNBHzC9RrsNOSJgzHXNa8rAdxUW+hPwNSa
UFgn7Gn38uGkHatLl3A15bsze/X7gsF8HvuxoeeU4/EvujUhld/AQMXy7m8cpPvp0H6cJRBmRSau
YfjQ5YwrfDklA/ql0eOzV+ny7IJBE8KXHSpg1ytmi+ZGWdW1EbKmxa0hn6QJuN3oBhLDhKh03b2g
XqpS2CJFP6YnDAiDJWfzzde06P88Z1HchneouPAlwFB7rsiCbOP4LaOpYBVxBscBqUlPhartl6Tb
srbrYxWSGcJMJH9nDOHiomYn+0xvqynu5x+XS6JZd4OZsB6ByOlJNmizuHdJaMikCW6fsKKHw90d
AD5UCoWsvQ6qDzfGijl36g5LTRd1mFL59I4jvs/ZQLNwk+Hen1VRmfBdGbgshvVPYgW9ReP8aIC8
wMiTOAYqjAZz+CjLbe6gkQlmbIn0CjV31g4bZYP8boDcH65FiOebQVG0q2awoDW4fTb29cVTO50D
yTa79EB6u3GdO4USzhakWd17BY8HlvwCcGe+aZSUP+ay/measZXMKAtx5vkkmhXbUF7IaznYiSaZ
IA+8mc5ep7MoHHLRnmymO6PtFISxpwhQNSgMNNaWu7etZuIVfeZGps012/qvmxmNgUcPEFG/LOJS
/Wyj1jUdmhEPIs+V9MKV4r41HZc62/oQaG8Xowq9PAGz5bfjoazcnsxLcf4BOSLj96pfS2LFNfgy
c64h5aiABQIrlGJvQmcQ1TPQBYHR3M9QfMROAcmGAIAQve0dIQwJipgwjn8S8iPlyuk82/uUDuZY
9d9T/Aw4ThPMcn1N6gqHbPgyZkwm4f1ou4381c9nok72n8I/kxttJ+3qQqlJAxG+hC0ZDxJvIGK8
CrEoRFIOLuMLHI7u/YOR3IwvqKiwv4DL/9FYTBygW1q/Jh4yjAJvMKMIwbhqNXvO52MCZUHYZ2N5
XEw8GMyPoXpuNkv4vM5tv9ZaRFmxr1RI7tUKgIVYZUVi1p2JeM36FQTjacca7rhttwsk9z8oQWnr
NsqSTDDSxxggvu0f19gxpT7XZqyR3kU1uuJjuimyk2aylkIzB/fj/x5mNEbwbiuM/BdEcJKERdOE
4Fyg582GDYgRh6ll6JCzFR1LQojpfoJg+RljEXg4Pu7c2Y7nF9g7TgQZU1X20Z3zaNFangAx8dz9
KLIF+YvNpEseJJuJdvMXtYEMSLCH6y3T2nDGuxkiIL1Ax+memFl5bbEEXjSDacAmI9b798xxL/nY
lxhJrycau+iGu/xGW7n2LGwF4gG+SS8V3n9nLuRhdQUr7qqsnhCVIEBHbSBVZsLJXUxw7h19+wBr
z6quR5MtaiAvk5o0O13S2UXjliUAgFYSMuYFLNT1VSBxIH6Cp930cKUbAsvB/YAHnDkUSZUlqtrl
JqNGYRQaCGayrianGcAiJZn2NDd7QEwYlVvGa17w+ditdXcroUXQpx6iIu8Pjj8HZp8RmtVxZbWm
pvScPO/pMX3hIrJaVam+B6rDgdK6PnTBAWy5IR/SneWDT58illbbXM/ZFz0E6UImAlrZAm8S88jd
joKZMdKrwPtLSDI/gXyOi5LVTSZu8DH4+4jARm0CWMB7yUJ6l0RELTpuq7VKbWL8QHzkgFAdbyxs
7q+0LvzVipeovge5IrEU3rOe0R9fesb96zqhmVIfFgh57BLCGxuXqvMSiDBGTwJ7H8YId5CAWXdy
UdCuQvMJiJGWjPbYYjnnO0IZtQxToki/C5NWDhdnO8w5TTNTzNM2u5pGxsSvMxOTmWavjBzJ7I1S
tP/VN2d6rQxtpFrh55Ug6BxcLQ09PdXQVFxi9FBxyXLG/0AkutO6dYqWWdZgoSmUS5RO6JCrGK2d
rvMmhnH9zCPisMh1UxnxPkIp+Byt/C7xVdGwulLk6q3QQQlazLmB3hyT8UZ8OGco+yhhdSjZQC3o
e0BFm12b4pzDF9qVkM/0TVL3sBpJQWbSJJyAuW1GrdhhLDGjcwxWrjQ2wo9whKf3joWuX/+FkkOx
cKanFsd/eYxB/kqn3Wkjedly0wp3HZlTBy0VZOHUXE8XrNEP5Ibg7F0scqV03R5uFjPLgDO6PROk
W8ywTF5G3d/HM06KFAmDQWFM3rmxvCCzS9E57/A1KSY0weE/JI1kNF3kBZz0LzaSpGho30I3CN2+
354SPVUpm3YcgN5FUp2Dnbq9vXf1FXhN9JUUuUgYI4VZ67cy4HdJBhBg9RC2fBBDd05oG77ZEp4x
9OAiwwtQT2yBi9ciqqS+pfVxySGOVYHvPmUTrYyZy5+6qrhkbBeHJGv/fLBY5i6NeoDx31XLg2Wx
2OpZREyeg8a8f8wp0cPTR4BXMBW4XLpgwN1BnDBOGsews6goPnbyRV2cVADOJOzTWBTb84AmikQI
q82lVaPMi9B08/hmqvwsfDPB8PxkUhwySMSt0q237VYP1w/XtQsrQTTxgh87yPSLPaXEZPFhbcWm
O3oDPF3YS/NJ72S6PwGSzz6FWMkTinTyPk3jDavDlQtqoqF1OcWqZo4Us+VqJi4C6BcNtu3cp4HU
Y4T83urIRTmu/ew++MW31hn2LtHE5I5bFHvThREcjBdjDE1gXYhOM03FzDJEfo0x74bW8PssM+gR
GX8E5ErtX+Z7RyD80VP76u2hmfilYjwCq+BbvKa/cnfgOwoi1xs5o3FCh2hoP29upoHhsHUfnG4E
zIhihvTBJ4vqZiVnlx+KCQXVTYHGZzLnUEqiVCCuV5bJKc+J7ya78Eni7GaiRaqRh0rdTAzeoY+j
QW2Thl344SNkRezNg+nD4O0yqzhF+ncWrNM09U5/FzaVhuTljuF4fvSr1oy3RrHWSnG/5yG633KF
eI5wlIDstEkkZZnsnU82KdQSAdmS+ef+MO/6bPeZfoLh6Gw79o5+3ppS88T+U8gJPivAM2+Uvw3z
cJVbqF9B0jUK1T3HOrH0wgOXbi3rPhXTKj0VxWyYM/LxLnb8dtigmt7On8IH5Vj+AbgTNSSxDbJy
n+NnSl0fokbh8/XjF7fvChp6p/T8yui2sQMdb9d7755eyBZIcVqThxgKOPzJ67A2bBeMAf0i7QUH
a0R0So+L9prwpDABGCYG1gAQZQgutDaZSNgXT/f9/oEwfsiftaFKIoGNbKVNAKUEkhO69kGOUle4
8E043KoHgOP3zX7BitgGs2otOyLKPKq3RvE7VnOJlDQz5YX3TfQx7IrsaUYQuVDnkga1qUFTW7ln
fc+vuh4lvYAjGWLPC/VCp92zH15NRc0/F7ZNDBYFgrU+G8+mun5+NHMFF6wMhOHEPlAvzgb4m26J
UDoTuiW/bne/DnzfrEjhijG4t+ZJ61bbu23AuPm68fbTHjJ/UGis8GsQmKE6q9PO0ZCyEaezwisl
dq9GYqM6KwpfFsURrtQLoyAaKZ4Ly4qzKmsqRUlWX7wU2eX4O0iicLOV/2kWTzapHgKMQ7aKDD7E
+QKtH+cdFhDgSB48C31wc8AK5umszyJqnA1YuLE338UagXD3x3kOb2OO2y4mlJho5ljvSJp+xy6a
9feF7IRzrCedKbbD3EcLETNJDoGv5Lxcor93xbmQueH3JWFepWfxp9NtrkpblUt+IM9/GFjQ9aQb
CXjD/tu5urxp6hnj1FjuZW3NJPeLzF4pMBVLdscNZ9FLYqCyfs/3XVS4E/ZVqb6Ckh36pwFTXISo
PY4p6iViIOhVHzLdQPtV7TLLuuZSIwzfRHTx6xMTddzozyN5iet+i/4qJRmF2x0iDy2CGEg2dme2
ptozz0kcsOKFqA2s8+WLFJjsLwRMNC0F6r/P4KRToqjy/U+02Snhbn0guHk6HjFIXaFgqNrPXQXy
Bp5CVxtsC4ss6phC5DQOH4xgdig3ME2qq0ofmKOsROyjbvz4x7WAvq/mtdP9QnPlKl9I84A98qFh
A1eGojXKSqGHkvQ1yjDBlofbt3G8QZ94wWiJdZzFu5JY+hm1tz4jjnyzErNmnCJ1qpURCnKb0oxC
l0SSAe2Mbh624E5+kPrbB3rMxPYb9ghPfexhTLyR7xjZ5vi//+MxJvVaC8ulFOikOM4ZmbYRWqw4
Pv0o9DKbrI43ZmLW8YdT42ydl5HGmFE6pcmCGRjAxovdTGQbUWZM00I7Yd/HlCHrme430mr69UxB
lSkx42ybi7IC+QwvrOSComybnMlwpKPv/XGW+YAjkPQJsFKSW62+GgWr1ciRlDGrQUzYvIUE3h91
1ThucPtd6+Wk39mdbHzK+P887IUgZAQbdSO09X6cETGCJVBjOxqampkP+OFEjmyxC68nIOeauzEw
Kz4m/em4XRA99QGlCnHhAyi/+em1TzkR2QgkGS/0yoVDZQfx3Sb0TP5X0D/5nM+ENpg3hzzTkixc
gLVF/w5stJ4ou9c9Y1hPKlFlAplKDUboN64w9mNzTL7wHgS26KHg2krIjxeGJcs5mSl9GiF4FV5w
s5bkyhaEZROAAsCMzlGc/BYJxe9WNEv6omrC1NdLppYuSOWCDAmCDMnCppKxnnQgB4Q3CD5y6bgb
5t0LfOL9p7HyOrDsVCyPLyl+EMn6kHAmxlLE0teMLviYF7N6flvA6SoEyTkUQHhBSTan4OD7WDkU
s5rPqCIrixozmBx6fCj2TjnyywE+ViUSMEvc9wJxJQyD/KusB8x57d31B+hTK3xy1Lq4KHNepQ1d
30LdJ+9W2MputEv8hA5PSiG4v3bvFLTZ/w2BqPskUjj8YeMUhDpnr+HFInXMzXjGP1VlxojpNxKy
YXiRhuNx5HL3XKWeIiVAwr6ymyqx53GdnS6Poh4I7+Vc2931K7OkfhYNgbuWq7WOWkiVt5p7bNhz
PaueeVZWAUjGyyt3iYl5cZ/ORNk6kQT07Z7QGWeEBbr01iIDLh5ecgK08PCLh3aebftfloaRtHRC
XIJoR5vB1EoeoPu4MznUL0qvPriQ7/1RfWVQej7kuQ5KluwOVjiBbQ/A5SAbXNrttz63flnHh/Sg
045IusrQWRlE94cFd5al42QBC/+TaY7X1hUncWhTETfkm6TMv/XQRONlixyy8YNjJF+OPjbrbTAh
Zppn8AIcDQK672Bv11jwm9JA0+QWp+/Fu3qSzl6su/vLiVH43/LWovCjipBTxJ5TdxHWrnzICM6M
knUxadsC/GFtx9WI0KxNeIorRYI7iIbrYzNjukCy1OIBIWC0eU7Ijbip1cavtNRXVwXfxszrx4MV
JDxgCJh5Czu/AO8CCT+DxjfXfKQjXideCj7W+27YFma0lwN1ruMWoVpcv+7j0oZq92BZ28VO2jzV
bQbBns6ratgo7xFbGLjnyK2x5hUWgDlW0CpR1gQOlN3s634ijyXGKXALfOh/8RjIqN5+qdlMVehZ
4oJO58N6G74LL9KBwoBE6N4YMvbL6TP+XKPy66+v5/0zcD2a133I2R3fgurBF4WoF/9KpnSKYOpr
DRJCwgGYbEql0KrGu/lEkiwkcQyckY3pEi2VR0KEKm7qMGMuhC6Wm2AzuHUxRZG74+f3clQ+ZLUo
tcMUKUFtruzou1Sy7KUDeRmptgD6P4B7Cla/OWgqYi7hFd2rYA9UHXs2gh3VEnFF/NQ/zSWQJkWD
unjF3yjEZI5aljqW7F9GU/GOU2Q1DpjpkZFu9mRDDBIi2q+tNryWeFjSwwIQvfcQ4px9M9qBoebE
Vli25q63bGaEtmh3sM0u1w4e1a+L1ii3oycIBy/LJ+bpNdXLrhgTMeecBdnmZG3tZd3J5UYqWUKA
dJnHB+gI/gD3hFPhudrL93woAyangOf85O98+RMuGYyEA9cR4NyGyuiNf/QPHMBiFsUKwyomUvBj
kQGsR/DBTNF7+KpBO3j2PoUomVh3AuXWZsBaJgmtKfjddBhVBV2sW5VVxUEUUS4ZGvMJyfVF6NFL
DNbnmkuONUvnKsAR3B1fDGFdpw9/t0QFlNx3n9YbwS5X+II5hPSXk84IXxyE2VYfOmjvfe0nct52
0hTQ2BnN++L0mTmlnPMZy+JA8nWa4byD5hUbFpRa6N66LB7UrmGF1E2gtE6+fiHqEO0VsSLNRSqn
tZuJ9sxUw6sq20GeFFrYdUj8ybT5xCYEd0ZEoCmVmG4fqg6oNj9ZKnuR1arn8AzPVhnaXwQMeVl5
YQTadLhUdk/xBGckbSwIII89GG0V8WWKtn6Ihve9Vrsx15aU0EHCzh9fed5N/T4H0T9mcxLzQSb3
HffCBd6Ij7CBETI0/pJ0wnuHmiPO0d77iyKr/gtKaOB4QmStANjxL3as7ZxFpdnIIYdjpH0qX6RY
9RUTkwaxqR+fht9LeqF1YlRaL6OplBM3HN+UXox3+mnlAGFsMHNaxlQ9B0lOn3LpcSbA/R4f9C9g
Dm1gYTlE1H/tiTQeh1DF3RLaoJvlSejRlBoB+lqc3Oz6IW6PU7AsdiG27nAHUDl2v/4H0R0KitgD
D0sYYalkhjFd91cldWR1LPobfMpEq59oHDxFxhBP/s1u2gM19e0Fe+Bi0981rxvKEiDlP8WUB2aD
AbXZqwlT4vnPhBeuSU7sqR7ooqMAsEfHFUji6iGx5F+R3nPYGRUxQcLtsrKm18RG7rPyIQ6krY1w
F/VN0/LS0OToNVegEZz6wfc0lP0fFyfS2eWfgdRGZTSVgcT8hBEha8y5yLyr7rUJbjxeEn/murnM
tnuFyfMbYq18t0BAVXifXS8zpFG+KxwRN5Tb6GzSB52kZ5Wbq8T2MIscd/jeyZwq45bZjWOSYQCx
/T+8xvv5e/BDOxyC48EdIbO3+HWcVuXyH6tupKb8SO2OnqdpDp6ZX0hpc4ymyhj7Ca3C1Z7AXky8
maVUHZ0PgbsPWGWF0429cRGURO8vXpqQlDGl0euAwb/4ZsFnQwwCE1+hNpWYIG/RHLvIeeyoj8Ns
9PCMdZk15+nFOYpav/ZBir71TRbRMqTj1MIr+pWo8aqV2P97Zpd5fPohKYb63IBBCUqhAyLo1RvR
vJZW9XInsRk6NaWHSPDSf9mDwlBlfJf2ywIA78Vc1htctfyEtll+5ISVkOLGLzHBsRKoGucoXW6o
+5wDy2PebZDzHk7cDgpGLIHNoEdYoib3BZyd9jz+nC2uh96FQRdkdCJk6i8oO41uH2ZZrI7ELc1w
TDeu4PDqRIKD/911tkw8SjJfZnMc0vfDRETWkqIfV5c7BGs1MiB9Ng8Ne9AZswe78QjnwSDr8EDi
yRtD4X4Ig/5m0JVpnOXHALmyvcxij7TtwbdLnv6/aLS6GeLsbxglSi+5i8Tcvqe0JCFckcusERZJ
MKW2DsDY6Dhw/EMAQZ6RSDcw+de8kaWF5RXZWS+d5X04SzsnD9EzACEtisQRrQH32+8J4cA4E02I
lwPd0od3LwPgrGzks7nZ1beXSJs8oxlIrrabcriR3Kl0uY11X8P4jPI0cu5OvJhrRw4ohU1qVwNr
QcGjc5nmXcDOODQYLn+5fDsQwyONj8oeGoUTRy5mT6KtL0vg7J1pHGJ5QJ6cuPUgVgs5EbudbPE9
j2kIJGdNBJuJRaKMwopqH+QnZasx9M8PMlT51RKb1xnXcsik4YRYmNkX16pmdluGoqQgNKGw5UwD
dWYFSGHhdIBYdGNZpwCfeUGxrzn0cwvIlUdEL5HAan4xS995A3pXvGe5tKbP+kjC+KJwEPMucjHf
m3+8oCRa0r0zqw2xZd6G5KAnkqGTICklTs3niwERBP7rEwRM+gl0sld6Ik4SuW5JOTPWVhKkcuRx
4Zfz9pC9taB3lsGEGk79+WCr9MfLfsewyxvMIJz6RcCULZyQsgXT0dH9HFxHVHI3zrXU7HEDZCkK
5ww3kjednX5sOrsMjVFzuEWxhK0LvM7aAqKDHTu0Kx5eKR/5OcDxp0p8MvbI+jvppOKropk3mfbM
62ghAFJdKAOqKtLBl6N7MzPjj6DBLfPsK0JA4zOvMD2Irl/E3v0Rl9+EyGbsLrczkkfkHR+nxzFH
oLVngzMon2kJGtM3z77rYPKVAoDXEtYUteU8peVNO08ftY8LPXi5qAEozjn9N1Rh0/Hkr+TCj9s5
bQbk4UI78LvwM2oO8Wm/RBQRePPtaYRmpQb5yCDh6aq+zsZVpSsteGrR3UgIlwyjJiLWZ0SqH+cZ
J7b4EGxwkGhQHC6JC8ZkXhHfbESjJ4/jwbce38/OwJ6TEjPiFTAtIaS6xlgux0pGw3toB06IX2Ip
bk2ZFmsoRZDW3O8v3tIlsBSnCrAvnSvHd8XkhjWMy8/rI2ekjFxCDw1UgkcuMviHwUPD4VgOAI2I
GGHFwI1Gx3pbTiGD4tnc8mYj1VPJRuwAdoJZGScwV/jLWDNTy+ECFM+zt5zPlffKh5C88TOnID/H
hyH7W+NN6qvmQ4hzEhGMAPMe6GrjEwVq0ACMKmgp3a5Zga/R9reXZxmaD76gsdcGSwwC/r/EoW94
jnfkukhWzSItQK/xeOMQG4lP/7K2R4e7LnajgzdH6HltNL4cLxE51kOZb7DzishRHwK6P3O/kOaL
domAAkg1UIdVZRemnET/5btZ8nhQ81j6SM+coexmPxMeojIQciCTdyZYc54FNLQLvk1/a+ZVJ6NL
Xm+O++m3AfzLYE6/rdlxbR6HIKvI/SassW+7DH+KTmh4UugXJI/rWljGkhW+8TvRN+3WjBUOjXpC
6Rp+PF6EO6TrGQqgm0fPWY3DZTo34uc3emPk51D08VBOF1ZC31GBotCyNsAKLbN2cyRNswWuKqbE
+XumIFh98JcEVLSHhQ4eSg7oItBiJL1ehqpGo9fwhEX7WLAXmIXBwLtbA+irOei0w7tG6+9CjCPU
Tw2khgyjXkedgDJSoAakZ+DVjO4rs3GLbFUZGEhayTYLH/AjEu+gXaOn31GlPyxeDvdQtM41GwvP
DXJaFSjhHJEE0mht14hCDq1JpvmjUy3V07UAFroieflXG3E8/VpnbwXITWGgMQdLC9GP0Vvrhozx
ATOj3828tjjLAuWjxOQEwEMvw/Zt8ZaPRlyOaPoOSU4jHbVybPmwsI0ge2Vs73h7iIE/m+KlP/1R
rmIju1tzx6fO0kwWfnkZHaA6g46KlRyb4BhWpBJBwxm+KCUveOeGRCU1sCR/d2AixweysHLva6Qg
Z9uKATmCrXFCWm+7vg7MZyx/Gf5AfJ73C5pgdriLtwOVTfphJ24Ef/JNoSOOP22x2d5yXL/Kzalt
Iix283CTe4pZrYUma/Zf0wScYUpYjbAKNC6a6Ui1chBMCZ0EiaNjlXSMxL31xRGEyrG/xMMPxtyr
nJTIWp6MQ8VHVVg9cCShumqLNKrl32mLOwotWyql7hr36wQKCo0xcMeWMtUzfcj8q1w2IVAGqc7u
texhnxDtsekBQOOoFlrQEXIBaYqyw3Ai7FFY0PlVBhUJkXvYOKV5UXcoOrLN38ocVTEhmZ3+UQAT
lq3ah6sePxoOsAi/n+G8vDqUlChCFM/qZiyOfeKFgn6TymPEAeN1XMc/mS7tjXoiHGual0MC8e3c
DUmVSqPmJJy968HvfUPiu1G6oEd7g6FCRgBtpbsE9H7t2G68WGkhc0SGOIgDpR6qWTyd/199vA6I
RGJfehm5KlFNY1ykY69Gokl5uJpQsOCpvhvfP7moc7B3mkkHoQusyooiBnUbz22MKAQe/GEWpd4A
BCa1NjrSfq+6Lzo8u3q+ZMu4P76vv0zW/QCLWJmSNh/TWVO1aYw2kH7ymABdLIaPfFNoylsnE3Ru
5xsoV44/bIse6o9JHwu5soi8SwewUcHeF49t//oFtRgl9Xux0qLBeQBX1obWZhNnnDgkndyZE6lV
T+OicjqPqvKiecAcXf9Wn7u+Vkf50vemIAbTo4mvaQ4aSnXEn6zX4ARmBHR2YgA1sQQiX///Js4E
eVqEDcwvjVcUG+KnZeEFaLMUGFb7+bwFZ9BCM//2pgJEZOxYqKyrPvNO5IeLMyD9jXRmQlIFdGPC
BDJScST/wExUCBOxqDUMSdrmxrnDSYndojiz+Inkr3XXp8sxE+lpnH9rLEtIwFsvzV+w7Zj6ZSCW
Jm2/DeJSVg831wCnd6/xnso/XXAuuaNh48il/W7sXj0QCnmcow4PyMML9jUF1XO7/TOeWqsjAoc5
/OvzrX1pQTgxA8fGdoLkoDd2ZFq4baC4zCauLc8CMMymgyCu0lPTKcZ0sz+LgYh9Pr1KQE1CKuSe
6BYNPHb3DYpSMhSWVzYYDcvJhhE5E7eLpzQC2xhdKrmMH+t1xAFBEnDUBdkS3kK3UgipWu4S1bK9
rCOt1X2MHn+aNTDPm9D5ks3djZSpSDG7z+F4khgqXiu4cbYm5je8iigBgtEhqifqYSdeYWWS+UAQ
xBlRiG0OhozsLdpvzo9LypnS2KDw81m3C4+pfXzOczMMF2ZvH53erNWwfHsc8LYAQ2Giy1CsA6wz
fVEoUQwzsBqQbMYzdhSPFxtQAC3dTceIxy6eUbc99LVxy0tdf2/RDgxW55E2gjh9fWARShyVmoWX
qcejI+ZP/WX+k5Ex01vuRUTU1CneXioZ7droe4kILYT9ts4AlQoAtRh3VPZ2/F1r5Nlg7xc36wdr
wbz3E7D6qWDEapEeCRA36NOPP+YB+CDLSBkOtaKFE/VLyMYBlC4kjTCVqLEy3yFyTPxItgUtNj9n
xLvaEjgnCchoYMC4HK0CPLcZReQ1Vq6bq76pfHNWiFSfaVTOnAIdiXWFJrZ/kVAd1rvw/zCqFvCQ
sDrzuY6X2sISBifNe5WjeAVIbY6UzFMh6IxTkTS7R9UtqsEYqOnkwQiNmK0Pw0kAYMX7r66lGvbv
3ZJsRVotO1eszShb2ebWvFIUnoIvHJ6OzfUR3I5EG8n+licsPnymhWQ0amuucDEou4GZDVFzGrGP
f/gdsIX3baUrF0P/vSXqcLv7UeOMvB4vS3QJQINs5hKP3jWY+25ylDF+NW+CfzOyj1z29gbXNPkV
nqU/Jkk6Uh31/eDlzA9mwZ5ov9Se9JL7n2Xfq4m3t0p90bdkjD0lNOYUXdLBX/09uKpZcelIVvIH
EBWzacMrMoHQ5b2kQGpihk0c3hzG2RXtVvmeSXlyL9HNs2AAvXLZwWetjqDl+GgridifGG9vidQ+
I1HZtJ0tjhRPEeVrnLUl4C3KMtTJfhdXybAWvhmQRM087FUamS2sRiSBltkPr/rNPBOavgOYH8qq
0IgJXyLVhLvwnQCFYbAQj+pqzviOILVO++pQcK47nc4YanVTco/AROoTKCWizAnxXUPxgvBL7Yk9
1A9pYO95sJDfzBF0EMl8yixb6ADRep6BYTGgaqIuOUxm7/88P29VemEbylGBpCwDKZ/IVRSMO+Ea
BKq/lreLg9IvsPPeoYMQwMnwNlMhGKZbhC6V+aJ30exFc9+fr50ypueBX/vQ4Bjx+mVKGnrdQZ6k
2o2R3XxsBkXeePPHDQrGkaHnR9W9kdZ4qnQSohF/ZGfQq1fMphDddKFh8ORMkHoatYkZ5sQA8iDv
/z0N8+Gjw/1M2bwgdbooziMpW1Z88Iw6gFNaCcIGVqZ3/jRTJWORqu+lRluqjJdpb3dJaJi/tEK+
oEc6ygW97rXFLBpxRaAd4D6vWZdXBz8+JdLymk6y33ZvB7n/Ax3Ade8vpTZqFIqDQVc7KOxCzzUT
k1wH/J9R50sjgJKSKQNuh6/CijHNNDPgYy3sPZ1skvrsnzFAoE0fNhAQxLKhHPfGxFWmQGxrl0Gp
gISgA/LCP/B7oP8qC8lceUsyqEELKsKdnqoa0BkEF4y3bA0hjhFseZsUsqnk3dGNPOBPgiZ/bwQH
lYM+o40VYX9DVR94frfTVdWdB9IdVoxvR9cHg5jtEqZkP3RjVvMV29a1RD8uBpjGdB0PjL2oVGok
290wlLI5lisAZt921jda0YBzGbWctUvLa1m/FvhKE8ycLYFS88qC0RLmT56yi+zVTHxT8vKIPReN
RrkBtsV/gpTOAXuA1xY6NB/gEInx9s2TDfQQRF0190eQgiMHuZuGd1A2r0aPlqgjRWR7vmWkW0w9
GZ6dl7FnX30fjCgOVf6Qaitg/pwRxIDcve2rEXwt6UxW9BxHhEVKH4w2LdgGBT0rQ7WhJYtu1Xao
BUxP3Ld89R1PUjneAVE/uqx5HBf1N3UuJrhlcMcv9NOdI6YqfxR5HnBXgTixj6h4q1lPcQWD65Jo
/GeDq2HDdd7c5f7d27K0zUf5pCHalhUhhbSCA5WRSSOHLGVsmohjjiSv8jI3vHtkaiamatEPqd1T
IeJAP8cmkKN/0uPoE1LJSTHanZHbKWzaWVSdqEO+yt4Utc+9rOkN/775+rvV7gKph7Jjz2jCkdb4
z7VJZflcZsYqPyyi8dqcp0UzXVi2ilLjMbyME8lhtWeo8Ab+HL4trs7gY3IUYSQ2ec65RvlbWv14
+t6EkLj8mEhhXrr7IZkdcqY3clWa/Cau0wlOyxgC5BRTonMh1/AOD2+exC56dgi8fo3O22f7pxOt
oieTiZfd7ePc57JKzLOM4DUh28hwlOjaOzJ/CqSeo5LHeLQASDGGnDek3xNXSySuJ6bYCIEEpkxf
liCizFVB44xmdpvwpfSRRpzEWIuqecvNeMJ4SwagXon9mk1PnUYPqOeUvuUzrtQqseXfnzWugYWA
a75Yy0VJJ0oKQYir8z6BBgwQVsTFMSIubLz7x13Fh0Dpf6ahecKRXXUZXSNEMirVmWv3CXBzOu17
0mFQk22bURfkgs/pU5g19cFozMVlDn11LQDwqJRwYL/UGAvfEPDL0oEZC6NZzEKPxMqiA+Qdl8b1
hPvUFm812xzWwgrQBlbTR7+Gi//lgCrtBpwND59y9dnhrYxjU41Ef+b9jbBjjToq1oo6dykWVChZ
oRm61NXpWeeK6Rph59I3pu0xkrpXVAjVlSCm6jG0hpzRiMlFaGFIfjY9DKr15RxZ13V7u5bgW0AC
Pd+HZGMQoMf0bmiOdmvF6N5mxL+iGes/O0vj+7TOC2oTeMupKKijaR/UsPiCqmGf++FdrN1iY3ZZ
E/8v5F+REpVE4xbD/4I/X5YbnX5X2/2O99EqSlbw/icAyYxa1Y3qwraieWgmXnS3XUc5gW7kvSr6
OHwPb+bgDhigD7+C2X+fmFoel8XkS2DUjnrE1RLsOnDUWUf3wMAkdaHH2sOkyyqQhkedllquNgFA
6l0otydNAQvl0cTfGBaLkHmStqmRWrier2K1L8F/80xzXippB3cgIdiaehl6vfSrq6iNJNzLpNf5
fEKqL+GPlFcmVK1XKKOo8Rlz+Yr6XLYGW2rnILnK8lqSKcGiyF1ZzGa7aOKpPHu4COBz+9HRP/rO
+ESbE8HOnmQfRXdBthmsY0YzVU21LUXWhb6YxejK/LU898L9AloPUyueZ/secDyStr+4+pBcfCKI
FvsUGscapPRahJ0Z+gSdSHgLi2njL4toNnjwtcVQ6r3s47Y6DwneBxZ5lu7I4LivILMv6lkvS+A2
wBwlD9YCsZk1iQ1k1Khl/GGDkCD/R/bxfY1sfkAo50SE6bkoW1UVj0Pp1wClDsH+eajEDNY1qzvd
NRj6JnoFZwuSTv2EYZEaSRw8evX8tge9h5Dk/SPd94FwZPjXcWHWAmxd/0D4oLAfW3vbFR1bFG3S
SVZx3weuTmxUQ3rgTlc9gFRamDT5s5yTrcBw9wmdMcsfJkQqVcmPp+KqH/yduKflIjiE+Hlmrc/E
lVdU1OpA8Xpk88wy/H/C/sJG/F7EXnrbkUdR/Ad1bVHm9Dm8TPF2HAAXpvj2jZOPx4wnsLsEKKO0
Scw3W2qZ+yWi4JdDrfx1anUEEmV2k6l+K2lnfpYbuSpKnyGAwmzfuh1ePOP1YdelVCqC1jYnf/5Y
cQ9RHE0FN3sh6gR7UwfmV+klD0a3LY/+nDYp3CUdPlLs+lbzTDtvNA48euG7qO/QT1JBbPFvakMC
+qdK4rquH1WeoGmlPUKg3CzTIVJJCXtcERiuzuHy6a2cdiM1bEf1wLT4bcEPgNU/UgNyB0J6VmKy
VywkBAQUXCIWNFX2mdyYBQaOekHvRawA1O1ES7OtS93De2Z4AaI4CIA71iAlrKpm6Op6+gY1zSEi
jfVImC1d44M7Px3eqV8phu4iv5PbGnW3YlQmzOrSKz3jDS0+GyaVdsq7VXK6jlAXkGmEGJpJoIyK
c1p4a2wDYYQHv7SdHHvPOkobFmXxw76U81clKqp7cdBdNIbHLdYsLFU2rw5bVYz27ocP/JeuuwAv
CRzB0zs+WxuxPtuPzA69s4piN7fFEtGT/AnkHHBmz8TbhZIHZ23laBTChBYwUNbZ9IROfPNVfYe6
R52AEQY0Lh1irJvpAMi1xBj0ACOivvxGEH+siyq10YnY8Ts7Bg4QnBtQYX6tRkdRf7r+1oyqOU1F
xZDjjJt6jzqNw7xaXq8ceh8aJHzcYw5l5+kdM3RUZymh9Y5dxlFsGNneTnrVoPct9qoPCVcuYmGL
jSvAS0JyJNfz3qedSh10iOu+33EDQBstfLgTitjxbZKyj37Itik/5M2D66hFAdtOvjhgFXoLN6dt
5DP6WogP0OWaFNzcFrVkqAbD2cHj4gC8vVkU+9SGiyh/pujBjQI+2Fd91jb5yM7WNxdsQ4jYCw3i
PLyQdAGG46PQ3onMFuzFIdtJ0X5mr1+ylTaYJr8yNo88OfwK4rfNSSDjZsqYRV9a1zop5y4fek+H
HbVBkK6plIBZWy+lL6N2/BMYDqECP4agBy+m5AqdFy1eW+IlYH/usXbh8OX7Kv5Ivh/lfPNHaLfh
qgVzoiMEQkjsG2qJ+BSm4H9LYRtsikaghW7ueT8W5M4D+pHtUQMKotQMGV0lpjT8w6tRkc0c6F2y
9CqD8zvEvbc0C4G8kAUPIA4Czb8yoYhDFb7uc3L8kIKdK8kHRwGCseYLP90rgW3LsyPf7FdzMDAS
zn7vbd3Zv4mjS0d/0KnASH6uXPn1/DLgJNOkR0YL12OG8s4J/Vlwd/QxEtXof1OCtYmYkh9lSgJr
gFiBABB6iumBSzp0t75NHBKIg/TR16LNrBHBZY7dKzEjKdZlkDgfdJdZO6mbYtf2tQKXzhr3YIBj
dwizDuB39CAsZov8+lyxe2kJjg1PDGlyD4bR5WTTp/a11MPy5CDNXScI6DjNyifn26LuHgR7C9XR
czqojdnp6mSTZEhZXdJQ69140xBKzsAaa0AdZD5Mblz0Dad9VtYdQr3txiq8u6QTSjNbxZ937XpV
RX7aKAb5DtIsJdUpI8iGOsC8U1XbLGyemaE6xJKUPPs5mRW0y4dxiRhhqRCl0wykpXq5YA5BE0pm
wr+68HztPWMptoTddQGXx/EoomUB2Xo4qjybxyVCy4GnvObM9xNk/xobIm78PJF3xiE2Tgj7OPs6
IDRIFZ+83ajsST4jMxFPNeIOKXweCmnrQR3eIgUafcFBXK4rMolAQaQwtP0tVswPkoEa1OtKcSca
1c0u1JHAs134kUdULcjI9jVnH4YlIMlk1gEHhGfODAGAHic13nD98rSM2mnixP1NJ/SGzIvGBjaQ
p5c0+KP414GVUlfaiKzo0g2eeiepQ8xbluk6xsVWdH4XLG+AfjE4cnqlEsa4O1WA7GN3jbtbRPNb
j7MwK2B2mZzLNpMLLsate+8Ysf/Zwt2q/CVUHE+mYBcyQ5vsOM5nfHVJH/g8e2FETDdesKFW6Pat
ZmDDrdOXcPkI+IgYXM4gYBr+VFQqsR2qZfbsmmeKJoboA4SUx1/+/Xp0DvZ74c7OOehNqZHoD9LE
Ptf+6Fs055NVH5yCyB7MOYRZPidWnqavfz3XyQSDKLhj/7XhZpPt5b+4zoIG6n3mhTZ8cdp1kwge
EgNEOggLCmrmTUxl4j0AuLVIyS5e5HCHxv5CzD21JVz0U11t37+j4shFvMJjmrjN5oL4lnHrKMWh
T2T2pGJclwPXpeSb7jrbdNjRdGa5vPDTuadlRZ2WG1ezSEfwPHhan0xpS7C/BYhyIYIbPOugucJ0
SnnnjQMFQoWmVFxM/ieNdoBxVQRnpnVnkj2gE8/0re4ihBoOjdHg1JRzpinkVLxK84wEpWLwlLk4
tlIrC8YdkSpW7IYHtU+s9xAlxPTfvcqUtnAw0oRRkFCErsJFYNlDDORnhhT0eF7t+bkadjgvtm34
HzkwwlwYNAQ+4w3IH0KhVXp/XnzkOxNGty3arATr31t86pOOsg+cjYjp6WhiF1BsSQjOXPBUX4qs
Jj1Dcgo/Fok2KnHq4jxW98EOztGLlErpyFOg4R8cCBX0wuldOJTMfJeoz3R3H+Yj47+GfKajszYd
tZsyNAWY3tgWKtG5K2fMvMHbsQfY3lqHRaEBQk+AKAbyk+DZOI4MmnqdR2Vj6ptDI+rcOeTBPWOY
/3TmchMY52hqrdOaDZxU+OndSmJOaGDCa9B3DEYjkfYkUa3HyLYLFmPaaEUXE0zzk2JSU+2F+e2B
IUO7YoaD818IjePX+NQ3GeOgIV2n9kj1FoWRzO93mp8f4ImBomyaMnyzh/2T6/e1NblRwgnmx1AI
ejWZhh0hnRaeGkY127FXQVTOlEd86y7UJOjQPPA161yuO6410AhZ+WGIIgWmt9PTTd2WjNR39mFM
cTkzrDYbKUlcGMrccPpJnKki7wlvXjBqoYKwJekGCbGqRDEiD3PZbI0PSaVpWdWC5xjBoVPYtywr
pvk1M+Nvppc4lLp87lQWlpWo3P8d9CdryawZ/0UpR6+GDizdVxfIDfcACEnesOXT45jomYRMe+/e
W7NNsJzQbkd6Z2RZvN5N6HIh05QtU2Zwmm/U9eNW+B9gJyKPWDE3zsxMlB6fzZDwrBOpAT0XvU1c
j1GUsI8VjzuxVXCHUxoJffmAAAJBFHWciWiIOXPASkp8x6rn8ql+WQ7CfSbebZ2VgfRhAFcn5Pe9
AAGVQTr5e2BvXEfUeWWAyYCAOcptaVXy/XCibW8cyGZ6BFpHE8L+u5/w7A+NXeMq6nm7Oi4t+xyA
MfuhNwJ8URudIhtLCptNry8Btab8FsC9KAl+QqpVS8I4f8rfEe1USAqqKoxsIRSEVS0iN5nNMFcF
MkDvpfzP5kS8J4ppTBqOYQrgSIGe2tr5XspybJneIaPxHZHYGoIAoeWJqynJcVcWN66zWp4gW340
oepsP9aKugPtk9w+4KdPGxJDL9pOFpokekCtZcvGi3QSc2ykhD/1FkZ2wLQ801p/YKJyaY+hmNRP
MOzTo4PZ0u0hMa0Wawt2+tswamd0TLaNMB0n+GnbjiyufPF7/QGlN8OM57OBoEuAkPRPThqkiTwv
xyTb9mWDBY/D1qhfyxFIBLd2K6tMX3eKnN7ntuftINXVB53jNKtT4pJ1MK4ias/5tfg0+M40O5Kf
RwcY9N9fksl9915jEk+ypUopZpxcSZ3GvWEG8aHKFh8KubrlD4YC1N0uWgD2nZoT7rbas63dv8DG
+evrIyAXIjM+KVQMIFULN5Qph08qLKjv3JRwiarD9bUAQE2zt9WjHJvYQsQ1yGKNsvMQi7rCctTL
qpp6BOQtXrD4w/rwo+ByTvp3H4pKh0W8iQDkyfiDYr0T5cGFk2b9OKvMxgJP0I7yFKZmUgHcvsyA
1IaoHlaXKFTHuRXgmFUvkjb05dnkHauYKTE238n/ACOb4K6Y07KdEQAMSomcgLX0bHF6JKHfFvo4
PplHJZ7J20kd0QPPCr/xrnDINP/vQoQpPKNaN+aYw0Cx+ooN49zA6ZbIAspNv1xjJbh5TZLwrKl0
/10uGhOFJXshZM0LtbGDDbeLaDv2uw4L8q11YFrxMVg4kcC/7NhsuWc9HG8LDyCM0AA8FwaFi5HZ
AXq3wjfJaupTOjKP2RxUQjVt3qgfzqKHbMy40TONm8VTNtPZBI8XO21zo4KeK8Pldbda4XS2yyj5
CsNGY5gtxIHPOvoYjH58bq5+YdpdIYyttc4d6Eat1DPjHPsHDXAAkBQqMlrvk+Dn3GTrs5O9tNfm
jwtwxnab+QkLlMCRENAS9A/tHguc6OWK6KwNwQ8ANr/iCTDxnlHNdIQtmCsjrGEwMhqFMhw3ia1b
0ZhMgkv4VoqZfNCFefGp7VosXlgXEUS9sRcSsSOzjO3WDw4eO+a85RArB66OGe9vN4jN7F4y3Ee2
7n+TIyi/ue3jd4dOLDVoMd3C+FQFp61I2ksX4mRyMdorgZDOGTgaXCLQmglVj6Mz1yXUHzBQAr8K
slVMJBw7qRd/4UcCazsCjSJdHAUgwIGZ9E5+NZnuIA88Oqmgz/+7u/PNxXnkRM0iBuWkSDJ09cfL
JLFfEAMdM+qmTVGWtOmYhUCFPHIL6DU8HfZBt3U4nXa7TxdnXTpakRomhWh7HQ/ABtaiIFK/sghN
PQuBwAsWF/mOgaaNNmdt1q1gYHOFMn36veDvM0ebmWghr45+225BZEHBIArNimlZ7s/AvnhG1cy6
8wJNMll820z1Ozz9HQibmeeN9y2KcEGBbllcrUIorbhcP2OvrNnVaiJ5OC1VS0vgreJ/dQ6udaTo
DrzS4VlMAolUNot0fZLLrb6XNUXALajE6BZDA7CkUojJ+TMPPcynNiSUmuvOQnOO9UtfqObonrd4
ehCn6BeuDKimxYx+7j407jhlWgkdEajCR4zFikeLRWYXuXzAi2WFlmXvkFG1AnOWMrl3tUM7QG9s
V+KaQHQLeVwdXDUg0EczoMakk5exf+LXi6epGjs1OnAqedP9/Z1NrEbe75tOQ2xPAi56TUVAIZ32
EhBeFe3EHo47u0X1RmNEqgTssG8hgMGEWq8dyUO7/jx1ISapPoNAt4APrLXI1clceskH7A/+akI1
3CIW2obxdIOjHn//mrLzalNnE/wsnrgKNxlZHeFZYSa7eN02LlOuUdTQIwTsYVwPGbiCjXAfKQMG
i9WE+87sUjsoQ+OXAGqXGfTHmDIwfglvafz9hsYyG+zRTG8gbQiCpfB5eqoh3+1OmiUEgzzE0mOG
ocnIpGTnMBujy2WNSdVmRWHvD23NDNW4u6TmvKe5hNoVW85bqHbAMHF777c4lQkpQgOcrZ33Bph0
cj3svffuetXFBPpJl0hzZjNIvlMjxjtUCXJ5pbWPE4Al/0ZdJQJAh6NmlxR3TJ4TFHjJGE+YwA46
yuEMUw+gI8Yip+YLXJTgZCu1DXcJCQUDkS1hBkm9CZT89YVeo5JvWVLrL3Y80c+53RmaYceKsUDK
HWiZx6bRpaQFY42eka0j7XDIs0aXQHmFmv1K6MIIuxpzTnKtMU2Ln3foO21/Z2pY67qjSOs+L2cZ
3UTgscbjTi72swqVgCc2GyZKCJIZm1yRqTO5FOm4h2oNl696hXbTOv+o8ofhIId+5MD7KC24XXZP
rYmBCS8iUmM7SVQBqKkV7CgX6ieqZwVOtdM6fKNQ8epgLibhRMpoKuj0nfXOeXDfGfG4aoktaWJ4
R2j5QqxL0wjFnnz9IyrssdyPXyWZ9c2QDrWa30WJ487a1ckKrHu+rUR3CwVbwKHCHKeEkniVAvLr
9uzd1ktfu9Z/SrApuxFiHKQVcrDEq3ny2RQaqDHG7QdXGogbA4E3lgQdfmFtFhW8DSaC9l6ehWeX
elq6Qi4BnQ3h5+GSUspDl/2KcF+jNZbK4UVHL58NjMYrw9jFxdYNUAlBbYSzp1Euw/6gJ/XLtyiM
BDcfMjPWZAAGflWS0iBFPRl2UX+kDSbSoinby2BB1mpR7mC7sRU75huCD9l9A8v/ykUbXlB0aQmO
UmT8tCFCwYLuS87WQ4lAHqYtN5ToOZAW+ZrPzjL35nTWx/tmH2gROiy1b9M5+adbZWfgZw1Rgau8
Ucg3bvfLakWM5SqC0LS02fiquVM19bRh6fzUjLGDZlOruUbK/wFKigCUU6TQUgpLxXvPK0H/y3T5
hg0FKsiqkwroJQlF7aajHv8muk40ro00W7G3rmLySKxEgpl3r6VnXEIB3NK0R0CO0cp/aUNh6Tq7
hbPARbvqcV2hwVumPqmQzMOh1rcdKDryQS+JFzqWNwdGLHRm48OLSlBF6vueCUO7S+RxUwgEYJBO
pPrcC0f0ueejewO47kXFolfV1T+DCvB2y+PW2b8IvLVhXyhEUX6ORDeE04IedG3uo/JVVo5r3ymX
ttiCj0VY3IBWMM1xHh+YnUtnu5rCq88QkQNT12pL87wUn1ifBFXIL7hAKW5ZkYDj8xRhqxsEUtjZ
qVs+Svn3vnuibA5HgG+0GXBbCnTLwAPCK2IERKI+yQGtR+v/ioNcjX9DsuhOZaSrx3ZOZq4B/Y3N
R6nnBa5CZs0svZSTPF8UrWqakyjKp7B1BByfps/j1Ls3hGBTmAVJhwrfecVaQPR7sUgFo5Y51tbb
4NavwhyHs69XNTkhwK6UH3shtAwcczukHH5A+KPe2ymaebeVPovgkBLKhJ/iEJ6m3zetQ0YbVgo7
fyyEXOiIVnQ/RcDj1zbYXOl+HpuLQTERZ5dgXOBQo/190YI89VqBITgaCa/X4K8bm9zpN8n3b1Po
SZrq82BvQK2QXux8kf44SWQq8m1M5T9RA+GzhWjqalTLaD4UuC3hdRfjvpsIpnLNhKm2RWkpXmQK
FZr+mKhiXnd8gqq/tACkGfwa/lHmPkWIta5f7nKsRbj32p7eCoLdj2jIVJlAfH9PJB+vW0T+1lqL
7l322aP/PX98WoXZJmzucoweGxpR+BNZyO6UX8QReHXFuVRsVKrAe/DxPaw6tkVTctsiSPn/+fpn
tENnQDjQqG7zGATRaCm1cbquHEzZk8zmtKm18ncVObDtylxFMkoF57ptmsR13DAN/jVMlqk3h4uJ
7M6cQOgEGPhS6HcAZ53Cf3KR5Bm4tSeHwcQnZ4n//wKAZ90PfEZUOVY/CIjtzMkcb0kz0bH8Jsai
CC5IR75QS98EjJLKpvpyBuFD54NdXmz4nZ0NoP0h8xBPN95j3PY9X0Oullc0tJuth04YcGYVLoxP
16vTTa9wG/JgwhmbaoLmqMsIJg4Rbu2ieqCJwf4GAL/wCshpHyuJfNPe0CMHZNkA4kFkYgkcm02W
ez9CM8ib0ttf/JVBX7+4evRgrlyH/Hah6vecwb1snVMyA3w0fI5BcrxJd/ntHBry1k+LgLy2K2cv
WlmaIRGVKml2+dRS0FFy6NahXxn7u/01JGNta6uudZGSZ0sbQweWOUqDO8qowrsuN+d5xUDXN/nv
x/DBJGttgwrPzQRVxWSHHiZj0dAPzaC5x36fAxpv480YdmHEYpFiNDCTKJssZ+v80fnPkLxfeKfJ
vdxQWA3O5DGj/4w9c61DLSfc4aaIuT2rYxud/NO8x4CwHeILiMGAIIOLwnMKlJQzHsCKcvGI0Kbm
sSZE6oA6ri8ta4TArM97OTGvRpTQ+cfSZlL7V0EJa2jqtblwwDQLkL2MfinTIgbLZyYvDFGfWNtg
nNoyOkKRzvEFazMo4auhK0BI3Ym6xsFANt1P97IgCJUPQcJFqlGoiRC5k9jRH7B96DufVGuxmoy9
KDcXMWQs7iR6DVZVeFPOgn2BvokNuiv8J03/W4JKh2EaC5UtKNSrWhppuLWD0Wv/y6vdcjDOnKrK
eRwMHiz1I/CxVZHq82CR7tHzejxS+aFbx8me74yOTpHz+bvUhKV9qhBFbbZw+Avdf0PHEpKES4jc
iRD7SDcrJZWXsdJhipDfCuD3LekRw/2iih9WRiC1vDxqyINLGJC9svFc0D1TabHiK9FgGr7XdC89
8vkZvc8hBSFDHY+TUtKLK/b3H2Ad39UWS/DrS+3ifXta92NJH9ZSY3HdBGy5FZNwuMGbvxHdQiOl
Z2mGBCx4xleDTTrYEpfiodG+5kZ6aEhN6j95lXMFv0VF8rSkyi2ow+5ig6rhYRi5cYKoL5Q5/kFb
8Lg9a3+7LORQqHR2aQUxWiweWgx4UyFdsolDEnUQ/w6M5/qtK4Xn4Qewy9qZBCAIyh+eZJD02H0t
w+GiSZ/roUtfdHg0lVRYo8EcDfvhDObwEDg/aFBDoQmK4X7KcR9qIazvzOU/jLZePs+W5oc9rAyO
6eMmiNjMlPiyMu4JTfblOCCIpa5xXjr7vXTs+DCf7XROPSvIxxkzMS8C0qyYvcNc7uAyoZmMaXA1
tfULq153F7YiDItAbK5thtgMo3+GKp74TbB+LHmTMMxpsB9IL14VBouifqBnZWfrt1ptYclF28ar
KyjZo6P7Q9siNeLdOe/hwOQOFoTlcqz/zEfJclxHwx8As40Uz0SoK2GgmA88dCum5nww9G0+0T+9
nFweapRE8M9ZAb/Gh03HQU/a3mPFGgwEJFYD3jec9qeVS81jpn0m7vKiN2p5J7R1UTIvIe720gHW
Yhm8FMhNRTftjkMjv3dZ0S2wS5UFo9luSTZDYXKIkmL3K2fIWhoRA1SNVbJ+HJZQBfLzEADnoRqR
ojaJBysj9nNIHWH4bKyelfznDrsXTBJWfb/Eed98AWy8e3WOSv8QnMAQxT1aAyWl8vI3HcRZR9pK
QHFpTkryecbb/cyfNkxgz0DKyxt/hMoQyClv6VLr+cRAptCqEQMIDLPQbudWvsraB0SW/Mku8SKc
pgbdLWO98PdwefS2bw06shtJDtKWEMvfHWnqkZIqQ57zcBdNn1sgIN7znpAyWRXKT+4ehgDfNfk8
XEJG4AnocOTIu2eJTgGCtz1PVXwFK7Lqq0HjC+B36sTIQ1/pJbpStoLDzm069VE4qmTheBs9u+Mx
LvoSL6ts2lsmBsVUc4CPCZ0TIw22ZWXI8BuvQvz9YnsoxWHIKiAqCxcqbibq6wpL/HHrr0ojaQT+
84aJOKRS2t8YPQz5SuqI9xmcVjMOU4/zN9o8jLWz0hPryw9A3sYF7LlezxzjUw49ZFCrQT5ADMIU
syWWTXFOW2kKqxr+wQ7eEZ8eTfhMIUdlAbcv9gwqulK09lKtka4t9hLJ3PXy/iLaw6Qc7J4JPY8i
r3KVjwGRZbS6jBLEXnMMhCETwuJ8sYCry/ylFyu04jY+9ofueU3GF1dEUZbxg/3l1rdWbrYx/z2C
/J3tQYcKHSjAWJkyZwRfmDI7l5sVXSEhwLzc63G4mStDsKxaSTUrT4ELc1G1QATg/RO8BzrLA+zR
rRfnJ0UqA1CmBW5RLxXnQUqRzWrS23FgLlOwa45+7d8BqVlB1JSSCHF6tuvo2+2wuvpUbLa6Ghyo
av9N95pvbBM31BzXjLkWu4mFe9Zn87Ad21k+02kdTcGzmR33S0Yb2CMTBO+M2uCaFUhzIZbuEezz
cq6U79vfBufZ2xGvrD3Q9nPdQeBmxdmBQsP3h2rzL/yrXp1OC1vmQtloqUS4UPzz2rojCxiS4HC8
f33Z3b4XMOIs2nHHr4qgtII8c7X+7I0QHO5nWM9uca86yve1mHOGyI3oE3XzP5ntcm+pvJjUlwng
0Hn3o9bVBT8fMsejAIhH8Dj+QRk2BkKtgIlcz0MwK4L4YqGsGmwKZRSW50WoY2/K+tZakhd+8iUI
2zz7XpLv3JBpMg1S8QnBnBfmlxKiY8Rg8lReajZ+KO5dNVOn4lRcdG5aJSfccH3bP1KQZ0VWsrh/
H93M33cx4zd0kdQWebQBxG1MVzPFOUuDyvZ9RN6MZ9RfEB0cWyhVfmV5r2xy0Ta+mGTc0oCpJZlj
Bio1KLDzwO+F2PbA3lRL9NZdZ+szZAN8E6aaF4Bwmu5J4X/HdyFVhDuBKxcDTe4qD+mOZ81HGV4m
DHGyRMZoJtuK4SSVpa4fJ9jWkXe521Mogu4FZLGGerYH/1V13j9ORo/W6QpWcDKkt/iOvjo1YU83
CK5cGEi7gbZb3HZ6adGmJPM0IP7Yi5PcQj9RfwHkBQwf1Una1dDIEFIYfgHyogwhtuGETCn3syle
FH5b0FHSxHmnZx6sINqmFssHpWF1FHp+tC9+UsRff0jGkw9WcWub4KokntJgCEfdfoHwTXvoSUMq
OXA5DvKAZH88BYv21+T4YUodNly+pcip/IEkHKtNwewQqX+b05HBwmcAQSbSzGG0rK92ywHunL3m
f8rDqSNcjoQeCNcjNltjv8WKwRJ9UXBT/lxIT35mUNpHEIJ+4eDvQtiuLBpE4pd3KLRKFf6xYvA3
wqcsY7YGJPfykF3akxGrEdElxQ07tRPrAndC3kgF99tXrwr/06egcGO6ZjA6HJvgTII+5cyllJs4
iZVpc1b4LuTl2fjLmmhIfYpSa7O1kr/Q9sy4eD/H6oTedeYoMxGt7rrVZSkxQgdPuoXdH923+Gg7
B1Pbhp5Fju82JsaimhQ3fN3aIYSTP8etcQmDHNBtMiG/EtYGXTVrM8KUSIx0sbDVAJHIz7/EM/Ml
vlCaZ2ftD8BrGAQMPahT7sUsh9n/anbbr8qVcl0kOtCv1g22EYao770zlLZTCXM1xE9rgVa0dZhb
0gXuAdh7QFgwgjEQdkomaeOx3HjG4RNF3Pppe2LS7BusHXI6QPku9Z9VMLvIHmWDN7FpS/DdUp11
NTZBosPDO10k4d9eyFLllMeg+nH27MOpRyNsUm3raZVw6wkwHzYllTcn8AIBCZldsW+UB1Oqpq+S
FZ6kJyyVGWSSCvoORO8zB6loh+/tmxOTndPv4JVxDOzcQlytE84GSS9tkMTn3Hjrm1ywQgjTVFQ2
27GeqiNf5zruWm5HiFZbQrbT4NoPbV/DACsbvBES4QoY4sdEctCD/QRScQ+7gITPwr1EOaKgLO/y
HouA3j5r1duYQVpkDOw6zMuz+mKK/c12sb4iwUZItj742QGbhZab4MaZszPklrjqIywiEKPvEleA
uRihMdj7qu4LB04RuYmIilhF83VIwlcoN3wc3Ape4R+2IKru1JPJF0cGXfJBa/aNC/tTqdp1eROQ
Yj3Y0nYdsTG+KQnGmRydsDOpPTAB5SqF1f/dVajrEkUwwhImdeOlv+63tvsGUglZEUvKeiy+libJ
wHff/FsxkeBNcPkz2xfqPsMJO6o6NpBveoN3WBaylnytp3+CCdpwC5k6pyHkB9LmWHq3pJo+2ATC
OhxT80cC5YvQhjn6OUhLmw+zj8ylHOEL6UPyiZOoh0rEY9Cm+pnGGHWWZMok1yVVNES0CHaBOL7F
YiI6zmxqBBA1oIcaxJ4sFXyJ8us9B18gQmsnaKet38AVgXDpDEcA4MD1EnisL5wG3lStwJ++rK72
13EUWdWpicR1VSZ3Uq2z5XIQgAr0Qr56sYsHgNdsqyowqGDSsZAIl4mlPOe+K3GLIB1w2lCSGEtn
Inu5Q+2bVmSmqYgWmI93VpGHUCiz+6QNvlTkc77t9AlTUSthhGRRplXhcQGIFJaTemZLTqh9fI/x
YdtzmXP94m8wMtus1/qvp+AmPWdpFUZmIhVW725iPzaVbiayE43fzDkjabFEZHh9PlzLcCqK7DUj
CnSxtbs4FEikIlVB03MOXYwJQHHcxpHnkvi4kHkQxoGeFXuHl6e/+w7FykFg8BvUMdHSEgHvCf2K
r+tESAb8zzEeOP0vIpiC0HdEXmQMYOoTo8GjEuDOaf6Yw0nEol+dKtWO47SrjmS7oiJDqFz0yzXm
zANwsdjaJ8JXvoCWp2I3wve+9wxrPzeJJl3EJOMMmmpuv888i7wo9xlgimiNYOVyNFTlD3OcQHB3
zjXkh6v/lQ56nt9y2UYWgXcoLCAUCHnTYPGW7B5qABFfNWGc73YlP2fWjBp9c+LkZteQgrAmQ87q
7i9bmd2HaZTC9l8me5ij0dAFnUNhmLPnvNgdNC2M7peCFXEuiIImPZm98Orut6uM7Axwqf5GkkEn
/XFSjaW+BuASxfiMC8Smh9RweeOyLnDXluCcLG2W1/Z7ir2yCa6njXUfdA5N5aeDo/4BF5deMWJV
J62qBObfUGKuDjHqD1lGd0TkKupup8IZgENUx8+6tAciRI6iGZK2sJZ6wbN8EG1kRGvBCe1ISF2t
ECt4M7eLnSUx2mWS8HqEd0IukUNYhtla2PKRcIGzBIrK4UZB4wGKXr4YG7eTvWzND6bkm5wZh4jK
WfRD1wqqsQ2TK3UYMnGJMD3jw4VAencwwaWORd3m1Yi6TZ4BMCZgQQecJPjuRqxD2JQ/XTacgPqL
nkEABrzeQr2UpBqKZbk8NlDAjpqQxmWWZEkNX899p/CHVL/hYl6Y3eXvucV9wyQER3FG2QzRPCc/
HfAp8h9AREBX2jG2S3Kr7v4GXxrKIqi7xEhOqJSOP5ESZWKY+LZGemHK/16O5Al713GGxgQtWRlr
KSkwd0tXKtQA4y+VAiOHuAspofR4oWndJQ1njRUvdLlqgiWa3o8juVIJbrRG95kv/ISXC2RUNvY3
HQdiTxhp8BPcvJBpHy5EjJ0O+hVhRamgfckFjwP86tL9O8JncUBLqm05aosO1mj2V3a9XHvKnx9t
5ceOU5VdPWgJ0u5vzgb+j5p7pJtrk4jKg/KQvXO3zeQbynrc+JzOW2fykx3qFkWsF9SdSf4c0qIY
7gw2kZW5qHgE2sVXAqIpwEh0zd/9TSK9mmmZnQ98aFSNP/BnjhkOipxXKRx0GdNXdv3Mig7ewhHd
d/5Lt3deKkLdvI83H6eLZ2yVepdHdwGhogcWMJ5w3SCgw5Hoe+Fw8C7H07DIOHxmwSUbUn2nNmke
570aRd3sXvHgDdpsA9+vIIAIFfV7c/21qb9+uXwZr6nbjSKV3pdnvfjNxxAFf+GdYS0M8jQ1qCXW
Q45P70X0lQEtE6YThfTOw91qZ250ai3K/+557hJa6yuTxYWPGGf7mq/DE9FOLYXOtcYmvuremODR
9Q8oAXrZgUCH9Hj5lDItpFp6H5zX/6WIC0nNMUGSjbqxDSq7SQ3aQordutpLR3G5kFTUwBzA8l1q
1Y9DC04S3fS/1Ws9zRhPJ0bnNMwPsHkTriGlrUdMpDUmoHkeWKUE+uzyvxa54cE/cWmg+lsWYd1O
STHcY6ScEfmOxPjZRJH8RpDh16hQh53Dynk5sM1F9ISz9Qvy24TSVfJY6heDPvSB6fNjQLlg4Di7
+PvzZ00B6Wc4p31yMw/+MuCW04/A6Hcz509fKxUhCWJYM4GlpoXTWyj3wG6Tm9HNXa/PBKtcQLNt
yHIbrwb234wSaUMB9GfAzvVohz9mPJJvXzrtY8SrLNCWESCAbJefvvFzP8GUOljLkvDMzMZ8tGAL
vevQNSX7ij4qXvDaBC8BPdj70JaxgmLAeajsvkDVaZrabFpvU/556wa96A9ct1zUsmfaCYBk+N4o
gS+YOrDTWGaRM3Lb8yuSVk/l2066HgI3wxoqhj/nd70cT6cbbgR9KQCch8bLEGuGrTyjCfwqkcJh
Pn6wv5OnsDcZ8E4DCovkn1GoD5I0M01Uo2RI8T3Axla9wcwFzkZQwJ6pz156KszExU2HRL8gEmHu
LUm5nec+QKYvWHGXatv7J8lNmJGXdwzuDLxVKsqaGtMRKK9YwSeAamXiCDDLDplHOknJO1zYy+H3
orcFr3SFVfVYek1XcWu8MhqQpHWY9WQo1zAAbimaKUh4htor6NnsgQFH4HWxYB9GYSMXtgC9ZeU5
JCrqpAnIRWVaQ7YNuUXA0qdsdH2TNvC2td1tEDdMvgywmf6p3aw+sCsPWNLA/WSpQMQhZ8hpXE/V
zclN7SB3CCv+kzPuEZuMrVznNC475N2A7UhbEZD2yepB54x4MSbHZBggxXe5ziazV+KAkeRxJ1mB
DjeyaKexF641oaFjDTKUQgR7BKYPFiXvd9T2FJ2B+ygmep2jeKdm9Y1SZLMm/MRlft60Lt1OI3Yn
tWK7At7N7iSjoVjtXbXCsEvmnxFhf4rrNKF4njCMhX+/I6MPLXOpSXSUlhIIVmX4QZigXCPn0GQi
/1YbMrB3/qIVzoTPmR4CeH9o0MhRghz6W8SsfR2ymyDzVOY5LSj5iUIxLrTy3gFqWGYTmZwCd65C
0s3r1PW9ErubXRjwQ7vegOuhYcHoXRl7vW3d60jrh704kLfUKt5LbmlcSeSidGaiMe4D9211bUaz
hRgcYTiu5jiSbnwEiIjiiJ/WVCFICcyrn8mUHhIfrEhMR1ivg2qUBABP1zs/e8+spi+TUnmhYlr0
2KG3hKUV6QF/FUyRyzp9AZim8cdIYiMJLKWnl5nYSom8otfQ8iqOJwa1BcbmEEgOGz9DxbGkCJ9c
AFfhi8T2d4qx5rCEo4O/7QIekBMk9/LawTaWzHd3jbqxxj2KeZpdIF75diU60o3umEeFl+EROZ7u
t/PpTbF6MDEDJfiTZzp8S+nI+kZN3+uGamhVGCUagNu0CKtucMpketJGH65MGdSCNmh5egJLTRY1
uRApvmwVuNX8Fvb4tk1tJJx8FR/SLli+ia7w+XKkfnoEDQxsGbIn0ddFR9h/lqL2ljQz/rgB5HzD
strY5VdPkHS1ZapBXTv3cjYVVBHSK+xsKzPhwgogiIqKOCkfpUT9Uwtl13uXQcXdr/XWjWPO6l0s
79NoRRUbHsshdqjTmH7uSycG+xlJgfhm5DQs28gays1xlpzs0rHxpKtIqxTAhoxM7v5rjtlriUwe
jNJelOfkUHrQhEnNZXUi2hm+fV6LpHILXR/+efJrm+DaGdfTPMVAjU3jVvWagNFvVhRcODYNJDjB
Pl0ESd6XA9b7spjjEOMaxqSHgovsXbnPjP9LG2m5UjdByOxsFSvYoHGa1x6t1W+v1i6aW9Czu4bz
Gz3Vw01IM8xLZIuPkOF4OoVWX7yu5vPry0jN1iF3rfvvusFS5vrfar8Mqt24t6JxhTTwmXGLR8zf
0xadrYhovgOqrrVSuTbzIAZfjvvLPhc8Y7JzfiQhxwPXBkncY6NNABaUGoYmQFm487xqlH3pM5bW
Bdg8CPxpyDDL/NOsTvBM54BMpYi3nrfS9XeSbjRQq1vUpwkzxBPHJiZJWzusFnD3pnxJr87sqCyF
KV//PNXIpxIXk5rKL4o9k8vwpjOYKslxHTYknMARo59UtAvUBT0Z927kW6KZLh9W0V1MfLLnbFAx
RkwLild41xc+aIXKArVSpV9hHR2mYrRS5muBRHcMKx/B9RIaa+seiUp+RwKVS5uSW5RLmqpDGHkt
Kmy7z/h2P11XMZafNfZEnLOUqfrjfv7hmLvlyG7pu5enzH1DUcs0EKQLJHEB7D9wjMHYnrzrDe6j
0bfZYLel/a3SQ5aA73IpKEACU/CKfpYRnrsA0c1o74B0xCHZF2t4PTFwyv3RTFMx6YQ38f5t30dh
gCtN3vIXhl4m7ku/gPsr4I6SyBHY4h+ov/p87jYU2EkocXKSCc628ecJNDpcsabOx2/1PvZBQV91
FvsuIyf8R8Cu3HwfUfc1p3bM257diADvsIcLTi36lXtPMA8x6yRAbHRgpQHKBwx5Yj6yQU/jflxI
/2eDnKKyZb0ockcb2YdZBN3TdClAT92jekz03plvRX53BZo6RSrANcJzPDWMVBomoE2zHZUNE887
weS128qt04zg4Kqb5atq8V6a+yi+aSMTi39aV12jrNpMgxbLGugV4b/nxNAoKxXjl/Juus6oMjJf
aXNFJtXupNN04pzrNMauEHtdBYPal7kkywgAKlx1d87bukxRputD4sWu7IWPFmDthtBMHb+nCn7x
MnEslAXgBtuZjloBj/Lvgo8TtLNozt8hjZKIZTMvY3vlc/MO6SCELlqwyPEUMVdcMFo9+VbMLAVI
7mlNrrEsMLexfSBh012GcQIFc0gBCuIjARhI+QTIvE8NJh3BrbI3vXqfOOURxL/qDy2M6HwDuz9D
6XgABY7esfBxl4J7by1j777ElVXzk0WoLTsn5WJcZ4aIzbOXtVyiQq9YJ1J4A2fI7+qGSDrCH9sP
x1eAIkfscmRNF+2XSHb9ltEDi7I2OGR8RyHuKwNFqMLyqoHNEkPitj785uwegUWC0539ublnyP8h
U32AX8ohktsdULEfb4aWxb3lddkSYOiH567tneNbm+x8tHBqAYr0di3W9laDs8KLAu4LpSfohbpv
ko1oIzK6QZulGaJkYN2QNWOMwhROHxsr/cuKmNmazraCxd8OFHbyXWRj0nWSz8g0lIj9XiqXueQU
FMrgZw+nWMOkBKWHgfNlGTi3dtyza45ZJYqGk+xVFEOUJFuv9MUq3y+PO6o90HKUR42ddZDVJfGW
FJahKbaDNNrfsYFZijrdvJhV4V0+GPisf/XyHcggLf/HKG6BGBea/Jyi/mn14wDGq2MS3RL3GKFr
Wv45uUFBg6fd1VaKTKjUu980dLJeW7OvPN59gyRZD25omKHMlLFeGisc62Xh7ZVX+EbnUr/Z2skM
91K1RHJ0q9aOp2pFc7T/U3GS/7ry8v64Nt2sxf3c1FM+vaq3MNUegR2lQrmuCIjxLwD0zhByqd6o
tEPuvqiO1HGt+InWNj462kGrcp+IS4b2bD6QB8SR0pDFj2eMo8TtyLQFvWASg0FmA1zt5td3Fzkh
3xOXjsLoedIBu/CNU5v0TvNR8O/hh1EjJbONqGw5aag3ZVmpqBs12sFgL6evVmzlWgKhlB+LzrWi
dqzY5xTq9iKxiYfxWizp/2QNcE14VDEjiNvFW/NxCJrSI1Gv+yRb7FHVUbIN7j9QX8wPH6VwL7MY
dFtvELLRnDWfEftrr53FUXaj9SdU1CeGHL25hTGOP6KPPuHKFai1vZ93ulLC1imWSjsEHNS+YuDg
h04N7jkRcQajLDeq66eY7Bne9UkTkTUS4SixwmF+sRXK5OWbBLbKFFTMnqD2znNGIEsTqKrgAEdh
Y5cwwJhWBkMxX3vBpq5Pc4KPRinDAglelV2o+muPaGyg0UuHfjgVj+QU9b2i9F92bLmcyQZMMN6o
3lJrNxz3y8Iw38SDy0O9G6m0YK+DT8tinb4Yx7ps91iyUKGtdczfqP4TSFYpwfAdVcdYCAw6BSrs
paAjVyGqX6CN4HAtiyQfCY4mTIqB+dJW08LL7h2rYavl2VTW84OkgjPkOZADR3NUsU9dkwuP5bvv
1IlCAvLik3Q/2fkVcdz66oBIwNi7IWvKfYbEZoavrGnU3pKqvSBbvh0G35CBaa9iRpU1B8mQUiKz
gNAgJHxtluFkIfHwwYOshi3O2vu5gZNw369jRTkzxZuHhWPRzF2gDnxT2HcmUC8L36nUVk+Jxq/m
N+bi5NDkq3zsElwTa2DD0JfSm9fQAOg3TG8FgUPeEv2vdPDc4Lxc4Y9nH1IZCixuvGyRWdfa8u7/
kFxNY2ECrPt3q/DcFP5yq/5BKSr2LQSUuuJqUz6fTwjGo87+D9xDkqZ3XL0gCQabpGtIkwqjFsXv
bV9U2rjb3wl3EwRvV09dBCJfRB/jq8nJgMajVVErKmJt55wvuO+zijHsEmXxPZBWbmv3JQhsNwhp
KZiy0GuLZNCJid0HH29fDO+ydu4XFF8JlJhJYFE79tvaNpP9RN9ZaU9tksRBW2yvizxvfrx1Mokr
TPSCM3MeJ2wIQiosL4o3pVENhiPW+FLt5uCrtvEB+8+lpFx96F9acxqpWqsH/5KRQ+J3sj9QjRrr
fQTYj8WMTE1hVBb5DeMLyYX4qRDbJspTXy97qSvm93nPHRK+iOg0UTqxnXU23qX3THzx+Ibsgs5W
4eJLR76YqG68P3Q+Y9aFXyVCH7C80L0cwTWCLfegEr/Nt4Ko5CAUthS2KTNuc7excXuafN9WTQI8
jmoEC8CYr4pJVR7kProUpOLmeTYKBNHHdv13uVytu0ikWwVfcaCTK+yAbk6O12YE+EidPgmTKVGn
K1nkqWoaJJ4fTYi6u30kd7parM2+bBdEbv8tlfFdd9Pf+8cr4SU6e1Vd3F+z+uDhmKOjf7NxrSue
2K28AzxeZKcLdMAFDhW5f7dQKSLiD/r6zSvUSf/ucOVo3izN1Y4XmSbiyKSvmKM76lIOnk/zJBOn
4PGY3LMD3xrExqT/q3KVa5vyUqQw6iy8D1Ei+HpqG30Bz2jLFFKqF5TC1FONATFcl2u5TFt8WOjy
L+hTdzJyky7Tc60zL3HjiJyrtFnYis+6uYndGuyEqUQDXGm128M1mI73s/yEY+R2pwd0zVpryCpC
jPwrc/gOKPC4r46E01RZU5PAgJL86MBDmSh1lxDs1WucSjOKXwf3EVV1PYfoA9A5R8z8vSVgXLZ/
/Xet4qWmLl3btgXighcvQoqhx62Mh/g+KheJs3g4zZ3e9w+3KUlr60wi1VetyK8o6bQ9AJYarDuQ
Xm/vdg0gi0vNmXb1jCJOXRO/flfLxfksxE03D/v4jxq+hlwrhb/sEHTwzbJFna2l+mJppR1D3C5X
b4AI7XlorVoVAxOqiIjfblwSvbgJgoST5nGLjXM0eXpgZfGgJCm39Xnh3taanbyyF/aCLuhqcaE3
F+cYshX8Q53lQlfMU/77Ajsd4kuVL90X2HxaxXyh6qHfwFYw7y37dtwUwSwzAy67gfN5bR3jIY2G
WHtSwrGn6ppSyqzwrOgUxWpuiIscX9TbNcdVGXRYxUl3lpsyyQ0T3qnpm9D/i26Luy/y2pcs55uF
CXC0/AJ66hiOw+3uKhEh/Iheyxb+5916Wl2XsUnigg1rYt+ZNvKFYDgCmkibRfWwq2XhOE6wG/B1
gB08B6TOd0WSuDby6J5hVvZsfdr0zpDfvpyCtYz8yKmNMw1e197PQ2Ib6QgZhos9GXx5/eFtNyVe
rDe7p9napsJWivnKlido04QGAjf9K6292m5x69bsh/G+Z093lx+XC7TrR+i55n4cmNFJG8HryFZu
jOtPQm4YAoTsb6QGyFc+suKMF7yHNIJZQ1aJB0XsHu8xaQ+hYn889F2K5Cw8FPcBVk+bVG6HoK3T
DEpkopluLDzzFp/w5n5xhTCA4s4uLD2dsxYywy+jitqc+LAmZbaJ9LTTWzCX9/LD0QQ9pAgSBQyj
iTtwaKkFQ5+mSHE0/5psCeNFXASRHcRBraiYx8CGQWjl34CzPB9/AKtkb3DkkYHghElt9KGFtI/X
zMFqnFFTLkbOQp9Zu2DVNZhrJLfHC5KvZwS2GRShJXQ2oEqwZyWLimQUI7fal3kOxdtNH1q/aW81
8LZPy9/2F49GxtBaXCW/EkjPd25URIlXYXO9ArphGsnGaG784km95ctXLjMheC5Opo1mMtjEZgMi
6Emq0jnszBMm1SMotP+Ge35BFvxAjPeXqHknbQdyXnTlFH6oIxiYPN0pbv1EkqYWA27abmWR4zf3
9lGyhPZdy0z3y1xo0HfMA4VZYLq6/W4MaqTYigNprb8dQrJByMTfMBkLxo8rFBn8ESbyt3n8SLYR
PIVs9AFLUjrBluz/vLB6ra4Q4D70yN7GgnIJEBOxKlb5JYypZoIwmgmm6Ezis1gH8/Yc3Z38XZeY
PW7ET+v+oHbH0PiFQFpcMf6JitQd4A+jUK2qNF2SJVnKArtUtZ5DYTI0GJGU3CRg6C62KR51Is+W
qYUVb9XvRkFFEWoYdABddz3NIhCCpao7D1HOm+3D+HoDuPG9Pvu44ta3leFsW/jVrOubH8/btX0M
ZqZsHGc57GwEbxHolLkOJhV6dHwL8ajkOKPghft9598PGPXB/3V92IU6onkpYUCryJyh/vacyn++
sZJ3K82+WFa/5blxOKEsblAl3ok+xGb81dMeQfwOAOUNCc6Zmriqg75sqMNyxSiVwE0Bv4sXgZVh
BPmUalPAugszfUbyaH+3HS0DDR9o5grJuWo71zwoPSMqV4qWVyqcnFtT7+OcfHrNGUI9y9s24YL3
aG3LHb8AWQDlAauB5Ob80GfK2Dl/OEh1sj1dxQ8dV8iPBg9/j4UtmUeEtdBNFMVogUUqf262PR4S
O07Z7Szg+3Pim0xtZfMnah0Fl37AuXl+YQ65tpiOrom5qJm/nwhIBXiNo4/Kjc1ceiecedTERabd
AFVVW9mnJT9We9HzdlLSpVoESp1Sg/cKYGiqB1CxD2ndPGwvvIBU0lbO4eQgMfIBUNk7LSTM8m7D
91YGq0eJjaOCsPrs5+0GsG62NnX6SvnBu+eJyq78HC7tIQR3jaqc+PhfSzJT9Z9oK0TsZaUyKDiz
UjlGBzlca3quEplvQEo6v9RjGlHlBdrKgLFt6m17GBD3Y3RNINp+Jh5BqHL6wo4yhfZzGa7quuk/
ltlbdcCG/j/Gg8oySPjWKZkShjBziucoH5pm+ulIBOf/GifjRAnhnT34eVC9jPfkIyRhkzYZ7/eU
RnIrypKRt+gR6UglFN3Ec4hRNu9OAvFFY8j0cmy0dRr7HKQwcAMZeqdz8kvEr9unTuJqhoniyoJi
oayc0jo66z6bkltXu1OfvyBBPRH70FQyLguV29Jek1km0HMYmLVihdzgfK6hikrMCDWIjQ6k/OvB
RwFMgB8IgCiRlCyEKkug+hj6j0XfvKpdWJusoefzfr/PIBA92fAHyNJL8v2L3+eT8o8uPy23bjxQ
5PxJOkaUCHULAl4wI4qzMgcLUYBQo2VmWS2SW0z2S4a5Fbvn0tGkcdCmH9KkcHWmquFvHlZP71XB
mFW8j4RQ+twKaEOrt192EU7wEmVpd61TlNoXokxSDynrdJE5OFzWjVpoR6pQxofY0EkK2q8zaNt5
8h/vBSQW6peELorYS/DwBuiHUT4/VEDGDUQTQZ1jYqmbyq2XrPpTOpxPfXHDgCvbgsPit/v2w9RV
MANpcKTBhoNCF9vT1jfGwLty6IVgoNIVF5pEsEnJGSuv1Nd6iaxmog4iVbWDSMJWDyDEhebt6NCC
i7Yt3A5PN0xICUV6w5cO+F52YhHMGZSt30zG/YpanvuADoMpgacqu78OCMwD6vzle3+/x+zNNXEM
sKsLioSKr/kLBMaFHhPo9wjPMiBmdnFQQkVFMJy+zTZ/INUoKXijx/B/vYuAvIPmVakL26q0EyLI
Ufyr7Gvgf0CCRVJ6cH99eb/scp5j9IGoQvSE6lmcY5B2z6RaACEYPogCyOUXj93gDcqKF0W5hSld
PQUM4EM8IagGbQsQV5RKV5kEDsa69CJOlgxuQ6t6mfQcLuPBpdOTBGfCIb/ZIU9Jes5/APSqrzX+
//FbMRBwfrHEgeJYQj/CYj8KDL4dyo0GZFx0s8yx9fz+i4EiVZdr8lYPCOlWtkt/PAjuL++805P8
HqPSXdpMrfBw/aKJNdRWU+FcHjIgpaBWRuNidKjK1sFlSJcDe4XQ/E7bXKHaXBB+H4Y80GloJxhQ
/cY98Qw4UhKAPjtiNPjulhTMY4PonCoN/GgQy2ZcDcPFf0NVeclNuDGBlzyUIGJ7zFict2DeDo4N
BVx+RlgmmpmH6dH62Uo/X5JDyV8BoFR18vcL1LSH7an98+gNq49tL5My6kxbcyG9YXW6HZC78Bjs
yosf4fThfy6tBjm/qG0/Qq9m5v3PzgH6XW6+ZkiN1Ldt3n+hWjyd17ZV9eAZS9K299cbJ2886A//
KJ4gVKYpetYMeOE2lZO9wa1oUCMgODesqVpYqGmd4yFdyMbE9xdxraiQqUjEZbRqLOJuiof+dXfs
k1gtWk4DzdALp+7wSeNoVWJvGPiyLvnt0xFvtuFkuJm7J0gFRLDfqG0wp/0onwgz+EeY/OUwA6ej
ge715SOYOMIxVfMexqzJreUZbqEJQ02sD7eDOKhj7p/ybHLkMUd5y2qPOqa3x6z+B5LcACec6GRc
wlrXF8xIsisniZQ4ScNfebxWIyeWtj+ryLPsw/aKK7m00tencuq9f8xDCfbfx/yLvmofdLX2PQge
hyYzd+bj6bs/gXxC/rM0GcU8K5z//p6jmwC6/ungmKc2M+c2nOUXi4ZDujI2QU1iTgWr1VzafG/+
0+VfLqXx0Wi+b0hZW+dIhv057AAix7DQFgQXX7+NEenIjjZNqWIV0jj8XWJtiKNaOTPhJKR7ZpFk
Atnv4HfJYp4qQinpaxIXy50Rxp4NgbSN2LWfS2DwuxOfxjOtWe+/nmAPML8OeY8545LgAGD0IXly
pxJVlRw9YBnJlyjpVmDBGuDOJ8CUnhJlyq/HepFLEXpHvDuHKCY3nb+na61LKC1Vino3E0hawhf7
5AfKhTpYe9E8ornyi+7XXOETm4WTno0fnxgkVNHGpG8g+566/110Jnoy5zVtKv6pJkLLNZwtxOhm
oHgfPkDm/jj+HuD9Mrf6Q0e6KfNB7DQoJnxoS7Zr8bfwQUx5TmGM+NLO91hD1B5Z6CSUUUsBtIer
KSroxnny6LiMppecwSFNbZtwDs/zBRXzya/c8qiB9JFKOSAJ1bjNd5MbLV522YZ4CmlDuwoA20XH
0ArZllGA11lG91LbRsk73y4++ZUxUR3Rug6XWwsGWAYJEbXYckM79tn5QsFnLFZducWKqa2TnLtz
W9evZa6usmUrSsdTcKVOPaXiOrwpIcb7NyUZGNHdXYLrcTF7LyKn9YjtG4QKSE+/yuE7Qo2XyygU
IDzGNhmV35TuJDeOLBx1c6ls93UfGllaY1bs725GM2hQw1USh3O+t62d/ekeI3sQ24Lo4XpyWdJ/
8FN3lXMo9MFvSHhPvnBpMjLF8A9scG5FyYmoBEwNpeme07pnhHq6uuk4hnppLPLwX3DdINaFQWDN
0meosFhfi6Lonq6X9A+XJQihNG2nxiMqwczjmohcukbQE3CLltNNAp/QICH6frqb34M6O8iaI12G
GSvekqHi00glxjvX3PHs5dMKaRhCzWZpiKZmzupgGMM+Xc5DLbBlCKwhsEF4+AbIt9+CJPfU/PDm
z2/ww0nY1SSwekED4GzNGXLO/u/nYFREEf2cVFSAd87Uun9KFDnuax/aHquEwmzQO1W1m2102adF
B3akmpgP2J6Pzo9cSM6GjGzzQ+j7PkvoSEOZ9CAIodMd8BDmzHVp27eskhnxXSiHHzqLGIcCZyTz
a62bjtJEjbdyABeLqnBZPCT/IcAfglhAn+xqavLqZynYNk/99b1Bm1FUjqka0vcM5s3wI02QhAX+
vgj49R9iPbhyF/Wm2v2L07U26914qCIEyIrg9rIEzvEBtJEgvb92pthlLx60b9QsJckujR18ghAN
D9JZ5LGZJtmG4gIsoSg81oZ8cYr+O0QuHydDWoi46cbSBGkY5qHr4qdHgvPA4Kmlz+NsxwcT6GAG
cPaWA0MIZWhQJo5Oma2dw3tQPJhiIb8YDfosVZ9NaKjrgZnuSUJxT0fq6MPGqX0EtMQTxFOTTFHz
96SN3Bs4e6eFCW4vHDxzmapqzSaYVPyGsfr+KEBQe7b/5Exyw0r+TQ38mbmOxhXzpZvAbcBruG4G
VgIQ7BYAdae5Y4MRS9QSwWHp7VqG4zMFgGOJHpQNr+doDj82m8UUbHQd1UC1ksdqTTi995hVDyWY
7jfWe8dqMy3Mo0hLlcy23WR2YxNIGM9SbUAu+2ukYQVrgvJh3F75xyibeXNX4wj2kUmI3OU907nJ
E7aXFP8iKfrIX59WJPWONg3XsEhtQQaclSXIgW7QWCmkKTKLAvJVz37yt2k88L8yPh06qQNGG1Wb
4jYRIVja8j01RH7fpzscN0lsqxvW/trkwfKp6QGiXe5zIRROtgi9KSwnUSOc41tL6JAmhxOIh2K2
TchBxNyhToNgQiJKdcNlGKjU9mmjOqZm5gK9VpWMcubUiMgYj+tlDDSrE/lzcZtrn/NJ/SxtNqlC
bjY0MnHuVmufZyaSSe2XF1zLuKbYzLH7djqDa9OwsOzW4cM7x4ypQl7JoKyDCZPlvFtoBNA8k/+4
rd4rW9WQk5wkJ03BXXg8NM/pQ0XpQpv0FE8I4wBQfAN83TUojBH6R8q/Pu0pk9NPMCV+/wrzOyUl
gHPoVBj8KF1xI8f47A04FLsgxuuPnGzM2Vwmk2E04ZAKKc0HVbKB/0+EoVGaSHIG3xob3uW8wUOL
VPgV12XIx93LAK9bituai2T1Bu/OEez8p9ITGou/DodLXEoErg9b+1HpiulfoIH/SwkcFWIr0pA2
GsOLPPu0n4wW4jotjv9XmYAermEmjGj8sYd9VrVqhJrtygX/LVtlVZubbAyNU35nlDJrKk4KSext
A0SgjJFDsMfYu34TQXMrTWAzQInhti2ZGFj3SGEFqL4XgWd2jUWfWons2ok3H1FTlBs/JadaeIjI
xNBW57Nh+6aFDFyzjCCABokEUBNDC9rwm0zImgeu51iq2nB3lyMcJfDUln5wNA24uwQTIOy/yG4n
hpVMQ/Sje+jRSs6NGdq+Y+4QkJ0wDKpUBQ5yKAyfg6EnEEd/20rUsEQXwRjzZIP6p3Im7fz0LOsM
IlqL8KpGB81kizuAc6ZuweEaUO9XKmZrIOngLMWCc1VTuueBFXkt8Jr6QGjEFSNj8VZoxUo0ihxf
qaPb2lZAS6FgLMl8AEjjOE/qUB7FpgNdJFeje/B3STnOYX2PBNYvicP5TvmkXNKfzJvlLRdTRaLh
PDA1gU9uHVYRcnzqmAyhoL0oDIznRbyHQZh69YqRo1R7bByQ6fytAW2nXS706J+be/mVb1J2e8yx
o+aOfFIGolIbjKEupRtN9KKow8jezCKHUCC7GigDVHvVHpjMps4bcyxpiSC9FhKvj6f67IEQUea+
xZzW2uhEtY2D2aXmwwL5YmOTZtA6n99RMKjyj3Uuutnj3b0+C37gjW5m3Qd+AykvZhMdL6z0pdSV
fycFl6remxqcrkmmIKQBbKjYCm/iGyPkInO00Fbg+9hX5TDeSHhHQccVCP6osMM1Z4ZD3M6MFNvJ
gKkyzxY2WZyUJha2cB8w3PzMcIME+PFn7Ix7q92pTGQsJ6XoEY7winG+u22Jetp+YEsygMYuXyBr
76II8iIXvj7kN/4IpLT4E4W6K6NgX3FMnHHWbepX+ZkmK4rKAEwJr5YYXSz9lPuq9exhEjXASsWe
sGNYRiiSqbZ9omLMAEVAu9EZI5/Lu9W/rDtWEnN4Mzq2B99PcaJYYGw7LxPVJYTPk4VjP3JcBOG2
WoLiX6byZcQrrmCaS8jr8FCwGPbnw7l8rqcZtUjzgApRvzHgSm3IQ/oUBLkqOnKBMkh1A28CAmXR
EHb1fn9jeMybAEtb5VFPfF29pkm044jKsi7PBJNyZDhbKBsQUV6rEV76GQVEdJ+uothHk3QP0z+5
8wK4e0fJKIDKivmU4T2HICW+yqAsbgC2Z9vOM54Le+b3SIGBnEMB073ltwAxpfLx7nTP3o3H6XAl
J0QWljeXcxCi7VQDPdWEYiTuIeuJssGDglTdEdKvgoeXR93sbFZ/fdGPS/l3mJ1vjIVyXSi7JJ92
ZcNR18bqJfra7WQTa+sLgiXY4T0l28F1S/GhB+DkLjdU4iPfwvDa71ys9nmHaDW5vy6lgHa5BNEH
2lkYQEL0cR4Vz33tBCz5NxC8UasPcbmdYcBJBp9frwnsvrFq1cu6NjiFWkQLvD3nD5/FhwekjTwy
12D/0IF1uXiI55pH8R7vvCaDvU5apQBEXCPEsyURp+o9S/1vuFcA9tnva/VfVX3/UIdKsKdGrUuv
nQjjz6BpJ6IVGx/VKZvPjy4L7FZAGDKsh8GpIn2XSLJ5laVjipB1Hlum81qVFFahO44MLObq158R
YyYRCLcxqR26LgL1tW/e12p6zKcgccGvyjqPZhhiPJENJr9+uHHxYB9vk/6aJ1OQfnZy9vsl60mg
bqpIdwR7OH94xzJcbRAjC2tMXwe87kx9aam4ZcKQ+78mj6y3/XMMPjHbTOnyxjdPd+Ul1yVUS7u3
S5tZpy7zv/3v5AQ0qYwINe5eIJysaNjEIi7NNzCtdu1XpZ0k0Yq3WyLrXILAajDBHTNLrYQt9Gw2
PdGAjrTQNMzyL2h5c9pzlhjIoxoBqWcBPm57WMuQf5lXxlOi6dcKmGQHwycM16Ff45F4pX0cuoTN
gRDavZuSkYtfE2QIzRxJVGbYCgve5vk2mfxlHYR1+Vtb8GKu80ZOzaZlgb+MzIqtiWUUT2Wh6wIU
2VkdxiNsD8uUvW3xbtn8aYcO0sViDLTzpSgrmgZ/zppRDg7XdVroROj5NMzuKPTxkPnXS233dRvd
85gAwZxvLa01oYbwFvrUCMhx5zwlMqpNK6PMpa6q13KsLNeUX01UskdKCPnQaacFCGlTk5aR6YUc
wHKsvl5t7LR4ACm59cv+nqXbYzBSJn9GnuGTA/zipReZlUGGbB51Hx+86f2MMhJoQcUq/7QBd64I
mu3S1+rzTQ+xlLrvNZ9pcmiPqnkV2R2zyjorr/tnWbneMtpGOaUIrjbE1VxvOhqhVhN082Mg7IfK
n3wfVFsvZAkGOrut2KrWn5kwfdQtf22I/lMpx6MsYlti/ZRAvQBjocpVy4Ru7m+Y2DYOfFTQpns8
reRYLNqC4TKDjVmPgCJCNnU0RsYMX1zwMPq5+xDAWMiBWPOImuyN6YjfCYF3DdsQnhvIzeTrUG6/
rOg3sKsnitig+4qlmAmQv6eLd74YzaXgfUnwy7gdJk/R+nbMiEBv0XDluPCgAS3Fh/ALA5aYwDz5
X/3FEs0UehxMQ/092S1PTNnl4Whm4e55deEI5hLEOOvt1ByETfjhnnpiOCzuYhQI4+gS+Mv9fzJx
CTgMePzhaf8eV6ud7gm3mx5GSzpHhfIe0Gaktt/n3eBj0ytchKH8EiRQGO3QSObiDpoapsbyoP7A
Fgv6bZHt+m8EBPuzd12Yry0omoMoXAGx2i5VcmhA5ZY8LeYB3/UJsyuU+ZdvmK2YY8ML2D0lYT0T
/4Rouy5kJR4Ho67fbHf/tphbVfFAlQ8oed5BSuRycskXggW0JBEe5a2ahQ16zq+JqgDxvUp4ym10
j6t08eyprhkIcW7ORBC1UUS7hruSiYbKQg7BYFyDPL5jZi9js3Mf4JIui+tLXAyadZOqK0B55WDu
XubVHbAJQooMkSordjhhLj6QzMOcp35muxhmfSDDnGgIvlvva9O1l7C3jTV/tXwwA83oNGTCflO6
RhIIOKvTrZB8ytJ+H0i2cWvLFTbCnOQzH8k4Se6/MFu9hdQhqJ3GrrjQTDOHQHO1P0CJ999/DHs2
KUcYK0dn10NKrqSEVJrUfMD69yMkSuDUvAmuImwwWVCmyDZ54C9KYGYk6D4eOf8neGiultmX0vVT
bG/smyim84n9LwhmF3MNdsYx4jVzxNxLTy4YaE3TbB6XVCOffcQtlgZo6LpGX16/Yaum5oN+DWWR
gi9D5+caRcbeukP8O95DWm2Lk+GuhSe2tNh3eJ/Ks1DeRutr1U0zLjBFbqckiw4DoLsiSTLx8j5W
JgR05UvOQWoshK6ep4PQUpjumbj3sUfP/JoWQUyJZoNflpDDUJ3mv+WsYHird7+ecFsQUe75OIel
6BtBWP19PUbIDpoZldVF0VmEKySxhGKu2jIGb5bLrte6ZR7bgqlfwWR9PVSwOWlIgFQN8FYZkMSt
2vnL3m+F+eTfAU1klP6wZrXCGEosl6rl+nhnOoyXBTlE1zp4v371kqMZfJCkZyrFtPILibPPYCc4
G6HqWwCG+AXGgSw410PoOC6ahk7tlcW6/ipJmQz1jdyNyx9iENHsojACDb0MIDzgZNG2mAUZVprt
RBk+T/Ym7ERDZvT+I3ACU5+WWe/AyqhS3c+gTCF0TcbUy5dMY/vMiPnn7b6N7WprfyiW3ETIZ8i/
0pht/UhI71bZNuM2uB2f+Rh+hpedorXFTqm65vVxMYrKnt6XvowOlFG6jO8EGuXwY5ERdnUjozOD
0cPlbd8/O7Res/JUsTi15B+feEJu5n9Fck2VqkjXQoc1A+BHQfVG2L9IWAOEVE5Y6CL4kxJclp0w
Uvm/Nde2gT63b6ULjNjscKe8P4oqMAeqBgNDsHDEZWeylrecUuSy8wKUBibCSqwJbWaP3+nKEPBm
q8Hf9DuAX4cYzshwlH/ABg/QP39HIOJxt2OhpzzpAncfDABAsgvjDItPQutrygMdF4kckkf7v8TV
vQGaQ3JXMG/KgmsO1Xccgo9luaqRJg6vpqcUYqWGossrL+NtaIjuhS1DUTp/GJ+b5g+0o3KyqzcC
rf0f0YOx9y42/KR/1Li6oLSjMdDYMwpOnvDz/go6rbMYaKoToSqm3PVeyQ2u3iyjCGY1EYzmAXun
nNLQmHNkcz2lqumJ7QdWCcRAATYNAW9PtWDAdOWIcfxlmvTx/MFVtPteXSEKIydg0ijgyIjHsXGa
UMdpoCV+d9bYitFfdkH0PC1pWF2rmgG36IudOnLdKGK7s9XZz7fMWZEFroMtdg8EBvkfgWgV+y34
3Qc7snVGjWV3roa296RvtIE2R9INbZjanxEVu9V3bZElJNzSrikNo90zjGCMCGr9S/LD5BCmdgLA
EKQC13HX30nW8T4L9akB/UWRZ+5uoS/FXu7BaE/r9uMMQLlP6e9W7KtJfYUwahiY6WKYqYImY9mk
vtKB5t3h+NW/Jl3nYcuOEHuWTnIBp6oPZgB23U6VVpt0dLZQhPweljpxckEPFTR65CgkE+0OtCPT
ZNlmdG47tgVXBLGES0+La2EwaahFPP3t98nYZpDJSBWFJcATlOX8jyXHvsrNIA11gpom32m//n6U
1rgwK7IKSiEap4i4HfwTQ+Miykgl1Y/mEJKXtNaNifNeSDEX+BTF0oE/RNT4EMe/AZ5r2epepOr3
EEpAU+AlWKY6NirlbSAKDRhaNNKLiyldTrzpaZ1Z6stSWcuYAiDOQPpsuL5eyobXHe9EGjPAM1zB
c10lX9OmrraRukckRwVPc1xPp4Nig1lLcOMDiTXembREqh5xVEcJAQieHV/3c7LYJYX6qWF8qRbA
GGbLkDJGzXr8e2Hoszf8sdlGxXMOAFIhvf0xOVhUQtxcM7twLCUuR//iD2GEr5y9Kk/B0wRJ4uOp
xmRTerNggtjj00/zhCDPZ2KF3mM9IWFRTaDW2ACFi5o5k6U9o4xOhkMh5nU7iaBt61O5NYlpN9ra
sqEWcZVSiZVQ44dq1PbcRkJP7CLWDa0pJRYj4+ol/jm9hX10l12Nn12bdkJeCKUHIpee4/PQ2Tco
QZ4xAVWnLDNGOcHP7bi0XBVF3vqjcs3XE0TM5jsQ7KGCduzj3Hwk370ns73UeGaeJvd76wvUci0g
S9IA6kArJ7U/UolgMwxwKqWkaW+OPbPHAjJ2Ca1GxYHoL2Gdmr56ujohlyH2kBEjAYNfPNyhQPhT
OxSPv48LNd93ysvrTTkH/GuaNUkqF9teTMdQKCC6ecnYJ1ZKoalZsh4rz9ei3JXZ/Lr3sRNES7Li
k9IhXB2zJ0yD0D9WsSVvNUr0u5XiZpKSRrT2uuH702VL4O9Uky8iGqZCPxtuCxPMJF036BqEnKPv
iOUMxnZ0FAwNEc6Zmcx485mQxwpWeBf42m9sHZ3ZOpp3rxUtgcvq+NdHghqbPvDmJsY4Mpe862tB
HA4RW5vuRkF0v6LUc9VlT/Jcp7wUz5Z1isKKNmGuW8xmDqESgzjtqNAa1/z0GbZlK0piA7wxWS1z
HhyEVh67e4335dh5K+ZM3o/CDiiRYOlwIVMpYX6eav4S1AMtZcr7Fnr0vhjm00459YIF6X7zJGFN
oGugrOoFPkto08H9/VAYrQVCCgC6Knx2/N27lTI22F0s8OrlMZq/DVweMHLXf9JFJ2UfK9LmIxq0
7spef093hiz+z56k30gv0n4wNiQh2FUiAzhvTIWyoZJ8toBJE5IIc0Up+15JtW155tNvkMBsYFAA
Fv5hmyWYyV4xIQdEY+WDaz6o8MWSrag0IY1xmDHw0iayIWHNWoMtHAUy+M3krujJnIV3SgdPsymy
cRQvMxqPc1f/rkp2jSyFb1jDqOJGT3NzfnCaC1WMAsNSGKnUaBSC/RCLZV47IbYSShNBHXQLK3Ni
EyRpYxQyA2ia8xfCEZ6FQt/AYVSUFbFoj3IzUJcLtvzb08CR5h8vsOgQGOQ1nhxFkXsoIjubEsJL
ffteplz9AOvd2mfp4WfG/es3S6XQF/SAoROs+DRA5+4KtIPHz2WCdid15YcSIRlw4l6XahjC5VPt
B7TaYOOsIvPopWNOlVqvoromthMLhVaPiG0WLkNL/kc0lCVcODBemj3o+ivL3B3OG2IkZcLdjxYo
JAnz/3O+efCZwAulPEwbAFBh+Dsj7R6aybu/4HuNHx5XPaos4Etn2ERxaS1dfH7o/PIFtqz47mjc
HgG82VnrAJ5Z3vL+4iBgPWSrLydL1CAro4xrtErwPSAyUAQ0iGvn9TY5D5NW8WYHzft9JiS7f7jN
R9Go6DERGu2sB4Fa2xxGTUXqBnPVDoA691b1mGa8220bW6mb+RUTjlPvoSX268XbfPU5hX0vYpNc
bluyzdO7moBseOzYhNYgdPnQOLMtUaV5hPRl6MSZKQTKz377ineHRLZefqImuC5hEOxOjDfim5md
ncgciszDFd+C+n5ZrB8HkweM5E6mWWVSiowKE+hgWiMSNNCptTpuCExUDIoupcrJ1IYy+FPY6smC
KnWMR9MW8Pi8LkAYpZDwJMJ7KVn2hmjNiKqqTPbOEMRnKOdGXG6hvmzEJMhTCk+srLOShbSdDW9N
JYjdksxqcTdzt41buzB+VnO3De/aSZwgEOrtbtTo1grn3H+NarC18RU+12f1+0V5SeQW5AvIfvPn
kdXr56XYjR2b07j6aAD0jGMAymliR6kDewQndvhTY5YojqCrR3oFMqKPNfDC9jowSylwMj5dqkvn
XzUnqVPAbc/nfyWi35biAVyNclhqAoxYb7VpXflYg9s0LGZHa+246rUZDfbbKb332knF6wwZ9mo/
3jRO68tEEa16odx4OaLFaPNz4KLU+yYwS3c7zWivHU0EYDwtLia9N/c+IKgB+0hmITM512ee+GRx
+GFaKa0Wb3IkI2L3iPvy/eU+BxYuEtBoJ3S5QqpMljBbl1bPdY8RDnXNSSqIn8ky/7ssL11KY4nl
ak2uWiTrhB3nSGOI7Ixgy1eVmrpQsNqlL8RmL1KeV7jk+/lGLLbDTf8AmlQoTg/D4zcP1ONCqMOb
US5G4yqEvO7BQZs5fxqUAKeCocFuIo/9whIV/orguTFMDBHXZjmQvax7Iz/oT6F6vF6Wpfuilzrc
HmM0wPy16xAX9yObIhkbZi7Yg+ZiYrp2f11sA4YsUMWylI9XYNGR/c0IiVSQc3l/WuKk4sR3iVyy
+NKlA6dgoNpNjwjdOiwEcmRivVjJoqAOzR5U/7QrhBdl+jHfotnYJY/zxzBEW04sdtCwP3I27R4j
eMq2JijFW020iSAuIEcbYS6LIMVq3Y/7PR5AfPlPB2aBvDRxnMyubgg59z/RhdMkbnEL97NQUw/5
dA3zopQQ+Fb+d9kbwGQa0t6xyOl3o2ejxgRzIN1TBFNyak30NsV+CsuSZy7GsD5oYVONTEKexIiT
vwkx2Vkob7Sg+uqQrM/RjBkDkV+GZpZeVB20jIeSaNc7diBo2KMhVPyfCtgsU6EwD8a+WOwCu/4c
E6Tw3vUjhvf/Zi7vqvIigJOT4AlNfRximCQsZFUkXY2uMUiyywkTUt+2J8XK4imCm/5u1SHChTiK
11q6x2dUlNHWDwGn/utRXbEA8FBO92FZzRAGWkNm28XoIGEx7bCGLj8dNWsz4U0ABpdvyvif1uCf
gHquyYZhcX0Lt4TRM90fMzrpeFvlmfZLlu4Hi0YQA4e7nnXtS3CspXuNrHz/mQG+OAIkXavhizD4
kGgFRrJlN941+4zodZmDau77HuM8EDbxhjaGIAPQYOW+4gLqroQykizrRDWK2aMy0ddEthxe7YES
i+Z8br6e5dK7UJ/2fBhBln+5JGPb78Mv/KV3aJk0Ae79TOEqmjgHqKdwyF5QxrnFCaSVz4DmxKyw
6LF+nWkXFPW7lHKYbqZ/DCNlEQyscUSPiY1bnleRNfMs9Jo9X5eE/WgL9xv/YLpvd7/+JtkAymQ0
0LFumi7V3gVLHs1F2K4GFNlB7oFAWcIgU2hpWk6p1JyTGfgrRwpUmPITxUXSKKLfKv6Mf/nO1hxC
mYlklGle639DmXrHnehXFwtnsVLTz7kf9EFDlMXfkOMIdeZKTtBqOHCqJT7pHSCb6bApbCWskRUo
A/lsjBj5i3EINrJDBf2RX3PE5Tj2C3gEFWnNSIlhvb2aPa38NPRinY2gGlDRungiBJW9ms8GQo+A
MQlFlrYN68GfNkIU77fbrvcl89gtWxUIADaJXiIjol0Ohl0O9tIEtlsszNbin5LZ1x3yxQy+xsc5
/j79DesPGGg0n0DGhFqNddOf9fQ3HmaXeRe3GbOo9qw/E8FCs/LrV7jEhTaFQ/0kuJtLMFhe/Qk1
HuShOnDcD87t87ls0NIWXwjvxseyB9kfm67xac4wIRlCqRAEgr5UpJwYV07h9iOUW/dlDZHis7qQ
Lt2fDUZ+3W00DJsM+L7G+8VGliJlrdyTFZLDZ1WHjpxICChdePSMLSjVNrBn9T9V96PSyV0XVURs
2DCIR7pPyZWrajEFmB/Fjbd7hh8xx0ZxdjHR1jj/A1GaFDdz/cQRm17x5kLPCvl9GHIDs+bXySvx
erKDo+HrX8avOtcYwLsC6TZllHtGtdF0tCapd2uRTSOxNZGkliiMJ//Hz3T5jQt6XmlO/Q1Vffm0
apN8HD6fcF7CJeaYPUZnvSLK7lU8eK7yjs+on+qgfMql8EtRIdBG6zj0hO/EB44R9YtZovPo4koS
JmyoHyQqAgzC2p6XNVEcr4GX7bIyxSlE2GXfKQ361loKp2kQM66o0kj5wsvw9P227vVGeEyUhLa7
Qc3zocfv3qELF5DfZCUN8NxPP4WAh9QNR455uFFbfXsTl3Sf8wuCXcHRmwI1DFCd8qwPv9r5TaNa
UxoMgE79gc3yTlBfTzUMeztoVa3XZX2u0/5uOyVzqh1A/eqFpDlEKK/QutegyLCg6+1hXnt2EoiD
WOi27vhPauNIf4p98LjKPg3oU8/WurDErTDihnOJrKfIOl5gjavH8OzAf1SLaLylx5QSjByMOMXO
c4Tbkm/gNkpUcKN/Zg5Q30GgwtHM7FdIsl5KOGeMUWogkYMzWlNqGNIBrmGUJr/X6x2rRLq9K6Cs
471YfoDZ2B2Vi8x1kiTV36yQ7Eg7IH+L7sITXRSTuRRiotroEKWZaN/72c43WFLJPKcmg9RGOKlr
6PlslvsDGaJXz3awp5UANbSGcheOwIhzcxilXxDIuOr+YmMmZFW97qKdH0vR84PRa11MJKUk+XBD
JVkg7my2sQpMxuJ00uX2QA+aXHUF68YZRzGFrQoGdVsIcu96q+9BRxmnakVHhhA36PsevWYlLUSK
7ESnOwvajICth3IBdoD2S0LRQv8wP59Ta/pni0vLaZY1Nz6oP73GYiCAUaYlHuxwhCtzg15hv7ZA
aNib4PDV34o0tyJ16GfuoLeQZ0gkzAntsSAa4xyW4BKi9jLOQ0sHF9hsAKxb9z+2aG0uGiREUkxY
Zo8eki64NizTEzabL3c6SXwcBIdroTQ7E/bIRtfxgXxqCboe1pB89dBI29MR3X5ixKUtJ00fbluL
BUSG+4WmudhoBVSqF3hl3kRWhLZxmePGZCExiywX9sTHNZXaJGsA3pikM4w4RbsOyjcSiKRSZY4h
N7bMeWymLmDmIQMJHJGsK5MKpZUDQD6fENSLpGprtXoGsjyZmDpYMsuvkiH4DJ04pAvO02bAeRus
vCpOga3uD6Djq7teRJ82zmvv/9xfANb7LivOVaCjeYNpLLH/4WW3LAe1MFoCvaGuzQhDI3IgVgXi
H5rJB2y3mBfuFjN9eMoZTNTAWOw6Mz/Ii7BfcMvKj5rZS8GfbZ5AMbd6xVvC57YHVOBb9TxgqfH+
tmTPzOYLYPG0zSVDcrUvek9zwBFgyKoQ2K6uE3jgAiMqZjtKhIHDHA6Q7bBk5VwfbHqIt/1/RemQ
wj6QZYfkPbPsyBfUVf1+tG/vK2PA1RIKYE7F2IdcoUDq4x7z23CznSueVC4vhlZPh/nKtTzsEI1/
Qeg1Aq+WWeE1rnj59Xs0qD7+EdvrVyzY/HL+T7BxOgUnUfRekGewVtBptkrFJPdz/6UWiou4f8E+
QCieFaj+/AliFftoYh1Sc0Wk4HlZCNVlZW5QtHvuUChcha6vlLUbZgs+F3EeqfJsoxe+aoZwksMn
x9lO+A3CKPjuWH9ckRTp8/E1tsjTSPE9hyKG0TsiqMKdSd7Bg6TlTcpGsbJ5J3+Rw97dUZbUiI1T
mtjEqEbBqm98n+elHvJM3Ujv8Kh4uis2cKc1rNqmrNOMdxbQEkYK/wuA6Ue9ufirH7VEDUgrH2I3
p4liebb/vlZkpHzpIqy4wer6G/7aPFSjkG94BSe0St0gbZLthdQiALM31UX2B8bY5G71NeatP9a+
5jyHIwRTCj/z8b6cJXJpBDn54Mix44lHcLYrFmYoXHV94TzQ+80w65iJZjTKPfuXQOJ8A4oxHjpZ
uP4ml3EoYf7r626ZgKslak6yiHuwVDKmAK/nw3A12d98mLyRPHreiN6XJz8g7ZYU8mGvDNu3wNT6
wIfhcsFwnZXMRGLhWhP6IHWXQDWp1QRc+Nm6UpFtwcDi+GlM3JFz5RTLQJwx/JlN8OzIcA+lvZYh
ZYyADFsY6wSkOX3PrRd1FF3xV3LuR4F3rI67jrqy7F9TYDonbcIclzO/G/wKFySBKUTJWsJv7rxn
22JqM5hpK/gWR6fECIwS3Ek589OZeo7565JfwoESwIgQpDZE3XAlporGDEMRgKxEHEeO+pMEhOuo
TVZ0kxeMFUYCsfSg+4PXMLaIaIvDr0poApQfCUb18SzBqNeQeNEopypkClMKUlHz2YbSR0XYMAXc
BWi3OIS9oauiloc4/+/qa01nbmT6dMNRIb+NAAqVMVcBtcwJxz47953j5JzRu1tSyXpYcfPkfk/A
CFjPvFAoX5Hkd1Po0gt9TzfUgjjyGipiQ8MxG4GL9f1Vanojs0efrOr+1nUyDPYy0QRw1GWHjCmE
bpty2Ugy4ScO7LBfsNGzWEih+VUpm+bN3YWCRWd4GderuOF3DIvUB0hoJehFh1fDbpnV2mRHFdo+
m8qHO7VbRz3qtFta12AcAW48Pz8F6Q6w1BIWSe+eYjnLoDWnBjBUGhO1xU+y1tqCePb6K6y+OX53
92oS5avYnV4Kq/Nuc11ix5cgMJu59xNG0gU+nwnxXUeVKR5Bza/eNaBnuUg5tyiON/+wDAUDHW7t
oM57WRDIViA0ODofpnBJSHBGZQjFAPePXYJJIsm9iUNZ70o8lXiOFaWeLgriXRAN9tcY88Ay9fBr
uZgcxu2U3Ha+bNaUleWUTTSUqXeUexdKzD4XsVtES5LMvIX2Y0zzexC6yJDk39pbQZjlofF+Fqh9
rnYlKiU8bFNAzkBvD8TSf5etDrxZcC5MRqOCFPmo5RZE+PgSnE0aZrqntHdeYe64yO2z0poe4gUv
i1vesfOoxOAwDO3DzCnfE8o3AZOCQ0zD0hHECSdW3HbUaLWT+mlFXjlncWNUqKuEWOVM8vvgxWKW
OPcN0A3Mwyj/5RwSRIXufUX7xPwnBMwhhbhdOfw2GNFw6M3bDZ7VHqoxrEYJRaKV7NLVQK/6o5z5
9oTVkDRuuPEW3LspdpCDTUibxQysXVjV+IzdTb0Fw7bDtf+mB4TGEB5Cn6tvCBSHtmZ9AM/GstDb
aey/+1TBfKCjkP7CxUkCHcMuG719zct8Ss1Q/lAZLaTlKA28/MTEhd1Fbj40yJKDdpD4W+stVAa/
H7gsbueW7WpliAI1OWlVKp0mQUG0ikZmVU1kNy/RPB1VqBE/ICK0pwBaIIA6fKjBfGTZ28ZTPl6I
COD8g/rAEBfNUFLCgzSmHTTDx6Rq4f+8rrIIhCdF0P37P7k2k9Tv5S9XLHPZRoi8qV7BFx58aXkG
395BAj3oTzIvvgg2FC5lxd6ImzibQpdP/JRk8uYJWBy0JcnBsDa2dDx6pa+zHgwGwRMep6JN4UCm
ynhGeeJBstRtY4vS+X3E3JJLMVkuK9+V2jL0J8dDA5BzjB0wVstP/BWVbq0KkWa1x8yXfWtjNojE
zYOrtsTvdJ/Mta2weIceM4p0bFcRMuRqYg0bPO0rwaKT5yIkn9XbMsd/9zogexWBUTwV2GVYPkO4
vPvNqou2s7DcAzvL37Q5ToEb5tm0uY6ORDw0k+T3IIZthvHR7raLYmPz/1nIyXa4NpTsmCGMGQxV
XAEKyrIK4MTjP+IZ1DukGXNjq8t3blcJcTI5oSW5QCwsoCa2fLkpJ5t5QBUYBpWFgIYBoflohpBu
zQH2gudbWzLQR0VAa+cb5Ao/QYjOYi1w/J/eabUuN7TpdpFTZtXSQDocBJdwhf2POxiLG1H1gcGw
mHIHZn5y/r4QqaWnFp967daaWjZ+bPr/KxqmUgjHbD+C0xXcdmttHpHjEz0AzoVr6c6g4j9weimG
DUNP0Ueo8yr/N3cbEGCj4GLguK2EVMKwR9sMa4Ga/OGRI21qnbyvL605b16XYdxOwM4HUI9vU1IL
DtEVNSttGRc2vhwDYK05AIRTfzn6oRzT3vwigOuc5lA/+9tpL0guP/NRF108QZ+BJM1R072MWfvS
nJNwf7dLGgb3JHoUs8NEospelHp9dkJtoiMPRT8wObb70BXiJRuiHuZkuHlC7eMbil+rKGXcU7Zt
7r34JgF+kQZi74jnh263DbdzZ5SFphKJltEeGlO3NTMgmNHBvQleiG/EsMEVVmZFkYnK2OL72p6w
m+pru1RrQg8nZcnrE4shu0ncJWjSoO1e1Fa42gcUUWZSNgWA+3oypc8Dp8gIiHEwn7oJGNvgHEhK
no0dpzmrYWHK4j8zSnG7+kC6NvEMobBXjf6Y77EfmMFS1ew7paSc+/xa4/XBkmip4fquAfx3Rk0O
bn9tilU0XJWg24/u6NN1NCPEOCieproCB8By3ZagdtdtqzCQFw1S1cH+KhVHXRGn4pnQUoEkCI++
m1bquZvrnJKIyKtr3ofrGuJZBRwArDRy2TJQjc+9btrocmuKU8xnH37tIdBPTfgjLHkHw+ozM19w
UgwAF98aygpJnkQRJZV7Ndrb4XOeT+eQpOHu4jXYnrmY/yr72heuOrTeBjY/dsktyBxbWsM38P2/
kPj+Vhb39EYT1RExq/Oa0RXQtBzvWZRYuPtNfNrWVV6HgLjWsa0+LK1N1Ny6swGXqfsSZeqT8LOv
leogQJQSNPNpQxr0byQMkc7kPqNJA2HCiycy61WIgONCPOOiZl7qA7t0DRTo6W5TyGqzyOWli0VA
xhewr1RxU17nGec46Fdm0xwYOXk0E0bkii48zJe6cMEaphm9+5vobPJY0eSO6+HjsrYflPDIc91F
Gb53QTV9+zdyLaP+IguFr/74QKC/vBKP/IiCdtwhj+MT94e3jxF+wf41iDJK0dmtga6Q6xFDCGry
HZVES/FAfD0ZA/umRPDaq1rY0nsaMblHw+X5nAOm3akp+kFzLtyWIQCz7OC5nULPckcrHOYmTX6R
ACk60DXouTC2Kmaib+jb5IAsxIZYwjWMM5plQFehAfosLKzbb17dAf4TBfycpLWKHekHAnnCSALs
SG5RLHEwjJ77gzX8qTQyvSgomVF4l4DkRyEIpCy3XnGBM4dMiXpSzg6XqQlgCSegpc8rcMFpW2St
+SUYiBHQnJE7MqqOymRr5pnUMu2RvpYHU6MJq7wpH8YXDW5/QAD5aAu1hdJ6lHwdFp4yTZao5nwg
vtPG3VbO3kMyH1j0bCCUzchbIqjhQB1JS1xYRyCgBPqoVabvnpZYgqK+eiK6yKSD4UTSXKD+ksGp
mQqQc+uF6S+QUuqy/Fr62HmomkcQ6beyQ86GxbWNuPjSP2ciruUuGD1qsNxsQavytGjQZ8WIGX9R
CTe2BSVH2uNo/Z3982pivrhcBwdxNuE/GJzCbgeLCDpHxKnUaoPijJDzo550zX95RhAEfE9TVmBY
NvKRsrlf/L5BsCKiTil3Db1e9LCLcXckG6CAlaj+Z2Bb5sb4SiJd0JmaM9oACVnjog6F2+oLegNy
7ORszT2HEQLMCSnIXxLc9/uIO/6cZ+cKoOyEWMh7UV5xWBp0Vr9k0JDOUh1y6DLJ3Bwp2IGNmnxk
og5Yvw1p0KrVHQ1gK9HqIpYEGZUctxVunT2thkq3dFAnHzKvQPoAQOBIWAmIvhAc9xsXcyGmPFUz
DIyG4IYK3JAnNnKJTvksn+wZbo2PD8VSRaWQcAwsgASnV6fQkBE4id44g9zbBZ+RVdqECQRHaB6H
CAB3L2XlUo22YClIoW/Zfl34/NYwVKE+NrXUHAFNnhXXTsv264IQAB1l/xKlP1l05XpJdK4DHRZ2
bRYkJpNdKqUpMaMvofq2F2Fmdh+AxxdDrnaHviuiCJqA1AQFUslutEGpQ5SXlOKaMzfzsjYDXnTt
L7LB0JFsN2ot56OGLenJ6CmNLciBPA163Gxxr1VxO0KombG+KWKunw0BBnrKkNPbDPxnBspkZgFc
XbRJLfMpM6IGQyftSOcJlUBuHpmk+A/Wwkzr9+Lf+KK3ZF1+q0kKUqxqOnir0YN3/NsKlCjtVaX5
7aXZe/lMoL/t2ami4e5GRqevUYH6uojkYnZ3pai3IUfo/WlCJ3OoncpWJiwrChN9xbiCDucHvSQi
HKUM4Ofu2JVttLeE/qcjNRhv68+XDPiYTSUqtoXreQSy9139xinuVc9jQzty7eGeSOY4uRTyYreE
N/M4wD88d5Rj2ihrZRETUWEF8L+qxZDHPBzbQxiAoPO1x3sJVJpl9vu8GNMzPOz7vBMmWXNm3Y9D
74YZcKdH3bRnogJoaPSYkXxHz4wamqrR3rdXZR/UKysCtGXw9xfHpQEeW2fPpPkkG59alhiClzIU
onKf2pRZX2hhw/CLy8dDO4mzJIZIYWiuA1SIrQ5B1D+nzYIhQdIuJeICruWVCBjRQEOAJE2Blagx
HN1/aFHCDoCHCSMHGk086EiC2pqhvHn6O6HFkWiAEk4YqjrolTEo2zCCYOu2lvY3eC1sLePDqDFJ
p/uZCIrkVqpICrXO8K5CxFdWLdOl7UadZqmfQfqLN4DyLCk2sHunf1YifcOHdu62xC3OGXMECL9P
hSXamQWj44r3gPb9PqbB0M2WVq1po+m1R5diQhD/UppZTBd6nXw08FisjvY3LYJtIuy2D/84qGPV
XqBIxVxxO4asOtQSHiVRdTCyNMcbWk/L8scKWu8CDhVEnzsEtcBGDJg9sZ7B+E4VxyB19ec3DE1o
0SJoWTdyHMpF1TpVEPr9GkCLs7TEE7dKNgbIRFAyrTbrmuogUi6vwL+NjyfH9ae88QLiZve81/I8
FwajxaX78IHoYPZBY38f3PLAiNPimDg6ySWO2DqHuL/Pa+athYCyPjExOkZMlxBHIOF2wnsvTTVp
E0+xgdG0dlZVxMqBAHnnupKuGcuEtPYOUl7pixPHhezi378/MtXqdlQr6nyBArp6tGxDfqQ78GYy
PDrps2aZmKJ2WplgTmlwYuxZTaGolm4qYNKSkFByhpFmqKvibmmxVXgKohJcRbaIzV66W4oKd3ek
UojTSmVWNw/EZ841oH21klYcDx5BvPkUHIdg5A4orczRfYqgClMlfly+L5J09s9Fn86dtiTy8VH6
4TDqrM9sG55ed09Lz4BaEC4pivWlAeUO1adN5Y9yWoiTodZN+KaXCsVuRl/mK/luauNzWOvGsfPC
+OddoMwE9eFnU0ktBMkUXlflvnGxLelx/20GkNIzjjXVfzol4U1xyt8bb5rBx491eYvnhNogcsWT
e4XMFF/zTRxUrtFWLXHmAV9MHHKXx+FLBC+SXTpZmTNYGIS0h18wS3FKNG8IDhOmfWGfEv+kwDp/
jykNmKbLsjc8vFzMX7U6IbJBhIT1XW2VTF8smt21b0C5aHG9eouRTz5T5wkILxgi+tYSlSnC4eWu
bfmAyIDkQt0SH/hOUdLeay3uVxM07m9hHkLMB9ArbvO4ZLoKZ+3Iiu63/ZiL1ECUcuwQEF+m4tt+
1cBAym1tz3vsNm21F1jWVXvKexR7FKCcYeRVXn2EkWm2Fj2YljLGEwR3ulT/AUkrG8JVJzypnFL/
IJQ7OTUfAVEUVAyxlTHz8kGmee6xKX4xLmhl9Blt12lWiOczPPPUvjUqc1pFlExHqYl40UuU3L5j
du1ZP5Ye9VFa50I1v7Sxda8A9RKGQoCtcyWgF2Jw1Y3zTIdo4zLuSBe5YlodUsfJl8/WsmFuWZR3
mbupPGURcluszpztD+Ta2p+8Glgmv0uVIy4h4vb/wMBwk++flJlEKhBsjbf2VIzqWV6iWZOncv/7
6xl+To00hfeTWjCwuN3QCx89U90dsusRqjTUrsMUakRPWi1JQJdVCJGsM2rtFVDdYh35ZOAkwHyh
iUh7AXaww4jadv2Tk9S4jB/cq44aDCIaX6p67B/+WgjRfnBFhUxEo1kCWIfU7Rr+lsWez+3kjeU7
rHOtlEsiFL45qemaYKjY/NG9OwTW12oCfgzqMGiwydGxFZq43mtJ21pZiJf9IG0/MS4JoWHTmvRL
L5RWE4mdOGsVTmgYkuqe48lDPU91XK+P0lR+O+ShqZE79qrPZcn+QTMQZ80Z3X5fdqlIknRFa246
jfmg5jYQx+vOTbz3ur+J5nv8qioxdPaFkxK3zsKnriREjtZvCSiEjqmfC42zFjVGT4uH6hYXJKSC
1Zx+JlBTBMvfi7gQRPU9m97HjwbMEvH126w206icDDwzD6tIHo6R5rdF3O12B7ZmlJF98dLsmK8O
WoS/nwtFmSCjEObDfIH2OB3wKLToz6apWSssxJOg8aoDZvNB2oC6iQknrEt3Y1FuixqNevUI6aTH
zgETLdFNNNB+fmygibfMy/e9vj+V5tVtPIPEyW19fnDKwDNMl3suFO3IIRC0Gt450A5dyBhTVaBD
6/2Jfg92TCHm+BkTS7SCBEqmi6BefaIqm0VagwnHOHlQ7tlQdItn6KosEoCHiQGE8eRil73Mmk2B
t65Ct1apw664R1L5rEjth3/s+VuKQEoDUcKdhBmri3TerFzDm9+oRqer1DxdhsATrWQgiBz9xPSC
dAvYVseeZUT5tw+UBFT0bYAyYR9LwO+fDUeV5yGcFS/ayaEGPHMvPV/Ad+LHViGS3D32wruv4+E/
VaPVk7OILyGgmyk0koGH9GsYrbBQxruQK6ct5wH6QXurlpschBR14bFkBtDB6iTEcEeMkmqGDEwN
nnqjvaT+279mZ8frSkuZStSneVCcgCWZR0UX8pe6urXhg464FgVR+zXe5p8rAaAcbScLSwLbPm8b
xU3oHJKay6wfWU1vXxmmym8wVEZE2Rs1yzheOjphlJh8h6eqw2bixm9pkwUV8wrKWl14Pdhxj/un
J0G1juhLCWq4JtOzTOjXImKHO6c6eOvXai0reJrPPFs7d71J1hoVoBq/iDl6j6cZRfUlvBEpgLDw
ITn1ZXXaEyPnMWZ9kRjFeWisn9iV8WdmNjoke6Aa6SrRX2YbHaGZRiecKCfHzvwEHMrSXot6sih+
NjKLVYsXfCKXt6wgET0K9X0wCKN8FffIcIlO0/WfVYJNKaUue1iIFDJAIMltfCwqA8/W+IY8LQeP
xuoUH3ArMtXgBMemzcsh1YC7BMf+5d1ykPIz0XWNrvc8l0e29VezCGXC+qSaHSVsxKjt5XQ4bCEa
oEcEfODnoeM5KmT6Kezg7KZQaMGi4MlYBXWaxGAj9xeq3q+DmgZMvl6o7v13XcUc2u488DA01Y2G
p0iCDqWcZDSnquHkFJvxX/T0BEfEIDrc7fJ/8pF11mIuKdyhmxa2XYdzKYARXIVQ55M5wSFbeuQZ
cj/8bDgUDr3WUcMeQR9BG+IL43rUBskCdLCDBeZWk0dsO63MTlko59G5yI1v9LH6lpWPqsHztaD3
y8C9zojGuY3meKCVZaRUNnCBKmE0xvVqpnO6NcSkPOhe5oCX6ozT0iNYUik+BnVt7eEy4nbrme2l
XhLKpvnfX91YyFBG2oFrfgf5Zibn4IN4RCaoxc/hrGuNsscmXMZecXwVaF2mZtktrTC1Kwjme+aL
Pq7SEDdYx6p6whizQWbeZqHlzJBlIG9QDMuunvTiqhXmBq44L/TqJgbqlJkGv14uRDczqFvs7/sQ
ZNglMMdwMgzipPmza+7VRCVu3/atBIAbtJ2pjEAFlFLEuoxns8BDf6W18g5HFDhIhs8Y9YCXFEgU
UrqHJD2LH56mN356+r4xOO5EZXsQOphVgpJDp47ru/lpKi1FmnLgt3rpElFff0+viSe3/dEb1HBg
6pvqv4vABPXFoHt7SUAJiTMwnkgqjuPhD1HnJSzk02GlN3wYvqLDhfquhQbIrs0vEoYBcyjQWWOb
e1degit/L70gMgCulQlyVM9T3BjWJUVzCZFo2PCicjCfIWvRSPFiGJHnk/F+9s7hVIkLGlQAkFhG
WzYiBKj3w7SkRUG58/3rY16WLhwJc/KJMGKKyzte53FTcoFRoQzbuan7pzA9bVgb/D2Sem/grF/R
Iw/GSqGN4Wzfy3nYQPFBw5fnLSDZTSARV4n8kdP0mvCbH5KLaKoNpK927FnCwIqcmr6rbVNvcIJc
vc70lwf0yQKjXpA1cZ3ZoWX8xlP3TotFpHZD082ONzsVnOZvIfVyIL8P7kHpBR7BMw0FM8PvtvJS
y2UYHuSHDGt2RaH2CjBRvZEvocsQuHGJRHVJjzWuax2VLDL95+FmgU2QP4aenl5bn8LoyaS49o1G
D/BI5xhVocNY1dVbmjjiapJ5jE87rHLoLaYmtoVPXgpJn0Kj/5+bpMK6d0QBuDmlKQ3eEWKT1nWM
9Ngsh5+3296pMxRWH6vzOKcSK2QzdDBD+LOxQmeROKJ59G9RPTBMHhORFEEex1Y69XUBT1xpxbL0
uxPywn/Zz/u0o2YLCtc3QOnONdCXqkyJR1zG8s13Tyhu4bBX4+Aj5/Oei1XGF1C2ZwNbe4Es5ZJO
W0FsDbOdRtwZmFl2+e+p8bIEC3sWTbJVZ0aBemg+AG0twHY51DGHWbPOUd0Kre2bgQ6G9C6TE9Q8
vxzJDRATXAadt5g7spolXYJsN9XuwKbKlzpVPg05H3z1JpMq02VDxM+sIC6enOCUhgmJ1fAkCXym
Cci/JMgs120+2z63TYgj0aLIMEn3ZbBDHcyT/eW4LlLURE1kzs+NjmM/CytqOaWs5N9LfoWgDuYB
B0lGZ31P5TOTe/7UcedQ66/sWIZgY93FyNCWIym5LZEZtlswT4hwMRNVgZmxiK3s3SmS7bUXGPHM
hcxPNvI60S3hPZQ88szIaYX52c6z9VpBkkQHBij7UZKNnIpQeinLrx5vRDe9G8mzbwREkO8BIl80
xUwIRt47mpFyKCz3PSdvYCDjOlnVMdY0ZobhI/kKG/gB2knPIZ934b0c0Hc8J2IAwYktdLKK/st3
WUBZImb/e92sSxu/5FvE8vNHofF4Rfs73kUHvLV/FiIkcE0LTvJ8ozJ5I693rqWzABzNCCE5aGcg
yX4steQtB6gVhoHstTLr11a4SlHGCOEXCcG7dfRzQqrvqSWj6WExgmtmTzC5QXUGgFMs2woTNQQZ
JR8hWr9poP3h3XwTyF/wddS8TDTnz3vsUA0uaKwvuvIvnHJlSmwq5R922sF6Y0ACjX2XhbOpR865
zcAkXWaislWheN1Wsx9BbOzb1mRV0MZ+ptMVXwp8sxRYmv8MNtR0Y4PR2j9jop7inXA1/X4nAR0L
LLtD4PS8wKrpCGuxjeR+eAK/BEFaj9SofmPAYUgFGcNKVVgai57Od7mPVmVIDRdDWpahQX57wxpW
w1zqBllCIOxN37sIlWCKdPebypDWInW3uH9cNm9d7D2aULd14TMXOxhr2zNxe9PKG80ZSyVL8duz
9ugbMFBHh4Nw+bCSA9HqoQlur2FWEGuIYKZdFKTeOFabS5cJhFYdQUMd+az3vF4ocq+dXRLM0huk
fNfuTBCd3wUK8nn95wxa8qwTiWZpCav88GBzN47GkVlAKuw+kBZngh7Y0qZwy2vMHcL+9Muy0yND
LgAEUvLLW8n8YYJ9ImornnxpQaG6Sf4iS/9+G3pU9pd+Rat7I5QkdlI1PfKtiZfDbDqmYtLGfPmb
BNieIfuBuMyndxic8GwiiT/H2OZQE4CpW1HX/p13gRe4BSAWGJlPqSy/DyS+EhxNSpKKAzvPxwbj
kCtM3D0o3Ty1lQisIksHzNQWpRltrz2gbWIU/ys+X+eBdLLraNs7CFnUnGxfjHsjAx0tySQMm/vV
fV48oktwal/Vc6al1e9xWh+CDcIfgCVx34pnTPTnZrI52lLbXkahpC++qf4npoZ0gwGQAQwDJK5g
WeNqBNVj7mJoi+emtf5aa8g7Nu3nDrYYcOUjfbkAgXOWBgn6fNENVWeWw4ATpa540+iXwMYVOOG6
x/Q7nyv8cC8rtvj/8jhIF5TsfXvG39wsea3OOxLEwd08nr1not6E3ZWUmLjHfK7pavdoBMbtmNhn
kE+73OGzGYS0f8FfwwCJ8F38lrjOC2qAEoBTPXTZvLK7xsbIOHBsKxWGpgusLfxO2Rcsx3v7mucH
BdQsH64xott8LFY/XbKltnLURTzoP1nJGLGzsaHJXJcff2iu9+4heBb/yMR5eLr2Gtlp7ps7hTee
yO6RUppCpecUVksAhAT9P4YfB+gUClJQRf5dwhvdH8isrG7NxMZsDVYnaV/E0KBlBMMi2zj5xjVJ
3pJC62o90Eq0EqAVQz6ZMi1mHecF6dxgEKaBKcwjZiOYmSaJtLmvj2NMDvTgenB2M2jKXx9WRDDf
AOppastEXs4bWIaPJmiuFTZudL7mr0SNIzLkTiRJV/RfEJItIrjmtmrw74ekJ8UFMgcKaKepdEbh
k1uqJt4v8SiLrb391TEt6jq2U/f8uA9zjjfkubCJ8QmgFKybzX9d7TgKH8p+Ez0jE9iDkNIB2GZZ
pRXq+95I/XDViLc2SBVAhGlFtE8A6gZQ/IWPhs1POvlrEG5v8JB8OHOHI5oVuZKJXkIY2zhVtknz
uuzX/J8i+xnLyHYPIeOC1sFtMvylivNEB0xDLdlv+Ut92UsIt7koNh9Ph6O1NPX8eKRXHvXDXs5g
aLRWCvgN2tkVGi8spej6SMJv1mJeu3A1hXVSOJgCQFlF9cfw/hdHhtGWgjADSxzVqMC+lLIOZQk3
WYMueMZOCwdyfVD5S14lmlBOOj1r40Bgl/J1f5iBPDrfgGd+Mgx8DMt6wAPDDDhopjnU77bmaJtF
EJ3kYxhasCpwgkTLe+9SPSSJPeHOnHqN3QqagoYXOBlH55ZGRuLh9CKJenKJvELHXm+sdTzmTO3i
03nxSCCVlp3KPpwn7/gwI39atLvpYpzpOlRKX4L2jk3olmxtM2fPvQQFgnYEgcNniiylO3mBVrQR
jjg49szTE3oIsaoqNYTveZxqxAw06GrlGwBJ7rEfHrIt+5w048fbWmfxG7+W5TixvUc2lL26+zDh
d36JoKz8imZHdGU7qqqdOBWDwEP0IlOH7F1F6ysHt5mkjzA2yTKlZ/rz8vy3bcDsp7qYzCajV1HE
R/NGF9DXMsyj2uMO5nz7xjJqRvzXfO656i4ZHN4wh/5ATITG4FwMf0y3c0FBFXIDgLKmFEiFKJRh
CXeAnpyKG41aAE1t+GcqKVwDw/2gbVk+vkQegEtR16Nos7biCMn0gClgWwnS1yessw2OFHI0+BLq
WScy40ouH//fFcLmJC9qoVmn42U33c0bnG9K/eCA7JTzVaAxZTF/p0H22C90f4xi62jOmkIeMPNn
I5vEvcMOmtnScN91DgZed8QC19rUpgyEV32WI8qMQzGgD/Pu02j7vaN579/PrzZhkyEEQjrmrYkc
+ghyeLtJsXyligst0kPktnJ5vTFB7G+hsvT4/KZz7pmrMIPsQRngT9eSgBSxpNzsg4tzhZx28BPS
JXyUPsln7CtId3pY1AUFCxxqMEzPUoUqLYUuXTkav82UgR3J1duxRhyh03M6o4Ys15QU+6+vvnpR
k9NHy21MIsodHeXDlulUP4jlOR59s4IRvI3FgS4sk4IKerBTO+Wof4QI/4FaWLIWY3ILccK7G+fY
N/qndJZ6i/Z1IuMZu/Vfy+1iW95Z0xccb0ThCJ8ahU/iD4ow7+6hIItHMjsQof/qXQzMSEGZ2jB/
MMLOnWhkvynolbZT5nwEqRLe6CsRCc8YPaNZh4AGi9z7paXg02tKp3G0lO/D6DwzRA/QXgCU2npQ
dXlgYZzkWbUsMIHQ03G4DvA9wwXbkxAyMBmnQnuJhOGtnL2kv25C4YAuGuK/L88rKCbYqqj9ACtL
GyMLHPmiT+81kycsecGoAGbaLaQhPQQSKso3dDo6isiWZVxE11Bw3Ny3B+RI8RdggVYlwY4DOK2w
+rLPilCWzpFhsHqPTgp5xMgFmEKuXiJMIG5lfBWSR9mVdYlr8JZqYczBah6IOI/6CoCmQctGE8C8
TN7QbzRW720r13VsgqW5mq6TlQ+3ivm69KRtS/iBFUfAES77Zul74Mmz3vT0/3DRF9x7a0g3tms4
Adr9CRCuGt9XpWruRx2NP0A9Xxge+vvUDYOa2FD0QPhMNTzfU96dMozsRR3Nxj2WDVleWsLVsbv8
3gaW6v3xqdSUlJixGXKYCwHJ7+nJvowqkqAOm+bOcf8cHAjNJM/kweYOh2V6a/Epd1e/VqyDEmm1
a21/SvIHfm/O47vLIEoG9YA27MExHHJh2Yj1yZJRLHOg/3NJijeXSndp8vOIbbkKyNJ1wGVNDPLB
arIx9hXo9vOimQAxxCO1OZ+v/VG6qhmfdKikqEc4b/05zfLYA+LSHN/p3jc0By/LDIJUgAT6T8hj
1E7BckjoTdw19yOQPbpjt5EjErGQ9YD4JVHa4dlQiGbFzHoJOowtjZvwhhUzXsMDcLYWR3PvCQoY
TQfwWa+KGEZu5hj3x6fXhfctE/Cfb9mv3UxO1YcAh8js4KAOjilQOTr+EoV3+xeMYdFJE9Jq7VSs
pI5doe4ePaR0WdkKlMTDJ26s7LnE0P2BGhA+29wIj1OfbbaMLSamuUaKEuZrg8qE0bF4gtEPVGtj
HmiM1HfJwL9LMvzeDTfq904UNyiC6A9kXelLwBzyZo54X4tvXoU0ATXwVzPhV4TR5SPsf1PIbweU
V5HUVHgI6/JGjI70fp/tqvm8sqAz8LxRt0/pXIOI9oK98ltRXtzavQeSI3gVpllEuZJy+lT6w0rk
uYMYgZs0fo/rEL6CtW5Ba+CXUlNYpL37z8z2iMhzpTAgfj2UBoWd1LJn/Ynomlq+ddmK2YM08lDX
PvxGvr6FT+6AtrKW0a3XK6NthZmMqYWjJyPi1i9nK9Umv32xI3PU/WHTIzwruxMpwOPyUc7RCFP4
mTXqrfbV4xc2GC+SHuobwlVDPVSL+uS+jliRlyf1OAkj+zijphAywI86j6J+rQmDidOJTtktpqaA
ordheGaPn/oNufStmGulwLWTPTLMSts0ZpH54QV8V+W0O6X1wNMuAlKk1zoHZ+e8yIn8BOIV6hF8
6YtysmFE6xBoEp1iDdEcSXAdUam9MCbF27APFTUEkmXpM51QklFh6H192v17276eh+HN9Mxm/H5y
5L6pg9Bq5kjvtE+Yzmt4lmciZ/P7bnjG2aVy7bl/GZVVdwpVivNbuJzcO/zyAfZxisRF7fqkYxp3
ERmItyMbT/0qpXX41MrxZboEJGvE22IKwW36lBs+1c98l3DApIANXIW4+h04yGg8RRJXXXB0AOXa
Jraz4LayqGmRER+1cNgoA6/Kh4PV7GI/DaioibrV8Yck9/7Nz5eG6l/Wd9PeOHD/NeDXXX+WNV0E
ZPsj+h27aprfQnSMDtArOGBfyUVrmRHWWjuJREKSw1r9AqIrSHhCxR9fwmRHVKC/P/m571p2Sqm9
FJp23eudI7NLYrLrjsvbTrRnmPNCiPozRSbe4Af05LplmuXaV61Pvg/vxXn2gPt7AGQEqA6ivu8J
2pfrsMesS9kk+EWhAHzVey7s8/CvllXSX+/l6mZZCSgW3Jm7/mTnFRTA40HXmLbGvznTPQGCotr0
vg94Tvx9uh+pXqLZhJoFDhKXFa8c6yJMcQkgPwcBKkBFqJHpkxQbXziO0I1ooensSgWidzPrmxc4
yFFDOAZkI6dO+Nqwr3vrrFIKOalaDHQTmwSwgDHGqJyulxiJmus8LAcpAlT3pbbDDLdTw/varIvu
wWH9oc6yEFKY6bQe09kcqsCVOTIgNa78ApFCago/ZoMyLsxl9n8MP7XUn/z1Xxz1OShjVKrh78wh
e74mK+mBTLAirxG/c6bBszkv1Bq1fAY8n2IVg+SKOmcmttD0zEKeEl9ORmMauSaslviUU5+nWWVM
qBnBSnfBV4Is+lgMqBMltdLnaABhSDf8d2ZBFblkKP0fTTBwT/mRVavt7VUM0EB7pCgdsQ205Ie+
JcNXZUyTni5brXimWcCey6bEQsFvRYwqwfC46XGXYzqvN3FgtEkXXDk38pBwKokW1wNGX6fp7kYA
oFq0bG6MMgYeOuoudFC0l9JfoZJlHKMYfyMRkAleA9BhW+p3m0kWgWBfzSNvificJnSqsLDKwupW
TQ01taVNcRcqvAnlXNflaUiXQ5f8qBWCebiOKOTRTxi9qyrxMgupHav/rkgT1cLrvj0v97/IZD58
uPBTTuB2G260KahLTL2smHOuZf4GMlkByvd+KaNRnEY5fppe8DPM+478bj2Uz61ITnm2XMvqiKXW
dh7bN8YhBjAcqLEmZgfssVyeOHWNusdChCC0aOMgnZDTX3n0YxOn98oPGpZfBRdrsmS6NxO2h/9W
uPaHeKt6upG+tYrvlkReHPEwxO3hEER65A9jJqT2J1/kbV0Qbp2GmbrzEyhyt/dXlb0RbdyT3f6o
vUkFKjSLcVZGGFXdHDufKWJxzCgFMRZcYqbG8WmWqicifp337vzVB2mC4mEcZAWFUOYeezIAf3FE
U0tWpHpXmwS83M1g3FdYrhgk2Q3zFMO1ZMYYBk7d73iZG2yWhEcazlRgsg+cgyP0feilZaYR89Zv
cL+5AyU28q8DE31h9t5dehnYeYJPjunc49Ka5SRXFCvlS26EkDqLrs4G6o86I9aFonBhx9dArivR
GRBnXlBR0rPD4cJKzz1rE4iDrunQzcMENl6oQBjlep54/Rai5m9SoQ9d0T8Gwc8jCmC0IvSlL+hF
vMpcMRCbre2cPBKQwHUCfxLdFu2GjUo9BhgH6aqABvLCVACJXBzhKaHoTwORvYNV2TPvdLPC45XB
leV7zO3/t8muDUpRrT8ivjYIfMLQunU8E/wAb25fgzbKnp9jzE/dRLdrFzcdauXE9BxBHPiH2HyR
u31L/bIXPJ/0dUwF3ptS03UNqd6kUMJkSWs1jcWJZwLxl8G0g5fS49VkzZk7Idgk/IdRbz/FAjf8
itmtupIajbaaeWp3YQq6oGHVgABFpxW9QGXnOmx9Qw88JG2n/axQrQsSFwLcTsPSvVDBw5N4Ebon
/P+1nfT3G1QWeCh05ue2rpWUCOUDvunm0Dglt/LriCD0hSP9pP+HKtjn/aCoqSie4cgyu8Tr5Ab5
jPeBbv5dqFYt/C88DH9Pv8FD3C2T9oZGIA9yeZemxCGPkzmdou8Oj0xtotmwQiTGE4vIsdX8GAgc
lf8E9BmfW4P/ZZ2nvyZB5+zj6Ls1NnrnZnNZjEeb81ssxB6b48rXmnC1DAbiNYyA/dtfgZvxYvgX
WSNSjT1xZ2C5rMoTqVDjgiYkBz+VVxKoStyoibPZ8KtKNsBfIlzPM0EQSL4AcaTxPJ9m2yawVqcm
l1k7i+JCMGDDt06V6c/u0bboLEjWWP1lCkVgAqh5N6QmoPhEzftBGJQRM5SMu6c2QFpyvVsfztBY
j3twdCXyKmEQINPIvz6m6Kxbw/EbP0Ne3Cquia7U1CcndfWcPDpj+jNn1pBOrRlV+AihvBLT9a/5
PwRsE4EdM6Tix3yBENi2cYSW12Rj2x8IJd1acGV2NBE2rmnhWNbECDQdiIeNL6IqzC69MmTRbY1Z
UA2PHvXSbYiDhNOYH5knGvRY6HbUDULZzXC+Rd0F8XlbWWqc/OImsLzosqXa0zilZ4b2wrjGyXeI
EF3+4foVRkYHFuhl5ZBlEpapnqIhjDG3BPlU7d0vh6IhRLLOcMhS1yuYM2cLMrK5l0IwjwD+3V8y
ovH8efwD5o3MciBGEa651PjEdfP/+4W46OQ3Arg00nyicykogeZO79oZzwSjp5YtjsfG5eQcmSnQ
J5VQtxLYcMR9iclyJJYZsLkKpDsKU0n3RiURhDmgG22WAYAdGUK2DVQF0ymmCuz4pknrkvsR6wjP
pXtSNVlwGRVBDc0G6PEa8A+tUItUrzsNzXVnu67JMOKWK1aREEiDvr59GrjDAswHfQSMJiUiJgTY
EE7dkD1uYL8gEJNmUMXDezPqPHxJCLXfxwFrwq/UuCRQbDA+AXusIN6FSQWbkzWUiVqW7t14iqtO
YDro0ayB3Sf5ILvYjPQQBluA7X7VRUGHf1fEs0zFjSCb+bYGsXIFoincoxYBcw1Vxtk3HQytYWd+
1gXdhGAQm063YdveqtdDP4a8JIwQ6BJOtQm3NyhcbyvHjOp2BSJgIdhDKRQdPtzOqrryzNsP7hfR
kcG/2iorTnNUjnA4o9A/syCCSpeXv06aCO4JqXxEBsq5oybLNgcfa+susEoMpzSrk1ct5z3QZkgK
C7xC6bvYI6WHs43H0AUYcIk4MfZYTmh7+XYV12HtZNVFypRapzN0jA+8JsXOU08wAT4047axeVBc
GnC7lk08fDh73f+jnp8LntEeX0yGhUjy1bsXjRPuZ9lScl+sUKIL3G8NCAQ5F8KYtKe4JLcWVE7V
ygsj1yJg7CdTnj+1pGPltm8p8yfoOZx93i4YN5ga70QTbq2NYIaEfhpBj3ZZzKctsH0y9zx53/YP
HNpnxMI0aUq/n0dW6Ovi7IrBAl0gH1qXxy5Fk25Uyrcg/f6sjA6mcs743hka4QJAeUexanFBkziD
ObZ2eTiLMJR7laPAb+bSHsvPjzroMbZ9Rb9WYRCeXjSIAVpdaFv2fnBwoO9zM2zG7SJjupKuw/85
+6EThh90xRC9gqelRtKYS0i+RFlmmbfdkA+1WOMj2gF+itR/a3QMqHbNA5M9cnSK8PlkrxnCM0s2
feAqhGZxHHTDHUVTSCxJci8d8U2O42g5tNMZpa2OoFWJuFGjjLAV2YZLAsmkeJpymR9bnZzHcUN0
o7V9PLRB2FXaJ5BZwrFt6GdU7bnJAZ3qGKuu3NM0nX0hg3o3o+6+z3KMRpfdvItVatcdlpRb1OcR
Gb00UDom245kGPx7IbNyBAdp21DAwrKln9EIfS+F4wpdDz2rpn2nNGFSQlNvWAWMoEFIlMJ6/9aN
iadxJR1SDC+kqLjwXV+CE+MHEzs7Kr9wGEMuDLxIGQ+lzs0fHvZ0Dav8Yv5/jP1JptW/poZa9HdR
AvNVhIUXo5NizLlvv7LFwTvhA0qK6RRVLo39An8VoTZqF/qMrfuvOUvzc3gz7JWCP+mI0N7/qGi6
THhYvzPRwxfXotao85cnHmcdTYr1yaMinWsQgTk25d+FSI52BQN8SyLxi6ubYkyWWNpiachQSfae
D5fxDncv+/CKlsBaRfOlp8/xIjBbD/49sC1UtHV4d0e9ke1CapvhsSKGq2WbVM3exPz608qY/2hz
IHgL5V7aZnF2Y4ePRP/ByJZRUABmaL8aG2yvN9nN6sfE8EWOWfAZIbhNovn5nkQvdXQ+ndiksuQR
gz5h0yVz6rQ4Xwh65L643WpYULWm13N0JnD3FETQnkTM6hPns1admmdcRLMf/DeCJaMKRTfdJ+Dj
dJuC9R0SYIb23w+LolLMrCJLavkcKCZebgctwS9OCi5bAl2ybYtZxuupTmlDuWO7xXQ4ISOqMTcM
ROqNNJFENTbT+GqBGBPSaj3/9UbIjjSzl/0uxBXnMOJrFp71MsbdG8VdfmBimbhBPhXMYQSts/M8
RDER+MBJpgx1k1JNVzSSgfW+bzffGNnDNCtvBW53lm8kTBpSdYC8hgh75DOJ4wcDYQs6KFEoh+vx
+WM3SNdhTTAET+5pMly0gQZYgrt/uKR/zR1NXBkeproa5gPoWPkeNaKjTAyFZccwFN6/jy6dMH/r
sykq/7wjJb8hBVryEzGEilofdwyOIPRtmXi7KG4WJo7/IicmZHdqqwTzLorba6O/d5YZ49IZ4Nbb
1qB45T8/qFff1+nOnI5Lh8gLEFlJQBrl8NbyTtqGw4BraAPsqOMm2Lgl6L5VoAfg1XkZOkAJMi+L
SLX+FiGTd5NAZC4Hms6iUT264cR4oYdX8001rAginHiHbR+nYkatx61BarQX3ZBBJ2g85H2ZTDGB
SkWKGUfFKjLzVb3WWRzgQZg65IAwXFg+r9jS+uiTvPKvMQyX2uvng3NMybzz4eRovOLAXuv2WyMv
onSiNW84G1a8zl/Av8rFL09HlrgtWSAlBlPBvZg5dOrg+Jrswg4iZ94pe5OkM+lbYsV3xRnPoDkQ
N9ZrVjAuCW/t/bpYB11S5YlDvZNtXY2+b/72xsbCGV3x2CYE0IUlceuK4af3U/qlpf02iCuA4WGw
f08NvcJOLNo7sH9ZtKdrlSmE0dYbMZvqOHqbAtlQ3mLy57P1OZYPhNIe7fQ+IiBhX1gKkJUViO9A
5OCgXcMrkRJ/r2qm0lzbQNDGNeR+3JLxv3zYKMXrRSPQt3TiwXjZCWBYbtiB/Wt8ZUJc6bFIv7QR
bBLsLikNZbXjxMwPo9z0DW00YiwohL7t8vVJAWEPPmsF68uodgWJFbQWaotEGGW3FvBsO6Vdi8Jf
qU8WF5OMS2uaRzzb9Wy58F0c0faeKF5Ub088UTb2RCfrNc5gs2BbCDADu7k+hTD/THuHX50DmIub
uRKc3a+zfuCcvRKnw2mCHTUhrKHgG0GA3IjFdjztMFd8mg/2qWoEhbVw8kvPmyo3mg5EBnZdBO8v
6AjuJLYbMwwW45qyLdTcW6SAPgjH7c8E1WiXHXu1hqLM3RbS3dpGSoStH7RuT8fU0GMpxqc+htCd
mMd2Aroe11cNpveEEsfTwwX0nND5DiS5lJHfTidek1wLnhBtG4yZYPC5+Zpc6t12aGVxbwvbt1jZ
ES/yhCx8PtI0gEpmibmYduDTH56XSmeqSMVQlXMVgusPQ4/ugaWJrmITJq1PRJS9Xg4aEkeue3pP
ILUi6kTUrBVjYXzh5/Q+7TE1ojiFzq6CFasUKwSjwHhXVkDGgJX3t0tH7/SyvJNAdbIkfnNwhSrF
vV902gRF4QrqLIiQaNCDIV8L1u25lj5E+qcP1eL++zZ4/3UwRQMwjDB3U54d4PBPR5ST8n4DHLlA
rrExVPMdV4KoRRxZ35/9eDe/e2MDtRgALDXxOdZW+y8POmsLa1DJE5Ex4lfgoLlb+aFwAC1GtFcv
itnF/i0M3+cJBRrzDSei7uZqXfk5Be8EXer8GzyEGjGRiG5b3k583kdw+n+VM0NHgTiB5eZ9p0nC
GLHCtUai3zBeg/j+kZ5Ee3BNWDVMc0qasNYCYQJ7V1vXslE+Diyg1hNz095TEqA6zAnoCt6cKbTD
vHyNn9nb939PTEriCL2vBMZ4y8T9hj2qu17SWw/AWcRcH35/Ko1vpdUYyOXinmYfu04EHvQOxy3r
qIB57Al/l7jbGLqjmZ70HRE29kDigZta+e5QxAK4cotMv9L1WxI2+EVK7h2j1XIPThKP9FpbG8r2
28F/BInpDF2AaDAE81cCqTw/eTpLY9ixVcUHvZ0rSe2UhiaEnOtyb6QT9EM2QUWfyppijT49wnz+
zURriClKzQLjW1TPX1vI2BeVAkGOeFS660x0njZi23AshX8DFiFVipAR8/AacFLfsHDG1jtwNrCJ
MGWhm3uD65J5MoSCx68U2Z8diQDT3DII2eFJA/50ycCJ7iyrGV1u5iPg1eCDksB8lGoatRYsv8r7
UqBfQ1jk8NEnhy+PFg2WIPGba0xouiOz9UD+c5x50H5+r7BAUH0oW2wmd5iM6rT4eo4XvwJE6MHh
wPchU3UDE6qwmCf0BrrGeERYIZwi65XrHcixVvRxkQcT7jYnmY99ht6Kg0s45A/Ivi4Wu3bUdaLG
zy4pzlwwL93USZfcG1Wc58DBbxZtRLr8yox8gkG2aCsH6GHmcm9Gz3ZqiB8YdNtbAurgY6yi2GvF
L3B8007WK20dFcUbekNHZXN9t9J0braPOpUgJ8x58iDTjJhbdSMa7Em7orOSpTHImOzG24kanqpB
YqGJp06ukFI2KLYewLdxxWtpG2pfrPDTi2XLlMYjiZPXoLcH+F1cXzdIR2eee6q8NpM0zIwWHtia
4Ek1z1nXP5wVuzWI4MLOJvB9c+iM8uXMgVXoFNOXn1t5f6oR0rRBnRVNou/o0lGOcXi+uOUs9ccJ
9UgUebXwK/m94qgxEwqRpuSK6Tawm0AkQZKhrSOLd9IMx+RbATIPOtjO0zO6VFRpE5oNp2fsbYGl
pLfSuCHirJbyQ26P7FYP32wY4slq7m4AvY93aJzakyau5sWDbhO/m6+WFte8aFnrbDwfTurWP7Sx
uKXbzt0ndJuygFuE/cKi1gClzGabnbqwcjC/OjPfFvRRkwQ0xxaQD2BDUZGNqr5IXHcjh2UXY/fU
orfEt1gYSDp1GS+XeP4CW8xCtooY7cjxqOYeD3GzOiNBau9NdUgsKl/VgmVoac5vFJQQb7yBeNsh
MOfuQ4Vbx5g3ArDYMXtTKKQ4o8jO/+PF/2pGwo6tL0OIbCxH8Ov3HWh0SltPf1x4ZRE5k15nwUQi
0849RvtwRbTGSwc/+GwQSQ0giEXdPi4PIuGBTIHWwmqZkLwC8W8ywswLc2EVV7N+nU2tDB04X3zp
gAN33quwfT4+nBfPguMLCYZLUoRSyiMa2IbLAWJjwwM2RXau5GGzQvU0wKg128o/LeNd1Hz6pfME
1R1UHPwHv7duDPasYfBSPnF5rHIfdSeRhTCSZ4nXCJSravPcUMbqyZrJWI39BX3L3apX77QFJTOb
mnkpqKfiNxhiy74Jp5upNSq0PTNS5QN1sSCAwhDHxLIhMSOTpsUHEPQluVKlknJiItPVT7hMa7TM
HRXXs2iOjVg59WXEEz04B5UMuljaq4aU+TU3bzBzL//fUl33VNBrOPjuVMMz94B9w72tqVpwwqHr
ljSqrZfaFp9Ig4WyhCDJm4hlkDvb18LS+VjA7MhuuXje/NQKDFkqXIAWPDebPZEwVsdg5Xa0pLJb
rca6H3gltRAArWHkqUA3AbZqFDl9ayW3lplXx0izmhWda128WWVcyxdkAltzCwBX4qkDgUYOYIDb
1uhLeqUWkwGbqwMmamaYXXczv0LFJyRBYOyuuYSTEAvrOiPJzCxrakHceOvsXOPi9xOTeRoAHLAu
YrzEkQXB/swSWtObdqTlsy0FbIevTiGPqL4KCKRPL6m5D24rdKrBlIgXlGHUxdLaR87/mjM5Zc69
U1NL2tCgusOOU91ywIsUT6ZmQdS/nKerAx4L3HqLm37mULfXMccDGCxtS2e1HqJgfTvneCEyWEh9
+ny91y7gBSg6lOcyVProvyxP19TNvyLDrSbm7xmk4oA0gI/6gqG4aS+dXpYY4K3+8mFQEQK7JdyV
flv/lBmZaep1AZS7ZXdP8BDUOwRD+sA/xAuZDGxxMqcM0OOX2vl/k2c8XsTwlkv8dHN6RwIia0nX
tzJqtHuO+O/uXlHqBfV5KhA/eKZKIhE4TKr9hgAgb/GyHyNUaLxUWFpyh4eCcmYcdvDZa8rObOJ3
X/2FnU4E+2X81rcCM0y4GN6mBiuPpp6C01QBVsLW7uoThUUCenGTWS9L6MXk7qmOBEOYWTxxUdKC
6DixaQpxrZzqxiyVSl3oxn3Hpw1w3n3z21C+Tl93tvFF4oGsWlKLyfbh/keZnenzuEgMV68xyo+B
qc53JpQB7sg96j/+u0FWu0poE6CXODHALXBgzV0t2fnp71/IxkxyGxdtAGrOavaETgQRc8DcnK2j
PrD0zQZwyveal77FhTsmMqyzkJ7bzXgUFHX+5OGaXUwLrSx3QQoSLCLlaDkWlZ0MZTCkOMtKaXUH
0q7MXzPDeOGkwNrtpA1SiwGUAm2kiTxr9Ufg9qqzsU7/2P2w6Y8iCxsZft3/X+pH2nmNZTvAG6pW
yTXkktP/U22jhtElYmkLRnMCt7OOi4E9xXj6C2TDUVce/ezS2a3t5FRh+BuryUNGNM4peK9jM+/E
oTUSu2Ssi01ksctjSLETQOO4jRtKFDmokdM4DPGYXrwf9/+wqlfAHjKUelHfY1aELcHFNNDEEhMV
kChyYGqgR5Y6bAkFkJFGB2MMZ4o99SRsejZ6SLTYFVjYCIxizmLtiwUxjE06w0uN5gqmZgG5vHkr
qdbOGgtlliEl5PUUl4ORY41xKlLgVlZZcPHD8zj1VO5ul/v/R1XZpAN2l+SqPG9nWAeNDaRWV+4c
uUHRIl11hmJivZessPZPNE+T/HofNipABOYOIgbI7ixnsPhVv7fXDAOrKafnLe0LEhqew532OK7U
2/VLvAao5OPOizoz6hQrRFQMX296rqaPpS47GXoEOAuqGPTeptUuIWo7AjP5splfJVOOnVi7mZl8
YBxq571pGRLlD6gkA8kD2HLSCCmjxWYVhrj1NEIrB3ewELv3yiXe5dFq9PPyH+ftvRILCUC1z0mW
VbsZ/j95+FWuLYUcWOQ7EKsZ0hn8fbmjq3Umpt/RKYNct5T2qLIjZVd+d9+6kr8JR0UxiaJwVTQy
r5lCBx2oi+DSizmU79qATxJvw16S8tkLeAGT33CxW+nu9VMuWp1MymyyjtfTs1iykGRWSTKXw2si
nYBJSTZeY95H8HkiZg67AbIfWoOUjv7pphzyozHniVFugJTHbacRp213ze4BDVrZvNjtI7gThZPj
W9FkO7zHrVqf1JKhcjtX/rxOpoBgjRgkNz1tZ0tRoQXmx3xc6rA2N91AITKM0oIb7zWF/vY2ekAy
yyks4bn5svfoBP8ddWo21pRuxi8u3w+11NzfdCZ+u6MYT+V/J5fk1mln1Itt/hlhPDUXL4p/ddtp
ktl5idv4BzUjVWiWPM31rzS2EsvX2IeVpZTq677+hauhCX49iVVQNkdShVibsIdLXXord4zgogkm
GvQkCW5vXlxwvlSNNzi6E5D2R2kYAyf6CeVpXAzA1VG40W54D+MLiPlbMRN7lkrwfwAHxVShH4rv
WVRVQKVJAp81SmudXuU8xgiwBw6fY9U8THKZj2Toj2Yu8vpAgz5RHP9sNzumuwuDn3gCR7p3PJj4
WZTpCVyanXy1MgirdHYbzw3YKTPjLkWBy2J4qhhkU2QFYr7UGgfQ6krNXsf+wFs9P0vEOAXtUQwe
mbj75Hd9FYjqMKa9bP4hl5zXtQlW96VHxBNsSGtn09lHYn6Zx4RnfYLzYOzWBxH34jJiylaSRFTr
t57etrGUmvF/TXvJOEHGzBs3lvFicU6LyC+/35wHK8ujjdq4K7NEGStErDhGSxAxPw2kymTAiofT
DW4tDTLcOF382kT+0lH+271hoZ+lRjwnxu9/r863PVmE6IX/OsL8n3q1/CWXEwsLUaSiQ3HCzI4W
ojpuC1Veu28QrOF6EMJuHLoKjbcersrfrX/SOgBy/2LJ71ZLjdISckECWiBVqKcPLSXFC7cB9/0X
Rh7sOIT/0t+SfqzsmX8csL+fx0AZBKE2PerkB8ZWEAChyz5gmdWO6oJeWCA5jMlrnGovTNRO1skk
9aCqrzNCNS+jZqePNNTPZTGdbelq+ZFjp5RWWSryZP/oAmuVNmfCgu0xNt8o87OrCkxm0NAHDnhI
+ytzkEpW8PonNl5Mn42PkRAua75Wqf9n1R3+ABiW/gCX+ZwuaYJue7/HVaR3uFcRa4CQYSF0UHUh
UFORIecnBumGjziVyhpLdx2z6z+bxujc7RPU32RLZGfdsDX2W/dwngeJxsIh8aohR4hLTeEZfpr8
OGrO17mv/2RHRn3HRDnWSMcxrp0F93iAyuGwpHrY3JxDq4sJ3+VbszkgfT+oHCyi7YqVOkeZGMoc
p60c0lgwMwq3jufhYVE0GVl5jwWS4BxvIvVCJBEe/ML2IMvsT903zSAHws1rvngASuCuzU7m760E
2jyQAGKWR82+rSmby0vFt7NplO05WA4vjkWOUZiROXYBijoDbBIyrMNEZhHTykyo4hpHRjPn9Eiu
OnplHZ+eyvkea/Mve/Y2UKdE4B3CpixlFUMFmoqm3H9s1AKhg7mq+m04mQxpauwAI3mGBTze8nxz
Gi8DKKRKgfSFNZtLQIe28G+trzNmYUU1SzyDJQBpIhu9Rlua/bJeTRDkBw+cEQVMprQ78zvqmJ/F
o03S+GVPBpxtsemGLoIp42itXsd6beZ/0TkQ10dwOYqbWTWb/MXPW++oRNvvnt7w7aiPAjVhw4/P
YwpejZy58XBBWbVrfTeH6GE84+CIqU6sZeOnCttRpUCsurOe/uU0b5nsAwWP1fzF71M6ZC94kING
B509nm9HonxkQnp3q5OnTId5JovTcpT88sBFNb2R+tbHSZG5Nw2MlRi6ylqm4cSM/Ks/BDN+JDWN
9j7c2lb9NruGlm4NuzXiUMOGr/Qj5dn9TwfrkzT84/3vpwo6AQzEFPHzF2eWF7fE+sRNYj/aygC6
lnIyckWea6n9Yq7gBKGhG7p83zmkNyIlY33rAmGw4pSO7XtdnSSYxw0n+YDoHVosaM7E06bb8qrN
2ADOZwaoTtNj8FBUcu69RZh3R1uhP8SPjiY/If/G02TxRUgLViSclP4XMeru+eI3Sye+rn4/DgQq
s2btaA6+WGvqxxpfqBEl+uQum4OMqFxYP2vM/zdskXZH1nCTPf65cm8smlIPGWzbzIINbW7o52yW
AvQL8aOQh/1mXmF2MoT6D3WWj7hocFCH6rXeAudf8L7ReMxEZ9/cH1i4XnAXLrodDppkoKV8k/+3
3aZxDL6IowGpXT331QUjsb8KW3p801zSLF3AiJohrJwptOxRXhhL4Bq619VaWJ2Cr9a0DaSez6Ax
RvrCWjHX3qF8/TR+AAfb7wPxrKITtt7sd/FPxxOISuiAgV3i7jYzxhnNKwxntmpLwMchCYi5Oxyr
M3wrkiBOiEeAW5JlBdHmPFcUHafQ9Ml3DG8FU+AUEcxLDTbgdsPqloK5uzVBRpWV0r1+7KCpTI2d
XG2c6+X00lW5+lpFcBNwgDF2cCLB9OsTA/WOCVDDvHNhNoW8y+wXOBQZHMT+j5KP1TTHA77cb/hs
7wr1w6z74FzqYeZB+YKwYGizpAEmCxOch6kpLEIuutjA/Jmcx1tnrNAYln6EpoGsoF+tGiW4N6Ga
geAciUU53Co2lE1w9dAOV2KNZHWKL2npAVEJt5LI/sGQnCyIYNCP2QHYKAaI5lmJZSbgrUZSkp2I
WfoGlxG1gCxgAS3Z8tTw2Ltlwwvlage9pKFwefvXv86gTNgT8aQbERwNHhM2w/qcrhYwxrfvssyG
bcjsohbiBcSqQQDQjAz9cIPagCU+UxVcmsgSlDdSIQZW12FE9BHeWlEHLhzttQNG41jUIdMC8ij/
bNJzOMsKQDbSUs6CM3RovyyREY0pvcKktEEHhXfRSUW9OycOKPg+pE1rWtJp1iXwbVBbQ1fz2NfV
m/M1ldqTGudb7qlrG0rInxXypV0FeVX/AvDBzxOcsd1fLM16uN3hXQEbrqALFem9xS1trFQKUc9O
S2j1MQjDLgvPqb0JXFjlfhcJwMXvJZxzG4MGgpNWMrAd2U/8kIM7Ctd5KhBGPMOUxn2HvFa4omvM
vBQoJRotqzaqZyfr61e3JZmW2dnXnKfqxkbFHXdfTNb90XCY/fog4wKUQ5Q/QlH6qdiVG3PTgRev
pLCMVjLDJ4KsTjrjyiBkEmWM2VoBgyyTgCbGzn2x8qbNCsM5j4zWQxEYNNT4A62gYP2wFcIttBi6
mWT7Hvmj1b0ZxK5u+k1takwe6m9Xo2faNVbr5rAbWQCKoVcABXew2QFIAbi3pV+x4vqdpTg7rzIU
PtgNGDKuV+3TKFc1RQijIZ4h2FDt5vPBwVYC/v6IG64t76+wwSCyDAbgSWKaKAan/i9jOtfGmisR
pR1Wk+OLZbkuU86L6o51wSehKANkKkpa4/IuFe/nWOryqSayqqlVodQbDsIwC1PyvsPD5uSQT9Es
2NuEhjUjMUQ404mQ+RQULCTJeqTsE5+lTgcsWTlbRarOizPX0XNxXKT6ULk7HYVPLDU2vja+Ayts
nH4YEsrk3ZxEub8sP+7yQuSY34TI6q071ibZJadSR1hel2KHDVYG7CfaA4+vSEQvQds8jBwNFpm2
XYIGMJol8J9CthEP2y5+mo7WBnCpUkYx6OJ2HEP5PnPyVm67IZ9zUwtcD1G+sG3JoeY2Mjj+jI2M
4DuHumWdgnTPEDk+Xyd6eLkPA5NVDB2pvRGMiXgrfxSblnCR+Ehmf6O3CAuG9B/IMI5WNmJ+pLuR
AfZNoDkDcOtFWu/Z2zND942F0FboQGxteMp0FseOJGgezoh3pP0FK+IoTohuofV6ZgYd9589zGXR
UaMUEO30To0eEF4gGuB1T7+UKMwoqim6FTh8PwzhKG7G3ymRDeVgGwGVyHuReo2tfCF1hMLWN5np
0GcSdIBlNQXJdHdh94YNyP2a6zgKy9nwi74V1nvlIe2HJA6mr5OOSRcRL+uG96N4fA4C1/atpMX3
Vi1KZ4UiMIvV36h61lrctypH7HP+NS/3OTcPsXBwkupmtfjmoTcUddpgBNGtNsnHQ5Jym+07xaTt
VpK4JPsYSIHJDm787M7BxzBq1TDq/Gwh/jCFq4q+CVM6UQeGxvyc35EExr12hQ8PyheOZ5CV/OiI
Keeb2ESZkeBBnOxupdO+ZT2rgAhT+V5F6mNzQuzC4wc9S4F7flmxJHhcVIYL3TApeERnhFEYK1h4
WyGrwM+naRGSgjhwQve6egTBN2P6/maRGetmWzxUrCp7UPGiK6467BLm9p5dN9A1YXxmE/gcuVMK
OqUyJRps7d/K9GGBbVjzXBhuzCMT6dT/u0mqWiVgnv/KVWwW7DSZu5tQ6uPLxEsPl/QWytCxqDaq
z8E7GWWtsTxEM6UQkpGdY1W9BCtnIj5SwNJEozcnzBHCR9DJu6/a8JPtgIZLOqTcnRzmfQDefHQr
PXwxq9KyJ70/XTg0hPODr13wDaboYA23r44ykOZBluwpGKY0B4S8IIUgATrWnsRxT3hG9QPCq9+N
8zbeWMZYrDBiXbSZF+3GoapWo9Vk0lG0eoVThLYozWLt3qmdWAQBeuDXOgSesdiRkLkE4gt1t6nI
4glNek7ByeegSdrxsESVcj5G1GtGo8rZsRrHGwkS5GSzTV1lDRWtV3BaJHP0SXaN7LNsetpC9+9d
/fMhpjmgD7jrqQ1l4ebqCATfwT6PH9j42wIr58eF3S2UD8CqaQ6aqb/STOqh6GdZwq8snT4Rt6Rx
kFOFRa5nJzzfPa66NVRKooW4Yh3bBBPiEgWp4icvc2D3VRR9WpUQ/YYPkWIPYmnKQRjUy4cSTuEe
7RJP9wpNcNOcvzkt4Lwm5WkI21QzMiICSzN0728dMhkC+b4Re28YGjT+gpVizMZvhH7OZTfgiPlY
v7+VqytvClMhRGgka+8hUoMxMMH50B/1TBK/cdfezlQjdMeM+/j/0KUKtGapU/IWHZVAkmMEqQ/e
+SOJfiUFRdVPuEDr2CFXkmQnbOcd2oJitmUApqIQfvQnluHyd8AWEKHwAhHINzGXaNuTmjiZ9K0B
aV1s5tHbRRZD+a7TTfp/9KDPrdFAD5VCp2x1vXywOBgq7zZBsGqqN4W+kXOo/QpKZR0f4eO170yZ
UyG8qKIwOkkoVWBTxujTPdAmU9cFokJRPI7rxVwURin/j0rbAVlHB6aRUmPgmHZ/FZSCZfcG4t8G
OmQkSARpv5IrOmYqFh9IZcQb6TM2cTra65E0opE3oXN+/O+LqU2EiKtcUx7iLL8lYhnFUlwuiIFn
XxDLOAD3CrbpmUkepZEBZAP/rLRiq5b9lBIOLyhn/xUJCfhUdHfkD+brpmBFEBioAd8RUIWtSjc6
ty2Vjq+SpiQcn+hH1SQohZloq3f4XL0EvOC32AKPiC9sfSG/PiOLxoBdw+n7DVxTtq4dkSrTEV7L
oV4T3EPkD6X2lLUANA2fiM+GuINbUSetAnaAcOTJ4nZux2y1HumtuRIdiqyOsQbDETNurict9cCS
X9P5IcsSiZt0yx0cYZsy/vJxR+VKCMGDBLlh/u2Jw0DMYNR/wWdZaaaUTppeCfkqOwlhvH0h6fh0
WGab6mBGHo7g40iqu4lBFeeYuKy1u6hvFzOYltvdnmo0EyZA4tE43iOkmlUBVwB/p8M40FXEu64j
y/vD19BLWJ0sedJWFpHSUY1XgoPdQWSlSdvZD+RQP3p5lhpSxEFf1Lk8AejvGbfC+0vWzMRC1kin
+Wf7NApA/Ua89dwC+Ig/9Rfj9sy82G7SPOPuxN/unTHhx08IH3+eAQsYqi2fzTr/2Z+05mXHK3/o
ce6JXG3soZpUPpq8loud18centubfTiiOgrx0jNEtTivoaRE8yxu7lmZGK/hB/arbCUtJKTlwB1I
GnIeNu/VFeKMv2DYS+1OyjydCY7nwq7VgVzySN6MTH9Hjh9BZm53apRzbczYx8EiHRT6vbBsxX9o
T8q+ISnzXWVz2nFqyhu/9rZuOCt34aR3iKbTa6hUjzOblVdNBLPPPDqzpTrDZd1A0fdXVhFl+Vo2
3fs33bOiosxCmyWQwzZZnICoDOGWkU+6UR5UFtq6l+bY09nT5SgbbKvH5k2r4Q/ZYwpT9Tm3P7dK
6/3DartjbY2m7TP260QgcOSAJyB7EIhRa0nupyfsc18iCmaqm3xmSDRZa3at4za/1Xem6BjFYd+/
SMtusRXSQ22JzuAlnNtlmuW11ASgd5VgUDuRBywCH73jV54bPZyDYCxgOIQGUcmL9khwZ+eCDtyX
L9dQdxfPoi17DhiLL1KN8LZX/L7MqvYTstCYxUhkbV11EJNCIHHSdPi+A0wGEXnGoMbE5w2gZn6o
ZVQAf7t36oU3F2oxGQvWj/cAWqnIs6Lzy03Wdz4QpbQ3EynEYewBtDvhCmOyxxpjaDXshIUQAo9k
qRK3S3UxpBR2Spov9GS8beCW3PeMIwGuF0BqpMtQo5B4MDAOoMMzzaoRscvPnLEZVIOd6ahAa+PJ
8O4+Ib7dU45VDPU+VoJVq2AzJFwpET/DC5TR0mymyTHK7G/WUTW6KisHr7wmTHchX01234qpLZhj
H8auTfevjTQ4X+VCTfSd/nSSLu2Trv6n8k1b/JCaPTDuh8pWaSzdFN8Cy82NPFjsuKyjCGaTlMpk
ztoiCnR7ThiiUVymmrTCVFzVOX8pAQ+S+bsTa6R+uDQpfxX/23f3VWCwSmAWyA4TnJCm+/AmZtN9
ZJLeZ/IsWYVzzv+AfhjNiaeylcr2Lf40BfjffRwer/UNpUXlYPLTaiWI0i2DUMOlJZn2itNvGDxv
kKO/o2oBx1PARscRsCLbaFU1QhknVJzEvqcG0kSqHFv27OvVe6SbZmTFwAouEhGsBMfqr0FGYP5g
t1FP1m53VqT7NoCO13h76zKciS5CQJ01J2ezILFN+SN1sOAj9L9JURmNr6SmaDDUwnn0EjKQktM7
PUNMwFqlpT9ClYltDc0q0oxu/crNx/SqpC02OAsLlJCPJeOwLxNp/9xGww7n54okjAH3fQVYtcD2
beEA04b3tlJia9Q4tbm51SJBKGKcsotwS9dyxNnxhokA3sjEqYSWJLDEbQYarhne92Wnr7zt+25U
w1D2U3yi0gb16toS1n9Ko9O8quJLknwEDdmZuCRg9oNM5KWelq8UbfUenB+cFaxDBjGtlrkzGLFQ
bOoH8A08njaZ3/+K5psHotUiBPq++KsYmvBnQlH6E25KcsI9aNCetdNbJrN7+q5OmwraUtqscccI
FRjpO5CywTstuDbv5SJJSxD63i2jaGlA+iuabCnr8DoEdvJJddnU5NwvgAwu2diy4a0oOA0auXcE
MB1H4uj80OxGvec7TjbvuMgFHNLcsDnaaTo8iUtFWKWx04AY75+oloHFUfrFCexxl/V79lWo3rwr
2l6EUjmJOUnTXcGKt57/y1tncbONi6RX1w72wcewil5oUzFXy+jBBcFjdBe7GMKNvs+U7Xq3ivAA
yBAUP8VVF+XxUR82cJoMkdexFfshb2ckUN5q9EXl3f7X+82L7aR5wn/njZr+EbuWfQyYwKArPtv4
d3ZX0Vke5ReWSoUm/HI/BWLv+ADmPU7CY2FD4ApIJub0hh8C0vMqHcIG4tqUga0F0aUsMsuj10yF
xxrNM9hgibHRlrRS1FyJLry+0bh6q+bflaQ/LNYQW+MLnVgDsu6tFUoTzseTMGqOG6GcClMZZYdN
VXKcjRb/aHtRoLNZoR9lXkNwfIUi0b+2gAwRAqtBjEhmjbEAuvl0oVWmJEDI0ED2ZIE0d6J3j6UD
ojd2NPSS2JOSBoMYc1+oxdZ7AW+UJdEFehnSYndFFa9YaM/bXMUjmAOrTPvmZ/AgCHAkzExCXdYl
dXJEKdJTOezNGIN/AscLUjSmq3G/ev/D7N+6pEF9o4bz/+upI6kj0bffh+cW/hpKGFVVfwP1DQHy
kJSiV6onBJW+FsFym3FZzoUp9bCxH/780iEGUsYzR/AALJd73peVj73GJpJubtUESmsmbvKAvJ1O
Di0fB06GDpztP4RDUCrEG4sOYgbluvzxaU3IpQNz1C3OJhU43NW4lJ52Mk0BbZb1ktn/Ewj1lls9
lXs+WCCuwHJugCdmwIlrBvdmwjVHy7QdHr02BLuYnowBe+snN9+mpVxYInYw5/XYoIfPk0P4ia12
7hUbyz7O1cjjBoBeSSeIYQzL/k1vBQ0Yh9Zdoua+8ltKIVNbxCbsvp0DPXjrhW5MQ3BWatDxldMT
DFi9YYOpFDANY8C2vOIaOSCcDGTvwFkBijfJqBkDrHLIoqFV461YxjkGIwt7Np+wjfEBt6nXh1+E
SjqfRooJ3durEPRKIT4mxk9eW/JNYXiyl3CEE+o8ZoPJgGoDTg3wXree0LyR5NonehGQuw9whSBO
zHOUeR2cj08o/gizWGQ6tYA8rUgpuODohjHdHCFk7ZqGB1MAYJTeYR3xErDd60j3cLy8+QgzgsLv
tvs1RfYxCf6jC7tbie7fsqMWzHw5YoxgEvkOAbtk7OharNstYxIT/vRTEsK4zW1xKRi6AdxsoOmN
M2mvDsbFxyDC0tn5uItFS7pPMiOb83+ybdW9FrZoG6eTglihu9czVP/b7if6XtdC4cmwUddqrhm/
It87gC/gP9CInSdlHFZGmEaxXSzu1KUKlJxbg7jDyVbBKhmaFwTcKep4oEX8gYbujjkfuW4JJA7L
SLYRnQgJrnX2kz32EMnMnioroxB/CgXbuLu9QHxgUYgysS9z/csG2V8V0FMAEB8w+h26GqKO/bgL
meC4o29XrFoV1eVJstrwbNj1f0TJXWxwiyiAa6zhktr2nkHlRFRa6ajbVP8lcWj/haEq5oekwG7f
2EZRFcKoLduOiyoZx3CCkagUSt6GBA2YYRm1s9n9wJE0I+ZRWX1IUp8cz4kh8kGm43OKQxwhZdkj
trE/E4I1ZbsklTJKtfHRyHDQX/dObb0qT37mZFqr06TRGcIJbxQDly93Yew/p0WF8XIGM2Jq9Yg5
LdgsRD+0BGAmFwskemajb2XDjAwFVl0ndSZZLLU3x3tIWnC2Z08bZsZTfl0Ya5ufvxJRsGSZdLmv
2Gd8iyyhID2XrHTTiW33nw+Cvrf/M/iut4jwlAHMLsN8/fTOWez0JrsJTQXgfWaz8rAOitbgWZfT
UMejZC9LhP94xH7u2kWJatpwEtSF1Z9CRd0FU/KnYFFHH6gcvy1zmgtgQRkv4+EVOT8wCmhK+bNr
pjOq0Q9JX96ovryT77vKXEBHCJn+IPrQ6RvPkr8AvYeiA6B6ly0S/SFng5IPUX9wQ0JgKJwap55x
ewJKv/+YJENUNd6DKL5/wLrgXj7CmkqXkVrvnjzB6kuIKHHAkQs6hONfDekJyoWgaOHdAKXlqC+g
+a8Yi3sRvF+K/iztpOjbxSpG+XXuCbYZyQZntAhE5kPqKMeJdJqnkd3hou/6+d0Kjk1crQcJwfls
+dWra9CtW5RIpMBtupGihxKf+ZC87pg7a33KzW3jMdiNhIRZOPWl9lVG7hXUCGC49DAx/Jbro/6P
dOl6lEhT9Mx/Ns5ieY/fOzuIhVSfD9xbaYez6WFkqLX3IfpO4pmkZ0vVDk8y3qUhvvcOTLmhzoSR
PYA7iQ7Y+CN053uIN8TO/UGuYmESzo7o/wsAt2zveImDuuAeRmuxr0JOS3kq1efSqgwFrtKGAYV5
F60zIv46+LGtB4ZOmqY83GuwnccVjts4uvtpUo6q9HDbKBCTiCkR9/oSyB3ME9wOalER+bRT3lho
0AF5Y7M2qsvZgh+39l9vTdu7Nf3Iwq14uNGqoYsnqc0z72XpCuYz5rGp58qLwceNbgizAkxgI5R6
a9Q4y8YAS+S4usn9w401/fPtHMjD9Kg1lADQwSRSNCgZTYl+NYemjKseVTt950IHOednoTRUwxT6
4IAX1qeY6K4bol9Z5aWYRRBUSEczkEmUJNfhgPC40LGYfhGr2WIkMq4NIg8l3FN7s/ZoETn2xaZE
+pLtE2N3hkJAxqOr0OOpzd11WSXctx+M0S7SsCKPoiCyT55kCMK/UbsscVXULURd8Mip72tzq+z1
fPtZyhfW0zVmLz2wrc509mEaXfNLLG70tuOfsls5cIYWp4y1pqWzD9BCmX+RCyfwOMZIPD26PdIV
FidMYSWfcuP39Qi/6KRwOO2JRyB+ZgQBjscqqbQJOWKtZKEwMMQomdO7/d86eEFd9qD2m9MTyzY0
TPsIkVUVejuhRvuyntGPGBTv8QSEly0wxmrLQOYJDuES2vx4QEWg3ZkC35wMuOVob5HijeBmLfz2
rysXfp0oK+5Gfz3qERiaLavGI39jDBD8cSqTETPi5MjP2MnIvwXjotDZhaLJMO6kgnkZd3TMa972
Mo9IuTznpIcUENt6iyOb6MvDlQIJlX5ptWthBz9ZmVS8Q8ShpvCOT9vqyK/TZBJEJGRtOpyK5ngt
Gy4wUcL3Lb6D/bOhzC+ic2h3fpffkvZoY0rqNP/4w2u6J2m7xRSVWFdgdka9nhJe2Uo32TCgCX5f
mG2hCkBbK/bcex4QQcPtNQCJdpGN527GLCPkUkCXQMhq1ttP1mnX7qouclu3r+h4wD2a53u/AXRs
0xZ2B1uD2vM1oWR2ualXhXlcdFUchs+ycnATu1NNySuWeB/WUwEEQTSPZukfKUkrSJmIgRSDpkhb
MbpkR+JHwhl9RZ6kpSPMlYjfrs62tVGGxj5siJtOT2nDBjpNi8iEnafCsJgupuN9mNoAKydTADJz
3BZ+dzsO5TWG8zRNlVxDI4fMEYaO8rCycGsIz2pOOsImVY3GD02NJJyE43Zk8tRfUcvpZlkNQ4nb
OKCrMUiN38IW89sSALjqwSvf8LxTrnrgYeozx83uptNFrXcrU6JbRQv+H9dPF4l11oObpjrB0PmU
0GZMpxj+hUKaHKkf2sWe46JSOabfOBrc/RGeWSBIiBVWoAbOFwesNgNuzhwrSkWMPKqllwpyUcPV
EI2KpQcp4mRdRhHq+arOLHb0KG/iua8jWKUsci3mlQZck0wafNCChAuQOcej/Z66a221pSiidI0R
4b8OJj82HJzT4QQcFfqbVTelZllBm2hz+W7gNd26s6HgDRX7tNBrqcTj8mCH0gcZA1YFjIQaIORH
HtFpZ0PywpQVlC/W+nmypeV7aKSFcz3D8oM2E34r6LFjBTZ4SIZLXeEOOriqDNxgCifIxMQDJ0CM
7QcZXhY6x7/h+zNlu82cOirzkC0vJgSlhOWlhY2MgGDbObAyvb4e+urDbMEHMfFbTlLB81vduLsk
uHEhp8tK/mfIos7E1y4YXnpDU1f3WNVDKozIPCCbIpV81LaX6h3tx4JolmFOi38R4LezCQHf4QF0
oVW86vgLVX7L0g8J2ALJB6eFgdtgsdg3SJYDJUpUvo9SapifQr0DIaQIJGuXnCQAl0O3EA7eDjPx
7Dc79TZtI45+/SMhMPwUgpnsVCNGxsnYON8K6RqG/KPrf+vWa+xnEOxRpNokIIoQ5zDIDoJxmm1l
cmIFHPd8FDYMH9fGjdniimdUm0ZGBSKVEQZUylY608TajAiCWRTV4DqsSlqTNtJlAI5QWENIfzZC
i32ba+OwivB24z7TD4KH13SYi6yODjSvMTocv3UnF5xpkwMv55cgSt/d41RVzCFH2SHvinzPMpL3
mBJUk14PHFECeUp4KbyTrlM9gBd3ke90lttn3lU4iHK44TJMbkgLR3yBHo/0kssm6buYgj5j/1fU
bcmKxNoGdJ+wCidAm0wTG907qdn4UdDIHFjnQpVuUSjgofqRKDgcTHwcHv+K34+D5iSrzEfGAUHz
Um/0oATAthTrASFhBpquOnn6VunIoUL7EIl5GfbkJNyQaHps4c8lu4/1EhILrEIdWnWculbUgL7w
w4SLDiL1uaS/aSkpdN1U6g9HVVAnZb+zYTSfOptT2Bz3439D+cyaoK9n6erF+gDo/OBebfjeTmqb
wO4vF10J+KuVlVa1eC9XH1B1wb5j+DmL2GThhZET9rk8STfOnvGQ8+WXNBkVM2mjBBMGll009FHq
xwcaxZabgfLDo711opiq4ZgFLrk1TvnNMuNngTgzX2vKZETV6m5uAP9JkZK+69Ca8rfGrS87ViH7
VBuNh8kRu8GFV5oXDNg84mDB5Ilf1LutKT/BMAaF9SPE482Owr86RcvO0ARIucAD9+apyEtPnlTy
DBIJpIbT/I6PpTbbWAPJin/is8buzH42YNlS1WPwjkcIQt3/C1KEsSdSB5VDuAO4OVHTuYvUmY4i
JdCQb3piDTrzavEReFTAWCnYeZZZOLAE+UE++oeFFGHldgSM3OrimwWTcKgCqhdFuSfxeVXnWr9W
Y1QRJ+R6SMJHEsjN/L9ih3R++vGN/hpOHof7HNYmJ7axxR3qsd8lwWJl5c8eNPAGyQDtFV0/egqO
QwjJ2jc/M82XL7zIRs/ZfoQMM/o7OLi/M52jyGt0qNSK0BmAkNW9ADQxMIw8J2WqkOds65S4OkEl
TOp4aTNW0oRIjjeCcf+aWGXst90T4gd/+bFysdAMVnXtiXc9wFSGaVRVyn2eqeI6LeHwTqx5WW5F
MRcsJOaY8iADzxULCLaWMJfLw6tQklfcIO9dWzx1w0vXjnDLfShZF49VxlzwiL7GOPx3i3IS88+b
mMkAKcKgnqZav/f5ONjRAIxJm/3ByJIxp0R/2A7ucBTnAWSGn6ICTBTto5+xmre97pCS+FulJdn6
t79j4gsU5cDFDqKOWhpgdRYZuvYFrbCjtnANhwdmfbLZXdMv4lExyfZHJSpXViB98gWMVktiKEbl
iPxcSuMHC4xBU7tHk5BaW7xW+H90ltyaWx2sRy/18g6VCdzcoMAZXIb0JdLzSo0=
`protect end_protected
