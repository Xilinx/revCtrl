`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9072)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/Y3
LeD+qw2K3LM++tksXDWlRgF/znF+Jw9c2JQAPXKM9TKRvOl/czmCOhE3aNSoCh1FUwlKG7QK7XW5
1i+Y/6fuS/CW01hotPrez34/+2hYr87se6GBDorysLqVAXMsLY/YV9B7HhDUSw8jyNyknIEmI3U7
WudHo8vhLWlCkMQkDcMf+Ivoy8TEGZRjbwDtOXoE24Tpyh0y7Szqp8vQqEDariMqKoVn6oTmJYLq
2DpWhIEswln6tRI/+zBSleCqwfAdmXyYA/Icw782kOJqC1rm3rVrW/fPVK8K9QJVLjxlLtCOUsdW
MXHfW8zBcf+OJ6M5Ps5WfxcGaSo9F93JhZJwtp16qQc943Z5uL5S7F6uhx2/2/JNEiZKR4nwO6YF
9lApKneiqiV4lMknv2GfPf3Z0yt/epCJ1D6rwzHUxOS1WE+QGHCe4rtK8iJJPU8gdqWBAV0E38zX
DrRSC8OcTDpaHRsM4h45UtUZ7QHuncOnjyjfle45UXlGJHuJmqtQtKoBHlkWLaWs8IxPTRJdashu
kUk0S37b7qinz8QPzVNDizIo7tt1mrqBCLYTAlFjqwSpg+Q2GoQNpEbhhjJSmvYKPuGddRJZO7Wl
OSphxyLgZzVvmxDSH/t87kHgGHsFgjp9dviohojl/U/zWNmgRey6ALjcz02ZkQE6vzh/zBsU36oI
1XLzZdPOsmsFTW+hi0YtW4QXrws+XJn0lDvqAm7a/4zSUan/YXPqgWJAp0UJnu6AAEQbDjLTTbka
rmLtzTc+KBM7Qh/MrR0nLXOt+vB6+4vpyFW6VF57FxmXcsdwTMv34b7IGNAHXV19xTd61xcwO0FS
hYiDkPuuZYyI4HEIp4JXLUgW5zvyHVNvmOFASRRNUBRiTkDYHnHp7Z/O4tBKX1n17fF6v/fg3mwS
2JeiK4If3PXvktkxXJaPGyiZmPmt5A4Bthy7HLbet//JHNLV38xyJ74gKq7QU9oEASiPXGEAhbM/
x9I7SkQ7MIJFc8uqyxac3MnFNurIiDEeYdHyaMERPao3PN6xhb/2oFOdOfTFP1ukLGNEUsk0hPd1
LgkUtfW5A20Gbm2UqEhuCsZlhhN713pRuj/0GuH8RmIBQvAjd/LXyOWfuP01wImCTKOjz7332xEc
vYTB2ZLyx0dZNiESt3YthzquQ30BRv2JZ/yMS2L3RICN8EY6volLZIQ9J/ZWNZnto43SN9PZ1A4d
KcVhHcitoNxEjWlorIlUHZeWcgjrKzRKTms/5Qvq+XK9VFq4xnGh7Oac9iup4UOYCOq/mhqKA4j2
JlpoYNdiV2q/qk1GYiR9lF2o5Ecimhm4F6Qr/f/9tQ8wUUD6qfkiHSEpOGq0Z+43W/6hQ3pmdtRH
CP6CKYahbYpyAC5P664kR3KSyU3BSn/mcTnKBa/6NWGyfV/dwudwQZYVTSGWPphViyNhg4NXBZdW
VpNjfiNyjHV/WD/NL12VW2Cc1vUJznM7Ohc7WOPoxL3rTVqMbdkgPi1PL7rVXfy3t8gZU9LEOkRW
PzJtI3ekd0GtH6hpTLnCd4KmXpUwUPsqehrqFsbkKH7YNuki4EFBpsExEHrPqDWOzpH/kcA6Kdrc
YH3a3yqe7rPGOTbbq8kMXtkWN+YItZVlgy9BxRaEYkXkPwPE5k9IeceOrVP1c98Iv+echFZLGGt9
j0QBJm/V8zqFl/WSHqF+eE2suXsp689eqNMH9JYhg2llYDoxhhS7WHFNPfDyoEWMj1/FlOG8ECsl
8hbPn81Rxh9ZGPDmnWU1rLYxp70uYzLoDW9knjjlU7YCZd0swAJvYRhXsXf3VpO1kz3iv6W+nZMX
Brg1+/LfOSXBphl/YIzzMLzLBGrPVYuVX6U60QduJlfeyJj/jsupLa0YCq10Y7+A2WSQXESFHfnp
Oo1bNau5NhQE2DlB0tGBKT9+EPIslfIrUiX61m6Dkfx7lrqNHGsqror8LWJv4D6YsANdMsKop3y8
ywyUOABWxCDeC4c0Mvj7ZXbQ7mSXzmcBcrunwbWP74A7PloqWvI7iteJV7lKc7ctjR9u2w96DihV
W/DwvdUVHlOVlxCx01PJRop9W1LKbTZpY/0ZzTe7UocPsy/89bc9AcwM4aV8BP8oa3Tq0MJrZOMO
mP8yNtdJbBItrltMSYPKOFrGF8h5Z9v2p0WPw/sstYnkE2z48Rw+6hSemnVMd0wzek9T/E1AS1oE
ZrA3f8QL4jIonmJyBqQNSc2KVR9ezwV6djyk6MGEmqbDiHCADFai9EZ365ggEep82nSHyOwH7e7k
WAk5TUhv+Z/kHNdp52dLfVakxOtEHSbneCdm8hkeGJ7HytHDkfG0EsgZqwM5A1W/2scrmPjhfeMq
Z5gZil+FLHuqDgpnlqk6GwlHJoOLR6TnOa32UQ4VybJP9TMmBagp/su2C8/eaMBKHBuRVk39v7FX
8dhO0ZLg26Y43Dp/r3gPiA1p/bUv+HokNtQflnLHrnfgcNwAFuo4ChGQr1suF+/6MEZ39+YYcLQX
aZIHry63MB6k2POVKN1jUp6i5HvsZkxmE+SYqfeSDdTzqzoy3kdlF3NsS9UON2EiPWysa2Qu1opo
tMApEFghS37Yp1yaPg80jFeZRC2laiYChE9ZVjVUsteBxyUf277ypkGtcghPr72TPqQ1zQtbODEV
01nBZ4KzeBhaYwC0n8+Xh271Ug+NcvgaVLmitcZexDBHRfooei8SXKptlrX0Oj+5f74mAi29Jmga
Yl+J4Ze7y68N+bzIJgr5GmTFfbhcQWOQtM+BOeiDagj3eW0qeSPaLziyW5Otu/hbEIob2UQETk1p
onrFt1MwZK1hw3fcZGOjClWT219Jhfuyy3lsb9z/1Y0t7kkhyoXH0NKDKRuDurkJ0bKhY+0GCyGQ
H38L1GYASu7gN5ku/Zk7VkFeHIldz1l6oisOIKm7UGg0hicb5B93f2Pf12QemWqxMQgJ63mSrLMV
boU5NveNGoLsYDtDnaV2YNF+CNcyA/sJMBZrLAgN/9Y9uAUXs3U4HPLd5x0+voXUhAbX4JvYJBIt
lCVF1LiQZRVoZ0CoPFcTPy0oqZf5t/B0waoz6o3QOXzVHLjS+SJmInj4IqzXOmBxM6t77U7imk18
bLYCgkajPq5Q2BsG42RmIsu+QPpn0N4hg+BdsyTRZhPEP6EAVaqRoVBNIdfJ8gn+tTTv+OCdZ0fP
wJmNdiPolTNcs6vK9TbANpZeWuI7a6qtgKNBsOCOdc0zhjb/RF52S1BKEBqc42VuGhh6X5yU2mGb
ruL1Fd0poo8hfojdBetT9uzutJqvFkx+1xuUUrZIfuYOY3VMlY5n6iS6tCuK8VerRYRMRQ1w3ZNW
TjZmBq0MOs3B64bLdjcA+Cb5wKYCtVDrfS1jPXCYnY11vEYxa0lbOLvnd2vLtQkTwluYDygDt8eR
Vy7ZGhDBf2KaHmfrIu3ziboSQ5DFEaJ/98YCNZiiNFKkMhf7LI4MzhlYsZmfTO1rnyW2+tHTEJNb
Vm1wWgpcmdwKzr0Rhxk2U5N9VipQYIGLz3fFUPlkJLMay5qlE9EXxZm/kzHYu3OMPoUDf48zkJP0
4xFWXJ6SQ39+KeuRog5MN4xa7uxbbXarZf1M9+aT6CRIcVU8gQl7QL+b6GLf30nSN1afBHvn2ElA
yfIB8krcFI4oFtsvj6kwEd/5eC3Sdn+Iqe3wxumUc9BXCEWjITfrpla4uxtbBiTUWFatdfSqt7lA
uf9zUtEqJWCahpPEqJC//ghyQvyDGJvjgLnpdpngoG3BC2eE8rVJF0fXWzwojQlwvp6tVUVdFJ1P
jwlTtMKHaHZ490u7qik6XHGn1wtx/qgL1lU64nZ/CM7q5Bk3tqZrRcmljXruHkQfujV/a0xziFg7
wiYc+NJMMTV8YqDPyYP/7ZaPLwY8jxyqUKv/dxLuUlkhpPgEpQZCTURVcN8Pu+iCP252vAvejez+
0D54NWttijiwEZAtZkz7SkLxBttHCRIMFv0nZPTBYumQ7QhjbmeKQe4sU8rcfhawHm/ONLnz/zlO
OseQRJ4XfVzj8Rut1CbMB19r65UwOSWKn8GSvbeCSiJIcQKX2SYsCiUmzqS6YuVPnzK9n+u3jUD1
o55n6QuiZ4uSs92oPGJ7cBErGi87lsMjdauFQVrS7nh/BXmP2rvn6AYsdvO8V+mPSAlURqCQl89p
S+xvhZ4zxMRuRWUx7/49ru07VmOLMvoVCl4hoEY0m1kzB1/P03PDM8evS1hgRki96dTEDnFXQ34/
l5Qwpup8tIfPVpKgQcfiZ1JafZIYkd9logsqA6hwUdEkVnrceyDFM+Qk/TIuqlwHvN64EaCCrnne
Fis2w70NBUBswkbBgdjENmlCqoxfbGRIok4K1LaE/eKXbu24EeBeHKedKNH7dbX53EaraJX0hGXs
JojOIb2c0gE9If99xZuDuPKaCTy8lE/a/X+UEkGosFvgxMNrNZEDkmKw7anEOlyeyKC9fRb8JMkL
vLAUcbCj5IuWfsfb19l/pVGTuTYOpAPfrUbs8VwzoUWKrnPaFETqUBlB009rML9lIXpr6kDpTc0+
UFTMLScIoV7jzwQIddZx/MzfzP8c5k1jIzosShmZu4oWZi3CVYsjsGJPSQZL0SAd0b2vjRKQFEet
FFH0H3iIfOUP81qzj5IR2yIMg8l6sQCMsBRvXYWI/IuHvhJ4uWVeyIgxbjkA+OJQVbqUcMjzMW91
l2CJszv4SwX79jmfAts0RllrNdLUE7xCxeqF9kpKJqUuiZYljpII+ij5YH+Bd96TzpT8oIhzE+a8
XTznyiHLfm1Oc0YqQapF0OkUtnav/4keouXavyasCU50GzzwoVNngUCB9hBTtU/JePqap/Dqi1AF
5eb737mEfatCuPuXvVFgyOsjf0nE8ZDzvsrJb3q69Fq7rpZvt1kUfYjM8SAm9n6xkSb+TgkBqsSd
YEU41DSanAlix89p+HhEm4grzKvjBeFE6WILmV1d1vL1B+XGB7HkBtJ7DjHG9xdaSopg0fcRf/zI
7ly+nWt3I7qGaAwgTmukBhMGmszFbBdWxweS/jt5tUkwDQGDJTvUsjGRTjU3R5umiAhqAKxUZ2wP
FaKNC5RN0YmfEKghzXCmaBcb2WEZfsfaIRrpV/XPs+scWPjuZ1c0f/CZTdeNFWxJgRz2sufcZjs/
i1FOcHmYrlzR6B0JkeEtx2g07fMtPNUU9hv7qfFCVkAEa0CtUl9QvzQLKWoi29qaaUc4jxQ2X0sj
UDj/GrW2XrZQum+gCFmJTquvtgyt/cgPGbIVRSMmK0KZbmr/B+YIzsuwoXKsYOVCWFi8TmXsyGnq
oMOtTAH1v6o2TQJxhbOCRLGNSmJtfKrywd2yXrgfq9UesFCuufiHH0D2Ootd3LILtfoN4h7iaxoG
2tXQE3qrnTymUUJTOF89CoDRBMG3RkR/DCl6OHdHJSuzIyr5EFA0WSkmvThVQZ8u2OFCW9GCdwqJ
eagtyyYN3XP4eH93R10px8H1gH6MPsGkmDNku1qvMj6xvVD4hMPcY5yYkvm0N7EBTBCBdqLCpLaV
So/eHDxbV0uh9PUFz0mjG2ZPJkaJoECBZ9tA0phVDdL+O3fnE/yACE7HH1zXxFXOmoYFxKGcrNU2
8eqUYKVX3s8aO09iGMsGLjc1CE+R7+RxLNDV3KbIOYzhqkFyp9TcMySHbpyDUkPoxbSNjuc6fQYK
OtWtyIEqQrk2NXD1TCZNKkQkJOfAbA1ONzfd6OGMQIUk+iY+pdTn7ry68w/pyqHU+YyYJM2YeBPD
yl8W6cpyrb6mDY5s+6m8DSUGmrHyn2G1MIfMZ8e/J/jamXhbBO27zI//qenu3QfXCYcHHwoQasco
caMpHG+woF16Ac8CR5RnV9ZWGYQrmQ5/4enaPN6iPBjBNf21HcEa5QcCXiReawrQ12cldpRt2ZcL
FSePlGIbkpxq4hEloldBn9ovWjLFpYrCzZAU91ihvEcL+6Wos7Q65oDg7hER/fd2LJ4Snco4jFkO
ZJBaVdiR1wpefESAwS0R1N04+1CCbDS0tHrPkLVBQbLenyaOs/4SMj11RvHznTnSV0cFfNsd4FNK
/7/Jnh5CJy86+/KgjhjiJFsMV1eKSOjLm6wKDnPzGpGHWaDkQk5bdaUKimWmmu24Z9mh/GmLQXMc
oToxN7aWnDaPgRWLmRiVhq8CFhjHJUmoy02vzc8IVeRHwkf6kshAyf+kzPj734SUftDQvh1ZHSkm
gi4gi9TW5349WpmMpIfnSYm0DAUz7TAF18i21JXg+OmreQSQcMTcyYOOQNt4Z8eMn2nebw3wl3S/
FSPrHVhQrPIIOudXta/9zkUH1cPZHKQru03dL8l9zxLl7yu7FvK7uCnwUEI5lyRgb78op0s9QNVb
EzAAhjfMGCGgqXBr6ytml0gETD8hBPXg500FbqLoBj8MfwhvVaq/XacMHcK6oVJJa/6CDRfgrTyY
s4CS3wwCAcM8FQVHyRuIboKaiKIT1He9ptqxfbnA99Hfg+cikbrPEHQuM+EtMDmnzN9JpJ9wjXNd
TAlegXdPvdkzvRKdqfQ5ZjRbEPwA+anyq9SS2o+e6X7gvOIf8UUVxSCsi3W7E58Di7WJMJiyS7SG
4UzJlM4T+FXzNWmOquPpFpy0XzTDc+ppEp5fQJdymufOd7h6A2OFU9iJvuodSw7iOf7sfwZJBw2u
iBApPiNY4E6VAk53XfMrciO7e2/XHP55Rvp0jrFEZcrEH/ORijyf39hadQw9rum1xDd57lw5bz4/
Y2Ca+M8qdungEyEQ+yIJbEkwW7WQgfM+27t8WnlFmBTkvJ3XB1iV5lkt+7Xm+eSENZNjlz9Lo2Sd
2/o5WJxR34M4suZaji2eTb08qExif2/ZgabrhB9f8o24ACtZm1vl/eu4q/f2rosV4D11lCoOMrAr
wDJLC1+hikHA0Lnl97cXVrYY+el+GMBif4bRXHv4/pUHJ1zWyIaj/mAyj9xfPRQPXEPLYF5fHxeB
p8kQi8PepOeFBGnp1Ny94w/huH3XcaFq2PxH29UT7ezHXNdihh3Y+wI/8z5MowIv4QkJNzRkg7di
Pg6Kbrsay1xPEjIPgYQkqc6SkbNPtKN27ZVA0fxkXz43UwX1791VbB+Gr8L710RsZixnFY9pUqWQ
wtwP7LCg3Mx880rUKL2FCe2mYUfKV58ndvgFapDZQtxsIcuNb+LaHU425SPJfRpnVAHQ/1L35Khg
Dx5V2VXUeJfil8CTdRvyk1C33TL584nF6qUd5ZtfP5zwh9ntokH3SDSUa2gYnm96Q/hfemzw1Dxr
sbKGFszfTdJca44HxDgdcHKzxxOAn5+Dtw2cxAqnabYNsR+/rzFJntFa4juw7bfFOdk6XX8yOahs
Qzh/mvJLNAexnXcHvonWHYIi410b3KGa48pum5asmI8DukwBYfsK5UH3xRkKMJlGHePnF4g4TmbL
KrhNIbQb1fxQSvGE3w92/8ZR2Sdh9CMO2fkUFS1h7RksXgYC/JZ6AzXpk79kwOjtefOYVu3k3tqZ
cUYnS/dus5LTefYxAm536EWUXRSaVwzdt36dtEoAK1rGRgob0c2MFwt4dt2Y1Yj2ON8LWbWUu19M
+FeWD1owjDecOSiFnxjBlFv9GVpOb8TzgNY0BY/W5Rar9gHACcr6FHAWEggep/ZR3akKicB7Z/eR
KkWzGlh+0geV/Mv/jXmCzn+JSggo87eWvDibEzvnv4n6cn1uvXc3HsZbiDoS771IdFLhm9w+Rp/0
hnS7ZhG4d+V7RljY6bgRBwui+rO6jSJB5Ll8Sd2l5oZemXtSW2SzgWh+RinK/d+fwvk66Nw6QLtJ
G22+Lp9hGKaSr5rj22xWDcDesLzsBwvjlQECVFg/OOE1FmncLg0TVx14yQ7t1Tvwa2MRHkiU/Gb5
zHO17zok8GFr2Ftrvxn5Acy6DZqgv7iMqJj9aZAIQTC2RABLmhERLIgpUmBZbmSqVvk5i0oYJKhJ
wmYMidnRNtZjTdHqXlqejJNyTBlcKuCaByjn3RSi1b4QGou+rNONUoSlL31e78gDR4FGlFX63nwa
75JalewG55Qf0yU207wrcApw5RgZ/0tN6qs8VeuyjrWPGlEIkl7/k6xrKKqbU/FQS5Q1ilhyQmp7
jDcUtV61bKN7Ea4rKNPgLP9zqGdMgRVRqhvp6LuUQwfz5pbZa2pp55betmPz/GgS4FEqLe94bCz3
9LqlPbAPERI1DvGZsrzEvrH/SxUV9d5HVjx/t0SDhVff+j+q88TncIZBtSh4Ulf/NdpJZG9Rb63Y
mjIcJ+aQ9Bm7nupjWfIvKS2cuTUX+eoy+lr4Bg5hWtE0NM4VcOQq3AmkDF7NomZIzIBcBIS3HZCC
U5h61ari8/V7h/ZQ3fiA1hhnYO4LcpS50uP9QaMEHvwH4spwiVQIx+bDGi1q8ljaILlLIIpnNBI1
oMMjbHLd8QI+C7E1Y+hHj+/8JpS25Yi2XqIXAEojM3KvZqD7LKcwyPdy9CH+AVOEei82oZuuIBZn
JRzqK6pk2L1kwXRdp/dXPAN9o/13PUvu2ryWADiGlr6tT8xEnjhi3FjUkQxzcDxiZY+vOR68F/Iu
F+dfTcfU3ScFCIElONCF/Cq6OhfdCrJtdPjoQNzaiiiBWtbsL7LqBRltjvVXwZK43OWxeQysUU5v
P3JSl6anQSOfrMA34cWh1XpvB4s48X3g348F/3zNLnI14cb5Q10fp2sDtm0lHHhFym3FmplGg0lQ
d2Wwr5nvRsc9ugaapeb1JFc7YRrTMAGIKtM4YZUGurCJi1VVRk/LAm9ZLdI1d+rpeKeTYG885UJs
5jSK1H35N903AbnQT4Ikl+y4V/nAMIRy+g2RcNaTlAtFGjpUhWuFJLGigjKywO68AGCJXoHSTCWq
cn3MJG6Ji8Z9k7c3RgbnorINen+0y/hFWI/zOp9ttbPEohB3PuZP5TOaK0w/CJ93lSFvl573FJQx
DYGj89Kp0rYqi6jz5fzXezTZeArADx2DT5USKzlRVzBKvCfCH66SSLWFQCjxWepp8z4H1GjdDuUc
kcsaeZRdIMbe3hY9tAjcbPzJeHo97MHwJW/uoRPPf9d0Fae9kNE7dCJ+Hc6XV4PAgJMwIreAqdXK
QvlGc/J9p9hZEZL5pv4EJZ3hvhJNf05VJubFUlR1LzSNpMsc9uBeegHdJ//TCWzs7/xLSlikThiY
KaLTryxhD/HNgO+UmtMzz0fSACbVeo0vl1veEDXjmZwWcTBfUq4+jqG5mjXP8PjDmto1uQiU3Qa9
V1Rbuqi/S6aTikzYJHtwGPB8OPxlUBuOEr9vKALkc+CqDTMVz8NqPM695C3dfbZj2jAj3dsAbe75
YUxW+svYFDJSQ3ShMPeA4yvfc6bOEywways2mqvZQ8SM7bjFVt/C9WCk7817rsOSpz8QCOV45eeV
FoHVBYvL+lM2XPt7XLWKwJuvkwou8UqDIzqErKY5UgWJZndhWLV2Toh7Vp6a1Qxspw/NDN2tnWpu
gHTQxFaBDoocGZfN/lY+0pd/qm4eJDIrBf048kYdiv3iEpDw2K3otoR59gzx3bFws6bRPH7FFM99
USEzutU3N4MTBv137P0D9pY35bqIZUUofY3n4+6M1HB1K7aUzr/AQIol8ybFqvd957ZKTwO6dSqL
pyB+Wy5jaYHPxIyOkUC/zMekE8wZ2SHSOewEcNmu5Qu8psldN1HxQiYnEhMRuLmMVAcDSa+GK3eA
xF6PCIT44TyQ4A78+BSoWxR959SFVcgag1EpQpnLSQci7cMNETMMpxdVYm2WuUzx42xj6cV7ogfT
7bBEeOOjb1p9eWMNhPkyIAaGtGKajUx4EeR2WmMVPrk65MNkgVZuxkGX3JrDx6sUFlUjnDZcKKcO
RitPomdaTYdY6Lg3BIwAy+3RAzl5Di1fai0JRozERXXQtAprNDqwqhtIz/2yMdxe7a4xS9R6QLQw
Q/Uw/9HeELjw+9So2Fyq7Nw6jr9TLw+9osmlnK/p2d1oSrJ6z3jH/HtGtpVXkt9kV1m5afgzmQhO
gz+ZWWgofUCptjA47hkoKc3B5Nip2pwwtzuT04SNxz9YMXzLMV84K5O6M5yjGoxMHonTpzkcI7b5
nBnF8PwIeYRAhfACFbBDJjXhbmNh5A58Z1vEOC4ftpr0IFSLMZ5FONd7tNk3peb3wbsP4qmJHPhe
DVhp5cexkAJY5GQwsFOXR37pqSvRWrgLimG/KrsICfZY3GtuGjlMez8SXwXq43gmTdTXOT9yTAUU
YzyNp+4RB+xJMlJmXXWVJ1UOp0CTBHxJTB2ufzDa+b3ysGY58uRi7Lpvl9ovklD/pDk9oq23U7Rn
1oouAce79qYwPYdsfxK2HwggnBusOmcmD6aRAvpHYlPYgnchbeVYkwbI9SzEuRadk5radD4Xb5P5
Pju+1XBpBpE1Qd9bCTSl41C0tXnTg1DSRi0tnR3haz+u5tHJTMGLN1z374XFjZ13HpqSDMoCip5e
UxY0tWXdtZruUUIkaPGcysSsLQ/UwblSY+dTwYwCF3CcEWur1VdD3jyxsJf2V8uL8fdbccZ22RU3
URs0pKET7vNTERyv8+otqoKsoixeZrHUw570ab8HD/XX3WYZZMm4fCUChEwOtGZC5cgLDHY1L28R
mnOOs8VHXsNp2Zv7un5kcuXj1jJcorEcFOn3fg4T7Q+cZFVHhhDkayWJroA22XalyANLb8xNWnR4
N1bw1j217I4DAw6GDXH8/3vkdta0yVASGcMd31N8PjUY5V8HWRcG5NAmoncmq9EXwTU/N0VcBdwk
ckoqOr87L7hh+1J8sVm5A3BfFvp8wvjja3sDoi/3h2YvCGkdS1ikilTawXwzJbUrMYfgnHxWDDAx
lo84ISHae1r+La3HvhaMlr0ZtMyZ246Od8zfkVGHuO3MlIUCzgcXeZdcD+yOurWZD70JAhCFxuJr
0C6yP7/pzHWGcldJaFAX+5Uh2eW/looHNh6F92NMtW1/4EVuqdCENR3UVme28uWRXd2UQ+T1IydZ
mn51KSmMzeJflzB3s8YNuEWTPNGAeRG+n2QgWYFH9CfEFzDKvWup2FQI5iylympmk8mgHwpPd2ox
GtKx1P2nz+7L1SNfp+A8C9/pr1tG6ZtbT4PzRGQu65W0WC6AT6aW2mgNP7SsMxwfGo1yFGv0fBRO
E6DAg7YK9VZqsnsS+4U+N6G/QwmplLOgpkVI/qzH1o7qCvvLTSFy6Lno4DFpQxPszXWF+TEtFe0l
Q/MYJEsbgKgbkG4VRBmuzyxSr+dWmvltbJWCFeIG4rRWiCKS29H+oQmj4riLpEhvh5rYkStjNc/h
8uoqLD+sMBuzhcfcSQqOgC11LceRe750XgmHmWXZ9jhEpxU1CZUwSKMlMnk7F0zDaotJEj2+sPkf
dsTDY2pCjT1etR5qlif6YaHIAe9WX57k24N9MwsA1Lg4MdxuOsahUbspPvCWi06gKkoO+LlPf9bG
92Rs00dvY6VImNGYCxWaPELVYBkbsKoBaBG427QxrOHq6CBJ6jqN4vJhYEm1pCZE/NJZp7SiM9B7
6+aEOxO48BcLm4+O9zV1jIqIEyk3Vp4d4i03Vwlt9+uxeRJy/RLdtUfDuCFWPYZQ2cnLW/nhzZDw
lvN4fUX6gF+hFx/xOuB0QHp58UdPi9+U5eSn5ol7ouRDOEIJmBzyH/+GO6cHm5txvRuVtR+hwxge
Apwtg6dZtFpbNsaggZAPh+jXF87IgLiGh2dfgBSCe5LQlh7XxanRDtXtxQ2EIO0ByBPX3WSjENfv
6vkyevcY1qhAZBZX/DV3jy0eUi0PlTBFaXTCCJ50jdxmz6Ho7BYYBVEblUj9YpiclocLybRQqQ9a
6kHfLcSVaTSUBIXmrsQNjY6p1jPz3wl8+GufyNbZ83v5pjSXf6gNrMFNxxM481uyneClOmyijUC7
BI2ONhH8eC1c
`protect end_protected
