`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d5VJXu82JfSwswDjhvbEU9He9tQ5/1Rw+4/2nB84LUuT0wfekcnbAADJNd0/JtXdeaCUlOw7Zwks
Bp1VvQeB3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T1a12gH9+o/WCd/uq6lAozrIbwFwnflilDyEA/rZKRAxvRmKOSqBXtjVpxVSoEgX9El2BLPK+36k
Vd8y/iFx5HcwlteYeuYuGTvgQerRA9ycH4Qwt9s5DC83MaSGod9ecMMI8PPrmdJ+hCOX8sXwEsN9
IHAKBa7h08XDRsgW0os=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZE3CBd8eugZohbo93EvXvQkUxCnosHfYT2eG0uuvFgW4E1aUdxFin2hcHpeAodvxBTyPhYz4Lsqw
3nsUxnz9hTb8Lhj5XnlqKx2mVFP8Z35n8lJk21C09QHBGoSukklDPI8dbQUv/KxN+k1qsLBHfCBA
FWz2UAwKlgCaoOPe87s5MUwwDM1/P/D4+XgEQCRDz/7JDN7p8ZFVtltMEx51xjJOCvfGoEeTzG2k
908lkYgt+B4pvwsuFOHwC28xicC9lqwuIR+OiqTI+hvqIl3tijnK9dhEHXmlIo9PqdVp3p9K5niF
C0wKwI1gK4zk+Z+Qv31AV2g5KDXjXxSpUgHlpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1K/c2Exmx3hO4tktdfNX/hsUCqBDw6bH/vDRPja11f/SX2mhefMgy+yYp/XXIVeJlyTPI7AwLQ+m
jPsm9qUsxInkPzY00BDkxz+XjPmDvPZhWK1LaTfp3S2KuDInJ2AYP1AwgClVQtpRFpipBFYqQeNS
QrfV5V8iPYsCh6rtCZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z2R2Fz5uoP9gCKKJ4H8ByaZdL0II83JUVbmmEiqboGhJOssYqqghHZS4Xla1DO6PE/W7lUbFZBMN
taobe7WZ5vLL3z9KT5znQ5u/8vqZfQZBnNTCM9ij+NRl3PRmkUPrtcd6xURukGspBspXFvJDNTq6
HoC8rJF2dAK3E2hXtQ2qzFXYx2JspRBZw2ARE4ENjzYZSYK5AhF3nV89pEvyjDlChnkSNr7Ec2sz
zSK49rQXLtbokqxvvzCHRCEs+NoMqKlklN93OyjJFAIzYffS6GiGtNeycU755Cv+/fAQynybNWn5
4vdHnb+JcudvHzAJFK7/azTzKOJrOSm9uJYTZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5200)
`protect data_block
mvi3i3MBI7n8zvuunOT1BDhfZ9+75ngvsPXxp5+0g3QEMYSUqfdm6zc+CwjSUXFsRgLaeVNg0vh9
KTzQ7M9UvhqeIJs1RJ7aoXCOWi4NjuDVIH3MyIK5EDd048RXQUSK0FLX+6lFHyT5InJGYSKGf9Iu
f8lkfn6yc28SokTMFCEMrheN0NwxFip0ReF8Ee5Pc2dKl1uGrdF0BXJ7UZ049Mho2D7hOHXsbhP6
/RJLoyVr6nRCr1a1MJmGX0bGEWkJIs1jSJ86pFMVX03RQSM9+EAT5mT4E6KDZYm9N58GZ4/2TYmG
Le9tMXKnU25gtYdk+QeIwmL9YAkqW2cizT3yFzIJ3GJOxdwKQQekylFiP22Arp0YRD6jdTCOSzD+
qLATb2gd8+u2RJPU1F7ee12oxuNMYopqiD8YGpo3jPw56RybU4AfbAWDWWx270rEZPGJdfLvZOLg
diuudRAHBEhvT+AZg3FFYRP7Tv3aWR5QXPOh5AfNKAGUYbEA5BqCpeg/QQp8hd4tu2Z8aq9U9/0d
gSO+GZ+eH7ucon0OB1imnzVUu9hzawkdHCN3TN1GCnqlRyvh6zHg9r4E8i5X63lw4kStqH9u/siq
byMTilnoACbmTvEVALnfoiA0FVh/KHbtEbG1o1aj1HpQiM+TVVvBv2sa0F8YEdUZS0ex5GCVcdOV
1op3A9yOA0vy6Px0Y17qEdniKeebhFGDvxIofOWSOieswyb1fX60mudpT8IhaKRBo7C+Y88J5o7M
6yrducftSO1WDEnPR5oSOeMdLrTLXsx2huvp0/WiYpzSgepGPNSuVsdrieda42PXNqYwr+wd7IeM
sXzb89WEG1J+w8ff8HkZhOSS3c57sJKEgjpKqQEfULabc+KZCQ1XEFMjGWfw6ARgR9uHEMkMULx1
SGRHHv1IWl8nB5xUfuRA8Gs93qRNji8oDwM3W6I9p//hG/pGlMZ/PMeo4ci7VskgSZ3KGHPi2iZd
FLmJd1pCz7XiREKT4HP0qFOe2kpRLRKRUCqO2iqtzn6f9yAHvf/Jxim33bjhNE1MEiF6GN556Aq0
uEIvFKYubeC1fjYnTTuhS9CDJWp5gJHwPaCcANePSrOBxzw1hpDhg2n1msRSjmn0i4Tpo4noovcz
+98T7Qc78zayn2hIAsCgEmgbgstR+MnhnKQhNQvjOxFm0/q02svAv191eTZ805MduReZ5MuiSfNB
K8lGH8fohPn1BBMmjNlApthySeZ+zkt+HmdIOvrEgmKAJ5pGZ/x+2jGT5cYdJODsGBabXUWJNSRA
Fl7Z2MD+VYo77150Vj5rq7z9dCdN3gvFhD9QgGa6aY9eQ3Ct/MlxhAoD0gYfzyAqw1UNszpTK9ae
Dqad/TS2d4mmUbt+cfmwjTgvPprD8SP1cGA+y8Jm1+wupeLaHW0f0J8IbMI5pUO1C0JFHgwnA5cm
Iy54+GHjFR8LThvZ0pIDnDbi2jp5zlc0WfE4a2fgsM2/si85hfxbGZ6XjSim+cSf62QNdKzuElB6
pkuOTWDI/BfT2L2GastdVyUVDrHT0k6BvrFkwzZ7TgNEUKm7nvitmbbT67oIumIagQIH98gaPk0y
kPwKnmN0xucw3S602iVV/5HkX6SgMuvPBAZOVO5/3ioAfwWEA2EncAzJ/auNxSWarDgGLtWhH6Gf
Z8R5YRIpvpbc37UFSBpJV9gBUO56xtbt+LVoyKEVzQ9OYg1Nhg+F1a33F6hblxgJD9rhgdBxX/2R
/3nxDtrplsP1dtXZiGy59+p/kx5Ao/iXGqnSA4BwnR72iGSn14mDJQaDrM/22u+mf7dlEMcQ3mRG
wgBO/vgH5RsYvPTGxlaH5XuadkpKIDKGArvQ6jLImZ8gkCzO12MPp6xeZzNWilhMwDWhxEm3r/C1
DIS9fGmlD/gsxlxi3MZ5A9lZMD8LM4S/JiK8x6V3N54SZfY2RyioL/ClGHEmCRqbLNRTyOwDsP31
jCTFphGPrv7zsVs8+ycQM9RrOpMkTZy5ZUWyVHe33VPqFCgtG1oOy5myS9lV86Kfk5MTxmaGA7Lp
5bTLtRYzcnn5chOqx2OHVQgufESFfpUngCViGU1erBX1O4HH8budrblP1vUNqTECGn93r0G4mzB5
z+8xFqSAiDbmHrdiBzdavuz4Uu/V97IJzAy5FZUAJL3REusdrSfyL17G8Fwin75y2o755I8Oa4MP
Fez9i5MFEBSUfr+LKnX3bovKiB3HslCSIY6l1OUPrKsb1Id+BaQV9D68bk6qTq9i/ysJG9Z4OV9j
el90lPSGpe8dQb/LfMLm0lOZphyr45Wg962WEQyfMWD7ofJbSISiEL1CzWglMqKPEPpnWA7mf9VM
BYGBmMYBXE742BUNBYB8cbn/JY4Zm661TH5A4xHuvBSnI5KvKsjKHVHpSAyxDj2ISIxoNA4Rdara
3GOGs0z8rUw96hUQHoAHjeak5hmKQ4w60D2xKP2j5ZueEmRliR8ezG3kdPDNEzDZSy6xzm7+093a
S7vIgzrVjTdsrdXrm6xcn20gaB0me6GLDTnHWJcOtl3Vin0LSFMHDt8ieOWqGkTH+BBLHrX4ieGG
6chYuTsl+8xgNWr5dzNLHn81YM4ONShwfgGsTMcQaFDTzHC67c0lq5sOij89lpBVKpsS0at5CTut
qI5rGClhquVeCTyQ1gTm1ZvFfj+FSd2KPPxyhiqJL5NT+3XT6Na31Y8rPYCM8KeZ7aBEUarrvoK/
ri76pHkoKZk8hR/Evm4kYfpoObi2UNyG94fs0/cidfkLpL+w75w1EAaopHTCTIzuSxpd/yEvArIA
0UKrUAmMZgukqEszYOy3yJvcruMb76/h/EtBbidpEzHFNkzluZa9/qwTEaPMy3N72fwboDsc05rb
SBuSgK2pLbVtv4CuTEiEAyvfrVTFVGTtVmuqMHDAmhabPsb4wmiWhn3eGEoAmcxxCfp49kLbrTFz
ZVWRlbx14dKUOe5IzAlhavtiAhvK9JtGPYYbr6M4vXSEccdOiA/KU8LRtB3xSeRPGhQdwQfkWm5G
S0CMdpFYul6WrP+DsSJf15sDX4ZRMaSGBwcBig4lBgsPrc+EBGwwrOz4Cp4/oFTlYwMZLWUU5l5D
owYIe3y3DHRuEGTSffWd3wPXOz+QYP25y4/xB2fpFlEyixY69mqZPjliq7b5Cy4F2hW5ywnO9x1T
ufGvGY39985330Z9fNcXamBTP/u4iirG0zdWCqjD8rWIXNvgth4tDsTX/N4wNCzHMX5m/u8TJgrf
lvkj4XgU7ZOdou02Z/Hv8VAchP5+kVzWwn8SmlE1cePg4KohAWNOtalc8SLYK7Q26bVX9d8IvsY/
20uoBN/mm97QTHVRtMRPtNuZzuK0aHNbdsWlV1jnMH6yaWiDkDrkHokvvvFvKj62oJ4qKSuibv15
f9YqvxG9jg4D37Mu7kBrhowhhfqb9jO7H8bUtQE/rZ7kxI9HzYTXLmBLysvqnMf6XlmYK7E2+0Fo
nfPczUSY8iLYbThdf3OYcbOcp4C03A732ZE8f5OpnxAA5zMXZl2Z1ckVyhg+ljXUoHfRXV1RKq5Z
ktHd5T1JKWalNYbyQwmG6BOz6KOIZePa/DU0rqyo0mRYm+FfKbViNbvYE6/c85mx0+3TcMAaYOVa
ro1g79wd/2M9S9ShhosTIkhUsKj7XF4LKGQzAqzOhTDEGGyx8FMRfVefs5XztKWfUX2WN9nb4Jyk
c2m43Zrlp/qlqKmdnNuGWJuPc2pWGiLiDH1+1eoq6seceJH1pTVH73WAfuaV3A/Six+jajq0AFKV
B54Y6kwkbDDLvztOq3Ph7Cxw0EIKQ2HWHOxrS6a0yEYVxa3KuxM/m2j7TJsBbJQrHIEp3W3oVMTg
zjDB4g6UcgGzMF9vripnGwqr8Bc6cxvSSCW6cPfcLVGLAL/IThOfkK0v8viXXnXmz4mgtHyPtjo7
cvJq6isVmo7WZlS4WNlj8z/EPJsVyQ2+DdO6i6vQQKfmJ76Lj7T0td8dS1d2QOAeXNsLQldl1p9p
wQy2IM6EdIjzbdOWPppblYujxdVruHmUdIvqd8MQQtJkxIUrzgR07CWdt5NSojEmNUaEYU48SZBG
dQ/RwXcYg/6j90gXCNNf2d9xvi9IroIXeiYuQNROmW4WTv5Yo3pCD8kKs2Oz1BMFQQ96J2I9NXKZ
1Jwqtxj2gwq/4ieb4Bo7n+su8rR/k3RaQbMAVox0DINI04XP5WmuxDfUXPc6MQRRy+/0ShEnwzUU
lvMCy3B0gvbuP87/7+6gC8KMuqGONGYIWwg8tJ+T3tOfcXNTaGuwco+kLnvZNDjLTHocFacdEG/4
ykwjRBaA1POuDHZUdNTaIcAs4lPUbcVqkGgh69GmO/+ouyljYkaNPnagRZVTQE6CbKVkygDoE+Ve
kZdI2qwJLp+n3YSgEeOSlZ3CyWaZqTmBV5Th5lEGtqXhcejPkk7uV953nSNsuoIKZBEI8QenXgFx
9ieY6dvSiMu/YOQ/IRGs+SBalunKgOlGWQOKVIKqHgvyZh1E6qdXXJbRlI8m3/V9NHq+s9REzVSM
INNSycQzoX5BM8z2tybXu0FHr/SE/3/IivX4st169A6lGDQUVptQ9FyHi2J2XsQuhyPbuJutco1r
3QDLHPnj/yD9io6InRs2d7NxrszoI5QJLq6gpotFdRQJ84RRWCTG9E4xnPMo9tLr7+jeOx3Lq9IR
R579ftoTPpL6djHQ9AIPpJzmQh9Xm0lucX5lfAKnjX4o2DJeeUEeWWfAB38kHdghklpwVgTw/BlK
lCoLfy+0TRYL7PUoGDQwGoIhzg4iKHvI0MtR98hs+v+PgArZMRgz9ewWZwzsTQFUR0Me/9XV8DVk
KMIE6O7L1AQ8KbII7mgbfKJnaH6p3tsSCDipqHT/Rq54UyW0JYSszamMLrLK5mQtRkk6FUOkDwsD
CGnN6luStr/1BhRPlAfdS72y4ab2YGMz8F5Mqdln3YWy46EABHozx6s5+isX2GsG4bvXrzgjwDWh
uTrCNAgv73428Q8YDR6PNr3lKV7zCDqg3s9LkebfYWOSK9XwWTZXR6+7drShmH0iMUPwEzklg84A
EOJMc70WlsMLDAyBBYv9jV8UyMg/fZOIN/5BUMDNYOfaEYW2S86uv65p8hjcHt2X7Y+ZD9zkVoFE
l82RH1MLqlZjZIyWdYOXTvz9tzKboX4xDlQpQ8ZFoeBR7ktZh5cBHYsl934h1owp5JvkkK1mpmcO
PkBl7wQRZWJWmbCa1RVvm/ENibMCkS8SVBek+n9z2xwPlVfZ01WwF5ouXxuz7uajx67FO9At+VsB
QOunvN1nKfIMdNmQgV9BWMEMjVpYl4Bt3BmssTe54PKbAsE7yMqM5VBXGRnMSDY888T8a7ktaZkI
2WxmOAHJ98uklK4s/lktAH9JnyO8fdAQ957hT8p1xgnuhWDRGhitUBWGoFGSIcnj3hl9UcwwrLON
OIUQ92D2UrVMD/aWYJOA8wI4vpVYT19m3PmCAF37wa2y9AQRTml9HKA+A9IMkwl8QQGkeBtHMNea
V/LF+7Q2iGUV6lq2WMYLzh1bLQaRZ463DoU6eJ3MTSf0gwHEZggS7hTDB8g/b+i6hy5U3RUWmdh0
oM1OsJmcBEzs4tTGCIMljl1ao+nxWOytdfw5wdYTIBf+pr8SyzJ0sBw+4kin1IQGbqraFeeMc7R4
xbNsj7ulhw0msM6+9yCYuWCu8Pi7V7jhmixgB6MFgRLL3/N9aiCiXyG4kaIp5DcpETMYtGvvfopi
9rxnutO9AftTj/V4deV9kjtSifflwWxBDdqDq473lq3DxJkUJO+uCHHvtvgV3jaUayC1IfEio8RB
9602qRS3eKhYYT0UgxnOrdsiipALwPz/G1gUB5QwdcRaVXzFTdwj2jozqOT7Q4WW06Hbg+gSyqPW
tw7E3aOEEh7IIfIe5XbYwOoKXD2xMXe3xnzeV2AQ/QaVClzoVBGWW8uID4amRgZrEk5yxzM+kfZF
LwCiAtCajfENz9wTESSyp4vbNpyHdlJWGyHCPYzapJordoDZz8I+ldLaWXf4/BxynVBGkGoI1VJC
DsymFWeK7cc5HWyxKwyZX4zIFedpm5+5YNOTZ11f426C8dJc3R8CJPqVZ2afG7UWI0X/gQoFLOvZ
cLRyJD9cgSINVM5ciyQpt2yAtpngS4WGTMPKlTg5YGLxNL479xw+TTFPFT2ScuCN/3L6qfG1oGSd
hgsNayD4fqHap/i68xgjAgKwM6CwFnPLRQrbB1HbXffBr9+TVNnefVWfDmURwyLw9nJE9VlNI3oL
NTPvq0mFShwCqz1zDVlKy+Eq/UiGnI09rnTWYh3Cf2KVSjEvL+p89leJFJth3A2rgPBMT4DV21Mu
KgindOdkfPOnbeBQ6F2ISU2xEP9XdxSNyH22J+I/U73ZwjKLA1Qu3Nkt0P7L1ViNShOzpU6HJP4M
jqQqG7BHwNttTH7uNGvgMNh8lqO3YWsl0TYp/LjtQVmaWD44NSI8Akt4L4UhbaeBu8Q8SdfbvhYZ
PM9+VffZiavkBpfS+CI0moFbjKN2RKvql+0EAvtNcpFoTIJY2fbkMLZrGS85WTj3mX42Xj6KDlY+
7CHeVL4+2+DKNLFMhuzerMBVTCDu0zfawl0RWOlqTf/sVfIKxb2a1H9XU+KXltSIhopyXP/ZYBtc
INzxfiBRDCPl5TcymZlHkEmXKBJ7KOISUwZiL7qFNTd7YwZxFhpdA5PQ32khivCAZjAkb9KquaXX
O7XV9o8SnY1Nvh6ERgFRUagplJj6NbufUkMZI+g2AnT/q+KIBB5+j294TnjUZoIPqKvaxmjZE/JQ
/wjugKvApnjopI4DhEbbZgJAd4p6KTz6rTPaV6M4OOH2crIcZJ1vg5pHQZ3kd/z6l9W5zuME76x1
PBnRwpc1ywMQODdX1Q==
`protect end_protected
