`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l9rLb8eyF3AgALThasPiNG8/4BBm1wwJaB24bneaCtyp/I0xi7SHB/t0Ctv1xqonweX1MzV/pVKs
tQdRNspPIw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X5KWlL148JabgR5weT9wBUkHFWddJA7h4OZFLd8bdBf8Kop7kg1WdkOhUDgmpNTHeXS4I+xH4Y4Q
HjFAExnYrGUC1wm7p5WVL3DFzD5WTILYoEImzLFNcK9/mSAIwCGj+Wtr+9xrMpQDaly5jC8Sj+rc
Nr34z/YYnZpZdFjSjFA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XOX+x3GXJVQTrGGT75+NpApkQTW6W42cmWaYkzqsNsDYv4er+FitAoIemlb3od3AsSf9WRWhCQnT
6iXQilkemT2DzV4Xsw5A/7I/FZ1E441abMpjv/w5Z3kwpJvNtJvcGvjcX812mAAPcXsPvrB5LXuC
3JiNsCaNzfl0IQulHvHCqzDHmgFxZRkHPXNoL3EbdAxxa3qQNIHMXziT6TfG6V4ioLwZkfmj+nFw
X+PAA+oZbdjyO4IF/qvCl2mnZ/REv5vdMZsnEZ7xmZVfOO9rMWwJcGnuuXesJxcZqnyEOewdy0X4
g5x7ACzMTBvW4JyAsNl6ipSaUUNJcxvmP1Z95w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
umhSCUCmm4WZMMJVCjLiDlzFgH/9KhaxQqdvYM2gFaFK/BSZmXwKtVD0oGzsfgEnaEnfAZpnMH9p
W4FaTz2HfMA8FyEQD6bKpLwcrFDP6FLYTus4W9auRkdWk6MByslYcfESnbPd9BplDCjnq5X9FeJm
J+EfUISXG1WULY3BqQc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NcJ7q/waCn8/m5wYTzYlcTzCH0J7XhsrCXDcbP801wBgwPzwk6W1YaeEGpz6w5sg9/BVkYMZPdHy
s116tGvxEU4yIAoLSq1V4khC1G0CICk3cYOL6Am8EnS97sHVRnu2owQQ8/o01YRhaorvw4ApXGQo
FWXh1RTAkyoxms7xpWs910xGCq+5ztWRsH4I8eissSMkhuy7owGmA0f/OPnBvz/16ynnHSqeTcgH
5zrPaJOgTZH9aMea2bstTOpguVDKDnDoAXUHV93yikhxVZbDx6GaPXUh5fshHVEaMG3kP839Gx+j
prw3SfsWydM2YztaOjt4rwHOeUOZ19sYd2Gsaw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4032)
`protect data_block
GMQYRLdIBu3cBPESIImpy+xilfncLnKrvhSWmMznyv0ADj17ArV8k7sJt/5+kB3lDxZe3EQ9LAKs
LRseCEhmBpZq/WJhbEk4B+Dsr8KXINTjCGnx2aQgJr7M3WSj6oxVbLErFHnnsLfcC9qteWlT7o5/
VGi77WKuHIzp7dNvPZ0y1Y17J7YAjocvgWEAk/0p0OgzPpWE9BYJrvZmWqkGpQ7pMYQxnozDV+i+
uJ87Y5frDFLBQwoq+iTysNUUWDoP2nWI5L8zzNm4qufWDBLY2e6/Hm0wPDM5wqmYP0i0PANREPYx
fm8pLluzOqhnqRJD/uj5GK9V8sDQKsVzACiEOlGhX26FPpIfvj9+e6kXcwUZ6I36VfnQ4wMinZub
oaEW9laMrY0p6snUzqGEMzm7lcdu3HtsETGnWsm+Q7y4+TMy+yNw7eSoGJrIv34DvE+Wrr9kM4oA
WKvyh+se7a++GB2P7iooslOWw4doPuNZaWi5z4qQuh1/nPr1tQPdIjShZzX3EXdwcFW5YbLrb11u
m4FhntPXwhzfE5vl+REHF4Bf02DgEfrjcktcmjVGrqsexeqUu90eHFqNv9+kmPNSiUQFWtoE6fve
7irm+vmynTe+ZWK7y6XTDl8BUqgFdeex+wJv/SifqsHxj8XLQOBKBqMy8Bg95pICy+HlVDr/4Jtk
zdBuGKSyuWXtd8vuux0jB32zjKRz5Tu18sFanLHqv/Sho6C/jZfpjbhZowJMXjc9JIHkCTFAmhkc
C/vY3JwTI0hOYseQYHU5Ev/cBgwgecwUczzZB/OS18Ks9Q+lR7m2BFwavPoTLi+mUXRjQFSJjfhb
KKVnJzy3ykG4xJHlcGf4R6PSeN4tOO56e8vs6okWWV/Ql2YWI7PiOi9wRDgKFN0gtgTiZ1nFKYcW
wRRvjFkgje5kyF7yOjupXH6l1E5a0WcgLCVUINxxAkRIyJDecDP7VY6jYctawqvhnHxcH9YD9ylV
dQ2nHpgZ1hyQRYFDj0cmcwOMZ3NoKBfpjJU+FKORNfXjizB29gA5DtwGrDD4YRoNGvPANYF81S0W
Wecb/MulwUAppFNv2Ob4Ium0cLymfCNcuxE9i41GSBSQT/+K51De7jjsUQhVV1vwdAPLMZyD9hKu
QSU9wR7j/yPo8LSn4w3s1sP9D/7YLKHrsOWNHMNoaab8clP7Rx1cA/ngoGUdGYeOyrKBjrzN9/qa
1gu/nSBHyXxTP/tbdYKeTLH96oHuVDTw+brBkNAmGNU2wLCW6yUVUaiu/ZU3Pb/yYV3tJLcZNpnf
PJ0vDh9DJMMHsrJx/tKYGWZKajedfMG8h1rufui3gXfVNlD6cxMV9FZ4LNsYfRjVut00+mR6MkJY
ZBhKq572OcpgRyeMQQpsBnfFnRoYQTE6oczJWbcIuZp1gzN64cm99zeXfTuQ9QlJGkKbBcASHc54
P5yLwV8WtAfyOlUZ/Ksr29VOmhICuyRRhYn3zxayNAduTDermB0nqL1avg0qSIhew68uRGUlDnR+
4ubE0pk4rVd/MdVQOCswk8IHarf2eWm4MORMBuSdZPb4P2qUmliHDk9wVAolsAEBKQoLiFSKQmPV
h5WWlcBsd/py8424tFpPh0t2uxWRJoH+BNMA1Fo3x6trWLO1NU7GF2aD1Tsn42YY7Vhbh4kNekZb
JfRipkFfr3MRMtoHbCJEufkKNrtLycbsA7aX9arNzEIW+BPFm6f7GoNZuC6mQ+aXZBMye22uxyUT
QoYkapUUB4niUINqcHINfnFQwFTtNXVmA7qgdxA6KlScGyOR7oRy3+PEsI0hGfodDPelMInUvVHM
TwcoMFxwadKj9MKSlUvlrwzDH2/1No3MlZixET/cqNE38onWk+8Xr89BL2ReWNd5/Gzi3rI1tpKP
5EVfkohfXIHDYBGxEL0BIaV/C/idbNlbV5ICymNQVvAJA8r6jtG4LNoJZFTcd8O0/NaJxsQV73eY
AwFVlSpDRuNZDrKhMdSQOPzXFXejzZPYxQPEvydPa6raxRKF8BSzD6hDrNr/Q6lrXRqHbrlrCFSu
RmH3eDKOfY0qXgCzpSfp0AudalWSAca1U4aZ7kl3SniGX2YdAlkiVsOa+eSwKYoVH+JRXmoMQNDC
r4TRC3/+IlfpnzsBNmixeqPTfykLnr6TZESSRam8mcLdqsY1+ogzRWMdz0QrJnXxUtBLbF4D3QUB
m116AUBE5T5e0+dlhqx7gan/KBjZcCn4cL84yG3Ya5xHXsEx2ysZFpeOQ70O8JUoktegWlAbvJY6
m0o5eWCO2/0Mz+TAtQOSHh5KK3ODaeSkGLb0Pa81XC/xUQgIxqoGsoEczAL/dC7R1dSTFfPCbJIu
Xc4AYS1F3tdp7HFvP5rV3j4DQ6AbmKyQUdeihy/Z0/HheiEqoXHU7kV5sYsMHnUo0IW48FDabm34
wHE+OpBZezgp38Zmg71AlEKGd0A9sWeTW/wwQn5+ylaaeMCA4QV3VSEaSphZDU3BegIChOQyGygU
UP7KpmJ8LTtqDf3z23wDu4ESg3QDBLps3k/QZixZ810lOY7qESUbcVOlte+sMZ46NmLUTJ2L6U/H
n/+veZZ/bD9QIKXz92JtY8sIx7xReavOsVQ2QKksTyKtcQTg0G0jCJNcjQfNOujdiCyY53+HIYet
ZyDoyQU4M2tgdCpITb6gQDhPxsS3NrRm773wuV/mI4UCv4JDbyZYzzdOjmap87eR4xsDUNLXiZ7K
rjW3KgJWXoDZbCyKE2EamtbNCEUu6KJyTuqwCzjt3xi4sxhhh27zPBgQQk8bjEr5qZTK42eTVjFK
ySLR6BFw2wXaW/cVZS8MU8mu+3/sRZNy99Ryg2MV3WBUtGKm7g86j5vUvj0kiyPdRNBtx1Skf5bB
SNwrbIZX0k76KzELKdumcoei4U67UQByizHhz4QjJ68HymMBg5T+00XEBlAP/jJWIUm6eMY3/AtX
NWo3ltEShwgqiGFKG0XZgLeYOTrj/n7QJF3/tW5La95CHQdWPSIlr84qhgAXamWpm4KsJHzWCj/6
D+rWm797qziQfUsGJuXGhwISlcFu1oBof+rkI0j5/Kjd6+SklZDq/Uv84CDJ0mJZ/LeIACc9KVTq
has5Be0otRnbfHqvRl6DsSV/IAVLGqhrJr25F9BVjzkho8tk2lPyT6SLHY9pgr6M5y97TQpowJ25
T8ElJBpBPCgitpFOek2ru8B/Kwj9v59/vN//gTLypQ6AISWbTAhyjVZy18VoaE0qhatRO746AA9C
UtVqzLujugIMWj/TIjjt9kHe30W+IFBzKyTvV77fQYkbN9ggt0bYeP1Hp2lUbIo2dq+GMhcB2X3O
rSXpKBbe9+H9cm3EUQqKeusXOE5aQh+H+LKGG2DmfTedAHUNNUEEC8QckCmEo1TOvK/UY6K4ysgT
afkIDXQ0ctoZcrdckCk6QmBJ1l9hoLgx1PR27syAZJUGiqBPKKwhMJSf93/xkGdjUOcMTK/KDzxW
PcF3H1OkPP9Gxr0rtVjvxXrBHPXhxGTLm2RcFa6S4wT88unwiybJ0R0SoMRSSxysURERpPYvzldi
dPKrBKDYO+G/59VHwaex0aXdhB/l06jcUa+YG5AZl+2BlS6pB4CzI0IibGZzSLmrAApNuCmqzPCM
2FChIoO3h6cbUV/1QD1QUMzZRbTzRsHXzhf4P6ht81MQ98cHfq+CIMm+i8Jx6l0O8LLUM2tFjJyl
jjxI3WYmvPSpNG2Kh8m9Rssrqg55rfWd3FpUbds/PXqGwsqZCuNDXhmmBSPob0Yz+WzjOPGYtF9z
xnpmUsLpBv6v8AGHpwpYwC8trBcgXg5S1sQQwal8yRJC2irxINk6tGKZo3we3juiWkL06u7d/RNs
aDv62+iFeHhgDYqnh44YqIqS0uchsE3RJQLQ5OOmXZ8NdpLLDu8hZDY40eknPIK8KwDDcYtQp3Z+
kQj/tGoXV+BghvP4SJWr/nq8qKeUXbXhSSQluug0AjDBdqHeb5/UhblmcsUPWktADLRm+AhHrbkO
EAlfal1QBjyPivez5JfH8pZnU8R7IHINqhr+/cUbGK0FkokjriRgRTiLB3WuNsBAecCcThKuqlPo
qCzHBKfO1EWrZf0XCbPeAcbqzh+bEtl7PBXCIrej/K/rkJ5iAj60JgMh5Me68lbXNtrADb1JQKAW
D7MOI/l+TA2zROEErcbzNj9CEXmnuchAFJglVhbWMjGNTdRSSEu2VYawDARGLHt8veQ2n/zmyyz1
yQJlKjVe8Qj9iIh3dNQdpb5+aggKZ4sSy3qU86t2J3MCxbdprpYHwMyUV4jurTeM8ziR7Vlqu5wg
9iiw85JOmsqr2PkOWJBO2cVYw0S5GJ2zbg48qIbVPVJyeMt/deOAqpeAl6Et5J3RhKQkwfS5KHF1
6XmAia3RgOfD0XRaLi+Ohe7gMaQaQHbMbzXShnrkKP/U7r9PElrBdQZe67SbuxqfzgVp6p7HGj0l
FwBX/MEfafGnsTTMl9oMinDeVxG+1al6ayqCdnWMbT8cYlbetneaM9tRYmMgWniZn3shWt/hURoT
cGwKm4ed47S+oPoSMv7iOxGNHJaPGhslCroHQyIx/vu5ggcbolYxBl50GEBU0AbZRIqb6TGVTi/7
h7dxNeI2tL1mAC0FSaEFXeDj0IehTV0PKK8U4AMn/Ox4Cyj9vv//tYoOto4sWg3TsfAO7YDddsWP
GGIMWHg6D7TD/iZSFiWh5YaI11eU9qJVVhnJ9OG3kaRGsOTZ19Vst5CiDMZIfulHtjgJMQtT17JK
UsZSbSuzgfTlZMFiiXDm1KBGZkSrK10OR+pI4vMuAc5EuOCO1Oj3nYhmPE8gGRwgm7sWnFY2DCBu
D9vC0/zvy2eF5Z+pBEm+qve/6YNGFgrr75v6i0nk8ye0PmLTHvgN/F1Df/YnAMmtzEn9rejYrDXd
ZHEKTlMBMwt96tsAsvbvv57t1z8+AvdjYRBG0qXsWrFA7MrwPYj8NbRUuJLH3UbjjiQysgNcxovQ
dJcUN5cRjEVgJq0qQ3BTEYigAfZI1vaHUQyZBEtSovhMG7NPAbvw2CzUY9jWKsGf+2j4xI8WDvyE
3oTyZ3vkgp6uqxLfigXlHVI35WXYGhbIx6glQwsYqfti2th6HiM/t0Pn+xHdjVonVtn/dS3Kavx8
H1py+8uPMv223o2htvxCD+w+SgaSkOKjK19q5JDBznFmxiGCvj/9oIK0N20JyQQqJLNNbFqpdvht
sfJnK4l3Nv9WS7BnGE5jSdH+9HACIm32ogScEkOyX0HXeeBAenKAiSAH351NUJk9IQ/GyR16CXMd
qHJVk2i9Fs4wTZPnLd3F4XiP2f05l+PGHDtY//7Hkb4DEGvoUeHxNdmw
`protect end_protected
