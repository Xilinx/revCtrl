`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12896)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9TaBM/i2ZgCPEH+TSdpehCfiyRo
8iKS9ghH4ejmyvQ0cRxfj/4wEwjVfzJIVUq3M98XHpgzdzbp709gnnYBhuB4Uk+O2caXlcGdrgxv
2tM4rvseQ7XUCDkVxwvYSwkwavaukRHgEEpzgRnn0cQlgKtIxFT3zaVGPeeAeiD3YfMMANXHW9Nr
+/2SapGPwwJUGV/gH7UiOMkc5CnKwWkYJjKizXOH3f4J+tXM39Jw0/48qFmr+Vk3qXCsHW9fwEaT
YXa0Nn/WUlC4d+ZKiP8gX11rEHVTBfku3aMFBgeyOAhpCMwbUyUU12l8T4vauddhEIXiWIh/7jpO
dDJlE1K7kV3reVFr+K4GT+Fk/GzkPj+OeOhN6giGuPdJkQi9/GYlqn5g88GrhrT3DSFbDDtTFNnt
HVLVOdhPikh/4DXFEtPl78TA3VJFYX5oSoGizJrO7ZQ7iS+Toqo58ivFhfEiu75nHkJ7V5qTTyBo
IlVJM+aJx67At+ouf2L3MDm7j6NouIm/VM4RqjuRKlQmTeNVXOPd1MrIlaJmhHi/1I1Hw0DWiwaX
6aOez7jPK3uMCS4Gt1mkLIEm+zCfZ7LRi6Oy9hXzZIfmvemYiyVbq8U3f1+jP6fDydnkiOEW4CKU
fLNrOnTLfabYQ6WKbGpWoPzfj/sWcoMsoBaLf280UZ/Ko97KQNCK2trD9f1OmXPeQO4QenD0EA/+
M6++TqtZYeKGn1UvyYHucVDO2rKxEJlkCmO3wa6aGTgUFszsto5gpRIrubwlb8UpL+gfu/sPIq3A
/MFz4nKPS07G9In0FAW3+5RT1fp2nYju69MSQeT2z97DBO3vOh3EUM+fgi2qLFxoxZLT/b2ShqI1
ofh87oTFX4bXQTp8VsWMWhmAqgmRyTrLS+VVv8bjP/KKmezC09TxBR9sNaDOfb6dI96HqmW/dZQ8
IGj6nVm7+lGrNDCAnUQ7LTB5K04GWatD5Ge7NjMB7egHisSKsegDoXp2oe1VurVBEp80H6MDAO46
ZObqc2rQAd0wB1PQCpRVJUabqV87GXJ+62/GsvK46UmXIGDAksKf9p6jKplajMRNC/hn8MN4tffL
/DVV0ntK3M4o+nFMWlIafCmoLsxv2YLensPp+oBk+p2hpXUkEKXhKoBYeLRzXWSPDLNMId7C7wYT
HelbMOXZO9oDXK/JqkMTDCv6QXvBtWsor0kZ4PlHXWtzNc6VmNmMrhuXNf2hlu2mwTkPqlKuTgzk
YKGfrAmFwH6JgqIKjxFUD8/1APREgveWYU1RRLUnUjwWtqZK/EtdfuT+B3Eec7jigbHMxWPXWpBn
pgTCJEvviy00jMZabACBu95VcGvb+TsdSn61RW+WG6J6BrZsnXOAgBrG/Lno4F1XspOQcbxOWiu1
8AtDySErEAFL34SBiJs+N1ChVAh04I8aHi+YXxkNc5ndVWPsQfcbAAZAfbZIGW0vsrBGAjT1659u
h6lgG0Ei24OrrLo8J4tQHuQdToX8crKRjkbqdZaPP0b85xIGIs90PnoPRx55ZZqsmVrjAK5JljZY
kWJGMfGhVN9KFQn6KmVUuDGLTiP5SAseEQpQ6YefV005ZtxGipeyXIbcWDRRSCswQWx+bYSpI57t
Ku/EssrDfZZJPxDEXE/Ctu6ttyT/U1Q9VDFP/LmHEBH6cuM3weBZW87rAYJOMz06P8j+cH3jGxs4
LPUbZNrnbCunn6/K1zbgtUmy1l0DCegEKWS0bCht4zkNHjBkXBJWG5M+ORxG1PEi8SVvfNMafMGN
/DK6Mi8I3tIyCn223f5SRfXUOd0PbgYxsPNSgRnHyvyfVkYYVsz2g/zbshxwwjw5Zqe2291ARsEK
czvTORVx14LLsGh4Tdszbo6bAEWDxQ7cZf+PPt0W66o3Ea76clFFegCzA1XwrhiCOqGbZuBu7OZk
EVIPnKqFZENFq3yc4QtW5Kc9qC/GFSz6LiGzv5CCwNn2PB6urb+L5P27bup0t+N/BKctVzfdAkiO
7ytSqSDPTE/wXe13H8hACx0EjZJsDpMULOoQ9sJXQLSwTG3hibrNoJ0s/t3Q91IXLiPW8vdCwEfE
VhMQcFzZ5A7Zf7YKXthMdv0fp2ciOMUJsqUip9hO9M0pu6Go6k6FeGOvpP4Lf7TO+10tXf5MHBib
XWgFX41CLzfU2PoENr8lVYZJPCykDLCSAYokyLL7EFFgzF46Hpa0SoNARp1KPO2OJ6niZwvovNoT
LUWLItI46tlfMNOmm+mpBlhhYmEUUYWxFmXB0P8eglNlX9A5LJpRdXzqvlhyFlXm4BXhDyNQg91f
gyoaRAlimDFOprHw05sqppIjmwNld0aR00hJ+K62ZxsISu9c4K+dUtzoW98CqW/mOqjTuu43QQUn
tKc2fTOv90CZwJTAhdVAkMyJ0LtC1x+GsNPvV2i+ELqn+pL6n4ruHVOACwHesrpjE4129EAn2pev
YyleIJQEpcLrg431cGfnKeuETB5NgYhEXujg0NWMhbEtEEiGYPzsZyeaPgWL5kgMHBvBakjTgTHX
y1QO8MHF9UbGqs81wah/+WEe8JV88IBnZ25NnG2okKDm1Ws3FRCGFnjEBx5uYEiDRZuo6nWxbtC5
gWav0+cX66FwqiBve1zTmAM3sHSGhQHn6btmUmD1pfNdvqbATGMD59U3woqC7YmyyJQd9pKXjcSe
Agn5oplulUijcN/Rr9TFbNcYNKlP41LrQCpeXCxgAQdXuXDmtdP44oO9t3NwGtld65i6yVr32fXp
De4FweFhfm5aSvLvJ3F849KrxW63Ba8tZmsiNb5yEx+nUO9rNy+YKiUnYlKcKeYPQgcMwpt12bci
oGmeZW4YvIoJEA0BCKIlg6kk311GFL0eZkby62uP8FGQehiGndtBPma71U7p5RkUpKr7y2eD7cnm
iaQ0PmkH0dF4/rgQM0lEoSjQlALGFIRIbZq7x08Cet0xHvTHNbZpSfNh0GWrMWiCju7ibCSRiHvp
c5q6QqOu8Qn3rbqvhzVAtZP/Wrv6KWsJSegNQn2jocO1CYCLI4HddRDOspj0Aq1GCAMhLLSTGBLq
b5jzWcecbL/HWknMU/SuxuDTDWflog/u88EmK+SVdSy+lRQmMNFhChORklBJBnPEluLs3NSnOHB6
+XKI1cfNQONMCwf5Ia3E3wNegLBqj8h/qWIMnlnOk7szvAk1hPcAZQlccuxRYlRGIwRuf2a8wxNR
YGJIYOyoJtldBsKkZH0lW/4rdNR4xvd7Vlvgux9uzhs7OR+svB1Jg+0PruJHnzH/fBNulQb6ye4/
NTI54KRZ1Ve4lLrk/W30R9WNq4wWFrQenwS9SvmWvo+RAi4UIhcjC84h/QtHkUGnp5lROPwxq+hL
FqrtO9H9h8IPPjuhMTpgGEJ+4x9j8jRAOLVuIWLvNp735hwd98gMOPSNKsnK/4vhBpZ4ChSnjP7P
EH1qeAbRl75iYjstlbefpEqXrb7Zx34N49uVJ/lumRYqeXOFvX69A+dYk1IKYzGSVi04Es9638Sx
vT3OPgWh1mxvjiKJnIhGXcIAkzJhQ7YOEthggwrKlX3dkzyVMiLUymTknUbcrvsTVMmXS/dicvF4
165+55hxOWC8+WkXRVipz6A1RNCz3ggGsjsa1KGNfcmdT2F6FVeVWX7osHZuMLmUe6lVOKVn0988
j2E17Jk3eDLxq+NAqAdFTyhWymQqz4gudAckOVroa0cEKPco1OM2uag3hGwrnex3qzvssiB/5dtg
V8/PcFWo9sj3p0kLg6rhSmpur+5IAnG6WKcICg3CF+5aQiu/AB5tpvI/6wTJzMIWbt/XWuNU2535
6Tm3+82YP+MgrEp2gZ2vd+BJAzW2saSz4DZ2OjeRDFFrnd6SQ+UX8w+oXaVG+s/oUbDVs9qMkjOo
rfqnIDUye0hGkxdEfF4VYvRlsLY/sUKgZCTkwfPZazXZSRDRaCpN2Q3ywCLdJvzMTdjug9SKe0v5
Mh8uE2LV+dphfbTHu9PlH7JPTT8ElN/stsvaGVqQGni2wzdfS+PrTBV+qxfB8Cn/ehgIAcnwASlL
oyEp/A25yC8uoaqUON9HZ+Jce8zbvxj4FWzxAsGaOEjVfbjyP6S/hZqBUBBkb4d2tfDdMOUV7xRp
0+xx+XoYR8gfWhodpn6XF6cvksu+yHYAW6AZUU1Qq1RArn834+d+xFxISbezQphhVN4NL6p9x37u
+qxdb8kv0uk6Wb01gt1oT2k3TksFOPXNDbMDLxCs0Y/eIC7t8tN2ao3xdS9jpQ9d7TB6gPV1vjDI
btgbOvPp4HPjWILhQxsx2uRRpxCkA7uD+XzO8okzClmizW+AUe0fmdgIMUq7W9PRoB0rsgKGCfc6
CR9eLt20++RXDgbnMxa0gTUtBijDCal5X+w/LUBk9uOfHM6Hr8nWpnseieJVMX8w+B6VRwrwHR0y
rXr9rrCF6ARtSDjC2W4SuWkkR9r/NuE9KkwCV39RCp8tI7SNKFxJF4ac/bi06D1j7xIB1TkKht08
kLNNvdKBvPfj37Vhh6OHDY1RUmH+WtKI6s4MQ4bfoc2Z8r32mNX9Rh4QfM7Z/xLRNLu09xKqUwZ/
SYPK87iUGa5iDggCxyvCI0ImfHsrjBue05fi3UZb3F8MIaCU+nB8/Rl/XSmVeT8u6BiFMDQYuZnA
Y9BFE+AMjyS6mjhXaRm371lmYMCTK9eaWhhc/au7/rNWQ8fZWBuT2/vxWi0DWxxVOeH5C5aDQ3f1
pcZfAiImsSF6a7QBwDFIe+kE8vgrJrM/3k7RdzZvgBKPl/gqPw9B4z0bfOngDgMRWOi+E4QBelfL
M7ZsKmR5wNUoXaAfx9rL4pkJ/XgYiLAU3Qy+ar2i7lUSC/0V6EmxLGAuAadPtDGUbWmTMEY6Y55g
eN86QPCwzxF2eVUYB9w04VQWRSMOHUYsP/9PqD/T7GRE9M8wJR6ymW/o0hCXXI6JIKiVy78RIuFL
jSSnVilaUV+2h4FojlmgspK/AOMKec6PZwiCe9eJf0rnfwZJsn5/pK+SMDIXk/jUHqw16Zs0STU6
K91ohL+17O9PuXjuLLXOy5Lma4eANa9M7ua/cnDbsdyZVHd50s68npPhmsUhAf4dE1+GyppyEpI2
OV9E++u8XjhzSWgkw/8NYQOejZLLngCEWTPEjDIWhQmoZfvCVfpqr42+HXmN2PMjcTMIiq8dRlP8
MotBFLIFI5EqdMToxL//wa5gaKyDnFz7jswLVIvGzgrQaz4gk7zcTJ4xm77rTIMUzPFSGatOCgQH
8WFl7sI6xtCFnGlT4Es0bymLxr1XZ5HplsgEOLPFGTf+4CW/W90I9LzAxXznqc7FTjermYC0ZZN7
CicquAIB8Yy8sfcmSEgwc5SJmEYux7kPHGGWXIagevzZGolNfxQ6GkWRMf9Tctlq0kS9BkzCP/Vt
qPmZJL2zxpIBn/pszN9QNXyWESVMmBzYH8pv/gCR7OlMFb9eS/Bv0odN8bAjrTYcZ3K6vW2OLwn4
OgjNAICC6nyuVUh9CvOwFdp8XW8EWTlhaPck7sJrsabnV0Zfihz89MI/Id/Cdxy4mcZ3n3sAhLdr
44f1geahWLOM2DXh+wo2ofO+wwzESCww7s/YaFj5rY9S5xXoDxrkBgbML+YzzC4AXfkA1EyRwQB/
VG9uNdYct47SRrg0c6SItfY3NfR7Ow/tOEEuQJ3HmkEkQEXD02z1OhfdTXdgymNgp2VLcoNw8HOC
xRU4bGZ8jhCufisMDbKahyyPlwwIuEmR+iVJwI6XV5JvcTNCyJ9vLSER6XVSkSH2Tm0sHDTVZC6I
FJxT3T7XVZ+OpobE44nFfFH9xjqga6k+moaHAWYimnfR4rnYunZXxcsxrSL/skSBsyc+ztU63mA3
ZywMmwcI3fAJStI4vt03Reowe1DyZXXkZntogTlUVWv7msEqKuHY643bTlc/owUzFc5E9BlEyFzc
bMCAF4BSVZPWkUipMt2L4ufY2rObVhLV38U80pUEJlIXy0PiEpRbvavmvSikEdSm/H0beFNs0PQi
apgmj7QPU6Fh3PUbo1GiLb0rH1h/8mtuxXcLom9Kter2GPChRFLYsoWuP+jBAMMfmKHJvPO8OvCD
EPpwgW8pwEozWMMKPiwGRBFR8h84zJ8Fm0rlbyzM65lPjCKt7y+wQgyyuyeR/qce/lDPHm3JNvVj
+R1llCo3dhKoOGFacsVNFhehfegxmxoqm3jSgFRljD1s2gkmia6kReKBpYsrv+1oS0iOyFODIbec
+mWtAEFj87/frlD+WQqqVz7LXkio8UaFIrCttdS0YQS78fU9M1LMEiVhw6UN7nksBG3e5+f4Fbwp
p9QVUHDbLnphQWbvOe/gtmx8DaXYcIDNQKKKpElJcT76S3bVJ8w0G0cBWAJlP8wpc6dnGeM9Ut0F
FpVct/DLT5tXUIe3F9hlUfv57DhQhFm5ZuPKduCGnwLWoI6n9GwHbwekJaE9tXVlhad/ORddtK/A
YBTQqQRVmH2v/sw/kw55iOMwFod+0Sop52KlkxLtNvk9WWVAQFCHmVbkGbzBd1siSn2+aHTaofgk
CvnL89XFTj1w4HoSZN/Nxwcoy6vB5elsB0rfuIVrUFwFrkGe2/Zwzd/RxefSe2K/g3Zx2tf+o6/y
z4oXov4DVTvDiA9J3sp1omaMGPo6Niu20tje+4PT9vqQTUmNolD/lrm+axnC2HlWRcr+0HjJemSB
C17WLjJCN6NGFbgJTsxfhTUa9Iib9BCbIxIreuXLCUlK7i30k85lSstWPQnlnbmuGODO5pjNSehd
Chch8qZfXT946pbicNrDo2r3G57lM/nEi9ZnUSUzpQmrNi2HaScPsmlSFsbF5N91nAtCp4fRtinb
IN6ynonSEKQXuu7GjkQKUkCfER1+vrspJLr/11FY7mgiPQDJ92NnbvYh/qJpna5FKwjMxBAyAYa4
zpYlq+WSfndS2CUs79kEbCCAPORHGCDAzdfoBldOOLufxJmyQvUPRnJGwCh01sZMyKBRU1zRxkBi
hI5KoVfcAEwAqf9nPLUoCGpvJ+hOGvQJvbgY4V2SQKlrIJsXwbMfBlQlsBBMDFJ3bKfz06Oilt7m
w3IK/hYQCuzp1tDSD3P9b7XRv4fvZrSvwej6i2/2T07SI0NrX150ZW8Gs+rYE2OmrXMebZ9SL34r
/Iw805bYUxwyMb8QGMt0EutKsSMp3tGdcyHxcf0KzcvnlqJVrycE+x2HMt+df5AzG71sYqiVV5OY
sL9pjxF0UqrpuEdJoD14WqPzlyaak481ch1k82NZAwiP9zb1hxjL3TSNbb5TKyVyMVghyEz7KO2I
ci9A8eZJx6iaMw9jFH3ADZkqlPIbBxqmnZvpTBGspsvxktDJSzTge8N31dtjZWFdLrE89jaJBUxA
N2r9fIk+UxyxluCJN09rup1An8ay30aybwhY45ot4qE93kqmXAzNwShKp1vYVBSI8TT9hxp7aWhu
sE/g+eYvK9EEcICaqQoxWdREhP8IjjbTgrbSilT4PwrG/z8VYORLMZ9EsL5GbNYmgFPFBXIoNZSZ
Eq0gF1A3Cyv2Lbv4ZMCZftQ24p9jDEwGTajP215JEW6XLSiZ/u8+KUUAeFt268lMTM0NJ03Irl2K
yAQoVYV0CltO9+1ZEIyw0RGdvN4n15PA+U8xA4yAo0yObLu+kUxDqWS72Twj1s4OgixhRhi1DH4P
Eae0k3PzBVUHgu+oaRK2prXtxiiIyaPYvo7iv2R8fB4p6C/HGXAiqYsxixH9Oe+IaLGmwIX9Er71
O1oEL1f9i5qJVgwc6X9Li/c2Qpy/X446232mKDYJ2fcDUjrEbunHjUi64Nl8649PRDVNfo0Ewm5K
554Kd9fhpns/ouGlFgZKdu3ScS2qOhNMGuxYNhp1MwtV9oJXrnxHzrQWsZW3xfz0DKzSNEQPe90F
dT5eRsrKzNW5qaHp/FRraVxqFTp5/ZGvFd3uMN67UBkTl2X5CkTJooXsjRl7e5V8F0iY25MC1L0K
VidM5GOJhN2QSbQGCbstft6i9WTLQ8/ZA7aTinayQ8hc/JkGODfa2Q7RoLD/Nwr3zY5E0GgV6ZNI
t6PafwU6Ktl99IIoj1dmteJh1Bbi69fWyE5wUySsICUTL7VtA+JXE6Cg48wQ4sT+hbBOsTQlmVpz
NyDsCEaPkzQCGKjJmF9326Qq9PBy1pcZycWWuqYrULZUceDaX9g9i7bMVe0XclHbh80R+OH17v1Y
GITJemV7DTJW670TiIoJykaV88kN/vQs8jUS/9+3uGeZipQjCz5M8Vnf+llHsKIKzQIIwASZcbSt
FQNiJHvgmS+RiVbbPgBrAc0x5qGKQ6sPUobCZsXbuZCJHEpwimVkIT/xQ2Ff2nTAR6flb1zzAyVW
57FT1XsB+fo3YfAzLHKUutIlgFCUnMBodO2Of3T4UraWOFFEtJuesfjEoOQBZLAGGDM8DzAJ2Pi6
c7v8hXgr7r7Ft8nmvnLedyD+h85oBHjxf0LAUTmfXwwlFT3l+P/q3kfBjRJ+3vhNGcQtRivV16AU
8CGQmZb6ApmcFs7Nab7/3ARap+t9KZ4oHutbtuc+J2PlKeD9GP2b818AEKin4UIp10eXmoq36ax4
3HIXKRSdKNJWJSkoMqInZ+0FoBxYnMoWgHRa/skUaKEum2+zq8SRfv6L2IaUEwB0vjxSz2llBvVz
mpmyOvM4Fw9QzSEGpPHvjPe9wxZz080tKGjfp+oLa6A1eMCP9QMm47dINwjknP1mdWuoK+knL+z0
oe+oG+Bh9ULFgpyvOx32dS3oz7YOZgZJHPlMvVFnKL3yCiMs/Dcu9VmTaoy7Z/pskkrP89NbzU06
zTQOfGxILxIOSLn3yzKM1vzjPJeAW8GuhGA1qtQY5nRQMU06JZGvI6rPrXQC3IrJThCU+VlqN+BP
owzN+nhOD5cNJ31l6FIvocyFKWM1huM6XqxQJbfTgBGV68DqL733PhO+AraEuabgObeo6WOfqnQ7
BsDLcMMCARcvTiqxXiqV4NKgZM7LzSOW/pAzlNWg6G3YM2pB7kdYr4thrWpuoNEt7CXDNZldxCtg
9s/hyWcOFXcX23ph1X6hOIZGr+a3ItArzj01QiazMFjDfv7HwaVSCcSZwDBJQfBCWPU8HP3Ge2lH
mzUJ9qYVpb7f6hLDkiK6keuZvx+xybBTpP3EIiPCwySAnEAygmFqIqyKA630Avl1izbGZJINuQNB
teSFnoIWJOkcVoafrY9kb1by7JuU8aabhZNLgmBgaEBA4pf6FLuaaRhpJPGleQNjhqjSx8uRyWf4
kntlMj6CNqb8H79KJ9qriwkygMTEQKlQCnFR7mbP0S8uvTYfEkrboilrSvwHfrIfsPSl1Tsr6j/W
IXjXhklheGUAaA5ZPHp7Ya4ixiunIlGlzWXUKQVGafZfX5+h8AMzSklHsvzPzcrSuxSu/JlCZFjD
P6T4ra9P51+Xi4z9rIkcVZwtwzeSCz8uO+qw4l2PGcmk11PTFQ5tSrWydarpTv3balcHRU637kTe
NaE96myu051XuKRsRNIg2+MuBQWWTrhlA5r4w+DD6z+4gpi2IJzF9z9IFDk2bQeXQxP569kCG8Dc
uKHiXP6MjYmcqjhTduauyQRU2FhX1QRM3yLz6Ww8Cu84ABKx0pJnTBV74uhGjt7GYxpNfVc6lMZI
qMocZ15WeG7o47O1BCM9P9DcdlslklAUKYgrCZ4rFznk5m74jdCBazcNQao5L4UCKaZ17lnp0TvH
XQKHkCjyV3T239743HQP5uCZLgQQv5ZAvdA9snwlu2hRHoJdCK/x7UPGxr2Go7K8pLS2PDAfnF9F
vtFYbI9pZZiQZbtPB4iTcaTKylaHt0QmOk8DzfUgIzRAz3pwbLAmV18Wt8qkTJ9oJYnfu4VFyFUC
2OyeFDaLyGj9GJJudxwZ9UfNYU7ySvmp871Is9rB47Gw4inr5wdEfAPH4InchXBmWuvNHmrOr2Hi
4JhOyPbFNh6/x5iYV2SdXt+J25zb3oKoAV62eI25E4lyFsdlwlN7yb7rU5jDxCvTeZHMdl9mGHwv
lDO6yRl2NADuYDWYHvhIxN8ELpRQcFoNVi6sGTvTDW/5aTkMZ08oy0AeEmNA05TRMbOECs5HcBI+
vL0GJAk/k0HTU//dDhWCYZknfpwyjbM6fc1RRFI5Ka9vjuvVailKRGIV7aiQXpyCclBe8462AKSk
SZnrZxZppUTRhZCaC1A7gNr+9WvnxdpQGC9QruoGwurwiv6OihZPg91r/LZdwpzonZpTYV2vM7VJ
Z51Y0YF6PGoqsi21EsLCch25+HOTu5nEzotXFdydZDKqEARpysxYzg4nn4AtCbDhOVGnvWcz1Lt5
EX9RpE+yeQHIgTsLxOa5D2IqY7MjtEhOZoCTPXjCz7BmNc6Zrjg9cQFdPPlh2VZIojEQPSIDegD8
40/H706hZNBMK7yh3TudgkMJQIwOERT3STTZD+G0m1H8GjZl3lXfyvXtIRf6iQ8fY2ESdxIWU8D7
4fMAScn53Z6F6qrApZ6heXaoDMsAPMCfU4ooApt6K6rl0NMDV7bNbqNaDhMKhOITgjcaLhiOz91E
eLBu0y40F6YVKT9JGQQs0l4N+TWZALVPag/099h1X4avGGOJZUJ+FufPLlEM4YVKjMXCkkBNTaks
3Rl0UlgHK2oIp5mdnu2NDhz2pHjr3yxGPoJv3xjwKZkjvcuKeIIrW3TQl3/qGbY86PAsz6N/xDrB
U2lcArRCwwI6B7kiExK05mGFkO/xWBzXrCpIX84M8MPn98MUFSLH0C4TFtCVwfxuWVChQnlKeWo0
UZEOIohD59zIZDAWU+KFHZFTS0/9sF/OrHLydR+VngPiToDwNV0AbhWKKMuqp2rZK8ucHLyj9nb5
mTFDTyKImXxXaYn5m2yDZs/Fxfh0DzlnkFGOdRCN0MsMG7c9gRD65MQowsLslhMw6h+Iv3P72ka6
ogA0QWOxFiezY09i8P5uXkIogwVEan/qxSKnel8iQd+dTiJu5GocqwYB4vPQLq66coJZK7uONIOT
mncW0L51GorRsk0L4c6frlmyZnifyEJlKJSMA1VcOT7Q7MaOQdxCheOQQ8boDj0OdTOwXu4SK/3e
RSURO1Lhw4HLVGK32nXZkzvpUlVlDwdynSfRRaQE5f2gz5Iq8aSRug3obIRIgNNxzhbh3F0oJUZ6
OIw4JtTQF7fSUhyIofJkVbZ+xTZfqwpRYtzfJXRSnLhhUcYXrTloHvYNsz1MiWG8s8GPJ1XAST/X
Tf3fhva3OgEzvWhiRlx4VO8ulO14XN4s7ecg6MEHAMRjCzZx2YfY/LiPUYoAeqQ1vRTxUlBdFJQF
NkkuMzF2TH7gjVD4CxHr4H73GTuSg2C7VILSL666mh6Wp46sUrsVyhQPxzJxLkgydzBEmqW9km6F
lg4erS/VOwG0erbi4IxXPSg7OjOC79a50cs/CpRYnTBpqKYejPDQpwfoJtv3tHlff5/zVzHfTMSb
ML0hfRWqO/6crI4ZT5HMa3z7Kv1dGYNyVJHyMYhP7tas5VAPf1w2uESqLd++1+fr+id6V5HCO6iY
CUf1GSwAzDGzUYtrsemqXGUnTJrNqrSHPA1IcBIfwXfuB76q0SWQZ3N7Il5I9pAF3/R8N11lv58q
X6PE9RmoxyLt/EpUBqHeYlhvi73q7qDyXNA3/ooUvikNJhdMLecsEJmeZCrbcDUHM7tEfFkO82g8
tQ0tErH0NNQddBSFGACvg3AeWY9erbgQMmo6ZT+N1ruW7lJnv1ccRz5iA5MTuhqr3PU5g4iEsVom
VekF/UoVF1j6ELzIrcOh4od7TtE23y9ldXt/sr0mTROhtsqCG6K2DrWiPzkggDQiLim9NS/fh8Kd
5Vz3IlAyLHrf/1tvKr4sn6/UQeQimn+/65KcD2BQSjovXDFOAPAD6V2H2n8ODhmqgKEDVd1CsWup
lLbesUnhTfoKRUohNGfdT+5JkqaxNi9WY0l2TICttqfkRuaDgLD4Rae4KrIAj4ZoAnfXP77AKp+D
mviK/8JUaJHu7PAYQ33DhuOmdr9V31s1uwJb7o1DLvKqVAyCeyX/XbZgJgjiSE0P5bzQV9cAvBjc
mzD/7sjVP3p1yO4OV1/L48M4wMF88sBQXvFOmOqSQLgAlgNRFYkFINZpo1eyWWnr+P4q/L9hd+jZ
pXj3LEoN8ZJlAu/gTGj2bHxyk8NHWvLzZQYMuNDpDIdQidGMeY3wDa01dAiHAqaWuC42tqsPMJ87
PTNfA0Gl953DqGvqJ6zVZV1nJN0QZ7p+0TpmIiOtEiaaaMz/xItuLI/f0Zs4h2YXrN/LMwV0KdCl
269Hm0YBtT8WOv2nY984N8WlGmBddWKigrVBQmjA5zzG+KgzH9HeL+w89JpR6yKeovteuf9JrX9q
l1J2aebBkEQ5MFRCqO19Dchj4S5imG/g+FE+Ih7X47kXIRKzOw31IsCAY64gliDzr4A0D/A8ITb+
qmY2BqnbH+T6LYTntiNmiIHjBJkexPq4Op+SPxf+OzA6jAaTAfEdjjkNemd2kYgGmHlhE4ljp/fV
kaHr0bt80ojA/94PGiufBoLMiiUSsR0++FfIcI4G032CDxG1brQT3Av62mmzez2px9Un+WTsJ/sW
AAjdDNryiSJ9IRdnUdXvtdYly3ZliskuQNPXvwjiQkU6stB3AwaBM0agW67Wv/ya50z+hkq6vXGl
JzH1Px8uA5LarQX6//wyyGPN5Yv7hRmJBeZDGX8ZSAd1QoDLFg1Ljwz2YF8v2wAdt9VaSwNNjK1D
mb85LrI8Aegfd7b2CowxoNWAODoz69jpfP53Q0tfmsyqfhPvsNRIXOR3omuuSZn7yqqgpPvsNUkT
gSBbne4TO9grPB+qDnVEvM8pGoU09saRDH3+qdhrZrEltWpEKSOjh4H3j0VdB2DFkMCuSMSbOou/
pO4moS//JTuBkeSxt2pGOqBnSPmvlnKsTGw8KTvvXu02Gu2PO/Pe8XA3KrcVxPeR3bxe2De+7rza
UFDQwWpDowUh5EuBXAYbaPZBRL42yiJb431g40xkrOc0Un5CLVf9fcRKFezFthF/MLfQyQIyiZE7
3u5oJOt1X2Ktq8kcoO4HsThHxS09wo6/m4y2SWul95Rbox+H2yYEGuYQEO8IjrTd/8e+Lxg4RoP0
CWHk3+Ze/BY0AuCdB5GkPQICuMYHNLPAlcVCH+2FzfRHfzUezD7ANIwGmxwqRdOjANeKzaVOeWck
h2ojcuja4z3D2YtyIUkvPx85tdZbNASpNVulqqZ5CRAPEJmxhwRRYHvfG15m+SDBe2gV2XxY9TVc
k2BzpQzgLtStk5xZaWVP0zReKKDRgF9Ne9YCkRfvqHIe0cBo50QsLrtFO//y1+IlNUhTmZCYtwFH
w9aOkOwuIeYz12X52IT/nEVCVs0AF2+qf/YcqVPwMKprmeqFkmn1BmOequRO3lWy02g9KoWS1wbg
VUihQs+eShKQlydvufdMEImYEP8sGOoQYkujCkT+9XuzSlIYsoWjkswycKAWKtAFi6b3BHewNE4A
IcPpKjFqilNYVGQlZl+7uIz52uiIl3xqIGN2EF6yOg34c2wsOUKgEatXjJ6YTT7NtZ+KMv17Ea+n
YzuC876l+yj94gcO01ltUx3pA8VYJtyDyjj8EiUelKCShZ1TsY6OG+jeSnsdToXYOgN6CIqhfQtC
Nkl0lB3xuySsx4q3Ve0ZaPvdsEG9nchslXuIEYLPCZ+/BfhHBhReahI/welEZSfI01+B1zhyuMtP
WyGHHWCmaPJjlHm7jl+Dt8lrjfSaR/B6ZSxghj6je0C2ItDVpDAQidvbYrxcvofIjZgHFLdx5i7q
Ue2/F0jY4ZqD2q/oE68tdFkrWc6UAJloF7IzYydainUxSnvP7Sr43n+My2cNP/gIC/QjFwxhM2xr
9YyY8Hzn3qQxdkQTd8M=
`protect end_protected
