`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cI66OANCJw8fIIQbdpCG1eUZiUrVUYlTNQ823416CUh5RU0Z0lUSscJg0VdsbyeOG0GIlqnKKDcJ
g+441OyZKQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UgqPJ9i9WiJwgzx9hA1QFTAyJQbYygHQhueZLDtbtfbgNYIe9Vf6qQf08t96mKA1gKActJ7BeV+K
6uNMiJfx/3aUXCSX1zJ6wf3n++OQDmqvxVVq3gnHpb+740+sx3yxZnt+NIQn5YfqgmEXSODHM65H
T6IlCQG0Rk76FUmssyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JffVUoJGoNenA9JkXMLk3KS8XcomfWAzcMGUl6pS4bKWUvYmY13D3pemGWR5ICLizj6/IEASX4qM
MrcOHNOZ78VNNGbrwydnmhep2T8HUJ/34A8F6RlIg3EPqaoJseDBIuA+1YYmvMYUPXWmDmWnG1uq
4OVHNHuSMmViCS9G0XZMw9OZMd079W0WWlGjxgCIsCbTxgr5NySjw/l7QR6gLw2PWlOAIibLSL/6
FYbf9Pq748eBFOa73RMaFJULQdNMNcUKu7XbHElWwAbBAEQETSA5PY/T0Ovuh5VWjxfKceXk9gE2
s16k5nL5jvgzFecQSuS2lSlURIB4qY5hje3ZOg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6n3r5uCHMurGEnMpYNf4UX/MkeElsrXqvd4MQdfthvZDOuXHZxcs4tSf3laM+WPFVbsOKpN2K9r
vOlcg4pO3R/XBxH8buk6fx/j1Txb83yD004eikrbAzhD/XMeJoB+vwnOXVjryL4Tq7ewJGiuFj3j
3aajz5Netn79SPqpagQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ux6EQpdIiEpdxg0F62ecUw7+0Os42ovKYC5a4J5nt6L0NXwWYNruQn6thnH20HG3CkZMjYPVsVdV
6fsAhKiqralBKaBG/Ej9eLWDO0kqJYBDBHDr1KxCmmsfP7tgcSeensV8aAfsf43ITwJDMIO8VHys
LbnRxuW/uncBTBd8BpuuF6FOlCwImGuVwEh0SYaZjLlAA/zvuQGePlYAraOXp22pKz1CICW9YEbL
RHIga+6SQ98q3/eoFGq1j3ZXVJuLYcvW94K/kJlph+VD6UU5Kix62jbW5vyq5E8KMpqmJr9NNRFn
j81j5XKXBOZlfp+VVqMs7Hlviysaj593wan5HQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7200)
`protect data_block
td5QFuuLITbKOtkE3oI0mLzB/U3OEn5lA8+gSvm4NzDgr1xoKZ6KXCYimdZuYcgLb1Oo/1ycim8W
PFfdiPDalf8RhWG8Bm3Uye1fGmokMIeViJJFpudOlf2QwkH2Q9nSjhByWCvm5V/7FzruOcyzJZl8
uis+1q6Ca3nhUQR21H8IcHbv6Xy9XdyKOtDQhDkDGI8SOYvdtcIlVOvSvgg1PlHx6usdcjRT0U4H
P6/B+j6sbCmxYTaRSW+MrSFDCMABIOsqlOFl9PQ33XhNbwlnmFyLe8tBq6nfliNbidO1H1QObdnq
g0XiRy+Q+5bmptOPU4KeuKsY+CyWe+gSZWx7sR9F1KCyGDcBFrT2VBwymoVYyRvI5vxdUB3+YBRz
FmrHBd85+LV5hWGDGsoNeAlxuoCJZ9a4xhimnhmPybEeZIaW/cwOYSsIySVmatyomv9KRqSyFT5x
plbY1EaYl4W9TX+eeoBSNPVHCHbXnHAycjPs2518RrFUO7ZhXGv5vru5yV2qNNGPMw8E64EndejI
xVfqT4IJ72rQGgWyn2yK5gzLwHmyRO9sJ2u1oGUwTfGcAt/+bNQruj/XZjdx+T/pCUTB5g6RI4SW
1sPPoVa62LL4trVxz697RlCg99hexVJwWhjRtX/gBmanEQ8qMJknt6HoxQrVV0sTY0lIbrnMl6Fd
iNzNmxiKPcsuRHsnRlIm6sa3MR4RkV9S6QC/sljwL4YWPvCM1PqQd7GVDHw+CFokz5R9E9d9KN+P
czUx+HZm2tNSEn9q1JxgsiuqQRzitEd3EZc8W24OTiLm6WP6Jt/IodszaPDob+2ut4BOMLOWQcsT
mke/SrxzWJXhU/ZG63YOaoix2pjzVFqyTNFJuxsSppCeZIMHH1z4xtNqQb1st5nkgP9Kh+g6tXWw
dTPI5+X0B7aET0rAOysqiuprTrnSq5kuC3xjTCPygJZzL/dFMqUklhfKPj64S5SdP2wbN80H87FQ
nQnkk5OlJ6zm6p3GXNDYWMSouTrHZOm67mpC3LwWnH7T0/pfAdWmQ4rufIAQi+gM4qD2jOAQ//QG
slBluOWzc7ywEgakNL+S2mJpgHO9klPu/NhaLe5KIxv3JXalj4en7fCcwcRsAY26sRRcw8ggn0J1
1rHBzC7bcBA/rALNhqZOV7URMYD7hxwmmFa4ASbgBu7PHjZ/MoUzKjMIPsBG7pn0qWsR74oGPh/C
/ILnX0iW+p+Ye5XvoDM3T00Lgi+lV5DVYxTbnmGJbu0d6eEvGyNkK+qU9YmXdPPMlZY0HxL54t6P
6Fz8CE6icnAUg6yUsDYYpI6U0Rl+0yfwhoCJT293Q3P39p5QQRmmr/wsehzQGQqgZfnKSqH05QiW
Zr1zvt14CQhz6LRtZNLT/iNVxjEJ5A0ARpeukq4qx5IUV1GF2oDbvb5Cxvze33zpPtExB/f0WlNk
TrfxwFj94kLwqOINtYrmI3fBCvIydCmjQceNYxL62hawYt/MMFneDPu19JcThYBtUygW7mxxpDyY
ePDekjp7wREEwi70Oml5gfLvxk/yq+WqRgRVQlieC5q/Nagn496nauCxj2lLVg35JDEGIDkQplaq
BxgoZ5VE0Vw4Qc+Zw52VPmBMFvuR3rZbqQ4CZHaD/3CgH6X8oz5jJZv89PRafCSDXweVRywMm9bj
/08qvKDQC5KWOg399jpbZeBaEsIM/ncsvwQSb5nFGcayxkRP0/JHeJuSEpVERH5d+6SL2+O4PuCO
qMtp0aGh9IkxX2QrgR0hzoFPlqRGl+n7TtjrOpETrtMtqjyM8RDGUdiIS1ETj9U93xsihAwnkJIM
7xlEfa5lOnu3mwssWqJzQl68UzHUp1Yt4OxCRBj3xFlDi2i1Q5L7nZyFtm4ES6AjMeyTFvmfjj/V
D/F8eqHYGFrOV0noqBXhDekAVJY6Xjl8uZ9x4j/mpRhMbcKP53CcyWOlIxF6Zmh6HUH3i+0qbQaW
GzBm+JE4bvaiVjqxL2sv7rAbM1sZQnqGYfsxhoO1Dplc3IetPgWa9J8V1cRngAYMzD0Bxl3khagb
lh+x+DAV2qrHRqiTcv1nnHCwndNUJ1Zb1qOQD1NiZIhbnoTaRxNTfAHvFFN4SSx98ngPDiUGR94a
qoW6r510ybjzEOKjCzaM1SHBuET4pQmpFperF1r9bNTJnppgQ1Y7u4OZdvVJltmW34qjqyXvntU+
76uXEumAb7N/e7EoVDIve1vRxAQR3UmLXZk1ddFZUNZsc8Vj9Sym55RgPPBGrpAZrMu9ygUiAY70
IF0QXxDihE/zE8A4NqBD7q+9AN4omVWQ01vc6mf/1pfrNyDeJoEijx4NLTfTnNASXUljfneM4OFu
EPlICZPhh4GO/BRJGW2TNZsL7kzpjQ3jcSgAfSLeAVoObqOBJXr/6GtDhfgW2ZRMpG63D0E6xiua
6tk/R81+i3XkJcjC8q9klZk+CpNcUvg0M/pXNPa+Ln9wNwE5KPUgdQK1650y+tyJtWueiwhSwTjc
z2Ds14D6ldjm9YC9TEc/zpzTcljQL3DiVhGhoSx1ANQQEHS9FXO3npq/HJIu41+94xQ2kVPrFuOD
ywzI5iUPmlnOC/CY2itRxgcBnkVZu/9YqBb3DMxbsRWitLFt3+BlPUFc9+49l7I1GbBPE6uK2s0p
uvlgXKC3eP1cVpTIxCBrEnsnazFg89xLaL1xRUnY1K/FNAUCTBJwmbmwOLB+y8FQRtPLpYsjmV/5
8zIVxvRDA1RfD+bp8YndoLwgj952WpxeKv4oQEMKKR4o2krmRLsH1tgGKUajaDUDPb9YYxZe+mGz
M0kMXwiFRakaMLYKVCHfjZtOy/WtCa6y83RBAggXC+tLVJX+TyjlUU8MRnvGGVxfUI2FHF62Lp+o
vzsYaj9tLzIERODhEr4ynD6LNBXmyadshJVfx9v2+Y1+nUGv1q+bIUpoRYwsx7S5vSbsSfvGADjB
E3blsX97LAeWVm6dclgpZQ+MVC7YsQP4mqUlaqrVns1hqZdZZSxBda5HhjBONP8/H6Gl/YyI9XVB
eCyklQ4w1mfkTrbDs2t4OTPveqJQAMAjKIvE7adSJiFT1lkl7nkd3PchIA6nDlb0u5aV04/Yj70W
qzhGLFLd/J/7ggCzSJ+So74/KKcT1QB61boroJbjZhJMGt2Wom/eHlrdtUj5jcje+BKVwcvVo3BN
wm0ouQbVyqdjwNMCKnxeiam/WqGfsBwgUjK34uEZ7xOD9u8vyx4dghvw9Zya2FjM1BaIu8I2TI6a
CT9/NGsraru9RdwhMSN7ceotzQkm6xNlENlV6dv6q3SDnc9yMbSxwpYtSXdWYLJLLuaYTXngQxfi
NrQlNQRf1u+CJNhNToCCjBvGTQjRgGvjj1PHMbriFroBwukNqdTDl3roWYs+MjqbUF7LPoyUPUnT
ag9CKgHo2NGf6yQFx5VQzQXhS0PVbUbzzy2jMKmInJW+PnJYiH5tcn6LzKnRLygxCTWffXyZso0C
cAaO5KrUQuwnV7NcaAToMfLNWKmN+OjLA8cDC5AS7yRkxQKb8muHjF7aPMzbyprlSssoobNphHTz
OUCTsl/ZiLJpmnlmRiL87jgP9FhIMZgtYTPRrFmHQsyhg1oO7NQkm5GykPr0kqsf2px0VD1eLIrd
lSSKgLluAUGFvWz1XqP4Vlu86D3Z3CV1N+DAu/E4VvMW2dFwwleVsNWuAjy6FueO66d9MJ876jFf
+ZiFWI7EkGT9sAa8epuKbrwqXkXHHANqHSJAJUrT7Lets21AiM7HUwn/xK/XMRT9n1lPeY8FsUNr
TSxBIZ95RbDS3BwH+5qTXaQAgsZ3itulKwVcxb31hL91dYkLhbpSINANogSolwHQjX/r+yeuCqQQ
3HiFwhx+D5iBcQ0T6a/LoRCVdD0erOHwYZtPpnERackvHWyXBZWfHoyTsoB3on93qwFrlxqajyeX
FGh5JaRLevkzyvZNHOoFHrsJ+Fvl1v41ou2tyJ5N+yPk9dAFmH74/TtS4KXPSgXgp/QB82uEcg4b
Y+MqAuN+B/KeJuaozQWKBvlr4AIQlu6L3hAudHOdb9CIb8DkB5D/KtKwp17TTd215AIX9DdxcePD
jCS5MONWjn2cq2bRXVjsHAyOAu3ofFWSezgoF7tDXCmazz+lSF18/eAUDwsrNzbOgqPLGdBCX36L
sNs57oNEKEZx6bNzkQMLfT3GnRgWrLDY0dReY5gZS8pJic+o4UDtyIg3frLvjsXcuJZX+HgSiLSH
nrpYHJODwBphQFl6UROn2wVgUow2V5lQJmpFsr11u+61bkxoXiht2O+TILTg/QXAwphRbge97ocC
TQQQQUyuTFGdLC/QecArdgfRlSabyhrCTR9fW84+jFHwjOwAi/HuDME/uabxqg3TEVdVPLAJiJys
QmNuQNT5pJcHTavSXjsO3NnKlSwEN5yXj7zne1APN7t42VbX/0OtfnS7u9XAdiHqQ3VMIfumlQ39
xr/yg3WBEIBYiqnRkSCNhLhvCk3gMCnoGgqdDUpG5VqpvGdZdm4Bv5qXtFtwxb+/rMQhRavxxc+p
9MO/mM26icg/Sf0UtOhDFMYGW+kLeegvJWcDzZrwvgQnOK2ZbdTXOnY3ZcHEUx4k2CTQ9lJozKwZ
rawM59wSZ+a/rjtviVXkB/2OC5rRr72VFEU9vBIBoOMPYanQTW0/gJ6+u5Ly3TC/4EDBm9F8DwyU
oDZkBFZ4KfZzEcMIu6AR1tiwVZ4CgV+QXAmtYzIYCT5Hsl6qLFqJu/9QNqI/2jK9zJXfYaDweZsF
sYltNGFxOGKWIT5wfrBqfbAYnoddJ955oCCScNsQDM8myqBW3h3rRw5cC6CapFRwJIAn3FOAJdKL
XlwmZzpdrJLpG4ECUV6sY5C7BsRGmN4X12/A8Zwe7sX28p7lROLBglkuwQyK8Prx6pE7BgbYsi29
6s7RyhC3LnS92fENt5KZ57M+ykCEjQMpju9lcJm0+NhLcI+Dq/jOmlhKo4XAJNibQgjRnf3k3KJ6
n1i9kNrJxrQf17QJ574ifAvDRxvTnvqVHeiR3bedOlZ5eBPHVBKpA5h4F3x9TgPKdDVtQDsRdq1X
lN/EAtBztS9vgCxwd3z2kO+h2//a5sOvUB+4U53+sEI0UExF1daJ429ODVXBf1WtyVlZF2nxct7d
wyIYr/pDI2ol/feVyNApmw9U3JgxGJqP1Vv1jyfVGecWW9ScYiTCCS9LhMIplQjpKEpWhlnF6P+j
EjitKWwgCxsN+ksiuGoIQYhlT0mla6pwrkeHYgDMeLKlwUNqhHICP9FT3kWDjjOmwcuTeBDspcdw
FJabp4fOz0I8OQobgRNI0meqBEI7ix71GRPNMIQHnaOFIj2T/A6qHxxkg8m91MuvPrpc9Zq9H7kF
nooAet3i7V4PO0/02/4j66W2moCaAnS7BKONuesuIiV1YAiNXuriDnmT+Pa/9tmU4YiSoMThp8i0
DJb6fbU+77Yw+srz3pzus5JRz420IghKN3z/iyz3Cl08CNK4MJqeKN0mZVXa3F39pGThLWHVB8lM
2ID7o7yyCyYkLiFVq0Tybv+e0JZY1h85rJQ1PFN8HkHb99cvzONaeXtMAJ3XSCjUFw6wQO+S/U8/
UK95PWggZfFhVXDLwWnnUmL00acCyFHPYKBqO7BaXZlaqQ3dYMldBxCgZYRzrVcXrJe4Zm1TpVoc
TDZCWOYW+bRa/D0Z7bCZXPcc/wHZBtU0eHrmqOOzmtHrz8maCtn2s1XY0xasUlLZw/RS/UNGVmFk
p7hX161i8noRKoNWfupMxOhOYkKm95lmE+SZLMIx0KaLc/f1nnq7AbyVobbWJ/C2sX6vg3JmUmR9
veJv89TsbwJCARNHGCYgTgr6lH/FbetxcCtx/cG4osDYi3wsTpd+c2YQsg8DKCwxoAQlMPuiS3Zu
VhWK7gT8v/CHa+aiTrGc/icCxVax6LOFKwmtmLS3+7jMeDvG4Rc7fjCGVnsL7UXxw0vLAX//Gjrl
07CALVQnmebb9DlTlEGoc/fzm+w3uzXeZYftKrblvAdt7cOhIGcmTEVdqv88cG2KaJMrCj78UDgX
WsFOlWOksJWd+TR/KqpdehHx34kPmP0LEVaeSGDD1mJ6sYHXdqonQdGSHILbvIITTC4RBfcxYJNY
+w9632bFxHThTETZ46AFvbZc6AMg78JoaDEZ0a4sEWRGpIXr+VK36jlGFtA925jHzWO2sYx0wfIk
esIWrBmJo7ghYoZGPJHLJe2Ui437GRnbonq72mHci7kGgA3EOIIrEDOyIj3LJOUpo9T8MHQjxNxf
eOJMe5YthH/iSo3GvuIWwA0YijlUOR/BA0a9qPYQst4e77z+zaLpT4+topbmVy3j1g/S5krKsiTA
nDgkfs4iDSIZo+5eO85h4CFxOm+7tFCHSn1wUaMw0QCi7ExDLUfq10/z8eHNPO+Z7F1hTJxtzJNz
ktinO2vjQp2rnSikto+ASTLKzX1mXSJh/v4PWygw5LNVd9qa2kQG31NI3PBqgOKvykFTsONEUSdG
6BKDqT1sh/s6EB67RpNZ38EGb3c/tqnHYQnWpof6XNT4x8NiK6oBs1fVG5UhKPOKUbfwlE5+BQ+q
qCPoijZZ3uHPNCniiEg4NuHLRLU5cPhJ3zU+QgOyYxvK82aQfCvracfHa1y4UqrlFA3bYvomDXl4
LPoJeRKg3KIqNRw/XYRLVjn3aw1U4lekIuPVuD3s4V/whzv3sn/qerGDhc0gJ6wA54sW0IyP3v+R
0tESjJwHMjNUGM9u1nicsgE2m0ICwdoETuW3b5xG51wilZNwyoUAj5I96t5zlu0R8kaKgbEjeOUV
M4kTQX+eYlnFCg/5qhgaDs+aAmiXtJQ2dxU+4Ee9q+glvLLY6Nbl92CxHLjiGgc9jTChvwRtXNco
CdFbcB6RlOkyCv8TCs/JYjpxa7f4BH5yJAP0VnrdCN3k8H4WyiXP+Dh5q9NjALr6OR8ZOSN4a+2e
3G6cLQ+zT2PD0KGygepNNWW+RNVGABTMlwV1YMZOmjXIKVHTPkFwOKy81jTVBh5tKaHqcqwPJNFQ
h2xdGTE01jxl2luLgeFOvgPvx48gCfXtBzcVsTxEcCRjw3Pn65qYJjl7jo7Gj+BTnrTNynXLmnzp
lrkbzDif7AAJ37uz+MhiqwcKXhuaLp4GdKPKl74Hu9WQDNa6/EjJWjPZ+iCO1Ly6Mzr1SUrU6e7x
vL+js0QE6D9mo3S5f7hqyznjvygp0RMTwWgCynCOfKbQxLIQpcbE8kZLvqP6XmcKLKZb0MoUTNf9
A63of/t+Y7gJH4WRMnNBWStL1mPnuBReTmnaKoft3A+TaSWMD6uXnGKLaa+d2i6B3yaHsamsyFjx
6ML263UCDk77dzqBicEyi1MOCgcyOzCpfTpy+DvkuxzoB396NjLK18VCH1Q0k3IQQFZP4eghATuw
HR7hZ+2h/YGKVFh5IeQ71HttnDgI6kIgitvliUVMdt1v5WkUzENTqVyV/+hdP4qPRGrjSGXBTWV7
PgM9c4GzzeWTsRUnI1jqLBfjVYu26rze5EJ9qGVLnzw0J1kOtYF0D1EjB4wA0ILoirEfilnf/z+r
ZvM0XSuFl1CnV41XHLKhn6vRltIQ+k3DNaohwyioRNVndUlILjxSqBpLQ8NaW2pIM25glmLJAJUo
YeHLHiJfjEwQw/21XuoIzbTLIIixxg7/waWOkR+v9weeTKPfL46j7MjXfe/eoF2SfRsDl4C+Z6w+
3biwrv28iyVcVxPKQQciib3iOwQRRNFDMXo2pXEwskBPHOE5XBOCZnehr/vVbHPAPz7Vw8V+XuRs
+Z2eY6p9VlbK4cg0zcMvOcjKtohPBCMlra0lSz1DPw3JtOm2XthjtVs44RhjOuu93iuIWRRkJrAV
p459JUK6tA7/XdXYG88z7vEX+ieH/mVSnAhkhjLm58YB93vx/R/LvDOQF5/sZL/y1zTKSJM+q6Vn
sUQ22i0uCETBSDjOpLtJz9LkRK8KicCZCpK4tgVDcrIHM4hLzuEX3X4d7zi1ZpizHYuoKFJ9fSCx
2EIjVS+cCWS0QWZAjIxod3ROHwRmlnsx2afxoC5C2wbzUdH9q5VQRLUCSPhpmcPjMel8tA1LxI6w
imIa5Bco6n6/9/vmJs+Kweqv9nkHeIh5zfQ35Bu63A6AresuE5/UvezYG2EhPQ7l1fpuJikhvEvm
+Urnbt7p/EjBbiUjRotNoVSjRnNFprpxevSIt7+9ZLXlEVTvPSFK2jV2n65VTiLlfekBkVqSKs2h
l6m2j3P5Qge+ozjeUlWg+ppNA20GFm85DZgk2BDwAUtOVyF7XWFDmbPHzAToYEw4tACKxoCSZKAP
3dbOTh8BDKZXGWLRpmgaYY7j9VDwGpBxTX4/BbwdtSng1x6+9KLLqFM0yJEbWidNNXr9HT7TWwP0
nusakDAsggBPPlI/++qdOdPpyMJ+xgMFHBI3jS6US/8u2yTsi/95cE42O1v9PGkHUNTANk8IIxQ/
FK1ifweHVD0T92uJDVhHsHEFzLpTPYAp+pOWRgyhkDmQLseHJRAhyVJaZo7XeCwA3OW+SdvgwZwg
aCYbUeKsLQ+CX+fpDOUODF1wdFzyXpG6UHlKLeTB7NWsU+oDm+PI8QK275lG7cCloPiJx2+nBFlr
cGwY6PkDMl1qGlGSlt1x0eXgoLdNrepLG+ia84DJrg1QfOSJaLBNs2wGIZZZJnr9gN/eWhYbijBQ
+0EFiZLTKODOIhRgb3SyIWvGAKSvq9Jd+znSFxBHqPur8ZgHDEhzxkxHki2XNeyAshXtk14wA7bk
rMYKo726Qejnv1PXtbPxSDOvj4EWTJyJLuwCF6ldP/x0JjTIHQjP1+orG9vqLDiDZplx4H02EYbq
q3+VYvoXRViJsYJ4VRvOU3o8mJpvcQf6YvWIKzX53KGjDegxJoCSOTZorCBFUFhuNewYQ14Hv/AJ
tEGXJ1gQmISFbzD6YAMiIi/3oicihoO3ltK4dwzMJLAExbzt4Xj+ne6RVDHdRYUSCoHQKG6HF0VS
9tj1DcHYC6tB7wHy0pXLiyXZZFxxA6Ne5WKZK6QRPmplxXi65vHEngbbE9UzrAVpIjJzA60oOKfq
bgwYXq6eHKM2Rm7G/VtjYwfXsXBQTxQ39YkqGScuJYtFcJmYspygKc5Wz0zk5ZBzoUyzKqQgHDpp
ZP7KKOqgdKpRyybd+zk6LRYXdqHzBOgq0NGblrJzakTOisogLGuSoUXrpkuidOwNyET2LLmb61Cq
vXkagz5/mdQH7brZ3zBZZYziBbnRzTFZ16mZ/5KOnxOcNKsKGDCmCMj9mtEU6muHLMhXCsZYLUmN
1U1gh5R9hjxCYEDTfc78lFe+YDxEU0rzMlLdD9YpCMeXvw+INMmJjC00nC8QVFTsnkpjlTGPtERs
zYngrvBX3PoJMPddvaRsZQleNBGnoJ1sBTmg711LtkOuvdDTzKQa8JDIdhrsawJtiKXc59ZzSK2F
DU/DP7uh177wHxXUcjLttWcB8kRk+3CGTbzNaK/kXlyKjuO0hQc0RPd4sBc1U4TepEE1oexFIakO
Aslkm/d0t2nygIIolpwMwbx/
`protect end_protected
