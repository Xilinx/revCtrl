`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 318176)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbB/zJnlY9bLi0AUFrGn2gHL2x2kzl
0IsX27FVgcMWfMmKRIhoOf0LEEz3jR3k6cGTfmwrwivKTB5aAsPR5ZFX/Px/CzYUDlXcU0vgErYW
q4eUuhRuLmTUD7N0cRxvpabx6zAP9Uq3dZuxysUIFTTxIePtlg6Y/tWzX5azEKUAwpEmR8vOpBU/
bIDKzLdfTb9gN9mEpHLZLDMeuLMgfkHNrbJgrbjKcDoF8Q+6fKCMltlL/uFnWB64rVqE8zRRHSaw
/LfRvNBik4B0bHadCtpBFTHpS9Kr+AIAbDdb5dKy+4XiqmEHQd+U3yTmo8dNbnGJTI3T5zUIV3Fe
JLTfZ3nppg7d7hV7HAUXw6pQrhFJ8a+VoGeKmeE7SjWS4NOZjDc6XmZoJzbidVdi/Edt0WY2KGHJ
A1Gux8B+5EqHqjqlXjfaJNKUve6pdb9JpmG8LYaBbD1H2KTZAxLqNqm23ohV5pPVn2uKCpYipE+L
tCjyv0EI3hgS7WrQE660Uw3WPB9dXeJOv768gAMh2kxyL4EPQ++0TPaFDNaLc4uDphsRVqQ0Nw77
w/bNz8HACwtF6hMTba5UmMnU+OyGbbuhszlQy3wVevV0N2pldcsHywa8uAyKjqtkJpE5TDL/ABjp
rI5BGSiG+JQESGCbhXs34fANyg10g2JB4DwGiQhFr3e4zhNVRvUBZE5bVYu4Ll+HsRpVyp/JpXih
+wBEAlQoQLQnfMzTNW1Q8daog6U1ardqCx4LxzUExu9RsMGOxalAAf7NsicLO86YjpbFOsAP/Ofn
ntOlATQUO+pgh8iGZHOwv+8rXLsmV2EFyt8vzLMLn+azdfqb+BBkC00yI0WOmfZwkvMkk85PpcfP
mPA5bSC7n9BYlJToR/xnkSMADVtxPST/jQDjkH/AAWDkaxF1aBsv7WGksKVln624124O2Y2SNDEp
FphRZcmfaAGtg3UWohn8SC3/wt85hYDOtvaA53sGR9bHoSZo8C9q4Xm18MPAe0Rt8YIqT0KrBF58
WB3hSs5kyibn1FjRLDv670LbyYIGzjBftFyS6VZXAWD5rSpmFqj8ZvYsDL9KIAS3m4V13zsY2T+N
Ze2u5wyo34K9Lo0JIqj6kl8OWLuLDT88o0qeSwqY7NMbpedj7vtUlTxE3t6Wj8GGApO0Cp3BRTKC
qyR1W4hbdLbEIvw0rbRUu8XT9EwQa8sCEm0nM+G2dbkXUd5iQGLFnHdbftxQ2fSJrN8pll2CGRnR
oFcGrBmTkzh59T1lJ3timc9jGJEarM9LpA4F0dkR95NgrRjfUEzeapJbP2OYAoIBBaU5o4fMUebj
gIadpK3AoH3ZiH6aPcDiI5EoJBkQtzYdSo662T0Gj56yw5I+ztl6435b7H1pWnQPsB9vfwAfL/Bk
8O5yL/GKxMbs1ZPveLGW9L0/ndNsDPPofDmxsunw7KOIzTjcANjdwCH+2AJclYt0ZFHG7FuL/Kd+
ePHdwhmvmuC6MyC7Avxu2I0zWwgCsOYV3chN95WA/G5XLwsm4O9BXyLs7SnsneaOoFzsw69y25wk
h5WfE6LVZyV1mk0RU2ojE7oJL5LPYHpW9O21AAbfFkGuSk1+blf4HYsIfwH3EZBJg3QaqBLj/afB
y/2EfKQ1W30aDiC6fdv7HXdVJAcvUZqHKkX2R2SrwhqsuerXW5D+J6QjKhIHz0ONPAsKCp7JR1+d
gZ+RB6vvilc04ibZK2g71mJCPnDTqr9ReJeoSYL3gIHqmwW8fjQCqfcsmXx6YkzDapBNGNdI4w42
iVpVADm61xiIEwsGP4vrChnhdznF5jFy00D9NAQUXrY8Hj4KMXU+rBFHpU8jYrt4YdRcf+5q2ev8
DI1xw7ACpv6gQ8O4FXiR7jID4H5c0kL+dTuRTpac/MluFBJQ8f/HDIUrLsXNg5pktOnQjSPaKoTK
A4PMdF/VcWX5+f6PZE1dB2E7v1i20RXpHFMRM+lvwqz0kj7aiP+6HefS80qUqj5UXOnPJY0cQPBk
E9YFIrJC6e05DHLCGgnWOoJG7ZuxoZ83LdgdXNBDMVxqPQaAIc+PBJUX0hce7uytQ54oFhf8vfIH
Zxd++FX6VolnMdHVz9j9Aby3mrNYnGpsXcoE/LYNOq1LQ7NBB2ZHNkO7NgdkDTNqwXrlAGHqGliy
mmL5nFMx5tDpvRpqy7dmyrs7y1F78zD5fWMixYkHVJqSgJ4v/CU5rDPi+2GbJDGyRAePoicwERP9
XNxliRNx2zwjZkLElaJkjuWdyt6ovwR7RxNncY4m03vCKfdd+0yRUtRdT/P5Bjsdo53mdoTC+Yw9
bmvHdnFqKTkGKz1ILR86YUYNrttgsQVqNi5nwcApKoP29aN8reutGZpHYR0ou6vJEEgrHAqAfVA3
Kla5o3c6cz49ijc0sVgbEIS3b63kpy0aReQY5dl2LRBMYnw4/MAHMbVvyE3OUFqhTv6PfTwCt5KN
SxzIKMHQ3v3NwWrrY0De5l/usOG8bNOqb9j1AEasyWd0rS2rTU85mi4bNLYx36JN7AfXT5x/0ljN
s4/1r14FeDPicGihTsTp0wRQY3DFQMogdHirsfeb4LG8Q4XN+mZi/r4zd0EveJiJLvyKrIQjheBA
MdWsu7w+WHoZM0freAwS+vbUNC+hsEjfElGIeyE/rDIJjj/rhjuFFP6zCSr2Y6goAd79WraBEKoi
JA6JIwCMZ5kc7ljgp8wAlhADpw2NEyeQgx1A7MglBuEciIn1gjAQbMa2JH4qMz0eFFgCpu/rgof7
lxOSrBvzP8IMiBSLxJnxgDNpYPgpc+nVBNSxl71DUEf7EH6wU0RDsUq/oaZCWep5zEkd+i7wCLZ9
2s+SyRoKek1W6zsXhjUPdBx6P/fdlo405c/uPIGg+CMDGzB4aIEj3v7S6r70/UoMSB6UX84go7KB
DPe5BXUwzCu9dHl1p/l1fas9RjtNBjeO3egjAYYokf9fgNtI9o5eWU0j3GjRq0yfMheopwHyqsv8
yirRu2yNaGkpXdBlD4sPT1XtdU7B1YKdXNSAeBMEZ2wZXwEJTAEv2KHFhj4DLlugHlxW0hVflh+q
a7AG5spX0mxAH36hJ6RHCy/quTClOtFHL09fpsEG41U7iuLE8Z6T9ssd/E52vbHQWsEZUwaIQ0hs
2/CbOStkhL7HD2ThQ3aY7RzXgA57yLOOYYt4nw3B1y/1zm3eJBxiDerulNY04KtW9uZZKqwk7ymH
Qh2gh1lMevm7uUnUh/ovYWO3Z+1QB845sDzRZcGHzwE8rJqoRDEyCcYi2Yv8HjyPCuEMcrl3aPmg
vpeUrODb/d8I1kmW7OgYCKyzbvk90oORbNgReglnNbHlA291H31LP/8baMkpZXK3zfZ1h5exa/71
ehE6UNa9Inlttz0XdWWDqVAz4hFVdBxvR8jhwkaDmtK7hhfAGJvowFU4+5c2TDO49sLXmDSWwTfb
c89081o69kK8GcFsTQGWQsChHaAnGi7RQKDY3LoGH1pPoskKTTmVLTMsv7OJzhq8ZBQIz6e2dhMc
a1fSUVxGCvummJgExF8uB96roydz4y1Vr2ZKvEedm4QnwuwPj953YdmgXRWTu5MrmS1sdjA2Zt9p
eK3Iu7uG70YmCasYePgC1Har3YIXpM+b2Rqlpervy2biExv1OY+SHUTLiwRBbYfJH6AKUR3YpauQ
KaUbKFEppVOFzYhvlfSA9NgKhRH8or7diLuzRGjSKA6ejh7PpNDxmH7U10N8QFVADnlYV/WVpECT
THTfrVgqFyMcYkbUV0wB3WlP7xG5WS9yzTp9TOyaIO6mUbagTQqdlSX33bRXmp8i8KvDicVUsuON
LU9oiKnZ6axlSXO6VY17Vyau8cE2GdKPdTtoBAqKCB03hfLanrEvbDSHP810l/9tuPHNvDg7X5P5
sP2Ag8FCq3VDjHwAZwqaDPtLDIpYD8+ZLc6HSdivct3rwrRkd35Tm8fIWZB6yKY+sbm6MLa5obXZ
VP7Dx4Vs52V6nhAb3mKm5q3fgy+fXeOaxhBZvIpx51eNiSogmH5Lf5shJUHtp+g4pZzfO31L51Ww
Aiky6E7j54yi7fygakawMVikvdbmyTYaF1kJDwe7QVsD+MRfOK2in1MBhZ0lQRp+S7ZC/wT1EoPy
AOA6lVXZa0muWbbBXmM9SsNl1LyxgObE4h0w5U2wKFbmZFCrflfcRM9V8sqgyZuv63uoNLnl6c/9
cvzRs6xNA5QnNZCL+rZi2txBV/848QTN2brce1vo3lIqO1GQPKbc75qe18a6U27zPK65z9qQF8MJ
6w2v6ka9kIy2PP85u7ZDOR3XKx+3LqCuktjKHgY9ADKZk0zXd1mq3MyIQfnBrFiaj+say4UZYsmJ
4wR4w1E8SkUY+62Lqlfb13jpI8mTPs7Oopl12EwYVG3oBVuFb09f1PKid00BxtJo9D4rF1Ze1Ym5
JEO+mnDr9rVAeG1Sg4NV/h5BUQIgr2zMfBlAVNZe6r2Efz6XVDyxom4F1eXpGVPuobE6vc1IPoxI
CQ7LviQZw8p2qMO9BWE+6g3i96SpTmsnEmIbCSHWvUdUU1EZIEV+2Fo0NG8qpMZl7LAmJ3kT7p4p
yHUExjIoxf4tjKPx91Z1fcXrmFI2j3P2tzkCsoTqUD11vDRjI/xv7Sg4y0IPZkgqJhG5aPZWTsgo
sZnJeGEtNkb/5G4p6DlehIdg7V/jq/j7sH0GoN1D2DRKdAGt2KzkZ0mnEOKcwSsq3TgrfMSbv4Yb
2XrmciTRglhYYrzKgSRKGkba+ywSHnKlP9/NSE0cfYuxbVilNKLuR2lkqiyj7i4VgmpvKIy6mbUS
1Vr1pOdHFAw+OwDuZEOscvQW0nt0hzasPd4UOsVd62Rv7/8piA7VZTsCAIjdTnqQh22y3v9nDIFT
Y5bWw9QS59QUus3zhD3osfxRJGAx9e93PIopJEl2P2cQRbQzlM1pG/fAMcu0JZVhl1QwNuh1X4b8
IIQZEbv6FE6AUN1cmdsSIE/OePULXIlsoQg2HYEaCcGQwNXJO0g2IjJdhw94uTD4AB13I4CYUBKv
XuN/3cVOHdGnigEjG4W2fvryDj/9Uq5ttiWulpYUCuX+lZcghRxsZ7urobuPi45oCvMTo0s9pQ/m
72l74XW3pINAyPH1vh3BNYrkYXSyL1/eQorq7iVpGO7t61VpDy91eyGDcmZUJVg2Y3OgfbNRH6nw
NRQdbCOtxrFL4kmT0Z3DoWs4CMrfRBC8HiwCuCTKBdblC7Wxhah8xyMGrP8o5pi0xWj7WGZBGKwE
xuKWxRZSIcXk7EPCHVXzYa/BWdZof4szihqFIZALOk2N2q+5feSEsJIRcc52wVfedjlINec6fK1p
ST/YH3ex34C7lXSsMyTsb07sJ/C0ipqdIjH5VVrxewATSS0+xOpb7E/LGpioiOcEomG6AuMezbyy
ultQaZ5my1aLAXOq2ttiATlLxSmQYDvjd/PcGM4fV7FhC95O7JY2tmFOXqSVeRC7iCPMV/uCZeds
wAAv2pZN2TmHf4wPFiMWZR+IxLm8Dnyhat6Vi7+nBz8M+fjylJ+69qfR5enn9RN/xixMWOHyza/q
lA50+xaXcAU4igvy4AdDIptzYY2gDuBDAwrm5erX3ifvHkaAf1oXzpmibJCMvTNE3UM97az+58TV
BSBKmAZUOv8zhmxynwFA3YAIUVwhkLCD31YQME4Et6UJHTzAXvSczi8TtO+WAwj2OH4yrqWfiNml
gRd9phwL+V++kMl6grWHEmR7KoIDW20QszhrhsKh2UU9lyxxBnSfq1UI0LW1hIMYYqOfsKeZNVv7
LW27yUCd9UP13x4V0eSLc22TQQRqzdP/I5L3RJyEG5L/ly4vbEmsGbBePBHPgElhJmRuJHQg/GqA
sbYweQYZ72u+nDHrXRp2e27K2ZiqlKuW7ffV3xF5Hf4LQ1bpg8U0m9Bj3PERsb+qrMN5CC7W4P4Y
cm2GggJm7nA2KeaCWjW+H8akP6rac+u84HRdSby6keZVQYHhsvDcKJ42zVOdUVHSH6noS/X1/rYY
25AmfVjDvK6XeBdFhlq3wWoU23lzmBjW8VvzcCjz3NQBKdWnINf8rtA8b3qvhenEKXoCeE/n5Lhw
OMzFcYr6ekGFgzhRv9US7+s6KxT4PZljz3qUp3LxyefOl+su/48d8l0nHb1r69HDTVVT8UV43ps1
4xpL5prcolygYFzreDH66mnBPjIJr/7I2JJM868gPmypqWavoOJ/ZDmCmalHKh8JKhepcPw1hYJh
O9LqQAt3Fj26mc5IpiyNi4l9C74VTgLmXEYegs4/q6K/POUSZE7dnGZxaIvSA/7U4A7lBN+4z3yW
05UhwgWArSxLtgntKTHhHgqela3rNoIL2V2REffrvXyO+cO/yzCC/wHsc+7F4lbVRdLoAu/Ee1QG
bWZ14X7+2aigP/a3IPTDwbTTcj/T39SRWLVlkKnqveEoCw6zXmbjYrvk0NHGuPYcD6sXvkOgQrDy
vtvMFheXelSbtfNNYcELWh9w/C5Q2cD0bWml34RHuNDIpVm8BVtZyX2zq49MhjXKPlYsTVhBwHNf
Soh22FvU45xuN0/gYHWng20MKxMPk8TXLsh9gddz79HH4kHD578LsNCaJahsV7TtzB/eCpz9pB46
spFQVpzFaFpFtEBT5rnFyaswZ4oeAlITsSe8GFZ2mnzrGfDzcuxapcdJHr/0lApZrXQv7sQOMY+4
W3Gj+JswoH5MdSJUsN0SoKd2qQPsW1DUKaxEY890i8/Pt54bp9lKQsfKEdGRmzX/2XvivcKsoSQc
2A2e7QHD9Kc33GERR2DC0iCpp+RutOWdMbpCQT4LhjSoSAcpPJ8htYI48TD3iwT6A7hXoGXsUT9G
ia28xbl/dhphlwnYiBD5pgAE60DNUCl9uUYrgXw/JMchngpmnyeYdYplRV+e4GlW/76m1lU8gI3+
WX4wrCS1xfjdhGOukdV83lwtGsyo1+tZD0xSt54vxDeWrrN6ZZT75OfYcBAd/g2MLPKJNTgTqkf+
zaBkryCRSEx53ZV73Ce792DadY5KPHX6mnqH5TQDJl0LcHkhA92GKwan9xuajmIt9CPx2MegWIiF
uCOsZ7F4BZgQ5bzDbgPY1ovUYI8mehnF44tgCgwNLeMhLCZF23/4DMWGnXgK5bq/ZZFiFljzmnnQ
5qyQ2h0t5GOR8m8gb5PKomxjwh8nvCDdmLOsgasEMOZtwjo8X3KPOHH4oOTvOG8PsnxCeZ1iIff+
xOxHV24fTpIcqN6FQzU92NeWgPxaqzdawBBlBpZWA66+qMrI6xyLim9B6LJ4UfeJmbmZvQkAan2c
3+V7NLOCdQTu9g79xeRjYsUA/whbO6dk1pJ0EHgcA2WjvVn6omspIvND5RgJ+2tE2/EM+We17y0i
YpR0bA+PNl0UhlGN0lYtp/MyV3TlcVEGwP9TWIn6BWSxWS2NXDRB4LqlRDG50F+VV9h8zQVKRQWU
bAGUaSotF82UbNeRwCY0ENkms2cWxc1k7HIEKBWJC5jRzfFvLlfAChUyJgACY7fzUF31/EczxJye
Ufyw4wdeUe+//HXkKDHSGzb3sPgYQwfU1aQbcPJheBrJcffvYrYJX/xtWjxjr29hNP5lKuLgQrwx
sB+VkxuSKR9ELrNDqsW24cq3y+87l5vuOAofXk287gtb46Rp4z6cMez+1lJG0fKA72kdCKFbEqcB
W00Zcb+ds+mo4NOrK3U15MmNxsnQThFhyEE/OwfdcwVcS6PU4u9AhT+IQV30rGxpib9CNOZBKI1U
nd5SqEPQsYoYaOep5kvM5RDJRmjdcZYvMzh7Vq0mnB7zkZQgnTSm2POiiKYNN7QGVwqV8+4ENd3R
I5em1qub9qx7C8L61VCyLe7YyTGn+4taM0Nf0ERd20lxDFvK/s2nRUsYS3Bt9ySs2zMd3LPmjPgJ
/KmxQQKG2Sd0ozoDhWyeA3DdaSld5aMOJJGVJvD3UTXM25CJfZ/Y7QOKAiHTi3kYfgnxBZWASn+f
UJSJOYPqRlkZt1UPwxiZWUdxGaSCIyPWeGHm1e/5IXFaYPuVWBCBDCIzn9JrT3UITAXx8OtgN8y4
uF//V2XFHEwUQ+/Tc3N6kiSgRKgOtYAArCnH74TXlxkldeMsuOKvdT1Bxjqrc8zR3FZ+SHDU8aKE
2gv9tlteZvPbP2YU1l75yjDCFeKKMtI+g6bNGTS5bShjRpXI9cTXGhPpJgb/JBpOIueNALKfhIvr
JkpO9nuo8SMPRK+Wqr9uSVe1b0AKH+b0Ty6v09v76FQYeAadT0zEMM++ax8hccMWj/H8Y1LCCcyv
mpkRScja7ejD4lD7b48e9t5dIyTy49cn//S7w5ZK+HY7u7/SpHHtBLOPWKhJBu6ufZMyH0XZjYQT
pjxCX/HD9pha1vEWTPZ0bJv88I+QZfOI3PR6/3XRDxmR2SGSwqmBckPmxyjGzi2rNKi8V+f9zHEz
Xx1QOacqmesgDPLlr/W/Luc8tuDrXt4WysF+z5x0YW1vFINaJW/thZcr8Wi+KCOKKlk7w5idEUo5
gLWfXmwkIfBtlkB0c/E4QOLLXLZvqmsLAzCmCNJ6WVoJ8Qp/Lc52ld5l+8CNG0ad4P80Iaz9MKut
ddofHgPk3L9E0cXaby2/Tb1Py58JENKdSeTSW4vHgkS+QiWjtKO+von6f53IOkFYK8MsF4zHTMUm
TlDSFV4b+n3JxKJtzKDrm97YhA2uXD09IsvtBODFtd6jlg0dNB4xHMeL9Ik0xzUp/zclvb1pE+Sj
XH6sTK7qkfW59JqGXKlGUWdundcgrzFGU2wJTblvSeTqskvBfRqhN+Cy3u60HsGaMRYl72lP1/qz
QCbkqNdmK1OCgk1IDrKrcHWB49e550EBGKI63FWeUY4uXshsL888Qsb4VYkS1D0TbQ4PCTsj8iPW
PfDJgbyjoX+nHKOAvTJNfL9UB55bBnBi8i5/DUMInzdQILHtBCxwwhBKZWdt7lbiPeoFJQFOeepF
ACerPYnpIQgqijQpHwxeNWTBKqn56fj+AVImCLsbJPJqw76NyP8NqNmRyKE3L+xc40U+KqDo4Te2
vj4WojM5Jq5Svya5B5FcqaVFfCwP1PLp9YfsPDJ7k3r0FkJzrBOvS58hUF5E1sdcN4hIfEJ1c+qw
bE4F+UM6U/G21/0blKDeBgydgYAYD5bs10p6xJusgXaNv6MO3uCuksaJsnHP6WijKzeIWS0Z8z/p
eXymkFnRiB9plTe+yHOTknM9FYZTnWshOj8TAZ3ayDt8b5D4O1IOrCa8qMFI/JoVYBm6alcHd+C+
LYkz+D4ad3ZvYSaVBBdqQHrj9LHEokq8+9vBXZccuaTeAxm7VdleOpKQb54U0mWrebbTa5nED5WU
CQCFTt7M9pIQQMLHM8AjR7KIrHoX9YosoqqCUaw9E0gE+/fueWPsvqE/9kq+kU2JGIHRpIsWD5F4
oEKjPhFYgn+9lqHIcjnhjVm2/AYnGjqyeWA8S8dsdQO13IGbrwbfAukhO+nWwFTPd3w6n3SuPO/5
6goI5go72VeZvn77gVuP33ErFIZurGt1eeWiDDOyvS8xb41d/3y3e2308jXbfMWi0IcCpO0oCK8/
fhxGOiqfrkkEEoQnFpD97riWmPkiNhVtLzFjN127i2HjlEbIJenu0TRpupXBdEogvXvi0g5fMF52
6T6NNTM6vRs3nbVgeyiHldQp7wmO0iAbD5uLBRbjRSwlGc7+O68oSEBWaXZIAkbQ5x+X2ZLV97k7
xJNfvrlWItLhhtsIqirC+DXDGacToq8PAE5eut4SAsB47Y+3Z8DsfVuKym8fKxCp0bht8B3pfuXi
HD889kh1oU4Uv8yws2OU9N8XpgOjBw24c2L0AxZxRP0BnQcv3DHdGq1ECFfGHENPE2KMRhaz9w96
0nxQKsVl6II2rBrJyLfeWCGOG8jtdV7ZC1Z4CH+3Yc4HHoF6Er6JiCNeQJo74owHFWF1YGaLRsFd
/zpT3s3UVGfrvKBrTvURKZ8Hm2bxt7+vVqjrz7LIQBrXHXfBp0vGByWc6azayu27bYz0AAsYUA8s
RCOiB1LOEkllrMonVXl596tkInmk7vCbT7ZjLcWTlt8oNCmx7wFxl2mHjgnUOpzsO4DYOwCNO7jl
TqbvGiMJNo+wkNm1LlyPl/k29E0sNV9XY4snQrMHpZbPwzfsRZ5bBP389qOQ7V0TadrYtbsZyrbb
Nv61ocU8TE8AqMP/q6RI+oHTndveJewjAZRZXgJQyAdz55xL1s8FSMn5Qk75GPzgaG+Y9/SjZHau
ttnHNQTFNoe3b6Winp6QJOT0Z2ReiPse2Lc4oJdZ32I/vANCJFrj9SoGQ6LuJZWwE3m2p7YJtFC9
5Ik7j6qidOGxW6HCUsyw9u8M9AskzXJA8H4QqFHuY4iEmXbVJnhmmuEO6YK/k5aVo6i5NZJTrROA
dQRi2nAAzjyc1KIkgIkd9gNvi8VuiNxTWtWlw8HbHugN7e2hzCDhypcp0QmAyS7XFYFm7lCMj82P
bOpkMmyN0ejfdDfTJuD72pKKZ0fghZ48pb8i2PoDhmN0iQcrdH5JPwCI679v6bbBitJO7/1UUB3U
pfpPe3EVLTTw99rQz+Itepo+7WOkYw7KlDHat7120Rgnc9IubF7DGDFNBFmH0AFB148gumgnpkxN
vb7yniRiKj3upZfWgQP2GlzGlpxG+AjflYdcXEciUSW32WlXuFjJ43w/wItmtJjcOGRL9Ow4nYuE
pv8L4kr693IknhMph2WXEfvnzvwKD2ogZeuq57WWwG3ceIPwQnPy95KGCQC36TqQUIkiX2SZqNzy
Qz+Pe3UG/nh8B3mMjg6EMCP9wy1y8iThuS9JmGZ9lH9E7JBEsKfj2qmL4gdzmqn/Du7i0dqvnFRv
RURiiMsgu2xNZCloK86LwR61ERMljZdwJxGJ9OPeAY+XtSMdVrSJ16J0xyLLjrDzEmZZzFyisda0
tOrHyLDT3AtWQ/OEPT6HzoRIS0JVgtK0rBmFgjM8QuyKD1UrfTMWl5Q6TGpOX+g7JUBseSFjT4Uc
JEko9UJanMRqZRvtobfjzfchhVbnGcoTomRcBvsHF53dHPMseWXBzXPWLSZlkzVJPAh2FRN161yk
S1oltyNrdKHGldXqDt4D1W6srttHspvTZ5zkD0CO5MWjXeO3X1xmORgz5du4uhIK71QZC7U65aBh
VY43xaeu2H71vAKoV3D5hpNtAIUpp4O3dm2iulwxaAYEvGRSIB6Gu+WSv9YxDsNAYcyQHtkaw2Fo
oOBWUi8M/LO63jvidU8tlS1glecpDKM1pkFHCJ2C6J3HBSYkpLnYLeZ5ouzaPI/q7q1MJMHbwdzh
AqQMJwnwNpomDkzE8QUXvLDoV5mwggoHN6kBCOLshRjaHSKwT3jGJDNQfli/1gr0ThsS7090aKmN
TuiIk8yeh173ISRRwQcpf8jI6EXPkB3nLKlo3vSVfxJzp5jLQjSjZXF6plq2YadHKXHGBBXghO70
Tnz3M84Ku6gUOnkZN1OIOCMaAhLjcvNkXQJc1IrzW2MJXLShSecOXE0RHWMh/zyJh8/1SivA+YG6
/lGZ96bSD7dhb4xiUifus3DLkuVaEb9cjKjQN1z1WzJRe/TdikV4k74609hx78NjidVeQrZTMfr9
SQ8n6HoGwaQ+WlA2g+kcrOkInxR7NQvaUjFhqbir1IXx/2L2r+aJy2ETQBA645p/9yVlaQZ2fM2I
7IDCtbNqN6PHVPGbeJmM+WJk5opRWaz1cIR+B9SFqnRcIjCJT5oRs51GxNI7PLpxqX0UavJSOEfb
NCnldKbS34ukMICUuCJiV3Xst+2576WcImppsVRFQ7pnG7lWMBU6EUVsVf5Qan9CjlM3mSpOxzn5
Hkka9ATnjaODMwZfZzQWvWzfeCqDKdOtx2KCmWeXkyLCraa4Icz6Dd5aEMgzOr5EFc1W5KSeNK7D
bfPt+K9pYVri5kezf1PCNVcgpzIJfFO/XlaAgY8eV65dCQ29GRzbAWhiLInNHUtK+LdRVzHRlcHJ
RNdBUw6JtPeJAWuVUKG7QjP0YdEy4lN2raHAJeoclJjeVlDxqbgPe8ufbh2yUo0LqWPGfhLe3rRU
ISmeAT5/vgtXbSsd9F9+5DrZpBPFlKQRJOtK3njxzv1SpDFtBJUH23SNWhPZgoO06OjiLYamv2tc
z4TbCpRjdNS8uCSjcQ5QgB2l6MZCYDxkQEPJ50300oXUPdUZpVH5T7ZYUG5GHoGAcwg/c2VzV+o3
jcxjJT0depenpAFXXoImLJtEdpxGhCAO5mYzCKKmZk0UW8K+O1DDFGtQet7osTMMZAEMb+8zfuWR
ASQubwwS4bln9nR1jVhunIueDjhUm6a6NkVZeCfZKoiti2Cv+B0dPJ2z6zXhe9orGve3faZ3DdzF
8x1hmeXiwpEuYBjdVT03OYhl8w4f9wP3zmLfCin19BN5tVSItdTZFjdPjj2FYivN387+nxbNyiUa
cKhgTPgLOQyAREPH5XGKJgfU0S9Gh1rcenYAa3W1raYYKaxtRXC2v9GbutvRvJYt/0PAYSO1GTPD
awb5RBxcd4bEtNjU7GN1s4uRMwumtI76XiMpXU88UGl7RD5daQpix1D5IzIszBZrzAquLlRfAOWM
poTkzTSR1OmISdGqMx7wcvYrq8EtmwJQEl67cN+8dgD5zgUDTyEp6YII/LkF64l4zibefJA0TqtK
hyb/+Ym16WH1JAFvg/dVY7h9JhZUVkwL0Xo1ziJJcaVeWJTm1RQ1AE4ZQeX0T/6zS7TRtSp0E8qF
BYetUQh0oSNSiR7iw6mLaMijxbnR7atnb6cozl3urV3TObz27ZElzn8168mW17JRC6Gi1a25oujF
X3gUA4UgJQDBxgHw2Oj67YuvM0qnoPDKE+wWCX9H6hpW0fX03dV361gEfI8hl+6nB3aTRJGD0Qzk
4t9QoyYhUJOTtjxj4kmczl8sVslhqdOY5UgdeHaH2f5kkVYKvsRPyCqn4lF+byP4VjR1rOpHPYmt
R7ZvOwxkUrHvJfgLzIj4hwnE5JXDNQgEzzE+HhlXvyejgMW9a3OUh101Q4kq/PfCq2LK6maTlHew
xwUeAxiMH7iS3LAp8DQ4YR9sf8rWqGTRdngHUp+eeYa+DT8eHMa+Hu1oPm0aQAwzBhLZtf3/81Lc
LfAOONFqsVOZLQz7roMmEpCEjwUWf+KLAWpAAV0NedVDd4tt4wSkYRcA5Osuj9OkWBC9IFg3idtp
q5qljZFrgiMKr93J3auD9zgKMM408YKE3YMaqrUl32MqDhrXYcozUTs2qa92HP7cTNZSn0tZPDrw
gvPooDZUFqzNLLxldLs28KAHBl1khUu3PEXWdEmuHyUTCzV/4SK7r1ZsP4Rl2nO4uwx21N2T6hg/
saI5n7s73wIz1HTRN0ph+4TsbDYGFPhnFGHgg9q0u4oFxM/guwMG1TLrhJNOM0DFws66MMLUREja
SmIgq3N4BtQx1AkS1G/awast07vOBmuU4fRdzU5TmPPSRcGhr7muutJxaq5tbJhjRHfXOwNg8bFA
y4CSGywWRrSMKB6Lrn2+ctIhB6YE6ptZ4rZkAuW7/3rvMVF6z6ru0Zdu8Nczdq5a3JpFkaFE3fVH
72Gdmfr+n+pYKI/f/HHTilAbsMrEyP6nu8JtWGzZYkOt0g0UuZ6Hc3mDf15AwtkNpsUtsUTGTpTq
hf5nffVizv8RgRDvSj0jR14fFhd6W2in3xymjgMQle3rLX5AmCgXGzI4/YheBjT/gSe3PK67Z6vA
8YzQLh/d4bNIkhlO5Veu/bRx3hRXhyWH9ZjLOrMVJnN9yjjmq9j9S0uooU8CgTFTHVEq9Dh4O2LY
1LH65/g4/EMvU1D8Y4T8+V53Vc7mcuRbsDLMJRHYMR8bIDfgnqCUhwexn9U/1W7imZ1Jtprko075
IE1H/qa0/nxRYF8QNfR4i3NsPRkI1Rd9pwlbdKedSw3gpwzNihHUQaWWXQWgEbbp1oQIFSTZSGQ6
/e/KShmG7MulYRgj4rAL1duMsdCRpAs8DL9gUibtBf7qoqPmoD89jtNrrjHsl5ETYt9y0K66bsaX
KPuCYwrR1ikJ202LSegfBec3UHH5GeYQWDRdxxhTlPGnIP29DtyxUeh42oN9892nL0NXSTsXiZqv
AS7ZT1VkML/UQm31VXFWp/gh3U8BnRdxSbpIRt0TeBcwXd81FV6k3dhbkmq2Un7a5aNKOVPw7m1T
jhpl0gkU8AKzF+R8J6Dhr4xjNjeHGhdejnxlU3FrYcrwubfNNwNS+7bQEnz4lRAIT8nic4mygTwv
52ys5mQbcV2uEtkU+7/Kt/J7x+K7cNF2DuG3W8EemwZR1CvOtWPuEfdpRIQ+3RkmCIrLEvTS3Wa0
EeeuwjSvB0ft0LztgOubhrqbDiiYoFZjhRc9l6S23N29U5x5z5oZP58t4mVD8NFqhOamHnZVS5HS
7jBC07CG/LZCusjXqPq1yGZnONiOtU1PQRweQZGb0GBJ6+fJGyI0sXmVd2iS/fAinit6hbfe+A+4
elbq2nmdJ9QndPiw21M1q6iYbU+qV6IJm2XqAj9Zh3HIbG89X++ud9+kagh6Y03oqTf8kOjYVL2A
o/A94KlfPor9g97Mo3GzLrm75p1aZjcevz8UYNw+C7Elmv+8QuBxOhjzsHtwYfxhow3Rmwt1QWWJ
LhLj2Oz3LwUvuoCLZQl/LcxuQME65AWNpsMoBu+doqkpZgoVoP8QRr3xhG2GKT18fThKKhrhowtn
5v10AutMOev6B/pX7gMTfakUmkuiTdLwZdfbLs5Hc1ku/rcG8cShv6dIeDp4mW19j720SOF0cWFS
mxJMQXW6cnOQkWU3EM4lLU+6CHsnFz8nZr5XznWcdTAXUPLdJncleXP5TiPccYv7Ws+uWAychIv3
N8mc1SGc+Tj1M9EsLYzoQAq6nIWQHhTeoJcN+inir0hlzVVnQs17wPM6gtARkfVddE/sYbFvICo5
6hER9rcv4cc+/q4/Gjt2bc7S5pJiouS6XqfLgsyFuyuRRB9zAUCPvZ/KpXyIiD/HWAtImdBXiNNS
c9uhEMruznvUuN8itkP7TJRwK3dN4Mh0HFuDgCxQBeOg59NmEwssgwiYsHfzj6ZUJU8gD36gXj7C
tqG3i41xfZQFAbg1kzp0VsYJwVMXGhCRnrUlLOWvvIAhXT3m/5eFTcs/lrDyAQLgLaUySiHOwdRd
RUnyGrgtvVAOc70KhFnmj26nYiSFbqs1a0tttWv1UJN5WFOYSZ4KJDOsoyl51+MDtuQRenDgfNze
ti2BiLLn5jPTlDWTkpzXLqDfZ5nmj3mNtVb6l+ULO3ka5F67xyWcIBYjfLhnklCBGb2GPdCjBEVM
WOFkQNZSswLdNry4wCz38NmMcIB+2L76yPY1cFdoLfiH14OMnvE3QStpxt+AZYn1rAv+mBezEGgE
nStdocsd9WHu4choHXID4sut+wViPmyUMaPaBMUH/Q2QFT/H+7MOiT3Q2P5uqkkySfvKDWUBufLI
rL6AEwrUafAEfsLUvGoEX57HiWSzxPc1cJD7qGAbp8J1hgSaEuyDKWg5El7/2iR6jWmHmfG1/tjq
aXfH4R5vYoaC+s4geP4llDMYVRH3IX3glz8k0jhDspQ5lgIN3mvKEXLtsq92zyNPQoDTYwKbFGNU
BubT7E40jWO/aXEXs0dXpYVaWieXA5yUBhk1eG63f7XbMXNm0yvq4QNU16RmybJyj03btsCnsnQI
CbetCb4vzz2COKntPYNXQ0nmwGaIJyddlPo6kh+RaX02nqdpWk3h8CVRltH0ZnBdQhP52qQEsRaq
BzH99s6/UOkUh5u9Dx8jvEfCh7CnBEuxpJNlniQyuF6I/me8GdsLvGszwdGSF14ZPz2NGVhAf5p2
6yDc7bhQ3no3q04GasX5dmLeqhWmwbdygFNJEV8sPd4w0yZHVeKVuF62TB8Zx6+o54o0Sfu3oV+0
Q7FjVxs+vThE0yKHvsKC4Ni7cD/iN+853lBLCTgOzAlMFE9xsYd5dD7v+6iDzapJPnPCAYixlYM1
h8SP/3khTJVjKwV0y2IVXYhnjPDNPDyqbXN/FTERBAcumhFsndZdLuXrG62VoxiHvStjD6RA8EFj
oZsVpN1H5q+STvWNRfjrJeHpZ+GPptKjKX4UZNMbOr0YS+ra8Wn+1ULFvbH4G0eq8+krgua1dnxx
88wXQo3CuWQVZsCZRyNv3fYT18EQBMTVIgZnzba6h0ZtTjWmx8kc2EzNX6RQcAn/rDoH6pInC2eq
mfw9gw66TMcWIXbaKhVi8pSJ8B4mThVWIGdhcZebWXGuUvSRQ/0KJmoQkkQeM0LNYKGCRGBThsrj
/0PzPor8TTzjdVwjqI/fDljt2loQV2WbFCSHrcSs4xLmvfNQM5/C8mbCbMe8bPVxm+yDgN/GoCjJ
v9x4T5dw0m+kghTm2y0Mi45H7VSA/K93Ln+MZsgvdm17nHS29HtVOUO/zhBRTrpTtxBI+8oH5i4k
wmubTf8P1FMAU6vgn+Pc/guixPr6TeX1W5+gPDPJI4+USiNSFQGlGuzd7iQ88oRax4Ogo7XMI7pn
dMpLNYczozyPMOYI23BN+ryzXyHrHjBOFQT+EKXmOdJApfi/QehOGnYKJXrZmO3lsSYQRwWlfdVY
FltnJPOUcprS2Qyeo47ob5w1TFeIzZQSGUwAaozlm0l4Ggl7lsJDjruEReR6931A9//Rz/VulPM1
OziEwLDSQb+FqBiLo80vh1eb/zlsihnAcCzuxa2xpF9qPX7GbAiwDObpJ9O3YGd6IGlKbkryOgfL
qLp9RqMCl25rQSfWzNZEQJwraiPNqenQWZ5R10l5XAKyKJZOxyONQG1TBYefsw2YDsrjV1SPd2G1
Cq1BfxsJb0cs1mI7vHKyRnAW4oGtnBUY1tCelCgmvzUANgcJUxTJ2F2xU/AJTUsjFtTykzblJClG
Dw/IKXyX+6/YG1kuEUHi5AQZLL7dtUMf1AHd/6JqQBciQzLP+DWs2SSYyFetd4I8WzHnqICRvBMz
B3c5nzCNgyAos/qiV0GEr++oU/3FOQFFr6CTeF5vAa5pAYJOipO10Pd4eL9Mbsi4mjtXwUJdvM2O
eKgJ/6aQBY69/1DFd3aMC9mug83cpiccCMDOI/4ZTdlmvMENtTGWCs/XNoDT8DSIfP+voSDRVFia
yWotCgrBuLJ8sfHV6Kc/k1jfMoQxpcIbTkEE4YXKwYs0U5dQ2cj7OA/7PouRZztk+iWDDM6qSxiB
TQVZiLGfGCtEBdbzer0ANAI9dVTHY9e/KiEwPUJxJ3aUjSjquJwqjZwWc9Mmtk2wbY2ZuUl5Nku/
10INFDUw79MzTEoclTDJLftEPHKplB+6HCf9fbEsCyzj4aNG6VOXvq6Hi/Y223TbFd2KXo55A+mp
x+dtJXx6ihAdJcc1MFv2NUuErRdsSdgSmsweYN5LdMNrb4Ooq04tyuxYVcYuySsCS297pPMimXMw
raozEZYghICSVt8GbfGP+SecRJJydqnU+sdDFdmfON0prMp05cf1JaEJxUF2wsZMV7OtAaZByA1R
QRkMXeqnhP4sIVS/8JMmLPfb+8kwoyA1Ui7ibutyPAnBsgIQsDkp1VUQyLBSVDwH+IXj9x6Nl0mu
Co1bhWy5U4aLA41pe6qgySZ4K6TswWkXy3+9aTdZ6OlGSYDGs6BYCsvz6UDUwH7X/nQvvrV/seuM
f8r2f6Sz9acN17kOrskr2E5IU5NvVlFU6kNOihmNodc3B914pWFkFruHny7sCC+HO/kWFMcdSVD1
SGypONGuto3moMB52UwE0xnaYRq+CAw9byDxq8C1R9YE72H2sprqN2T3aqrH510LYQJWZlzzeEMt
4SGnThslpxompSm2rK6vurdnbeZ5g9EfVRdJPRkglVjQQZodD/sBGTcrDtNYRPloiw0l3WhoVJ1x
HokSF26svpl/UvrYaA608PFXPSNNkG2oquPMLNSAgLvEM8BwD5ZNNVm9QqFG7o4N+UocPJz9lv+b
AnSONW2Rpwi7At/UPLE9KZrdLMTMy1DQv5WpdXO2cSaK8ckpTd9pF79UaKpQQ2VtPTo43mDEA9i/
UI5G2NVzX93rjarzXCeihLW2yjhDTrBJQbvdlHHYMc69Ntg2YH96ni9ss4DkqvbAP16M21x/9F4P
bIMEXHhNmqqA9cYfGDdFbseTvchaDC8jcz1G+mt/RQ0D4Wr2CDakZhh/StcBO7gkEkRWcRrWZidQ
S80l5u/S3LgOM3KGm8PmaaBJsuzii3HYyRX0De6DtLcCapqMs9vrFbfllmszB6lj9u2KBC6N6Oea
6v12AankPpvk87RbKbnddjQ6xw28NUs9Cano5kGNYk7O0ahgP4MpbEQ9eORbh4EkXc+hsrJb1eXA
FA93zzA7mVpc6Km5NA7mMUJM1GUzwx266kbxAftMTj8dXy380cpM0ZVn2G/SMSpLgdyEBCzuHJip
v35ZsiyEjFB3N27NejcgOsdY3nurfUB0vNBryR88GVig5Pth476xfKcBAD8GsbGiFHiqIvp07FvC
+bHnbcyvvtcRuTHcI7x5tJliMv/6HCKdDwnHoJp2Vnub8tBrFIDkkGvbF+fyr4Ikl/oHmoHgbw7G
crw5fb3RMoMdkDUylKqsilFDwuqMa3uPwu6ajC+ZFv/l6Brb9VrixulE4bR13VUAeyNmDHsmyZm9
TQ6jwy2G9nE5PA4cCHvIRQc4Lway7+iSMN6BXm0iKghKOfOWI8eopJ9p5VHYYn692135v45cRL4p
6RcZxAEuo76XI4voORRlIRYM5cywMWCDGXiAby4EbrO10Xyi4qgh8uoePjzuY2tl5eqiF2ZDcjfx
7dxSbabU3KWngstkudULy5z33i8l/KAWuLHU6AJLUF8rLUTh6svOgByD52b76hTqwzODom01erI7
5Kww5P0QJKSyH4sgY1Jbln/MfP4HXB58cvYKKFN1D7enHJFYsaGKR99CRl8iTPdi4zIryUz+CX3g
t4VD2jjUl7Yq2Z6SV6M2JQD/9dLg/6DISx9hZEcDDsQNX4pqKbTiZqHFgwY9sYuKTqusHZYPJP+f
avpeAV4rbYlEx37cvq/kEggrLbIxlvhLJ7afzQhtY1eL9WOTCvdv+miq6P5JeHW0wDnIEudCyTat
C9R5ydF0pKQC5dmIS6rNvPtD5FLsN/HGcu+nX3Zz1f4FnYTpN3hTpvzRmQ2c0/dqVsynL0M/OoQX
+flTooLPoFc4EcrzqdjS6dlK1altNpJooedwwO5r6C7j/F7X8gYfC7SkwNyuKfBzrs+szTHn8R6/
hRjHfvVDiQm3qwW8vIX3DmPlHnEipfFfSjheToZC3RHuzB02mNiCo53SviW6ZyoEhS2d762PC2CK
ijTeatJx36RcWq64Axw+JPk4fm+7Lzp9BC59c4g9jVF0ICD7H8yP8w2pXRPZsTu+Cp2L1WToOB5m
ByZBnVLctTBgdynbWVyFn9Kb/YYr3FGaQ+14YRezB0NnjVWQnd/XlATeD6vixNwgrKSp2eFWzo9n
x5itTIqHjCHmVHZ6iKoMyiVF1CbhicBt8iw2z16NNXwcuJwOZz7vpvHMa+0c1PrPTD0s/EGz1rnL
EDLo+FKNuOZCk8PLa4a1qezyotyg6m5/9FaPb//NituJX4Csa82K01XEehgptnvUibzS1xmz3Oj8
FNfjTdoGLpR1VAmTytvxb5dMOL2GeGxGa/PIYeO7nNAzXufmy3Ivn/EJTcLCVZz/UnqY+yF8YkOt
WTqELaq9+5YdSjR9lRRgB8Zxm82xVKeWD5LL44GCXQGOTY8UehzQtRuByd0TQ8kcBASQS3SISh7c
q+LTD0fSm+7nhlEg0K8IcKQJnaZpvP81yNO91tDXsvrr+CQlAxxHKyRgD/ZnT/oRH2HGTEeYW7QL
1MYndRTkp51Gp5ZrrpLVEi/smWdu5AggJI2W9jh8uYbPIvpao18xomQRN75wgZXWl8f7vl1Xzup2
4dlEwiDJ3wUtAALtvdpqHPq6cO9Pg8bZK6Tho120p4shjOVWkN5ncuaYvCYuyGwwsw2w7URFiOUX
Fb28vh1vD0xur5S8Jz5/i3YHYuRGkG70a0O2/Vq3mlMBUKFplT28J1oPPHulxOb1Q1hkA2VcFKwV
LeN9rj1pZEROVAtw+gvqtK+vAIIfrLqudkKPghJEu6d2bRuwTzH6D1Sgj/N6ur+vNlGP4z+BMfFt
Ly/3dvDAvuKPhAmYThiVHieBQCSIXfz/8fix3pWvs08owIGJS6Gt/8oqicJlbt319JJZxd8ze/C5
6FYQtZOlXPIfHBrrqS8h4SWoazEKxARmEysW5s+ubxo75+58+Yv2MA+tK8L7v7SjW+bLWBf8XKsl
63K//1BVlYkU2QrdYlr83cz/1hzgHLK/Mu6u95ksZ78SmOO1B94jz23dvsWzblGhvSKsKL6RJU7w
MNvPOoDkkODdfKUrk7KxfObu9GwQoP0rHxju4ZitIXLCFkSUFVPOd2TlCa8Ca2COno4FvB4RaYCY
HLVarkwLXANoatUjxFNPytSRL7Vgxny2voPVUDtvaIW9m1t2upkHk54lhMyuBi5Zct2JBDrdFVzB
eh/68hKLv9OQz4KtGyjcBACEUneVUJHs66vlTvfwicR7ddK2qp9v9AcdqlvN+5QOD8dj3uohv86u
cgG6yS/w49Uf6w5lVo6NtQHd0657teg56Clctbuy93yb3kDVM1Bf2ruo5Cs0/v0N9kJdg7w96anm
MN86GqL57zxUKYZGQe/8yc1YXQsWo2GVUEw7Iysc8e4kwF3HU6J/09iR9PCvwfkArxp/2HuAOT9a
z4tcuSDWNY/dw1z8akbLhr/9dhPgzN3b+rKD7EQ7GqEWfMC3w9HeVackvAz6wUvyA2eH7Omd1oiI
lRu2/lbiFng54+nXs0Y3csPvlHwznqdFHvkGD5mszfNoe4RLrtc3VEXoUDT9495AtccbpoFnZmTd
EsKwcbo3Uuxgiu15mLiegsiaINay/B7LvRtbcstaxPqLTt5UJAI1NTc56V/GZogs8GufJR+ahPFC
kD2UOKEdHDnQVT88Ng3Edfsg1oTc3JqUc0Fh+O8b5VuWVS7ra4JYHSF41G5GmXAkm43J8k/k0M9I
dx7j38dumP6ahZVmWo9aLygTo+duvTvBtv1Lcp6rhNzspl6kaXPAw3ctPVZLLl3JXbgIYAd1mKaO
1fladssx9sWi5VYn9zWiBdh5XFVTrcYLPKGFfkqUhCStCo43ZT9cqsZJdEeuAvEi269nGqhYjr+w
KSXxEojwfeASidm3rODWo3BTOoK/11x9tjGD2FT9Xu4m/lnfcwH9lxAlJEbkbjEldT0HY/8Aom+j
saqmKaiPTzC69RO6wauyD4/0rzC/VdXxndTI8hDJgjLGmf9NLF9oOsiLr7HEZQAHKGe4a16RwVYQ
u2wF2eEsEQ4rpnDsaAOiZi/vJENqZ+VIKoPo4XG4eYXARFTzrsnNdWktYFTcAOOoR4UjEMjuVYzq
z+1q2F1EFq6qcbAcCgDEoegnt3X8NeqNMq4+ROjQA0XVddZmvGcXgyrzz2un3I6oTIS1lxD/zeDL
ELiDcr7UThJXhElN7Cvh0wSBoTSN5Wbp0Yi/4AYKekO0KqKoe2LvSVJuz4cOOtXhS/yFw/DHz0OX
FLdgoF+swxHpsqmJG1BHGd1EJnYxvxQSxmiqrVlypfsjV1HhziWC3eztKSZ0CoL0lhwr7iEfIGgG
fSe/mNCyyncVqTmL4G52h8kQRAsS+UYIs6bz3+EOM+Hlvky1pac4PdiG8IpgHfz76nK/Dxc25wBU
XZXgqdztSMTrE9AZB01XFEyIWsZfi5bx4FHnH1XrtNBts+OKwC3Aj7TQGzEjIIbbgoWjpOdAuCMS
P9v+qwrExAQfztM/HcYW7ZnYhw6x9WyO1Cml6GDmrdKEvl4fdo6wVsMJigGFFZpfKAcgZNVDmZ0g
nMovlGydY6cb1KBkn+MPV4yAv9VBONI8uUa0mc7K9fE+5l3nJlO++0RXD+BiWMOxjeQWxo858P4A
O1Yh2S+CKUdyBQ+KMbmDjrlRf9W558aGgaJNOaCUNuVzezQ5z2xZ8fcPybJeXA1XDvk81yHpVX2B
Srk3tj1XkMrBEUvi3+LfNAE4b/F6QQvG/Yf+lRZFlcBQStcJ7AYpGrWBrvgdxqYD2LJTaxg2xqHz
wHZnqjdb69bg8z/SIrR/yMP/csL/f+ByddM2nF94dHI5t9UJ5Z16qeylaJ+/RSbc+IOkROtzITPG
jZss63G6bdlQ9TvcbCS10IU4jzCucuczHcRMhU8L1PGdiIqywOHFcnBSuUc1JN1h9l2cD5KQO5xT
hyo9bg5ixqMO3s2Oq1CtWmswZm+7rXetPYLmZWNFW4kaFwWuIymG3ynuLPObsC3Y8YO9eT5xZ1J4
pwmMvS6A1k68RFRs/kNjLgXagu5LNwNjLL87zmFMw9tuuzaJiijP57oKFH7NQoer8DUldTmEvLuI
En9IEudtdDGrMY/drgGMW8r3tR6DuTTgEBTUrKTEkxffznasts2HtF6G4xFWMseh5rbmhkzIJvzo
Tml6O7el4pkdxUmWm9MgGI2gCnlkGGFeALuhrLfZq5nfcNwSnEoQC0Pb3t0wVYeVxRB4IZ8vmGhw
6WqHiQW4z8cq/N8sreWgrX/gd0aiLjSHqubExnT5g3y8rEtamO/g2/jIgkrd5En4CBMxT1dzjxyT
+sW78pW/B7UJXIHUZ0cSMwHwkMg6k8mhE194Mq8Uva2blx7S1vkPcT0mx1jGOY03wQrU8X7GF3sX
jd5TcPfPkeAWTHj1jxDLe61O/FbLxhf7SApWd8+EP2ZwNQRKglv3xnyphAQU2IsKHuvHDysyMsAL
ONuI2Gm1miBUkcBra6ncNtaCh0Le5cYJFnPeMAeM828O6OyCczw7JQ4HK5ro4Sw9k6bqAi9WDOHX
H/4xw0cEalLOUa41QZCeRFpGpVq2ssjklE8XBMjzTWk/Tg9z5A8Q14QxhGi3dbXYl1C9MLDJJvt0
F+8ZSYO+Mxvyu49xmHMasKLXHEgUoVGNtPlpqnTmFd45kLOiC+iJJy9dyPqSY7bVdLYQ26GuGDZ/
MTe1HhrfJQWibxGOTKnuPMQZcTzzG2tM85cbXdWLqafyZxHRKxp5x4kRXTh8Hm2RNqiOglAYIkXk
5X3xn2m7hN5VF7+JUeM2amDSssIkBa/DjGlvORNYlmmMmOZ5g3s9Q0cnAUuZT9rLLJOWWrBKUuSk
u1l+ALyqYG/fpo3fmyYNdZL3LC6ClwkUX4jyOasuHYKtukFTg9qKwUD6jmH50LeszJpBUPaxAq/x
UtAN40u/RQJMgUYoEFZVf5Lfobh2l7buCJ5WJ2CoMkruw3Vl/RmYIaFS72VZekmnSr4gusY1dQ4g
XtfC1HWW9XU2gl65azNGB2ot0OS+wN9qoFtMcegEszs58HwCb8qNg4RNeft7J7JPWdiwl/fdE2WC
j5oDSgGJWJ+Ssmd9SiminjqY7/Ktq1ghsNiY5RhJa40nJyAqW4kvMusGa8djFb+RHbdE/XXhJl2x
t7xCbwWYf5iKahScrOJpOzDt9RZhNiaAWHjiHPW0uWa5jwLbO/WwSpIzilORHI0hldPue3tfhAM0
FTNtp3Bh54Gp0UzDwWFD5OvkUekKJn1D77EolEGmK+3U0mRWOcJ019Af+RFHg8P7QCeeqv6axgEE
yFQBbo0p+Cr9GF3Tefco/qObW5CdLHw8gbZYmYEqbqdZ/B9hepLdl3VqNvslTqdIzUXTZUdrWDey
YDJm8/bAhpb88TZsE7fveYfrcfmTIL8fDbt4JEfKdwD3nAzYEoSwKnxZQ7mIpFluUHa3VX59uD25
Y+PrbqcT8V6JNWD+eJqhLmaya5uJ6j8YQCYAm83ghPYARfqUdZwmBHY6Osa02dNvsKnjf5kopudE
L4nghZwDTws815ZFigOxIKVZPFCFBErMrCTxvjSSr/3P4lbjuwT1bVj/fPUcmSWgrMBSt4tJw2x+
TwRwxmIRvKM+Vh4xq+PX2q7rWP3DufyE9YvrAUX8dCdD1Ze4DQhc7UoCANrxqHusnEuSRTUzWjFl
FC1W+kb2l/jWjlLINO/Zy+RefAP8Ca90rxPIVsBAJx29hngrzgabmJlSVpskNvyi8R8fuVCY9EHo
hb89bxQiHe+t4/4qD3WkEahgSsVdbNV7Uw7EpohUMTu9JHgFcZ3n6KGEvQsRvcBrAFXPMDTmAsE1
uG+KBgp6TIKtK82AQBF9sVzuvmXkpHpx7TWPcsuHs7L4fCD2yqF/uYp+DgK+vG5Sy9QeiQfKq6e6
iEyVJqGsz0VgfMOfFKNshgTpTuDNaOytRX1WaIWOI9AGXqdVXaK0uwLS99r0IPFvP+K7ocObL2Gs
S71c4s3US+KsVAYDl6fFGVwocLDPW5m5xZ5X0wX7RbsoE91DLdlKJZBoGd4/NmNiYRubLmNAa4wJ
HqQc/yn3Cnqy+6qsFzwtDIovGYsdUSj+yOomw0Fkn9En3Xzebci9BbUvF3oOLPp7m/YknSRB2pPu
Y4JjgAT6awnP9ngl9u7yRV5ZuGPyxrHSlNLAm62eUgK1q9xtYs6M7vhCK/Vjzcqedoo3oZ/vq7Gj
jkIoDpx6prAwz/CPRrk5rXSMDOrlYAv/dKfHFhhtAMWLl+V2fJEQ6bPvdB3npGxGR9g4kD4SPPOe
mknUYdoFTCQDB/y/nVTbmSUSC9x+bYMkzpdKZkdI2PMkPeEFvuh1iYJI2J2QrHCKLjZzhDgKufII
aofZbw+XSIKbHaclpgK+Q1xPulebLRTsT3fpu+OQYB6FtEGxI1OrJXrS4aA9NbaCStio44XaHg7X
JzBUn6Da92N1GOJ/VMBoU/+iBulPp3siPRRb0ajmFA0LkFaLKQ5w5BaYU7csK/iGvDwCWVvzBqwH
koDP1epvZQ1+a/U/kOEAelW/rxUcuMDY7cXm9gE0+3AG5az/RaMCBr8pN66TPlbNXlkwoPpoOkL7
FW+0fTCzljRXcTpOVii2e/VLjjaDRpG44zGyaYXyeQOrzXvsN7Xnsx5p5dbj0n8uaANFDi0HTo7s
H6DwTktw7FUOkn35W+C3fk9qN7JNNjF32lQ1L37SGl0h4SQgbKZ1Xl0nfR7ZqxzI85xrx4rDLTCM
PncEAmUoi098YiqVEQTTClam7bcGaggWbEGhVHP9XhxQBt8CpqCEspIEKP0WASeecQgd/eOpJw8c
w1eYsWuuZN99dvNlkaBEI9d+2EgNPhGz2bDl6sA9QUgR/olP+EhF7tu8Q6lsmb2JjylzZqXtftup
HgwkCVFHXrcvlMQbTFjL1czr9RidixOMNU21g6pv/u3zQXijPEtxUYB94KE6uEqcUdPMr7RdK3Fw
ZDEx0lYGMCxZ02+DvgHVueXolqpELA057r3HCi2RqB4w7gskup34hwL48WJigQs6/W8qf/GAHw2Y
r4OLn6g0GOBtn5RemnCO70wyizqQdJ26J2SHfxMUQ80/Rtubl/c9vyo3Tzn0dbgo/nzaGidOBe1N
EsQdotq9MTOjvP6kCRKVyn1X56Xc0tHg16pT/cxrBhfUKj05Qg4juP4fwLQLTSgCx0JuEMjVF+vi
xJwPFkrX37BHVUgnOoB7HhEcRChK4ZebGK3IaFEPPJefvFrVCPtIxBlBUzx6NaOqucadzgPdsXzj
9FAWalIQoeHK75sdtyJBcECVq5M11A8hwqTer0LqsyEPSyi+m6JcMlWm/G8EqcVo32Fwwe6+cKim
y6EpTAMvc1io9lfcxee5yBdrLlOZvP2YNRxBG/qgnhJ/sc/mB1+xBAeW/8i5gJq2uTvqA5iOZN3t
joS7BuYcxHkaTApPDQ69hBiT36Yp/9lkTBalDz7hP7Ua8+JOj/AMaq/ovjQjG7wfcYGjpj5x5bnL
6O0FT1hikJEmxdqT1wrrGhxXwKEwzsSUf9uHzPpdw4hMT+5pppk5sj8PqRMviCEWUzpeDdPuquHH
YX6i5FVTdNrH/Gj6xBUc4friz50nULX+qpg0AzL2EM93H0b9B83mKgndTpT2mXUYTF5d6kMhSISt
f7PxqdgiIXDxNz1mJFGMLNsUfBpYhBhT0cm7YU2sOP4tRfC/foKGUGw7GJ29m2n/BC/kBxvPfep4
1NvX1V9MG/euKlea4pyyx1GBfH1p2ODvpPtglZruY/5GJHoHxJr2jm+BAVvzuHC9tdLMlqg7OsYT
cvESiGttuHVgEC7BHb55zRVRFsuahdM6RUyvIELdQ+M6I9UuTinBd7a68mpOqusa0uo4CRkZ32Z3
UDgrBo1VXVmanXOPJsx64S3T8YbmzdHEaFCBSITJUmchYJ+MJI4bjy4Q1iOjuzMrtJVtIAev2ciO
P2O3A5xDBgaIH2Y3PxB1m8NISvBdPt8iYxXEOxh7bCjLL6bDQMAOM/bxdILovq14fuh1IZOsYO1o
S3Fstw7DZiZwrULmbipmbu9R6u0ntqU398ruGltHHfXskZ74EMOB2ezIJkVI6Qouqn4Tre1MzU/P
TUxztDE745AuVCtG7lyxP/yGDlesyMDE0++MjZ0AZQw72OUiaW1bwwlrK76M91c+YRh464lG1Rdi
zNcXVi1sFVd1h0MRMqmGgz9IULTKjPyUSikk5c4WpKu9tL/6mgmfA4V6ecR9tP/LbZNPn3xBCSNq
1hvUyilJNV0h6IZd2o2zMjOlPq9V9HKLaVVH8Kiri+FCbLwqGDjEpaOlYxKf/epjOEOrko+E8yVC
I1+TB53LgvbUvib1S+XvXPT+uibh/5zhzA6569Ci9Ytf0BJUj2li12Tk7UYh+fBZS+WPa4QcFPda
8TmmRh4q72Tj1PpwxpnkgvdTb9c8haVCMXMhMH0vqjHNsrraO5jEZglRQP7gsyzFH6JiQLMZwx/K
E4uTcTQk5rlgiSOkiYNeRpCtdFMvTfCRY17wSSFS3h6lBIZkwtXwGKzIjaRE4Tczl6pkTHJRWstV
LdBKs8v0CISoQX2pJ0LQIlMuz/PRMl9GRhFvPKK/FvhJ1FyfxXtIBb/kzS4flX3YpZj8GCkNIzxg
dzVdLCITHIvV4Y1+bgUU15Gkxlrb/AShFMINfm7i53YyNYirlzqzOnXUmBSF3UPK+CR9jQmpBxWf
rWeKDQJblhgJHX4NCgcYmVDqzhACnJs6jDIBan8KuTsvmAgIENt3nMWTrvHuvP5A5v9psp+zutrQ
MMcp/V67CU/wtDyJWQu/MsSjSp9pEbOFC0j5RX61p3ovvTb4QuNZAyNQ/VXUZIoi6l/oYRYjauTf
8m4Gm8T4hoijExl7cZMFUECm/jUohX23gFUtVgFp4wEiEiQhDQ4nFeA/iFOqCX9rPALyKTkqwE0s
1E75WJVM1JAncB0P1FRC6AyKTELB8GQPFAlFlZEGUWs5x8jgfUWYxZZ09JD1wgdwV+5yIxM5L8xx
75Dz//0iEL1HVDewaGCIIXXX2siNPUZ6htyLN6I/pZAZtVXIzj6AWiJEawUWYMp1Rk62OxoqGO2s
ly/XD3Ansb/ZKEIFVFC/qizT2radSYJUZvWxqDUa1Jc41f58Fm0fUwEIWuJKm8UWsVyTzJiZZJuy
RFOQnHOBReURGYWJ703Bkr+LrJqIo3tSyPnfhX1t6pDLgCjbYjBEk5p+kNCPZBL0jkLS1qjoN8Y2
Rj0TM1a1hbD6e/PJVOUl+A+Ek6mi6fUg2TUHGsumYdZ83oZlFKQUwlyV2BfskW1wuDLCwBkBu0HP
xqcBh48iWIqxoAXldJRycCBfywnoO9+jgH534pNdlzP49gQgK3BgFGjy4kMlgbPQy/6mSEb9tqYU
qmDCDxqXxD72iGuKV0+XSUzvc4lQAme9ImVXAjBKCVH9BuBqzNp1+jHBPtP9B2xEatjeK/iNzC27
pM7l5eQbXra6+x6qmn949xXDJoGpU45DvNeEjCqwEv8ha1QbmzeJcch1qKhdAxMraX13Ud2OWQ8T
poHW7ftTJGLVDyBH6RoTuBk46ghCykSQrLEUxD5LeoMmpWcM3OdK6OpdMb9YbhYjWNo8Rz0teBl9
i4JNOmuvjTrZrDLN7hRH46qiX28GX66ifeXJlBsU//hWyi+5wG/jU/Q5Vtn+QIWBFmehCPoGWB7a
j1w8O5bV4b99NClSloYgL92MlVJ+tUuM7XzAEdbpaRO7njFmxotC+HgH6sDIePKMYD6W95zD3DqV
XV67pBUrtPOuEwQvy/5fwLn5YZSblUCn0ICdT0HObdBez5J4exF2CKFlwKCbZ1BBaMxRsYkTaJfZ
l9jz4brqoHfNgZ22zRMeu79mrN1pQH4j55fM/Td4IZXT0aGKY+enkP9IFLj/CSVzSGPNEKKIZo7z
U9pJN2WZzr6m1f2culKpzzGz8jWI10JW/4eRatANuKvuDs3q/yG1kCsxSVpvfnmaSOXrAKXkF3Ab
UQ/QUBy9rMUbloKaFlzcbVoA7IZXWqvu2GMIBqFtGXXnQftCneXb2UYkrZm5LVLMew/MzTlU/K8N
4KmO1WVUje9SpzvIZnDVW5hoKmwr11a3Am801PKXaw45UgQL0RCXBmwbwPifxEX9DrmvyjYMGrDx
VTtPHpA+gCbE2r7xHhvXLPtWyIo3ZSRj3u0LQINFeflhZmYJZ3UlyGtBg7ihDL08xKLKdf1Ffv9e
VOENkR0Hd6nvJjhZId/s5sY5r0PUaNX229gh7bg6KzJ80tPSnzaR+AEuc3Qllbwub2/q4BWnkiye
dMQ4SSvoAzTWKIdVCuFlhCSgOCIrOVfvlR/DvPHkqu5Dilp4WMLgqmJoZUn9o8UxbQiZ8cN1qrxg
aImHIObikijQvjU/YMcWeF8u7CDZF2iJjU5aUc0ni+kHUVw6gbRFp/uTpjjJknhJUgC+5NZPYDXg
PXIu5YDolBE5i1e3ag+qsXW4nbxt/yCXWWS8QB9wiVAqEs3RoQo+b2EnsXAjAKPxnbrJ60pOiCvk
yC6/pDI3H71/t/RvX0TgNVS1TTLZ4Q3wfw0kXT4PPD9zPt6/K7bxxBJAWX0Fh0TSZ/wVcqsyZG7e
vi1R/0wgBvA7U6xjGxZdaXn6ah6G0RG/XCCp+Y/OQ/FTRXF4gmFrLr4aQJTGvpIsw6sn20xkCOEi
6olS+T6NvVYXfcJIwHOLeJIgduB5DSF07McWQ8FuRsdD7MU0B7lN3rXM/FsnSAXW88gewcyNeDkl
Tj/a7YbPSCYsTuK6+Nct6z1u0cXpuodWgz/wQMUN3EiVsJ6791l4WuRmdXNr187r1J6OOt6XZSze
DRyxyuMMkuq0nCoX76R5Jv7c52NLlfi1yVufj4kCC2pMbaGC/2W4onrHfehKyuTfEskjXAmDsdMb
O6Jdm+eIMyJjVfzq8stYio+1lUmE2TKhJHFfNusIoTjWqmy0E3aZ/+ibQZhZkAta9LbX/XgsJDWC
/RewKO7g7BLp1LVt207QpFwfASzgoA6LAtTIi5bklyPQRmZ5TmvqDY0YBXFKpqNMRrQ2oYbsrI5a
P5EUkAx6cCnZwgx3Nc0X5MLNikQuYC24eOKcSEXHmoENP9cHZnwZJqsnf6XG5fOOVI2Fo27CBGfe
o3tXqMJ/0R/TT7VAEzqfNS2BpL+2JlUWXHNMC3HnZKH0A/yRr9urlmlIwvgbpur9FGGZq8X2q50T
Yd+fArLkwiN9QrwNzrnnTycvdsskcp42bEqLyBV1UM9/O5+SYsoY1FSa8e5Wh1LejzTA9QwrXpCC
3iz4FDDpmqMKjpZfssvsl/Byt7HHKowliAYZUBFHgRkF0CuHDUemShug03sQPn9/O3DbUca1k65G
e5087z8E0XMzTHUkR+VRXHaR6aC9RRiAplYHy5TlEQ+jdl3K3DCBWn3R7GzCZcgL16JzWLCkgmqR
f03vEE6Q3lz0guiip1Hf5QX28XjCBzzHhRZuerYhHs0OkIa8gHH1TzBB/i994pD4JnDko7rqH6tc
KsNtoxeQ38rJNw3QhCzUk5wxF3xLi1+QHOqsSxe1zLkEu0UqPyBl8SZPPxKYDlhlnpMxco7/8+II
cxrzTr9D4TC0zrpTHAZ5lt1fdZspN9nYv2nl+cLY4gmHUqslmLUmrm1knWqvkI+S83U9LpppSuNt
tALitkA92G1rmpjKvtSkR0qPp6ulEeJyXVRM/DnGtCP3ht/X3SlDjQ0NkyvOpTkdIdWFjOdT4NBG
FP5TJv3HD0pgXb2qM0HL3zUUbPMQYimsYkZFi/kquCBG8Fd4f5YOaIKK/gs9NdJaivDUfdgiOiqS
lqu/ZhjQyk+CQKBXfoxWG3YgO3tyiZ/X2ILVxltP1SQbRUgN02e58ZAXpUjTRFDhvpPlpechvtYw
eQ/N61j3KOdeie5XegngFrVhFrxauHDs/wMiEWBUyoBpqqbAi0pQyLRtiMIO7liXlgyxYgqf01xz
E99iBuyut6TvgZu7Vu8wt67zgkq117OO0Tf1ymD+Rl5ol6ox0XFWoP/3pZURzr6CzONfgubCBgQo
VGChunEb1lwlOcbBikOTK9tTvxbNLnjXVdYp9ZmrGTzvSdphgzMlOhJinpIx4YYvcXzUf9A7BsQL
XHVbREhyW6PbIbDabsMShgjVGbCmvHSoDBNZSV8gODtob9pJdiYiXPjsqWSuMn3/6b68SRQFm0V+
8pYRU7TKmqON9xuA660kvePrGmunm/jEeh5LXuC50j/NhtNtgto/Rn3TMYQuhyspUI9qtxa5HMBh
wLvKaSarsCpUA/oD6BtHJghZ3IqP5M5G3fCb6d0Q2x4Y7j9Xtrl7BHtKOFo20XfI8WDwoZ0A+aQy
Ttw9gZK3NahB+Gu0pIwdKNV3RBfyQiVT8I4uA3HGFeYRatG/IzNLZpetdRGDR0WAAhAczpkNPIC5
9hfQn3o5QxR7sMW0E53les24DtyxOnn7XJ09J33WjhZ9hVDNwAPy5ovTU+8fm7LsEjlwMZC+sb9j
uS7dXjFqnAFf/Wo7+RGASKB/fvCM/LaN6L6P0jKqCu3Vc3f7nKD0OCCFToWj7q9a18LGgqye6iHJ
ZtNqLbF1UWBqp0kL1lnEBqGlXB9iplRFoCl3Y2qORqJstVGOEia/e+fuwfA7NUqoI9kVi9mMRgsL
liHGdfZO+ZcP8AQYzLeY0Ka7bMrKbKlZqH2pHLCPv2sVcaY47WjQPv6GI+PYAt/8yADBPC0t4es1
W0Z4McH1KuhZEbQYUGJ88ti0OJXOO/EaP7fQDnmu1gYoM4X8Yc9cXqkrNG2UedM2YweTh8e6Eps+
VHrU+htE/8gMKk891O9kdIbEe3XjnXnKxiKibRXmnDwkjTmriha7tbr1pZNzX4zXiZpp1hR7WDGL
L/YeGq6dlwOJZ6lNusRVpJ9l7oa0BF++Pwh30YL5nx0zEV0ZSZ4cVXzXhVGN1nSBdmU5gPOR5ubr
GyOYV2yvkzcVgNBrmBo8pcyYcLylKwQQPu95AIII767ZW0UgjGOlBWriBzMq9EDmBke8aVykJJdx
zjPGzx6N/40bNeG9vEZ6qIOreogJhsNmUMYJkJd+zWj9557S73TTE3HtBce+FyyiEp/jY4T/TOOL
gDfq0qZMJxSJZZGzhw5ZBYsPlQpq1mxPUoU+T3uVoF8T3hfcAnX31aVPVC9WYbESXnsakVwV8xLi
ccbv/5tYKlYiZYI50pQyjDyRMbROOEeY7qaMFdq0I7ZyN3Fj5HHizn9HwQBxJGExcSs/VpT16QtX
4lyY8+UhjexK+zYwy247sDPZhKBnNt0lD5P+F28YayjiDWetyo6s7Iqw+bvaB/jQjbvOwGEwXC+a
B59pMAR+9rlrHmXydAGLgFOREH3WC2+Ib2hcw8gOXR48P/uI+zf+rjdJR7h6FqGbIucxfB1ZC3kf
ZCkbq0nOLPu8aRpIJIrvv5ejla8dL04D73/4CQBCjrpZCFF3aJ2pdrIt1FgeMvF20NcHuZZEtQJL
XUZqL5lrwNNqTSLqvDLdz/MswYk2LbBjWUX+YboQuPab9Ph3uSVtiTEsWjU15GmYfti9/ccocZUo
t5D/U6b1sRUGGx9GR50tsf36krJJCJxfnAOja9Vs3AhCOn8n93rgjl4t4h76DhCY1aoadt7TIadz
MUmK3+Rc9RcxJZ+HasDjTvJr3egjo/Tm7AEtQx1KfXVt8duUZjEEoRM3uw8pzuUfHZwUQ/pVnvQF
5uDHNr4YeSHH5gy1dqMTZxo7KTGd75nATfNSC6/2mGbQvVJiTasc0mSsJX6DpF29SfC8P7L/BBW5
u3DdX1GeK8N9IjKXSIYu/NvrOv+i3bmPcB7tZmq0E4rl8JHAdnqq4cyHv/ojVr9JsU1Bpc80h/dl
bfrqvdibeX/48NxR/PB8lDlqbM4dINOFJ6dP0VtB6BMrtmbvxeYIDqGi51jU+YoKa3Jgb1BzhUyy
N5UM5uuA1x274pNBvrF3O0Hhyy3q4FtVRZnGVhz5ThJGs8qXZawGerPkAdDrMhfgTJR/FVdn9DB0
281+qOLwwN/25sYW1obTUisvvWoUl1rYHfP/Dgvkz72EKw/f5MYE4Y6dzQEsaLQ981QLjFUKMMyG
gjSDFJFTwPq7ckO009q8rrfcG3rGADVHXJl2w1dacp6YDHLB+Zbvf7VBoUuN1gCipM6dmlxItLzk
9EzrjPJM2vWiMWwPjBwVYY1DLqURtgVL2sKDrTd6yb/r7PYiWt2j5zyoBWZxm6Wi6qY203SWENbE
YHUwsu9VWty+irB1dfDuBp8KzQsTYk36jEvV47YMZItPHuH0w1/CgCG1NKplZGhK4uohyds3k82X
+iDiVHoqJU9C5jfmKJ3tDpnqFr+kA3IJ1+3lzv6Bxm+az89UTzdWtU9KOZnIFx7uwdrpOr/1WVl0
4bgokD/7SGk0j0FQAgsYVpqaBshoxVUOwQNKAjX//L0a9acW/12FafP/i7tmq2TOg5pcVMFPGTZq
NgE3DV/GDkLWH5fLBYYqMivATp9B4dIezOZIemmq/AiKrwpZla3TlmZGA2Kf0AKN8jrL1CUd/vMw
pBjp3jrL7Ce9glVCwepW+ZhBo9Fp+2NuIVAh/vjFdRRODy3TYrkc2XNmRdXz6nyhQ9uJl3IXISBp
+ucfP6YoVqIQepS3b/FAD3vaxJjhJHt14e076YQhvq8OLXDfgt8x/iMXpY6ca0fzsSqZ+Oxg99hQ
pwP3v9O/gJGWoQVtPDj5pBFXu9hoC3t2ytcumRPT4UVeUb63ncluz04U3wOwSaj2zEpzYmJrFtsc
+0BHkWsP8eHVmmEK/B8/ENZ1g+y1IIKMGLReYxF9h+viGgNP58rpVosydERCLCrls5rn+SvZoFgQ
nNc1RBot2dmgllpt5naDjR31VlEgIub4T2fJ/rgo7z/MVu/7arUB+RANBDflj60oUGcngclGq0O1
lFJBIxyFkWxoffDbZthi+x/SVfnfxhwlai9ljbWJMOSS7C1f8YKA/qIXBJXAKIfXQRZA8P8T3dwd
VKKPCcsKyv4qIoqTAyMGRaqwH+B1j+mpB5a12II9kiCZvprLw2xYOoBUlD4GwzZuC2rp+lwJqXJ3
BslCTcVcMD01ccZ6wCGNuOf0T9esCTEuMMqGd3p8wM3r4mtTpFFhr04JoKsaJD15RcXd/WDGU3uD
8wmkQ98tY7QaPYlE+qC3QGlBk+Q1Q/nrvQzE2/ROeeB5bmB3g0NZUPeKWaQJ4x3Qtr78bPFXIqNG
OWeaU801Opl5ZPXSK+ug8UgmuU4wkZ11AGOlrbTqokuKYZlEF8ogDqllia+Gi3zuRdo4XqgpXa02
hIbJI2DyjMoro7kzPDkKMBpoFvH78gkmR3/DA2Kclepc/W8EVPGMwe7GLlVkvUpdADqFW9WwDYMC
hxTpbBbrjYqINo05bEfKwHsZpmjgogVNUuvJUUlzJHOL0YxslpBh7efU9Lv5y/sqRM9qt2EyHT/0
UWt60GdOu4LcBArbl6KhDD/eHVHR07xrM9B6bKyNuLGhxcQbrCfHjWwvygI8/XDoOzgIF2nS04fL
HuFLGl/6bM1gyZAE6xJbzatbcsbRG2XtERE4p9wfBamleurah40o93IEmtukzh/ZvJY1i+axRUCw
+faFpZqbogcq+GASl2AwQnRKP2CiyDTzCVU5mFCW66Jy6ZFyOX5yNXPXXttJEOmjpZMrWWWIq0uo
C/bh6cfNqD4IyyDYCJ7x7byolf02EXxaYhrdJ0B6cKxyZiVb5S+xw1oT3BDDuk7aqmH6ioTHA/+n
IfzlOJa2KetqAJlms3xNWvsL1VWYhCB3DEq+NvTjDHN6qHtXGuVvPqA/8JDViYUYuOXBAD5Xe1tQ
rdUNp0FulAIw+OuQmDBqAqQmqfBouEnxRIi6EwsYxdEKwFQpg1RyVB4AVak1bHB28AXmUUDbzZw1
GSlcGvAjvq/Br+L5NMshAUs+zQEZgpyLoFNZlvA8yDLa5qnKtRIsLGsLhX+l4XLIFQifnhXGRo7h
uSmVtJaxNFNeGRTszn2D1THWgSOY6jVDu2G8yCamqKyqwuzKlBye7BpGLI9bR5modEKE3SLmro2V
kNkIW7+VwKO71W6RQdDzT4s/cll9xITkr8Z0UuzKZ5T/mJkcFXTEU2MY4mzxKChcjXhNnMA6VGE2
nUjccAy6/9O6oLwTpP+DRE6rhgs+lccYRJz+SwNlauFfX1mQ6o22shcL3c6Ky0qWpDDhJlhjd+gR
xvlj/V1iDjflzszOxiUmwbwFdFHgk/ahZmF7mPpZP7HOj6eu+46K9CYn36gbE5AxFD0sBVEJnEbV
lWRm3QH7mZHlMxDGDVXYlRWpvGAp9mMsgAOVTDv0puQlpeO547ZFl7VO/hqDwykYW0ly57JjCF3u
hcci3B+UTjll0oqJpv0Q2UF3HoCAORCPIAW58r3nb1KQBn2v6qicAT00ahKD7s5soqedjRzzY/fe
NVDDNAQcifjd9oTtSVDFFdL3VoWR80L/aSgWZw6zMRy4rRHO3olKFQtRhZWAc1RFuhY/gvuSbQbk
2YKEoDU8D12F/0uovyWlisEz0Eytw0AgpqSoGeqmGJ7u3nSzLtF4Ithe8TcQ0/3LLxYaQta01rLc
lss79Ynn9Ga9/QIPvHNxkNM9HMfrJVhIASsZOtWOr1l1AIf2BXoOOv5asocfbrUaKPLuPD/MaztC
H051boq52IX+26tWSKN8C+kS6bgyngrf8zCLa6ff2LjcWeqIQXG004vd1p8Y1B4i7jZIv2thWmhG
KtGXAjYd69tbIy9MONjTaSKYco61NHMkk10Tu0KY+ny1f0Iq3ejvBaeN2YiDsd4wdCcxaOzSkN2D
1K6vPSCNV5HDKCCaW+/t5OImudfcSwWzBHunb5pcQg1EboBPxdKygq8iFaX2LZACYGzTh058kNOu
3+ihvUDi2yYI1KZyXc8cnPAedXviO1oCDL29pa0EJYujJeJEPrEBPdE5pBKkWKHyhG+BF5R7GBu0
4Ydhp2UcgrfcSxhSR3OACebjTVaXItk1WPn/kAMVJJM2VGFLC1zC/iow+gvkGcuTD8feFCT48p8R
Sl7mC2hPwaP1SyuI6IwGt84CWnjA6tfjiymO8WMIgY/i43+hRldMMMx9C8At1DjL9adXNAN2r12T
WYf7rmb4OGKpHdGLZhaaB2pHcym/p/+Qw0iOWG4Wojl4d4H5yyFDicdnWeMlvOUHIMjm8LXwimsA
OsIjGmazN0VIVAvXEwnbWkG+qCZLXTMgE4VnHZO9Rt472SRJ3OWjGQ8qMMX02HCM0+8hlAT/cII8
pi440LsLezCd3D41ngxnwmSqEQa6UPPqQehK0q6a5VxTidqB9rOHUflhCrHGCyLTLeLOHHkGhHmm
0fbb6IeAwMeZ94Yo4c3+0IvdXJO9rcQge04k15FClwzB5Tt5mgLsO/ZQVZ1NGEB99d6MHxun+/kv
ve8PJZbq0EMTgxtUauXCSePHSmXMKxFOUCD4SRGkn95B0f2DqN2lEHXXZKmES831ZWFW/EuIlf4F
N+VUYIVRnVNgAlxEYjH5uZDgCORe0jpxAoF9EC2LI1kGnQfXQrfpygRTVljuAtnpBxsY3Tdf5H6D
cq1+ux52tJhydQG24psbzla6hUileNlr/TK8mgEMo+PDU0qwaAPU+KXR7FHL24dx0Pqoq0l4n6zY
+mUKFQPhtEdREDaHNYgBPG10AHSv84ZE/VDhPrBFA35rWbvKabna8LtGB8pgZ1zHn8lzXV1Kf9cf
t33BPoq+aUXf8tyTpoC5oHBVynqEsxmSADjLLqp5iDvFvimTOhO3hUd7Ze/HXCdqe4Bi/FII0HIL
QB5FKr+htD45OSi/fUWZZLMKKJ1wtVnZq0erktAbwRxMTXSxJrtLF0ulitm2PfKOdOx7ERexXIuh
CyQDqx9QxEn5YkJUEXQrSLtLb5ob+RjmHyuQ+/OW3wmsuwEgv+qhiENafJAMNdu4yhWJO60z/rmK
IxRIOp8BiUqkkZ/gdkBVqO5lqchVPMudwHDTlHJeh3yn+qW5+RWg8ErpawZwz4CH3FpTtv0r2vyO
eQEaeRLThPohCGWzBVLVBMnIwBRW73y+rjdAH2egmAZOeLEhJwuqlHG3TlBMok6ZHHt9l4zoITIv
+JXg0WXHhJdxmdMVoHoRj0ehLfvTeRRt90+CLiBLTJeRyO04zKa1bZWacKHoFEYrua9HHYM1qWtg
cGL9MvGi4qfQ4ZkeXbfuYHnYzH16KN3BWPmK3VUOMSGqxf3PZSU3St0j6EOxNf4p+sBKooNYF/1/
AJEE1OSb4REKayvGvyHWe6zBtrnk5O01NtOp9KPuz/Ky+312wajJhYrpKEywIag+A4cyQ5iY69LV
e/KpurcJ55LLbNwRhNS+SVqQ/wdq1ShMzw4i5BV2R/EzEmJSKK6sHeUrL/X9lwHJkT2tLRbCh9Ax
vnntEq5p/mcLiv1+ZqjjW+jRQJIlLRdLTGCVcJLfx152K4OLOt0pDokPF9BDfQ0Coeu0hbyOKH8y
HrmVvZOLL2TzOcipd2opUk7rC4c/LqGXl7VFkmkbxWd9W68LWIRHARFd8nBlFBDl5khmtRtKJfiZ
vMiaKvjOVb8dO7YaqN1QQ132C8M6HAqkTSqtSwjrOBcwpRiOpRgmKPLGzJNcXtdn2pA1F3BxfnLG
kldMLkWGf7NV1BMIV0QEmmdbSEvK7xM5yd98smvXQDYMQG+xTnd4k9TXQFjL8XjVdKugk1xd8NqQ
0LI3eMtmaL0qPYe5O0G007pHiuXZP3QvH/CbHIkTv53N9X+8r6gVX0BA/VU3WBc5TAqRd0uz0QlP
MwLxcVSVrWxXdqLu9b5ksJPbnVWwcG8ST/wilpyp5nZHvNGN4DmQBYa1hf80rtr9N4rKP3ntq8/e
R1zOK4Wi3ABwWLwhvbvZJjm+WzpmPv1UxIwvm8hEf/VGbd17Y1/b7Ds81P/PWjkoSKlduU6+sjIU
/G+zbZI1q5x72f2+CKZCQfnSbBzPpW3TQ2eoZrxHW+R4JxHi+fRrlQQpPfFDJio3W8vW75nslg6Q
RzIWZDZHCuPNQdGd8MlEBynhjEGvuJ2bswQjtwPNVCUfwFha3o6wBoslm2k36EwVQ3i15ytS+0ir
zDgIWtcsim0feLk/+v5hVnYnPHPpCKvXmMZ4ESyHHrqgOKClVlUz7L/lIxROoQS7lMQlwp0kzp2K
pi4vaHyvhEDzD1wFTxSCs+09zVOZaVuuIi4uMNUdwvfNf2vyubuXddj918npo+qezrj4YJPQu08o
r3FYpJZ0VnQnQUUS67DMzx50kVLPoJs9VArLsrpH7wt9WC7Y19KhkQE1WPJ8yJ+v+hK7GjWp4YKH
+xq3zUSbThZ5/lUOW8FJCRFqzpocsPEvF9/3godZPsQEFJa202l+0F/0PGjm3ysZN1EO0MGGbeAm
VtaJzR3jdhTzVujnw+JzMHLe+qUQuOzas/0ODpzCTpgSKbhDFNOkr3mSLdRwPGuTOO4+FcKUVaE9
HKVtZCNPUazIxEGxaLwXYSzFpaLTgz8hhO/eiZ2TvZOkbkzH7i9ShDCGTiB43cqnBv2qSVaUZkHI
uMfTd5aHtgPrmbp9z4r7VwFZ6MthzYFNNCsI1lMRDPBs/nMe1Kw/gJ5Fp6HCzG+Yp8jZFc8F6LO0
vXOkYtP5S0NZcJZt1p0Zua9DSe3j9ywYSXOb4ObAl9eGXPjHy6s2MLzH0D5eJvp9iQPqYDERGZsS
5J7BqXYdS+UwqucgVz/DlfNmsTLNrxUtb3SvqWw/PPYnHSLFiupg+JeG86btQQ+eBAjqW/iDw3vA
7elAo1Ldk5Mc0c4qJrOiiu5r8B0RSMnW3rho4cClwzUusj8xmpkHyphVzP8HfaPeQoQnsgwgEKGJ
pxULNddOxN4qdUqF8egTnMtL5OeXaXSEcZLTZcSVbNlStbTfgu/1Ej+NaBkI0rIKk1MmxvbnhoBc
4OIZlgPefUm40iAU98EMemfL3+/HWRNtEtNCOGqyIsSXhbFOiqfC5JO2fqzRtRyxIwJBYsZcGpzf
xmDdhO1sT2G/Pf1OIz3I318/DBD7x5i8EKvKyj4cy3eT259mwhSkS5LFwGaf/EGVyIf6BgAXJkkS
97a7xEiWTCl5Tp61Pxoj1nIJ4mfqT8wv6oJLeNeJaAJTzNX6HKWhItUM9K4G3IYVIAKc2X00FTk7
74octyQCxHkHjQKctkAStKuAXHytc0XYa8zP/EqFxzb9BOfCLUPB+i8Tla3OrrNgBgT1qpdnTkRN
cNWsS5z1qbwf1JIMEAyUCWLOxV7jymXTYrbpNMfab0rzotSptVQCC3Cc8cW1Lc7Z35Qroi+XzL9i
acs8ersyH8MDY/T6x+eGv6hRe+Mn+p3GX8iQr27qjDuWZl+n2rDlEFWXat2sRIhITIF5ROJx6M+p
bhWOpO4MtJXDh/BCiqWk2bSTsasd2Pqt5WHd3Posge16doQa5B1onnre7m1prBZK8C1Gu/8R+MLR
DaUtA8xgjiyKXoJU5dRVNuSK/DSJSVXjaSj9+0ENfAyrq0FviefpfekiN6aeTUHKLvJDXyyioF1Z
IlPrA8IRZWj674abm8JfH2kBSMS9V4NXzFLp5O/eVUGOCkK3rV9xO39pu3deV2Ay0t3tqjX6Pkrt
aQvtTxlZorgt/RdAuWlJ+FatzAg6uhK7C65oYaO3Jri5T8CZ4ZNRhABQQXr6uC1VIO7AlOyWBPlX
vLzOxau7D6laR7uPUTNAjRkMgADxr+ydPpT7iWHFXtD3O5PFtykyLALDBW740mISPmLjhfZudjXp
edKGalPFeKq7jOUcXlT3vq8CKr0Vs0qw3ii7rFlWlmMQ2tsVtrRp+nqrxsWVBZbnH240XqFs75kH
nMysxAN94ESefb1Ac2Ob/4xRAdKYoSt3wyver3cq5s9xkfqn82pQt6Faq63oSpPXBc+G8XzHwB7D
JgY3UKfD/H6Se36MWphC7+AD1PSFY1wYzu7R0NuUEk8aYIw66f56xx4XLb3ecfNVgj05GZ7ghFPO
ppkQNPP7GUSi0tDhJ1M72WHz/FdY7lCb1yJsBvzlqYJKkNy6ogroPxIONKB/TOVKP3AoYbZ97WzS
83IUC16j4mm9gElra6d1LnDIxz44dOPAityRk/850hQXcN5M2Fu6apjR4EnQUKMT5rFGUGWmMGBg
yYavM8Pnw2rF4scObIzCOc209VEIL0mUP6qO1C7wqD30Y3ckaxu2rL+TGsosE6TQQ3G2GSUurnqh
puowtgDgck/bVhIC59Z8R4ta/q1bcIGRkoqFujZ9IIe/96jsr74ujgslAIDQfeJaGPjsV51V53z8
vK7dlYktT7K4AKOTWoHjHsV0OMZhYSzOIHWnoHPmRE85V+pjUNrxa77GuK2NY/GX6/3GLO9xCjU2
DzSTTW1UwmnU5WfE9SWhHqp39sAeLvr5MWILAWxtb5OWMUCvWeiXA+lccy/zERuM2F5QTbYgi459
4FgBvJI1O7HoAp9YZmDKAT7lRjy60lNJACEISSF2auK5kWXFq4A75Q2t+TNMqJzYpiL+BdJ1rGUU
V2D1LGZK3/EJrCHPLJ1JLhItiQ4CarUU72LEifHDPvE9tTkrILRFDURtswXA2PLMMdSaWwOXv0Vr
P7FQIDreAg0CPDrASsSW5Mbu7630Yxh4RxBkZDRpv4x7qbYu8NlCcr96wrYbtfn/JKrLwQFHGkJD
EHfRg8pop7WCSKdJ2w3jV/RG2LobNyk53lhosezJ6lTX6e81w34SKOJ7KzJ1OLDQ4JJ6OfNF/c59
aTvSIwaiSPQyD+cyyFL6Xust7CYAZOk9iPovbqzLRH+R3deXNHG6IwlVRR1vZJu04MHbz+VmqtvF
eDePPMar3SsSBvhy6oG1EJmFfz59TS8l7qYjsi/m8Pu1zqMv10lAwEP7SyhniYuqS9ZEseuISCIW
uV7I0rRgjCubL3suUiDL+rVhr4aKaX/Pe5DS/f/zy65GJ5Qi6cUtFtqmTWTUl20bWF8q4VVsl9vX
rAMLPi/j865Bnc0JOcOQsPPJ5LQlWAk8L1t/bfxc9HxJp3UGneFohHJgSY6aVF0Xe3XBOq0Fr3cX
mTp41+C1/Hc2HFqnmPHMnoONtGjTPEpPmEW7hXPlNm0Gn35bgEt9vnvTxP6lYtiU/FQdUAfrUEOY
V8oxiUuO+NDmCHk2v+ACVlsZSA428F+CB/bP/Mc6JI+gyBH69Iss3+weGqEm1s8hgfWvcVF98Lst
K5/0XEtTEkDIB+Rjz/tDwt13WJJph6eR0IPmUwqmf0EcrCIky0BnksjmrJOxpLi9LZWBQtjk6sIP
PV2k0NjNWL1kfwhH0ekFWzE5rD0sbSU6RFb5KLrn6UgtkZ8yX9Wyb8pn4+KLcYGYFF1E4M8RKH7h
qA3741lTngDd3hajUT0ZeLvr7dFFrn91JpBC5t74LmoKCUzawTvedhGUA5xTlEGb/Mlt5eFwms0b
tgrLB9I59RHIOKChdLhTrrm7/hrJD7BpsYhydT4ScPjF4EeeLZ8LEFTB+AJ8TsCyKaENAqjKcLxF
Iqtlz2b/VGlYmr9oUGL3AogLzjJwDsJ80wvADMKd1qYR0PyK8Fe5cluweuKvf0j1kIlEhba3dWME
sxvGuAIm6ymEeITRVt2XiG/OL7CAVH+esNjc5WPm2R/+S8KvcloiKvYAH2AcYEAdtLO273nQl7WS
+sGPvs7ydFHIRF0sQ0lR/VlT8sSdxMBt8kkTiKo1aN7fDWyYL2V2RZIRgcM5lfbKBGlZaALsd5nO
EZXMHfADTLqnife0Q5mG8mX9LHFulsSTx4DHlWgMOZavRKo1rs3IzaUVmbweNNTK81h7ZYLzoVnJ
q95SitXxiJzeVMs6SSYayavQdH2LI9kuCX7nBIMM+HDwDSWxlLpIMcRX4t1SjWuuoVYBkSeGXlEM
w0unQihXBRGUtraoY6Gp+rCjhcSXzQ4ANq9uuPKNzn7574NgcDNgFXfviIXVHNuCnL6GT4Rt2Xfa
bsr/lTcsTuWB2Yy/w7v/eRGIoeCfPAkRh2Ij9PxcHQreaP+URGGnKDlqjStQw4o2rq8BJ4m4Ap86
C5U7LlGb1CgdTTa/Xip1+24xormNz1Dd7KATBO+mP8i2MuqUStscbdzHuZMQxGSzszvAslDHt+1l
t2w9Qq6u7P+LWhYiRzzdVGRoA7E//GznMZzjqiXFUsZDNl3kwQ5Yh/GqNG8ojcf1q/olZV28FvZw
lAxQtG4EbFYJli77bNioQZk+Fpbs7zaXzzZTSTdEInYmmLUQ1n7ENFtdnLa4y6WyPKVsF/3RJys9
5BEHVe3dWeIf765nkd+crGM1CAofi6Km7gm2E4Ivlm8V9CEgs50qgyMJvuM3ccHGmgX/I9hMTuYS
7kRI/8SGHcJ1aPomnrhU54+0zXdt4+4VTHtwtzJnClXZD4EXLdqcZSVmTlBQH4heOdfeWXUOtS9R
t0wwwMbIJZIoxsYkVXRfy30wBh/rf5D+rQfARThPGuiHr6GUlVcui+0JK1WqmQcCf/UKKcSZWxUK
HgKr+0XveSGC5amPcSG8+JpmreEEzhUNZusd/BeDSZuwDX/GECDmjmoxcStkoroWBjoPZXK5yukt
dfn97IDmybFXoB3iEaKaPgWy9qOXyXRs6oIEvgNady7U17TIL9iWW/HLL9PhIc/8UMYtrI4k805k
QDNV39I75jDV9f0KWGTuS0oQolxvlo8zlvEx5Heo8yMOD+MNSCJeJ1hB7KxNDxS5ZpNkUKjEx4FL
WGP4Zjn8UXl4I1cFCyz8UEp3sELZV5vKW6NjMlbXV/iO1SFeyeP5FpsG+Qguphoe/gpLEze3dnIL
y+qlGOvIHz/3PyySNWdM+YM4jilr4R7w3pay9Nfff7xNVM48dwtshbUBqh7SUtTJvm9EAuql59/P
cp+EbU/BSTXUHTVVqePbBu0hXYTZaNdreZvVwF76V7hnuO5k4KP5VKP0H8fiGUssoltI9SjeY21h
4+QZUSxrrDJNHpwHHZETJH6bpBtYngdkFy+Caof8gWiNDgy19G0IBV1fVmZQnchAJ31qFefJqt1l
cB2J9Nf7VD9n0rmH94txreo2fmv0b2L7U9hXPwUCx4XjqOHiCudRYLpAPzlM04M6AzzKoSAOmX2t
XwqQqLS3TzSuRLwXmB6nRvL43Xzp67EXmStZMVAhuO+yUSn+ZMvL5SBvFzeancLDOkzIruQtGOZz
54zAmT308ETaMqOOreagbzBkjh2RsWSTtP5XySySubwR7ZCUOmiNiy88p/pNz6wF863ygLJYkJm7
75l0rM7fsDWBjVb5HGkFQyNA5FxTQJtb94VWCB4Q1pm58ek79UwOpIIdFnokhlrtXjBoS399nMaU
gbu/V8rErCsjY0451sQMAP4JUCT/jAGPUZJOF6LeZr+etQj6u6lbPTquaTkqPfk+payMxfLX28bv
ZisqVCGv+HBjrmi7QJJdqT/F/L+mRABXfSYYhM1mfEqnB3s3WYEXd3Zw8bG7xLi+SrqxFyuC+wtc
iYmjLUGl7O7fSb+1CLpwTHyIoceCqleDirUgVit/twTqv8TzItnr9bcbqkwlhfzQi+eeZHJ8DLr+
uETIJzf62bve5JNYvztHYnZvgNO+ftx7SZsdAyrEawsA2BQwRao4kx8xVPxcCUSwN3FX40z8za53
yrdFPg0dmpVlT3pyiNX3a/3nUVbXtPz/zgrsZWKCNojKvCMRUGn8jcSMW+ZeGTWGnf5e8loEyLBy
YxpfGxdE8zHHji6HjCZBm9JYdlnlO9gHiUPxqqy1j02R07VFr9aXCUlEArtf7dIpQIzIlsTLqCqu
cSEayC8TuftZMh7EicE1Q9s22hpdcq6SG5v1K0RafmYJl9NqGG/Iw/LtxxD4Ppjqm+bpizhTrhNi
o6Xx8HPQUh+iKfurIDFnD0AYGK1ZqTg2kuy7mRnIqw0lRzSGli2OhkgZHMWpuV4cGy19Ydm82BAA
ndqYCdv4VhiNgJRT/lcDasOFHLMMq/CsNYMvs2mrarX5d09Zs9U2hXCFf3+gt5djO+HIm3HdEXei
Uio1C4DPJJRsULjPdFQ3SPXwVThscvvmDUpDh88M6pYoo0k/vKF4x44ZbE2bmHI/dHtYQ+PCsi9o
JgCEz3HDy3Td4/Q4ifOO5euknRd6oBD/QZ7q9sE+psMmZIDIRogo6TWBbuGhRbzUixGaoY5Xnnk+
ry3Bdh5UWsDnI5JnEboj0/A9a7de7dagsHrKIpRcfILKvbV4qO78sBrR3wO+7sZMXXXB/k3bWhMG
0un5btpQ+27ULukGCqzo8JhJVEb6i0uGXXQ6lnZQ6WOECP+5M5fT/jb1PGt8HCmehzI82Xx9zLQS
UtKTKzsBL6/sRRIEw+nfSWdr5NmJujfHuyEzdPM0c61vy63Ceay9G0e7t4AEnAuK45r8dib658At
zoQX0McOBzG7Nb/D/JvfuvKxeLHAHoSxYKFDtQzI5zpC3OAxAvj8DxQFv6eIVa/ktmw5noAya17e
/hUJ1HT2+hlxTu0SG5TzF2c/Mk1jiYI5bCFXfR6hhcsr3Ewn8TGDz1Va034u5LQ1NFEFEokdiUx5
vNxy6hjwlSt044JaIEYsg/c8gdLXIvC/qGF8EFpIF8eXTfjLmGPM6AGIBUcyKT4Agihqt7juSJye
nOjZdXjcuMnhem9jk8RFBdHAUC5YvHMJQX+3RQ/JIfP99vsXcfVkZOyIZ7aZ/VNFflfAfiVHomGy
hi5Og6tkqJQES6h+xkfK3d+lNS7h0D5dz4bdqFf2qGv+F8LhzxLHZpwA5Tc3wQIM00tQl4uTB0tM
+nMx5Z/m8n6qGIOlv8wIdnu8YsBcKMmUbgPjkEdA2BzH7+9KQ9qHLvoqBfsFJsMO6l/iIt0ogejh
mhsNQIIIWtCzvLPrdF4ShPuC65EE4c4p4CgFll6djMQ7MqHqSnKz5S6v5hWAnsXXXLpD6h1Bax2A
cMO9Xq78yIU1FK5tpB1id3cpogoZPUFPwyc159oxwd88oZXPcSTnF3qJnlqVM0601UkY1cZ8nDZX
ZPzjkIB5123UzkbSf+hT58znh2vZPuF4smGC6bdWMQI/sSZuLHe7NKMyusmUrdvz0k7akidoSdgw
oKdWjfMCYJXdFoILzWIoiJLn1UziRzc6rlF0jIo+9QQgeQblCl6S4u4lntytA++IQykEVfelieYI
Vxw5+OpWDTVa+gSzytCArsT4ExO71vYjUhEM/RgL2Pj3ZIGpsxTbFMp0+M5SUX9AfOhSmmyT1Zjk
FyqkjYc/zfzloTXfTiWvNfoue9xiNJvu8D1neTV/zD6VK/BpL/JViEyAyBKBcRjpksAWa33aRVne
1kWmS12GNYn5yTfFbPklG1BBKk9n7IKxtmFfaD9j7daGR+u2gVAKvqsOHcvNodLLIHiqDxoR/TsQ
8Mj9e6KGrdJ44FlxTz844WRz6dZEqeQlyzPvKzZniY/L8OR8KE732PdU2MY12Smmx2f2Vy9rgstc
J0oz1qAiQnri9fQ/3xHZa2sSvE08zxuRah60T859cVWH7TNjwbs0p22Jmn3+EpGprmH4UD/gK1Cu
ududJ5LVcmcu6webvsbdH+5JcsMYztHAQRKq+Afgj/jtdGGjAjF/PkAqQKVOP2HlMSmDgJk+m+LJ
E/U66vffJw/j2Esbx1/MGzF4c2riWRoaeBEgj24ILJFCCERLC86x/+yhaF4AJzycD3z/czasGkxk
HZrTJQ5EC9KQx2hVcwG6Zo0NNRYa/h+FoT6JgPMTohq5cIxnroPHTpfopof88tMKRQRinmZBwjZv
aS/eAe3RJgJRej2n7NH1K+hqQW2unDnQ+YPiJZsFKHG4KVLZ59Eo9lTqrVW/Cag+hejLi6D5yZZS
Pu02IVzIGkxL4GLSBzYx9F872y2uuY/9FF6SNZyzfT4xf6BL03LBP7FYGYjc5b/moR4LVl7n5DX0
TelPncMl03mv2RMHwJLtTV959LFplqpfXA+z/fcBrSpd/e8f2TOwBHV+K8eD+ZkEA116iw+w9r90
qJnzgRgJeYeTCkY6sPWtOaTXdSifLrUiq6XG2daupuy5Mo+4P7sjzBnaVzZZOEFGUTITJYDbzo/F
fyW0YTE6jVps8nnbLbM0Tw/JuMlinYmXOUb2oSfra/aXgRtb9u7XoCJxUmkAkZDVmyECsm02M8Qj
YaZvyPlHlQbdiGxpI/16Es2ERWSw407tygY8gpjq7DMo0q2pp5RHQ0MFhb5NzuG9cvWKWgAV1QIT
nKMl15kmk25haphyOpUztaKYF08jsL5zgk/b10agoS3XYmSMmK6jtCHFqLXrqy7tAsuw3vIky0mS
dGPC67gSOyXft2NVdNDl25Oc96S3R7ox7JSkJAjdHC5gOPpTpEs6EKGjNutVqrG95l5ltSFirSYc
eOJvduY2aA5mmGRFOVp3QKBp4L7wUv0PfL1q526ZfP+9SYnd+EZLTy6j2DLkOD4bVwweFUI85Sxw
XUBPoT5o/Xw0wOfWUX8HRUqZHi0x/FwgUj/CHD9G53VpJqqkAsg9ajMFGg6BoWLpzHs7Qc77hcyg
vKo1NBs4uFbngcy748JS07q2nQrZ03qjbpNpvh8hkJ8fDuaOy2erS5qWFEkB02A4n7QUzAjkDU9J
qr0riKG3lvMJ/IyO3APEdIsmiBK9PwO2U8lo8d9yqMc6VEvNrC+QdgorAXQhEg+4nus6qfAxxAm8
+CvHlClUiPtzARe5WGAe31ROO0/yDjbaNhnIBXxp3jgCK2pC+g93bBQ9R5ZkeOGaYsqJlBiIn+tc
MJIImxa7tXFmM2f6jVmbFixaaCf1RLyZXU9C+8q3ZaHyK5UwT+yD9Z5M7+iZ+5pJEjGcjnLJiwiY
tnKMNVYrR3zkChEwypKyfcdh9s5+RJvtpQ5V9IYCYbRngyhGT6cLzSTcGaWlThpPGR6/71CUQZQi
jw6wUfMw6UB9/bnAPHru/jGbBrANwn3L6HAaqS3NcuKaFiBTefacgmI5BP0+VJYXVUhfzRniLff+
LhnsQ/TodBNeX1ldMrB05dl2IpVUOhwtaTUAjrRR0RLfFVjZI6bG1hg3uy6FxakEfe8BnoaObv5i
0+z+cqa789VeP/gbTzkjUTpWso6PcoPQjEW2t2OOEDyR4i3yJT6YNMs86IIpHq2SCUHaTCkdCihj
yROXS3pjQ9KX88uP5K1jahB4u/2T9sks5rfeIR9lTaB5T0yCp8Te36mj862VVp4gOleM2sEY1OeQ
5tjaU4eGjVmraQ2pHKD/3UtmoDijkngUzjUO/ANv+e9OGxoz2jh3QpyNsn7VICUXmEmI+lqe/VAZ
MIeKWq9WtOLrANKpral/K0ihUYz0qCNlMHVR05dixcWB6ivfSdQI6po2O+8IelUxEEAlKlpdkjmi
Xop+35qsIDeRo7OP/QvmCbrGQKYI2HcVB5QzkUQzeZuTRz76bys9ELIvZ7Yz6gubWquxewVbs6Yb
UCxw+cpUvjK+5Z6mg+Zul93ORgWpqZBwjjiYfdJ6glQbfCtMAhW/0/4ovJt9VL4dBajvznpLWsZT
6fGFTKWsOeFroUBh8WaPqL3wIyzKOfKaqMdAX0oBylt/K9Csp85mFTmkzmrAviyimbaLTZlr5iHR
IJ7C3OWU0YT1oAXk7isGj4VqxLvqULf3CRT27jUvAQ5LjrsN4mPTpK2xNkBLpsWLvV+YoD4QxSqw
JwT1bRMgIyGCHt29/1vuEpgWw4OYGHC308SHdvoU49IZ4xlExJ7j1Xkuxx9BRn9GCiqbPqTPyvZv
3nlzMd7eyqSzZwYnf+zw67QCMX+W7FIQrnzZCOLfnE26OUtLw/HnmzWrXw4JbgeBV8Uu8UmHMV5I
1+9FaDE7xGS2LLHln5NjpjD4TC4Ff8Q9bo09kEganTQRsOkDTpvQGe3bO+1ksWfD+Q6k2ryx/6g2
Q1D4183hq4wRH3s53dS/UikBfbb/1g8BmVXqNqHqA6UCDb0jphq1sAS4/DmNM4hxyy+avcbb1Dbg
l7WjS1oxmvsY/GIdrB6zSFDwiuEW/KF8yFHtTRQxY5cLE+bI46+/2zuWD8/yyvU72d/Fd3YHykR5
fqi6D8rZkWbrUhSDVD2QUdPLzG5dmpEg8jgCxfCHRgQa/M9HWgQrRn35bfIFJe/skN3fInljv/8x
aeSPSo1cMVjZvi59Be+DModB6Lk+tNFBXjMUJNDP+X3nD2zi5oOinsb9tWO0egIt3W+7PrY4lEgq
tQhh15pThbUaPoF2UIwtcFnNy12eZHB9xWg7vhamMCso+kmltV4tE5Nsu4AMLwW61hIOWRd1qSr+
JDiXszXW+O26s0Q5BmsGpp4DyHIlKxrCr4mQaDdC/ePjjvJMPCvccS0s9uLJ8EM0ZmFqTldG5KsK
XMPS4YButoiwvlUby386b5jUO+MOv4S+SwQuW7zs5Ce3RF7HxAkCsGV0rUTIBD2cBArrye+mEu1C
ZkZVYijiZad5qrI0xg1O2RfQziz1dK/cAAsUxgJa16yXN+ui9adBSFRlap9OgqjarI6dW2/CTnL8
/rg8W4ptcmBeOKg7Oi51E6VFPJywyeebT9qBz7eEvHl8w5DOGxzV1pdl3XSQ6AFgP+YZnx0EEMe3
SdeQIFgSBM4ZqDzL/JM4bXOnIlfA4ljEA+fLMef+RfpCX6ffeuSJB4eXmb37yt5iLRWdFl9ADpxz
/z/py483agdSKxc5MKowYZpxLP00a3TrkNNLqRBOQTKDmAPRRkM87IVibU5A3xnDcYdazqd/+n5l
l2cXyGJZaiNpLjFUWT0R3FegrrS25wCYSVIk4GBz1OMaT9qcORrSLm9oZrPbZKIXP0zNSNqqK36u
Z4VEqkz/Gzuyrcg9LLm4Y2+90d1chYUAovTm0umcMzJW6LuJNtnr5xoRDxYcSrdpT2lIzK0e0Hqp
Q+gPC37Wsi6Oe7DAMBLrQgtYvQSkqeU2y02BCm19A96589LBwbYQG3Bu3hCKwt5u/nFfilZUOYbB
iB3mjla+H1YVFXzWamnqrZlsgjqZ+senfisdtUnMsmVwFeKHCDxvkfot6TsJ/zOmKj2dQVl4izOE
Ji6WWxgk1ig1QEzeOLy2eJDvtn3j0Kk8MXLxrq4odkfjbN24kr6+eNpq/cdOI9FGx9uw87f30nwx
St20LCI6ueljMQI48bieReOYawo1OgmcyRXn2u9G3e+Iww131/xrY0tVBP6hqJMHudzlzYfWlbHo
276wv895xUzq8ngbExuRcOlHkRGtV7gAsjkx4L2SBk38IzS9/tW/DEMC/BKCnA1jDYhLYa41uzks
+T5IYQOUruZRzZXAx4Wpaebbt1YU9XxKRhj5uaBQhMIyIWfueaVBzl7LgdkwtI2t02NPa00vzaIE
aCwYXEH9eeissOa09Zt7HMGpbm8GF4yaggA5gxWwlWq1EzLZgnki+KON3PQ+WTiSE5czInakRKTU
if12h3Ygl/8dRK7E+IILVpBNtF7f7xoj4Y3GbPug2NCVyG3pgBij+amUW+XA1PerZ+/XcUTeCX97
b9VfOPfOyCh85XfyNgEhgVcMHHu/hJFAvJdFwXqjH7tGNyifCY6XR6WQIkuC7SpTMMnG662zlAqD
Hu8K6NQepPMiXgtWRHOPm8OpnKk0S1/WGA1i8AX/grPX1rQga+gs1kC+yZKfwMKKIEz6qZ1/RtDD
520XYswbFkfw6B6zJWRR5bOoqK/bGdG3+Hnah26yO6oBct9QWBtlzj49wAXgprm5UDm8iQPiGmDq
3zp/w3/rhtcuqF0vlYLuY4FHTqbYTAGLGHb0DSyceRJDJK/nCACD/mcbEirGxh2h2HB/tSACXE9h
U5Kx+ttNKiEpFdDri/0CRTQ2bthFCLS8dNMao1i4z0fptso5g+5RBjavl2X/LL81yO2Sxk5YUMmu
TE4qmaqG0bD0/8L6OaH2k7TMHeuw+cQnzliPOxKcSkP2p+6fobAmbLyFxukmUlwcXu1TlgaqCx0r
LcbeI4QPDeFhTOhdD6fpv/5xyoj0xfr35Z/r9dJKOHIPvQ4ArqyRntMZRaRwuDrykQaDCunDfjl7
rNO5gWivaPI/Ri37gdlWPxVYlHYCSEZm2D36shw7vEkWdu5WPhzcwH4wGXoi2Gp+gjBRE5krvLf/
KHxk8My6lSY5NNwUXufKK45U/E2RZHy9cD3yttkvCPg45EZ9xIWDFnEe5eXqgCqwYnFkPEan6pFJ
6W88gQU6NaYahaMcHKWMG1NPqbz7+UjWtmrKWuDzjIYFqhjJND9wjwt07ntUPlCtnlQ+BmsLQXTb
FV01ikt4n+pZuCHmSDnk0Rp8RoG+/JXYMXSwrW1BaS5iyDBGyd8H0HmmMLxRTpnzWFow2hnq694A
MISStfEdXplvDNEjaknlJSKlhh4wEUxnpteCFRsZtgdnJ9XbivVc0fLmx+Yws8wwSwTzGogqhJod
grTNQeGsZaGfuP6Nbr7PBmuhqn0rVuypmzX/mQRev2CbDbjHCqWDtUmG4pgB7MtH1KtMW5aFB12/
O7sSbTm3ABd2p9k+f69ZaYyQpWZkuWPQ/gYFb2SWOrqPO5yoPjL4fEG3J1BhkdWdsWCtjvyu/0qj
YU2s5Uc90KVTkPTh4Ranljn1KFlL7FvmdRACLnT7bd/u09ufMKlXpZGsdRQIli2j9I7wvAbdSn1t
tMMBuRVuZtA8tZhW2TmENWSlfHSXotoo5cGF25Dww9vuCYzNsvvk3CeSaS6kh2rZIzH2p4haujx1
+c5ag6GP5KH7to7h1Lut6yhpafHtd5lXzuzrY3uLeY3VxcZejGgGAe+gL5UveQV1ShBEES3f6nKp
2+I/m+EcwAavA23GqdWkKkLEKi+Lz+Td4K76cBF3EdnK5rVa9Z2rpuAT0nX5y+0AV8WJ9xN8eJEp
xFwlKTEfynb0h4LfTGTjz2NvrG4YT9yJYwTWiT8flg1ToG+E+UUVFXp4DgUl86MqyrLFd3CnGBEi
2UM49nwn7cfjrtUSeSuEuOGsQqB+X0hjOZ5sdE2oAiutMnnHQJyURxNEZCjs8B13Gi+VUKVzvywt
SE/twHucr57h1ihP/+Ha0O1xZqWjBEyYmKphlZvf6MEQa2S9vzuUJSD/3ATau32dJENvCNMzBtGQ
GV2yOH3Uw2jxNF+EQCsSkKqr4/BxeyXAxyRfcPlb52197lD9h8EJOor+lSG6LtSqIODLVuByxDwL
ko0+3zfEf8LcK8QbPcD5mRuH7QG2qsrTdOeFz23FcYxZef+A0Zza5Yxd+HZ+j3ONL2xkYgqWzVzC
58LE7BTcdVCXMAR22cSMmy9IO1MfIQ5U24fLVpTs5AeP+B8AiozxKheajIPu4bg1WbegfZm1fiuu
Ywd5qmr0Q4azuTQJHwAMJAMo6Z+fbwpkr2uKtiAoh/Az19PWesWnVw58JhG+DSj+U44OsScpX+Jl
Fjve64nUateBevFXspw4dViJBRh5uBuST1RtrBu97gC0WOOMI42L0eCT9I7oUbfQQkmTL/L5t3Ze
ValZBkkpWtySQPq3NSad77Td+ZcZnhVPx3UrDcwiqxoLKPzKExh+yxOtqSv8wg+K0a5Eugh/qQ07
PDLzZvk4MeOxdHCRxM/iE7MrQxd0sI1IjcsrU5CXtlX1Bqm7AEkAenM1WXNEv7XhGHbx+YJQBx/f
t3KIpxNvI0YcNLABeGS8YfIckCVRTTEZAjwDo0ueoGX6DASWt6iXC/oU+ZwaZ+Xc1UX+qWDey4A/
HD7kMYhgjNrXY4X4HfWbbGtdTqp4HLaAzJ732Uua9/7e5vNESCn4XUWkiMW+Eiix06wZ8R41kfIS
jIGBtLKKIChVxL/QS2TJiMIpAF60kRJ7spN0BBamRoP+6/3xF2FGVCxouNh6rLaoqAD3Nrw8WQ5Z
4OTVG36Y/C4vUTez1WMG8IrspQENiAx8j9GrKxRhRhDOiqcll2xQGaYjJ4vRLEsPDztZDI2JiWwp
pjHR9eXYHJyo2USKd78h7VGsWieiXjFNxFyo9Dkp3rX3julqqZ3xlWDRpsWPjuCUgvqsuBnUoiGw
VuWIxGVNUhVonD7nXRUjnhfT9hmWCqDG7UpvdYQYYmAZb4u0vpUI8mdTVF2lR7gYCtVcCCnmzvm5
Bdj1Y0AhYMdjCabXk9KtYgo4LKTrMkAFb4hb7P42AFOcq+KcGgTqGnywF2cimT1eNPO9VR/Vjvo0
9/jGRcRp75M2dmV2Gu5UHTfx1y6kosAjqFSjwEnUuh6gJfb7scLk/4h5CnueZ0kMz1MaBknKcw/m
R1h61zEhc36+vG7ncT9cAV1imRuC7QvB1tX8ALSb2aWo2UntVhYc+sHofQTpvYXQnuUQWFz8RE4+
KttWBozQORcQt3fVUhYURpE63k9v6xoOdx108Xw4Z/Ltg+PkNqslDjGv02pwuJEYpgkQXIWiI9WS
W0GJKzTHHGnf341noIiIc2iQKHyw4ZbR08ImOUnCZT3Pb925d16LK47RwdSHl3gnPYcmswiZAU8z
4eCdp9tAx0hOTG55MZ9wE1O0s17d2pMclW7/CY4HvNQS6asAIocG+sGLrrOGqjM9LiBHCGxwoW6Y
I6Yy7tiIO7Hi6Me5fJhWqXMOyEgwmtJ9/BbaIbFoDFNQzxE8c+UDXdO0pAU/ysFshrFyG7jxvAzJ
0g0afaVuGDV72HCt53nUgBhBHXAljDyPfslN76gEvw9qm7ZzhVCedSMiyNLI85t5A1xRisNc0KK6
qtfGoQ8YMOzAXpIz6voW8MhZTOVgGTAP4AnCKjBmBc8B3sqrZYdNlc/cm23ngCNeKwf6qo3yZ2Q7
McZ5UEg+4AA505USJpSjGOQSl3pElLq/1jSEPfOdXsx3Wqb6r0nnHikbdCQWmo8CsiFZhTp5/JJs
dk38JBqVR14qgGcSdgDHesXpma9Y6N2B6Wde2Ddq/iTQRY9Q/NDL+3hnxluJlMcK9t9Q6xADSXY3
wTZBIlQZ1VuKbjfCM4IZlr+EqsTVcsJgndWR/FRWAizOtxHE/YBx5j+ExZIKyA3qIl9pNMRiHsPU
SHbgioZNj67ZGSgePM1m2UW5wWQYkw/A/reZCJsvFyVLE0516vsaTg4aysvytyp4HB4dN8hEoOLM
dQzESwAEfOerTwqselayQeoBFTVNTqW1NY0Bruxj1q/x3CUgIMbRkaRsoOT+hus8XVo55/D5697h
Q1O6jfUBoOu9igtP8STdjedCM5dt8zLv8FJXgaedckkedA7pTYpGc8ZV9zAzv+Epm4a1NQa1kytd
8aLtzBc3esULuEZE/dQYUe1cmvqgY8+Dn5XNas2vxX2Plyc7+mRBjugzqJs+t4hgSU5coDPjRgLA
URNVIJr8qIzBCTgvL6o5u0sfes0d+3aw2LctAj9EcF+BXWTo25fJWNZ1RuWyFb0QYJYKw7qGTDBV
yLDG1j02EIc2pzT5kC2HQqi3UUIKilHmA8YtJ4VAAbEr4vo+O+k+DrHnmGyO0B9nQr4glUs8G2Mf
TnBg1g8dGM3MA1OO5fbQ+P593YJAAroafesKnXz6ToLMLkec0krMMUiKyqrAr7XoqXIeet9bTl1Q
RzmXbx82t0B//+HfdJw+bNke2lMlYcOraH3mK1TNLB/Stc3kH7x3Dk9ziH6Sa0cZmxxOFydMpkr7
0kR4wNDRTu2RFrkULCNcvnGnqvBZAsS1v4r8qXzKHm4cr9Z6NKOoHiUU6FPlXlWW+3JhJ7frBzh/
GnP/qxzEkTnz0ym5bPaKpaJly33aSE86ao7L+AzULEODGeXMyHRWEcstCFBdxE2AB3OiXCxVpzXQ
qwXz0Yyl/2Elni6tDJzNkUoHj8tlJdC2akitw1k7lwQMlWKmDBVlOnMbRBFeQ+duM1Ccm8L4M2W8
bHfGYtU4ZqiG6XmOlPASHE+GY6iUq7jWJP5dshMdaG8RX7JTMN572fQxgk3OT0G+BfyPvT3lup1S
R5aX7+j5iHmbkPPSA4oKe5DnA3W7MYRgnMPPBJrFiN2EYKTP4aZm1msaaH6VELzRr2/8OHrlLeML
NVQ5TRkSihfq9PlOP5hkW7AwUz5IIZKOBGanf+soHvoGbQzfab4icENyQZwszlN5fJMum2QoDlZO
V3m3HK+zqobLJ3OfGLDcB9SEiDhDXlqjHUufzmuhOErzzmXb22cXvWmOf17ttFFJvZR3U+q9Meau
YHV5ORGfzYBQniKLWSxVwAJ/LeXJyjc1C7jkDoUoYV3Xf8jtzLKqR0nDSkq7fos8fd9P178GL37b
+wVIdLRlWfpRq9i4xsXUXt1+hi87U1vNhcwX/tQSu9VKIW+BbH7UQvXGYAr9qeFH+YslPVV2Hl96
o6jOJA6RHQ3ahWB8Kx/gcMbOAYu3dnqq/xTdpL2eh09kt8ZSbQf912jGlIa+jyYP7XA6LKEjfkfD
BGxrb+KP+j/S0kLGqROxM97Qqn99b2h1aILJcebtequsukcuQaQkD1qwwl5wdMMQYq3rUP48kf55
/Ye0fhaZEWlt9s68kTRK5SHPOzYLIh2X5uzPyXaLX0xyIUYaDGj/g0bO2Uw7JhVXWukpNt3lv/UQ
Iy7SsVJvW48Q6cImJNI4PfM2/j2sit3BukKe/JtNs3n+C8y6ZJi8pbmqK3fikqsWdGb83y2qjecK
aNN8agCq35/ckGKKJh34ANFz/HLFFEBv+/ULEqXb5PadGebpnCzX5rECkUGbGzvZ0npkOd2DBk9Y
3QHoTFny8iOvbvYRloVY5cFuMvXc8qffmPADHo/1WyVrEa2nG5S64QQwW1kis/TNoxyFZpN0jdvA
lRDR1OeEK7QGmH3IHP+Kx5G6CMyQFgA/APb3hQoeE+2P4wCMvAJJNBe/BbXReqCsoJWwJ20x9Pfc
zQLY4lEgZUSOmfWVG6RSCh+lIA7lp1rIK+b+ocmBZcoP1BMESCtUmAjNE52ngW97fDwbXiVz/hFY
PgcT853lX5fA+EMQkL6WXYPfeXHpfHNZZk6sbpFPhefqNz/VlxsUd7CVtlTCBMJiLzPF2jzklkJ0
GDR6lc3FL/LrBwjHIk/o/Q2wV9Us6O+j5Qd/6DkT865uhFB/HohdpEVMtrz1SgEOWXCsrx1q/nCy
ejyiB1PtbblpCAcbPEij8c7Z9TslYhCwHe8ThJz6FLwwUVvZcLW/ACFx+BRZ4M4E/6OIaD8FHlB5
X2kT3W7MCBhvf9xIMkwzM5gOUooKMHBB3s694v1ck3kLO8zqF8Te+3UGT7EkkIF/IHWaYhML0+kr
u5g29672/06Rd67VWzvlvKLnwFVAgD8eppIGcnTQZ9dWP4FbVU0uuFJ69TYGHurYP4h6wIY57UdW
2RDnaj4PmNgO6GzlnB5hTzbly3YdJoVehhf6bFx3++52GYDKLAeNUI2SvQZmt0OL7P3p9xE1wiOF
sRAm9Mdu2VbeAmt9kJ9jK4obb9Uv2fAXKFeItdm0FgJH062/GwWsUVm4IKzdEbvFykqTmo17yYHZ
Ke93gb67MOnSouTjgvU35iHKYc/gXs/7xFZYEG8K9njkFwk53g3lGlIj+nt9ug4LSmy/SvV3WuaX
yqMxLXdQlet5eCCRDhTVQHkCFKkcEF9+0p1ziL3ZQcVYn+KVcTNFTw9zH0YubauZyxV/gewepcxL
hmPcfEuPFG5JjjlkKvtWvgrEcErm0WmBFDNIzafg88CjbEWT3M7KBGS7TwEnJr9rbb17928VBPoX
9IsYBpL+9+6PTsFYZVBWAbihPSca3AOZXNwG0Zb6FdHzj/jhTVOOsQiXMlx7ylqXsrKaJIV1DC6g
v+jprX+zrIsLQOrzTMcQoI9XSXHinSzidnToFaAp95ZwV9DNpea0hdgIaiSDqnpXa+ihr2CbW/XL
s80jmMCOy72WJDfS1+uEKPnmFq30uvTR5WJQPxCvDQx7jX3cw3Da1xYOQZ8Wjn1UdjX5WEvJm9Iv
Eh+0vrnJ6Cx85l2J1Oa+Fx9cr4TqyWcyo7n78SrAsQsYQYpA7dmrXPXrZPaVKjHQA6S7s6t4C3LX
ZrP1UZ7WbcbTdJ/5Y3pKyTLQo1j6GQM9EbphF+tfC/JEwKL8lVuDFuRlw81CkV69cBNk8L4hV7n6
Qvyklx8qIM9El7upCO7FeWIBBZBSgFs1DGSkU7Pn9+uZ+ioz3wbuj54IaELK3ynL1QWtZ5vDw/oz
ZKn0tdoh/jBVp2i81vaySmelMMP/WzzJJ9c4w1zz0YbLylMwu8HrE83jzyibk7/3bnwlYcamFdOO
wfd2fpNoQW49Qp+r6uP6R50oif0k7vCxI3MlA+SGQC0/SQJEo5Sz/6s0iB3LsBs/SsiGfcCWxxr9
4WnDPJkz29v8eOXFnRU0ags+d/wDmhI7FZGvNuJ3kzT2VPtNdhblN/JbaOWaIqzFvhzr6OfU7jZB
zVIbPOrnJsmlLH6qNVG7QBuoTVeBvT0npBJfsSzJ7RrngcpRKLAecRRkholbkdHWdaA3QtaLT7iY
R+bQcKcAkI6xtJ+mlkuZ9ePAAJ0d1GpmIqj1HUZR+bqIjnp6QzIqK/OFSXf9QMMO2v/x5NSdNZMw
oYYIXQhP6gIwz6XGymhJFM6rVNxX1BcQzmS9RkOrJ3GNWgaF7TbKMo2cqI+HWScxes+6Bww5pMhX
Ef4ccw86rd2HvsAUFDjb0B4whTBa4xwOCHVWAghZ+krQ9iMmHlEMVSjj+UW+5UBByz0WnAxnbl0C
Gz76CmfWcnqmaui1MeKdUk/t8D5RV/kril8sgknoxG/KwcTjaVQ6Q7RCAuymZ8wRgCWdqJAbvTS6
wO/QVOkCAHVAodxtgv3Qja2R3rkRAAOQ9Sdg3jvtM4u1IAJw0dJOEd1JV7bXTqrb9cYFRv2Erudb
mmMjus1nOShF7wxsVJpzCyHzuezcPZmz+JmRuOjlrQcPCF+/l8T6kkhCuHRm3DzCOn1Skjn0cxJn
q5BTrSn6bKmGZ4oFcBM4g3GsQ0DKjwjHVOPjrjsSB3XMKZkzOjXKb1pH/6UG7aBDOfYaNrDg0QMN
KgOd3YqndQ8XEKphn9fyl7wcWfUoXtFDwCJ1QsXeeTw78gwS0jnGaIPbUlJPb+Vp9G9Amm40okTX
tWUEIQsZPSjOKJ8f9BoxcanHvptoREiEidlVcUL8s6yGH2/086zGxub6HCa8tHZlTgf7UcOOR4Ja
zAINxScn67Tx2gM9Rl1RgNtcoAFcYLL7Sgg2PFoV9lZLPs++/ChOaUJI1k85qWkF+5qFsnbsDWt6
QdimKa7suRhCM9gFUulEF0wTddQh7XITnc8I3HGlvZa1kymN3ZflgpvNpduwV+MCkr3+j4JfWJ43
q+hkmTABe7AxM2okwF0bQew8rqM9bo1RN2OHS0+fSSS19RDN9+RYM3s20I6VFhqBKNnYLhWRwnYd
2NSXDzUt/JGk6jkBWYiKO2SgpLaYPTpFTjp2lTGj+MS/OsSy8Tsmv8VVhAeC6wa4MjynNl/GR40O
XaQWFzFxvNaq0iUBYvKDkXbwz83ehOU9PPDO3nqMmkcEgEzeLbCIvEQEfjM9bb19Hb7Pxp+3uPjl
iDtf9BDg9xH9dwCUYUrwrIhIOmk5AkMsVoTq8aVqfaYNvUeKSVN9stm9e04qvZ4B/zNJYQD1Tz8R
nrrywBaML+Yf7w4M/0Z5rcWhx9C1nDONBbJEMfcda9+unRDp3IehUPK7HoJNFK6ayJ+DBacYimCd
BcE8skBMEbs8CrtmxgkihDyQlM6bCmkYXxSfyH5eQalmhN4lq2sq0thZe9Xocybpm1c9ngugysuK
BR34GWb6VbKm7U07vCimjc7PHee9Y3xTrWAW9iGQ9XGdBtNzoYsA3XJ//rjXMVFeo0Dd15MnWMFl
bmR9QA4J5TEKGNbhxI2M+OJkkeX9rm84SKsjYF7KIz/+sbQ0WsPRHYUiLh5EyqUmOL4ztBihcJ/y
OF/T5uzG8MFo2/GB+wf975ZJBp0viWSUY2fvQo2h3lUkURvgikmk4dESi4nRUYGAWZojrnoYzCdh
aAUhPXpAfeJxBd0WO0jCrYYwLuQB3ph6XwQySKj7T2qt7257sYcJ+XmfMS8rEPkmqbW0SXp/sZvn
IKb8y5cnh+pDWxwYSjvI6CXOxZw8ei1vZGPCQ/CxIzrDVb1lUJaJS/2iiZmEFelca4G4rZxFNegE
dNTXfXeI/ZjTOGvZe7voO0QIv4Izbyp5CV6fpVMR5/lRmVjNA/iAeWf1YBSf7od7l5oBFE/3ma3/
xwLz5hKGTPRYwSLBkzQ0DvFUxe1G1DYqkWRWNG6mltRGXLsnxN/kMdP8dSRbmZOwk7Fnv6TANcrj
u31D6nK/LCxGKb7bZaIqQQjucJ84VLRiIgsRxn8LckWZh1sgKdRsnnEbWplqImr+/P6U/+19I/io
J92DSd7c/iya54UV2+I2aoNrFba8UYu3Du4oqTzOz8u+fL9A9i0gaXhynBEPZ1WeeHgTb/Hkh3i1
4awaYMiL7Ua1tTnum/zsnkKeVB4mqig8tj5mFEXDu26is55rWF4nsjxzEWQqBVwPoQoF3UE9WHoE
0WOIZKLjaxzMBgGdfzSlmANLBm50DtvCe0VcoD2XVXu8dFR1eFuYT2sAkefAoYi3k1DBN+sCo50Y
PznvGvjOo4y3PHwoREbxhRtcNSOgEWLLjYtTsJUeS9YFOfMSmTPt2bZMwirN8xJmFy+jcyT1mu8S
Na2F4vau+BKUp1fZIdY6lR2fHpwi65EdH2GmZvAHkMent4IlSK+N6s4sW13dLKo7oDKGUssaKsuA
Y4lHa8fDaIy/7rCnVd6TpENqL5TnL3z5zCslcuLq3zO7Q+nLPDFew5ZTxBVDARVVG9kySVNiPx5X
kA/C90g2J7JEh3nTbClMu3eGkVLCmBjAhoO2nnsay7/SkOxd4AS5VVeXWDOWPpEIdI1tnVfVlSh6
LKVipNnJ2XippTXZ1IWA/GsscbaIwwrWv6i1+s/d4Hx5z3yV93ewD9/T654vrTle+twYR0t4Tfls
0Rjg+M1ngQvF0Y9JmUdoFExpi6H+TlVsR2ZvZyfKvhcGTW5Id0p0FuLbA5KSeckaO2tiU5UBEpNR
FDyCqflgsvnIKglK3unFEdASZ6TGWgNbNcflPdZG9Z08tTW22lYI1S7MDWsa7jWlMMrmyofMDdup
pVfqqPblWFi4YhqbOIdpprMw3w8y2N7Hsr8J1jslM9kwAMjUqbeEf0tyfmZ2De0TJKrG2Ptnvi/G
VPzoXHc+PypRI8JEZE2sCoz71ZaIl7Zh3Z6zUk/ZmT5Ky3Xw/fWfLIkYACIVJhVBlyUQWoRCwYmi
ii60ZrxowazIZQrPgNM51N0CZjMyfK3k+wfBHyq8hO5qE5RwCirYbMDGCXs3rS6X3oGgxZs/WRCw
6PAZPuGp6QCQznz4oHozP4212HSuJVUaLVcu92UZkJX/FfnIc39mK5Pa8dUtiwTX29kUQu8D1IH9
E4QU2r8RDMigo7BuPITmhdEEJ5Iv9x8MVvLTWGeIdStfvcBNSEFduQXqfb8rVsl0oyxi9mpoDxrq
NAEAvNMoLY5ImFP5yl4wo5VFpV0vb8cPSIsT+SImZw8MimdBY+EL0kI5nMPkTMT70sSAzK+exoVV
NXAxXaR3Cjp3r+lIMf5Xaj+3R6fQU8zk+oYq4UXQ+Q8DwezoZoEWLGwQ39PsnsvHvaTApgLu/BFr
kf0O+TFjnM+O436WdXsCxZTetyQpQ6UVD6pyTy14W8Y7DbHPGqR2KEn9Pzij0WAihlTTiHZ1qbEs
TnBeC4gxnbOz3NCAmDqNrXMtV0l5GM4vA/SHWqRj6pZedz0l1JYvsxwbyJlrMw0t8Xfe/y4ncvYN
NZsAF8JMHW/5yBqMVbSwgOTZ0cy9aVV5Wayec/ViAWrde3Omc2b654qaQgG6x8xVAALRIiElK/ry
kLMJ5tNPnHKBQLZX7hxQ96JLS2Ec+FzWw0HYXUpNJiMVk1aR6egJHL1bUOj9vlEjh5deaqGIhf+M
gIth40hyY7Jp8PjYf4/N7z9BY5nLeTBu84+DPWv9lrd+flIIrYw7wcJzLgMFFyvTOP5hez19WPVl
GImjB3nNIWUOR0v2iwsuQ3iH9wdLRtaSXenuw+obLzRBMS6lWVI3SnS1xKjuzeFzv9XUSvisM3pT
uB6iM03qsiBmqU7IfSjBDeOuSr9uxORMypuywqksRAvtvj76hnxGTTxUNulAMC+jqzwie6Zj2geJ
T+QPM062VjNFIAA7DD43WXONkl7+afe11MlIqSe8+bdSILQ4EIu6sbboPP9tZDY+I800zIql3j+c
g5KiMYdDaWrPo39eTH+xne5Qmlw4//+p59zs31SKfKL3xypgujQeFo51eK6O3WQsRP+4AGdtaMGt
DF+nJ7NnKQ0MlUObqKQjmRDY0UQtB+vcnxLSqMuUAHLlp11SqbKiYm1UEOY7yh/3b1z73S/U7PVt
0fiS/hR6XGVO/PaxEdtZWGJLJGsbMRSTe3Np0LTDSVToEGux6hPnNCupKb+W6guE38JrKfXYF3ho
AM+dNiOCJTJxQmVKcCaE+e+6ZSDXqxDE9fGItpWv0sngsKg8fC4HkQauo5M+JHdruHyQMMKCxVZn
zMXorCNiYBZx1ZwEZ/jNvQa1CgBnW4ffHg/zR99BbTE6b0j0YFt8r38IlZtbakgTqKToroc15KUF
ENiW2JpUesU63pgH1cejn7j2Jwc3CtDYqZMDbu7y+ACKY9UVaJtKtPYaAiLp/fmFmUWYoyK9MiUX
TSzOxBmzjLd3z7moXbBeC37RwzOHDOYgGpbaukWg16WIiMT4u032dtOVgdHxlwayPezIZ/ENIYIi
ut/BKYt2wTyPjBRQ82o/2VHkMuOKJlP4L8v2mBgIYx+28UuJGgIFpaUZZt8HWE5T4QZREy34msqd
3TaJ7Zi2ej4WIgbMRS7CI9N6w4H1ZsWaouvsCAq0yZhPs87RPG4MYuNi37F9KRkhyvGaZxO2ss5D
KPb3ch2XVdNB2a7WFh4mbOUV+JkpabApIWWRUhCMT/BliKAyRnklkbB7ZqHxYAOYFlCBvIz/WOkn
uhPCidzNbcWz5w6yb9uLh+8igUt63fcsXPSHh0StPpV9FaLqFP9931V9eTIPC7aiF0noCXNBePeC
Tdc1FCJccon0GpY6d5jrFHAHAt6wPYKmgQPkgU62Zn+3iayfUH2gT1CVY5l4FhIu5kMqHHSrzF0q
Y8fO3VMvbmPrdB7902+lZ6K7pheRO2LGfx9Xl0Od9r9u9Q9Cbz1yAl+SamBWh15GpbD+x4GPQyNH
aq56csgVjaFCGSg4XvRMhGXLtcabqfsHNYVSAuhusl36VjRH4tLcZ35zosnp9P6L/rIbK24QVrSw
UoDwf+VKWljpjSYb+hgjHNNR75SJjncNMsKx89GyRxVNB6Ez2Lcyl9sucEXJzOet9dddZ2prs/62
LbfpiWBcXbsu/tAAPBKo4Aw5Af81Mm9W3eN6LXwzIvyzSCsi5HS6DFqaCtFFz509Zf0b+T3qI5vC
+Uz4stydonBDafkxZRdM24/0kIUzZNe4i5VDeiTZWp1hIj6Y9NmKVh5fjsH9SFLxpmNnNjFU6ZFb
k/G40PldVOQsbSM03m0aHx/ND69JMRJERjmgVyFApWY47dwn7dbFYWR5f44cJGC6XC3XIDdinNBG
jh2XzOSwyikBjxq871ogBVU6Pg6BH3XssVkrWDCqUZ8w5n6flhsAIwcKs5Q2Z1gO3Ibrs9GEKZD+
v95+4+wgUb/SJL0TFVLysF+Hweglf/KgEoKbJXt1iMiDDMKOQzlJuH1j49MQWUsTa0DECwomVNFL
e7zjNfZaVRSTkEgy/G+zJPKLBvzuDql2KVbXrmGapYM+XhDxTWpkTHj88N7mFyC6hchLXx1ZAKU5
IQHZIwAJ0cd4sM9nJPVThfLcinVxbpjpQpjMwbIKq4CZDPX2ZCJjivPvnf0CXgCsFlHHMw4Lftfp
Hbtsi/vhwMY+uTizirFEsMqA3b9bZ7PPD+qm1TjtI4DIwoc+ZO1hQfnXouNa+w17JUM6f8FBpxL1
A4KEik6Xs1s4+18uqA8Gl5joUofciKNuVGIcwMoKSVxyqLjXgykncJUEcga33jL/uQ1ArPyw/uEO
K89H4F0fMAuWzlh/5FkVCWX9ZeIZ8yV5XxuciwTxU92wMK5NqgG3jMxKQxVDmTkRwR4+bYWezgym
YHyqjbXBvcfyb+X6c3b0XgXDDsMG8KEfuoeAQ9DtV6QFCKJGi+aM42zSCIVyFV+fETUUsyCEtqWE
eKH8mwnWEs2wql5JF4NwAClZW4vLy/Pep0dRU/+CZIoy6bDVuEJl+ul7LbN2pmpC6XFIcMZ6muRE
YYCBKl29zk2aoLnyibsWkUgel6oajsYDrgbegbNFNYhriTh5emEEzFiaQxeEnozPkbOSU9lBtMX7
PiTL5wcH51evbjoXlOJ9XI8Iv30IsXgX6LZVAvI9HiDGRB2CCF96/uTKdogNdUBMRC/Cm6zlCY6p
2kLk//S1EDFzFSp8s4RbUq8w1Dx0za3oaXp+5J3zwNIdZAqeazhAezc9zAuwOKr4mLhM02um6eK8
rMFfhhrebpuOmGGZoJbN2NcjLR2mPJGuqNebQzlXGZtkMUnIqnpc7LPBGdtWrxDpKYW9S/oUb00x
5+frTbeM6KNQEr7320qmGVU39guz/KBmKQQBBHf4lfuiIsQgA9G1TpLQ9KbietR2ccm52zYciZkk
124w+otCFmhDrBbveg2QL/WbMTk3sgswqhCX58cqkfOC/FIBeVXiIBa09SjGf+T+42zdWL2TfWf+
0E4HVcurGshqPfp36h7dWJJBZRW6yvr5S94uKbOErQQJZKbhKYWoJ+FU7T4htyx+INah5hig/L6l
KluzSK3L9CzQEE10jsc4/18RgKxB4Nor3k+kNOl/94rO1TdbQv7my1DGUNhURtXOc075xrTzYiH4
8VPPgozOVERBo/zDK57gAs5MIAzjh7sCRWEr4YxzgaxaIuDl0udPa64mcNTZvDswEkMkEjRyzBvL
ANpphqJN1k8BkBPc5Lq1dT0HhLKcZtfq1SElxjz5+FwDV2U26Zdi+Qc/hIyxJNihDE4P5Q7sWz8l
sEy7x1oupxC9vC9kXVAGSBLZejG5c5L7CiWdVyGIAu626FG1AjTuxMkNHmE20lQl2zSOS/4rBY9U
vHXFWHtyZbThhJ8YsuafDP5AMqesEbHzoGRD7nVRyBsQhlhXEKst27mnGl0mveLwWnj8c1YDvo8+
/IzhuW6cpm/EOa/Ovq6IO4sj/EY72WB33JnXX/uHUF/UDcGaMq1q5O1/nw9QSBPPU4yyHOqVIyX3
8wLC8nE/XpP13Hcfytp+bXFOO6qgzkZXsakvSYmdBQHdIxmNUlmMZB1BPQGazmylQSJaOXBNXf3m
ntJ0yp/pK4sz+sTpjaBdi441rY25UxFfn7OcqDXUd1ICNCPRFChOVJEgXCwIg7gQONXtmnLxIRU6
9N3iH8rEyeaybnc8YL4S5q4aUrLi4+M5LL/1IDmf7ohjldRblvEPb90fGkNAfuio9JVmnk+2Lw7h
jNWUfzYi472MC7KNvgv9PQXiAVrJgvMKzR/yiLXofb68edMH8/r+PYYA1IwKqjj8+YX3SeuOmJEN
8ThGdgYGOYBfs8v6zE7mQoObTnmQ377RqRZzUs+pO1e3mNfUuyxB5ijYX8f3MXKDQAGftimwFCVl
1SuQI9Vvbfm0Fjirf2bQbB+Xvwh5pD4YTDBJ3s/6bk+6L6NJPQ+COPkmUWqA4AL4GzqAyZ3rXm1P
4tvvKG3DcqJ7d3Lz4WZyvPVKt8tbmzOfS+nT3RxsKuEusubAUjp8gQqpSq46U6F5p97UhJiJank8
FvZdKVxYV/5NJSqlT25Mqfwd/zdL8e7YDn/uYba6ruu4kDxN0i+xltULMNCmU6v23spqSQWV1m2m
Oa2baKd3RL1mTYuF0ozjMBVcTt2V3+N9IhcIdTsrCy5aVFdrea8puW3DBHiIrCW5btTBCk+kejq+
soCEgqXU7/xOoiOFtvAsmxqSn74PGNdIwQ9+c4X4MpBecSH/5Z1LxRsvl3MT7Ix67QPVH36aSBr2
kSyf/q3KAkT905OKfRKTemjArYbctS+vF/sB8E9Hh39ksKtb063TBQwXAyLcE/sA5v4rhQP53Zp8
YOgeHKQNUJ8FN//00WqO2WJgQ7kXk5NmLSg1wkQaFzZDbo5fJQt5Tccm56NZtUSJVmbd0FlLL+7c
KnBv36amyErkrqj+Li+mqJevU1gcNOd12w9uboPh3lQaEZ1f5bCD2BiYdW7HwjAtWi/0N+ClZDt2
QuSsRMWV+jJVGNmfTQZ9C/7inC2T+T7cc9UflIDa4RoAaNdy1hfsoDiGioCwAOwGCTQnCy0B+gGt
WDKxOqd8zSER55BK9g5tQnHj5fH/zr1tyVQVuXaW3sdLDcxG57p7J2YLg9+gsZn3QpKZ1ce5wBFN
2Qwd1HwGmlwvmD1NR37BlZZrdj6nS2dRmwHrI6vtEXYkmbct+0HBdk8ChO1ne5OwqPuVmuQog8LO
1Sb27pcnoN5xgb7Hli7tYSXPnIpNM0M1Bwa+r2uHSUYC0GbLBbzd0aTSsOO8Vc8nA5sk5mt0S9u+
kCLna2aZPAp6NlC/B1A/EobcxCQb8iRFDsR1Ncpp36FhQTgpGg4twWaq2N9TMM4wruq4yzjMpUzn
iiq+kVoV3q7TuyuFrq0oPHfxaZNPHU8T0aMjdi5RTnl5eKZFED4wFaok/LiOSltaYIH+yOV7xhnQ
kckMQKGzdSKO82u5JaGRSOv2VdrVE6wabrF7zjkMr/7w/41PY27SlVGR6UBDftUyEos+CTtBPS3l
02MnQkzaWZr7UuaXjhYCgqLIp0AVsgpVlbwLSkX0fjIwGGQf3OBjVL1tXWrUHKAGWhQlXPtlM55Z
Z3UdMqJCh+/m5yFdK2M5CD5IMtBJTqDbZ6ieWLxwAbxJZcV8qRgEoAb/1SRfQ8zL8/tyFENhgN9c
6WPpKhc7NfwkGXLkMDnTrvQ+x/gfaqKRXKtrXdC5miPY3oNAtr6YbcCe77flBdpQLTatDv9ioziN
Enb4mTpM8w50z2cO9+oIQORiomygZe+iyneP34KfXohnoIrm0ygM7vDPgLZn9fi5VPPFM8WfJbCg
OnGN6n+5vr7LGT3glJsTWyE6PoYoBs2sDjB0ZzLrF+rb0TYVlxv9GZGvx2NJAjxh8XH1/5+gEenx
Ro23013NFCL7kntc/Wp1RXE2CgNjNHTSQbttr4C88CUKCSidaquvziBmN+VlocQxAN9Fvt5jzR/L
9IymiJBFAAc+FXlhgCIoA6OYNqTJ9pbvqYFbzX0ArdoCTfQYHWmUMoIEf7UduUC1AXuk2jmz7RJ3
q7vL1tlPs1Pi392zx34GmobiGUUHB4R0cvqnWenrbA3S9KFYn7KQmfOZFgfVQCbRWRcM19BgncBk
8raOu9sy6vg9ei8GWFlq//qM/YeH0iXKHoPG9mFIwuACiQyHmJfhAvccP5dnM4H/JDfA+lO/28to
3hWmxsPCfCqUKTmkU/4RvaMf7Yjq++8wcbh5pnp54US+7jJDt5MKQhym21K4BClzFfVvwYPU9IEU
0DwOEzBgLEBjIaFptGxFS21gOFUS2/EkjeC/0440WRt2VzaewXBK+2IXJIppoOSO+Wpw7t9EdI/V
caqGvsDEkd3voP0Y+JCtzo2+arqzGMWxvJfArJPOHm/n69R4tad8LOK7MebvKZAIXbndgiwzIEV/
GYe8pF1zBCgSchsH8sOxRO6Nz5Hsw4m+AP1VR8uNKRt23udBnpKUvKXowwkS0dL7kv2Z2TqP0qfU
at1txHjne16EceojzRNgNuTbpmkjK3CVO+syszUu/s7nbnYfCID1Tge+DLy9Tvpf0C4sRwBIjHWL
Pm7yY9kLSjeuTeRnINfYzwB/V3p336cbKOzOtPhGJ2Lu/NgLD2GHrQFTHSz0Gx2thaBCfclEhzSB
fPvoOVwzA7x8oSuWGpc6muO0BLQmuYRrAqKlJrX3/Q8mZwTZ1tx7urmGJEQz7D8Ih1aQtRCURCDc
nhMaKPz1Xbamw5n3OIgZxrgC5jOXCe6Jwk09/DUlmHIMv0FZrW7I7875Bgg7C/zR3QxwGv37AwLw
FMbtVbiHOIGC1oFkFo/2eMs0/03k1R1lyRihAkEX8Mv9UC0Ra37+ih+NTbCLNdx78kCyy+GneKwJ
AnBNGcN71ipyYIsND2JTZZi8NPMALBMqPPigVg1x/qtMsYFyMrdhu4u1zoq00pCus2bA8ee8T1VD
W28XTJLnMepHpS29PeqjuRP2N9ouBETjmqCqWTWIRiZpuGxLcU3AmL1Sla8n5btpfQ4Lf1eKgAWL
kk4hDVXlra4qFQHvxm2WkAIYT1bTJnHe4VEV6M1G+2TREVEKOzZ2KGH0MvcEQXfSGpwlvF8MWBbR
7MVWdUW/KksF8TWKXbjV449mN684wTM0472N7NX/oT+Q4L+bnjmGedtSmL7i6YG4vYonjixCEfSG
HS8Vyh69/lS3hg5FsEbXzFT0IFoWeouBPXwmfSD/Ebi/P5cu2uZA/Rszz883lqVUQgrJfB1fjtOR
l0TOuvrxJw9PAbD5+R/rOxyO6HcJ7oqCDTAgtMDB5zL9l2nxJhP6sOkQdQ371FUDX7ODWYglIvbS
TiNUfNSahwXg7sxPQFEstTZISJtShh4BHWYY2qOc0NeYkaDgf+zz0MOJddmG4O5+l8KKfL6SU8ul
M9CUwzCEbAQtWdkSZAkpkWJuWa1Sh75OloWBn/5iZ3epAX67Iosd0g2UWQQxuVjvNU39n83zYzpZ
/jQIxNB9+f7PgtQDP/5Gl9e+md52xtkjOi/grzTG9PyJdLIR22YplrVMeggHCTsRMR5TiL8+DW45
r0mVAjnjTxmXmTxVQGM42Iu/ZkeRwTWVGLbSbPzd/OltJx1UTt2gEaja7WLMBdly5cNCRF2CgJE2
G19PoE3MDl1uxNVKXJT95tfllLrq7M7NyrMlLtt3Q1NtZu72SRB5XbKJCW7HvNVFujBz3KhTrkdB
rCSLLo4PQEUw1vKAwX8pbuMycyKgw/L9L0ke5WH+0MGUlIpfIs7m9miq3uHKumoH84Y1SfQdLuGN
rQ/6DmxmJ6KBSaNuTl7Kyfdbi/wJubM88GlqP3ZJRr84EUicvhxfco0xz7o3mCkpjS5BHucqpYvr
u6ai7G4JbYQPeGEK5CpZbjxOwNj9bMazA0QreX/bxiOPGQSqxqyBL3E0Q0NwIhUo7VPp6dhvPKE6
Jl3QO8fkFAfITbhiUjMW5SdpTCPBTxO+JFuj3ZN+D/h4TE5FFOZdRTqLRvKioGbtTsYtkb/urPJ1
mc8Jr60cYiqcHgP2lPUzpYo5t6YG6rG3EearZrpHCVf+0qObc8rNCVAolhlDa3R+OPtllC6ipXIK
YVJVpy/g/RA/x9BV3SI8onBQccw1T0dNN87h9VKMKfMLLnZAGAE/73hbgvJHzB4Ltd232sW2Ywkp
f/hBt0Z1kS7lTCMgyrI2upbZMqcsRlS+Eo7jo2kG7JldYD7oZBhknHYQLUH896+jDqMdcTm898zg
hqFUaHV4tH5tADtCiKE0WCforwmLNRKNsd8qzL0WJS3GKXFM1rysvv9MtVlZvmlBQPt+vfRJvmgJ
ZLucUVUDDEHkty3irpBocviQsPJoCGU6V2tLr5Bs339DycND9QZNIZ97/dCn87SbErceM7a8By3O
S8O7y9J9GhMvzkoiDfkNDMJadlAWPOHO4fYiGCKBIe0sIPN0gN82Xz8uTHqlg1qc0gIXSKPVF89q
OXX4gFeOl8M/fu/aeu/rjhBVavAOxqklcfTGcneqdIcrKlSO0rChsp/1r/hz8D+SeGLgPfKmXjrT
dCmUlnn0ktHgS/2DmHqHdOCfxe93jS8rcr0Wcj6AXCZqOgUB81Q/hi9WSD++6BBMgAAOFacmwrxO
MlTy2Y/Ssk87j9dhBXGyltXYkYtx47Cu9fp+s8T5D2yA1ojVhWH6Xj9r50Ie5E37fLvnEpSCyRjd
+eepEQ7WyP69I26BpwX5f2G+bzfMtsscOldyGK4l6W7BaIWXHbQIT1oc4oG54nbm+yjdBDjeAhfN
oIpULBp7o8vPt1vwX+iW+oceE/hjDROlZo9kQ12XTGtrCUATGlPmrZzeU++/9l/8tHGdKK4Udpyy
voqNHUln6uVhnOImBcwffSMcFoCbgZa0+kZHOy0s5/+9o3OrxZkncsPVFa5Te0wXb1VEGykSn91J
x5VOLRWOiSfBIVRfAv2AtKuQQSmspuCd1wt6ETX4w9P7N3qEOPjL+fsJ+BEPAeUcTth8yVOmqpOz
U0WUf8+NLOnzpNAbvtEqVcK4TK07MrtQCrvgfS2nnnedeCdm5Vea1yp7XtgZkV+pL6H8WMuAfLzc
yhfPO/hZdLNRxyOAEcazNyB6xdn8RRXoXKEcBRSJjMzR7udmCBYA56lT8gEdx9yVW6rzCA3iog+d
cJ2jX/Yh94FMPWeLrib6bcgH6leiJpwv3F/UwBikkzNqdytYip0IvRvwzTQ8Cbv9i23NTxiqpj2X
3ZnjBv4Krs3SPONe4N7M8eqVkJy7p2i3KfkNwzzEagB4PV0hQfjyjz4jzmUjNHmvwwq5DoSRyrmS
CQgup07X9trNk50StCpguNOjhNTZKNnJV7ePwZ8dskljiA/LWuIVojPjdb1nt3KfIf9EfgdeCmSL
Q1DHQQOpo6BAP7q9EHWpYEkejyoA/+QCH7qzR+vNz9PUR/e6T6tvs07Reuul6bivDi8S9aqkDmED
gVIqBvAvdn435NkVL0YWRh0A6OFSwmzgqzXs0LcC+COWEryvvjkIka5DpSwI+lU8YWizWg/7D5HC
BfyhRKOZD52OgQjr8RCg2sbCsdLgqxH8Oyyu5iAxxvauKqaj+Pz54lw8sAqFjcdqmb1ZsK6QePuh
JRNemI763OlV/qBuDX7721JesoDQSVBNADaFxVgbLyCZbozYdydJItekjpitdj1z9VnzChchJMZi
kdpfrK2hVcSO8WgA/xtqgNsrnsWT/VCxEHdCFtoyY6ogmONwbIgS7f0W91x4kJMujuCRDIx4AQVB
rJ8G7WVt7edmRtQ0eng6u1GLxhp5aQmkaaAAi9q6/M3BztiCW3rD6dPTX2lPo3vMDOEDVZ9HVcEM
eWGYWSCQ3DT8fnBTShbXLB/tFHboZY4uMNaOgrFWt/FjoipiGPNd6Ba8EUBUA6wz4Dei7SEltGTg
XbJC8bmMEaVbeIXVQ0jW7XgUyQJhcy04CrzTCBBl9avHC33CihpNt17GN9RBfbjVxVa9j978SppA
bq8o4Mkd/ydoN7Gk3nZWOB8cRnli9XdLGk8BwM4ez4DuHV9f2diKrDIrNQXiBbwIvOAYq+Vok37x
HFfkkyBXzGEchJka4y4wQiIxsG7zD/uAvEdiw3MYQwqyNiBpmOxSy6Bgbxf0oeZSzOZpPdcE3QMP
nunuFvnGSJGLfPYRvuO++REFCbBmnH4ZQ7Se5IO7LZXwTfBXOdeLPG769h29F2fslXQkSif+Ti7K
qYXRwHotTY/huC8U9EkVsHdLXUaRDIiTcxw3KP1ogy4sCW0JmgrnZ4B1tUWc/sTRIX2ha2rNYaLp
VjDq6+PvD8lfvPUboOmk/bgbrtyf8stQ9iJksLv0sIZ7b/VaIqX8r4sxZ40/hpxvdMXAu+hlRemg
P4UsrGpAeyIWEAxsfv8GyC5BZSixyoHlwzBlY446Hzw127QuTWkVan9EmWxCaSFiUOTjQd/CRPk2
tgRqOGXcNToD65Tsu0RBSWsHrnL8apb1Zf6twfbq860mWKzKpjW+fsZDkjdIVnGac4nXq/1vDJUK
0CYP38JO/8DuNhZLNId8wJYBkxD7HI9zmlFoHM6r3yReEum2jHDEOvnAC01SGO2OuVSqyv6ScKSN
lIb5upHMGwExbAhrER2ldwu9bXAOnwiu8Zfk7pzjrlD34GJoTF/T3qb177XMHw5aaO/WMXX308GO
4oZwE1trgARjwKuoAeQ4sKEmqYm4qVdfPXDJVb4Bz7HGzWeee/9jqsaVqjIj+3CifOo3xREOgILC
Oo9pt+TUaS2kJpQpVlJ8WWAytZftfRuBEjk67Mf+Z0qZLXlypKsNixJlgWJ5ZbqDouxOVCMFVI+5
dCo0FDGWOh3PdUihcCq3W3tE46UKXff7Wynj57FrnhxV116CERW0hbTtPgvt7Lfd0D5avr6N7JsX
dlXu/CTMJKG8tpLVqYqSCqUfC4QhEgnyW63OPriSLShMfUuHiOQi0q3r6RF39KTByPFZGeS9FlE8
G28wO0UvfB+MCQRH+wtYI3CmJPw7mG//ISoRXnU8jFgDvxKwim3q/mOVRvMN7HXU3IWf7G1AupHG
ZCkA8HB8q9QvHpHxFlfIIZWdBfwYqq45M81PPM2uZaCTT8uXUvn0FfZE3cT4AOyU/nUAsJTdQO0s
fMjf3SSU8e48OG3ImR08JK2gx3pj+GQLJCVnNFLxKpnYx3LO0VJ7CdBOVGCmgc2gYDXIJSFdpa+l
3G2Iyx01+kjrGhDL09O3IhFzbdseC613uaFwPMDxulKndI0oBUd4iLnVgc1RHmlFF5lZ51/bMPA/
Q2ddcosyNnYnRbymTnEsVbZIQYuzSDcMUNQEE4lRW68wwNZ17m/TyYv9FKdB7EYheLo7SPXpvdzd
Q6QSFmtDJ/apnLtR4mzeMXa3bB89WTYOkeBer/OjfHT9VipQo4gk9nH65k2WqVe3EJktdsJj96z0
6/W0sI0YVTESZKi7KOOLd809p9pS3K6vHuH+wkOa6UUHX2FtuGW+y71ljeRoDrpmOg15dX/wfuFy
fHwlMqjfFVHGcfYY1WMbcwlj5TxzCSxI3Fvsir2yfj7Od68t1cjMvlWy+wccNDKyYOuvL/jnfZed
klZNGJZx0MzAjRtJcbKJQHx3X3/tuqdPor4D5BgoD5vKDLtc8nONN6W3tnDgch4tD+FpY2vm+fjM
bkrZQ4i2XsFvCm8rJT4CDht6Dr6D/CjRbEkyqvnU1EQQa/7YnwZO/BaXZh/apgmrlkPSw+jPmVdh
CRhbZTqazHD3K4sz4qvnQqELRuYGQAv6o+3+crCKoSUvwr5/OBccCfel5woCstL77UBRCdSnMcKC
S3PKLqy8qamDrG/1Q7bampxhEnk2MbKPNS1p0Gez7GSYdUyDQG8XGkLMdApJ6wZwrkEPwyhVNCvR
HpsoiCVHcjRDFtAwX74/gZVA9oLWVUA+BJ+WKuzqYd1s8+VGUIWeDaOrrr15QAbuKZIEOjA9ZzCQ
JZ9Foel5y+gsI+dj3lqWKw+wqicfC2E5Yd4hjW/H/hc6pf5fq5gdKSHNAwdXyp1ojoxZ4fFi9YSw
6ZWgODB8wVGiC8pJAjItMAhrfiszm3dCChNwqifgE3OWEoeZXz+UoizPY/iox02y1wUS6I4v11E5
3jGctt6k4WnV/ce4w70+oh0wfJxYrC56b5zI/QGoGjUHjcu6RbptjH+JBYmWahixZGMZ/PAnJBzw
8TpIed6MdIVmku7hleA9MNK0rxywT4LJl1SGX0Kn6ioqG5futsWZr2h4J2K/kEGz55DEzH4GTeir
ricjenCyA5UWa65LGMr4YS8j5wPq36rGZaLsw9KUyitIy0W59ZSh8y6eUt9l9Gl25RuU7X64p3by
a4KVhF2enog0/RuOtSW2KltqaoAJS9wyIPnrzPmBq1NB+2AUMqzqFGEByZB+n4muwR4u6anNNsBX
NAzbqRhyk6b/MFkWDdaYcBthIoKoqM3fO/o51d1ZnIH5ykIgCDJRZnncPEoz3Ux22Hf8t2j3xoJE
0/xbY/+Whg3feVnExum4hN5JF4Q8XMAgN168yTvog8xzzpvtb/IFzsOsqe/+GZFlLOuP7/cRATF5
/wpx6tnzcxqNymthquG49ok/J/f72cUnJx7ChZUfFI+FiPv3hozZsirC01HERWIZwrEVH/GRi7Pa
UDxh4zE+uo5OI/EQPRRNxBJKsuOfs5OLtIO8o14yw0xuReKqNyz4W7I1eWHqTCuJyHaS87mP398A
SS2vvdThcqrymaqdhnOjbJ2zrwJLEj83++r3U5oqmOht5sdsocQf3movmzCfig8MQV1jq/jo4OB6
BYRPj3T8rG2Bo/vFBBPZNAO0MtH2JNbg0Z8LTqXZXGeWbQ8JaJwNlDBtZY0nShcdEqtnFwlQmwTz
9OMQlgbcxO6Q+HPXfCG4OXU8dpKRCOHsW4XPXoGggctzc4Na0GWXmqVvRxs9Z0p/gLI7q9keNp4T
DTJ4O4qkTIeFTOlBK7oqkyGx+QX6B5wcaA+EqZ53f05E4rkDyC+OD54Va+M0Bu32wu3N7P0CIN7d
B4SyC1nlEH4FQ7OvqE4U3t/BIOyrtLcCy1revp/JofO1BqmEwGhZa9TIg5bbI6KD8jq33O/5NqCl
J+MflMad9LPmZJnFea1XNOAoi7mW5nywF5hGqMDUkqKnm4aAeAnImKPaSWd9wtR3otbf9gi2ycNI
ghXsiQNdmH1FSrdYmTth5pb8epA7Z8S7JBIVh86d/tHuP1w5DiGX3RaI6HjddM1f5iM2g2sTyroQ
bG8VuL0m4be9Q6E/wqU/qhIEWS901C+T4RAHjC3YWL571tn1b4jbVDKYKrYhrkDmQn6wuHJj5Wsy
sAwDaku24CpDveUcVxYVsHqZCfOZ8ksva25A8JkPZxl6zuNIcZDm6TBydLo3x7IbRuyYqs/dWcWY
YtNX3VLYXWMLReA4Vr77xYZs40MMt9sMesoS/ERDCMg5rDPVxMdRMhn0j1am345YsAl/U9ov25E/
SHHYxhrkdmo4Mh5gnrgGQpePxmlGicHc8PveLPfkXvBGIbQhelvYBhM7h1v/M6+SlYnPNk/Uqp5d
7JMmsF3eSJkciuRU7U47KO8f+1x0B7xLZE3PASKYeK8TeSoPLGXTrYbsSXlev+xd0b6CftkFjBqt
U5cMvmGQhx0oo5Bn+rZAZTlSFu1nt62ovW8yxR/L6/FNE3ERynOOAfmVjis6EVpAZvg31CcaXiAS
uRwXyTzBLyjv2ujB1/DaQ3WSOLe3TNd5uYrFfnGisjtRwpM/hV4T9G7TGJpALNL7fWpBsMJv1+gV
rTT5cbGBunRyMtGWHcGxFYZ38ef6gSfeo1bW/DtcOlyMlZ+Nb9nXYVaSWwYRtgs/HQiWIkLLnYIq
U5mOln168u1YP8lg74tQgBs+FVnPDkIQ3JrNry8OJ2q1UVnFnZkHQTFlqRbJictbSOXCXbRvNELk
hMbNWnNlOcWNRqlRdrqAIFmRGLobaE5+imdrMzLVgNqAdVGA3bAB9mdNCRJCgSovn5yVfEVxS3CF
imfcySk/vwm2uCGxgQCFWigb49NpJVv3OvcHHiDH4q/Sr0w1qHiX6BdoBtuD+VxOjYBcyE2zZoey
eKrBwbWfWu8WE5dVcxEw0PJVaQuXwDNfugRJpw2/ciq8Rssivz+uF5qS3uh9aSGi/Xi8KcVZFGsE
shw/dPu9kxFEdTY2ETerk/R0uFGhaJznGJU14bMBdnd7RxAXnRe3gUGgixId3MEr5noih0b4U8/f
VE1WbD4uLZgR/WMHXonscL/8Jrs1edLAoEBY8QqP/BMIYtDKlOBjvBHnNmvRzakzlphgybEmdxbW
CnhtCxqDzejYWbFIG8Zz90EjT7+k5MfHndwIGGnxd4qd8jFL7MMKpfoxPJ7iGq5mJPj7xzrejz2Q
GmMGRejaX9ZC4YvQAMkb4EJIhp64JdiFB3QCwDcw/4+UDRYEspv/gi0anhUcy22c25rMD17amgRg
EwjL4FPsjABW5AIMo4ch8ebXT53+Fl8Ib1r/pIzi+PLvUlfHfBnqFQChrkM9FjIiv3ZZPwIgrMtJ
USL2rVygVkDdqDSXi+UtnuoYefABUrW2C/lKC6a/ytNAuTZa5KqKGnRa7nJ1DtnS8kEfGhWmV5Kf
A2c+tnht3EaiDWr/xdvrGeiNt4mGNlXIT9rr0AN+F6EhlWf0Pcy2m5oIIORBqeUH0OYDc6V4AkG2
CN5c/xYVCMxVOeptIu1G1HF/0UcGWRUvGFl2OirOWl7o7X0RTANvEyfOqLwlpSbLwDk9wBEGYm7K
E3SGgaLEUx3Vw9jJXU7+O8ZD7puJf6MTg3hVqz8a1idVdbUqFTJaWAz6PUWH3TUsXvOu/aiXAFqO
d8LG3GdPcv9naJfSynRMyn11DFnJ1vl/fu1Vg4znsZ2mF7EU2ed0SxjDS5MEE7U2FBrnFtK/5YbE
lqtGyZ8TyfEysR8x6SSaukRUNs4yfGOW5yCQbC3GIb1O+I5YhTh7w0kVG8hgpskbECK+05FqWr5V
rwoH5I2BJ2yKXyYPlWMsrUousP8L2whE5Ewb6C68neMdHtjcpXddvaUvUr8kxkvhSNgd+6zv3XRP
FJco+idMD3hCviJk78769WrHiMSqlvMt23AgxaysObuKLI8WW8kk6zzxlxlU9hpGSdPS54XNbwT6
TyHcRYWkBP+34uAtS3GXgHuLDbb0GTW7EvcsHpSGgau1n10BlPN8zTq+cfZH2pkdE6d3PI4Xzw62
q/b0SkuGYb+BmVn4ThL3AsoH4vDeAU329DnCoquVku7UW7F0s04W4Y9HqvsSAZ52WGOGx5MxZgad
5Cd38p6ZZeM8Lwggs6Ft5L+6QzrdgqXuQJZXjms2leXnyrR4mF/0x4Lv5cLTncUiiEKVcPTEVXlX
S0n+ijOini2lapB0tNFJupfLJPKpNc7AqM8O9PG3eJ3vxwubx8Mz911XMrTz1NZewuUXCKIPxYpM
e3WjRKkEOCpKlowiN4gMdLqMekDYbK7up5H1rH6p99hnwCVf7OOdLfkGF6A96QBu3ewAtnLSNmL5
WiE8pLTVQITBUCIYbm/bo/Xn7fGkdn9syaAjgckHhCXV71zgqgh5WptD+pME9YzNePEmEnhol66G
jdt1QcaXmjQoR41FYzhkKac+xKv/hgnmpCeRoYXopXKOKqbA71o+fqD42r6Jz5mH4yG7hDNG4To/
HxHCWDvEAlqiF7NvVnYaGcjt8FqlYYcr0e9lJcEIKfNBEyuNXCGtUjNY9Td3KWJWx7b1UxEw0Db4
9C5i4E83Buz10U7t85vuajOsNV7h7qjn67+eQo7YxyMwyRJy5Kf6KASBYcTjhBE8PvKDdvPdly3O
rD3h9t8AU2Dj/HH0g+G2+n/b/t5zBS/b7JO+HUJaj66VUxm3r9aBBNGm60O4pP/mJMTdP9YBPIFE
i4WFk6+UYSKzGUvAmNH4tPvp87o83Gi9/dvyvUoG+CDhkwjN6rG8CLreBM8oO5K36mNYF0Nh3cbm
LaqfgqSDxeeE+n5MQnXZWncNw8C1TmPT/jfTjQ8LbkYqAse5/Zo5OhdDdbmwOIfo1uu5ph/4ghO2
whefJiBMIG6lmCc1MZR45YLJgpr8Gu8HcUX1qR7Nq4HDrfvVQRomW30n4cHYUF87doM9PKgA+y2k
NCgGAv/NwEVLOZ0ZDwfgFKooKCLgAlsiESJydxsOw7xC4lIc1H7BIRquPU67AP5XROT0iBtoSkxY
sskXahMg22X29XY/IJuLzS9cVXiCbPcPU3ofhQdhNdOxdmxPNE9xNLuYHjtHNDkUdh1OTnqt6o4C
BvzcodohyWuQlP5JbsFOM44QiYN+XxokP6o+lMg0i2fVmzX6qpQ3fLANVHux8ab586FtMEclWYmv
Uk3mRwpigonqrzWqv1P5p2t2jqUVBmZFC5q0iibN/WGv6CbRhrQCbBwW2B6Do+40l2QCYOHjwOT6
SvT/vX8+WpKA66THzMZQfN7r78tr18IwgOZ4dkowA3WerXjcKNhuQk1rzAkPDYXSepVlX/blx4FQ
7xaJUfnanRaI/vMA06bP5Be9vQdCP5XS3cEMEpyYKkRBbvVi4v40AGmhkHUFcLbYqwNZEhii3HZ2
Fyrlnv7LVPVtphkhiGG2sPcUbD0jAkDtW++HGaDWR5/ePkl5hX53zNVNJ06h64C0ycAn+qkl20Ik
z+7ptE5n6PIVTKleuUNDE472tt3I8Zp+P1ZNT+TiZIzXP4q/Era8sZkhsmn9/auvKoqvBwbnnoJl
iyU1NaVOcNSTo45D3lYecRPt78lMR3LgGnE7stIrSwCHw0jiPp66APrLxo3PImMz4IFGDRrBW3kL
jUh66q1s4fIkyWeeIH2YAy2XmMVPwCMbgq1Zq+QJGOkMK/VuPX12WUrEPFUag24vbnh2lx3IySey
9QF1SOWG0GdqPlO7VW/n9qnAWKnlSBR6N0Namy1/gyQvTIY202WGQn98Zyv8baCB3Q8zdbOfTTsO
DLGiB0fhh74y1vSw3Or5Ko4VQrrdnzF/bM3JcHedmCWr3C5lFUpV4atbXfYiwA5VGbPApucaWoIe
qWeiRLQvl7EJXu2Zj16qlGYeKs1Q2d1ebkeRzA5cKfG3iWhthd4iFf+kNBUUfZUdvY2BQB18WC0B
l40aSlgbfwb0V70Byhxfa+TsgoguvgJ2XAzV46Zuyh1S/1UDtTrRz/N9EDGpw1Y28Uk9OklUDlrZ
vhHLE2wOlJ7oOiDxpRgaNZnkp8yeqhpPkqvo+TflGlzhW0uFLdGlEb/6yuTSVpqZ6bIo/FEF4+vj
KzYPKS6RXhnJKWKzlBFqSt8RoCbSAFSNQeVHabBTNSEMdkzQQWIg22POt642MTFwB9eZaiKk8YiC
BaoNKtMb4BUVzl4KbWKKHFOX+4RuR8MGp5yrx1uupLb2v9/zHQ3QPhcCIMDXCgViCAJ0ePcxxhyF
uSn/TRykA4i+/y/uMuDalL6rTuG+m/fbuxU/nd8aPPwWfcJvBOaZZQWL2KwEZzr2f97RuUVccazF
p+N3Lkpbj5VcK9hx3YEoaAeHSIB5hk+aYP9um9KdE/iaK7yYtOdeKbonC5TJkgZGQb2z6tuhh7MP
RDBtIKJA3snLiuyzcxjpXm5pwF0ke7zBvCqb9rHi10p7jJoMwm9SxY8MDcgN6P0pb8BijmeJJc4N
7Ec82jj9s+wwkhZ99K59AwOrGK67PbTFqAV5zxDx7I7XhgzqZ8diQc8UPvaQnrhI4/ImFdcyOnwP
hkLfxOBoWNZI4eA/Wtqi/xz6L2ytpl2CHrrlikWcZtq4ygKDiVs0ASMeINZMMrXycFJqH84e7HOW
2OVCS5BtS/7d1YAcBAEVdrz7Gp9jyNLgcYmi+NHqyPjuOiRJeNOKMfXTzS5aF4bnZd5EIhJ+r6jK
2LKf/IYIn1WAR5BmTexDISlNXbanyvE5M6igyD4VvTUAEdlvNWJTN/kVkpHU1vv/31j7mtwdI7+S
OnldYqbcKQ9gidV2niaMXohZtNOkpMyjm9Jfe7yzHhx+x+jVghnOSpm8aoF2lxBcyDqUWVM1MnxQ
I7gcaWpifwqDBcNCHl9RhBDXFHTZei6I5FeeultPBURC8JkO98Z7iCyAtmXs0RHw3ejv4u/pEi8G
8IdyIuJ/SbWfq0n+wza+VpKLimXjOguVr1lQfZe81jf53FH4GgTddu9pdHSBQM6Y1w9xF1dFUTLw
fDPmEBDCJHTg0uw703aw6FqrVlDKTLRKzu9qrKHfmGQuKQ1Zg8h+0Rk/Xb554aoDGIYyPB/QDvS2
x+ebkoYW9UMUwNAORLdUBV8w6Aj5Dl94w72/gagYnTXkHZhZI2Bwv9a5al6Qoam5vGZj5w3Ydw0J
Lo8rwArYYfARWyzcU/sd/Sucs7xfeyYJGBNJ7w8VhL9MEZLLM0MOuVm4DtQ4mK9/klCp8Ivr1mZC
QW6ukyF/TcnTuMd6Bi/QywTH/2apgaThq7fbIw4u5YKIVU17xp9pBMTFal8aqrifpGNmjwirLJJF
RK+STi0aFTTCocCe8nKgZ8pG4o18GhmNoHSoAI1/S68srUQ3bi1zp9PF+VS+mDL8rqvwADjVnuSb
xB9Hih/GMhU8uhvwpqw3xag1n+ya1Bs7ERhKjURaYc1V4DS1PL3/xTaoHeqP2xL3M567C+0ZNX74
eimYg32t1AmXlGBDoNJCTapkCFyIxVrjxJ5mESCsySYIlk9/8PD9IBYKI4OBu4iRH+AtWk3nl24V
LBgCz8OiXjF1HdhgItLWOGSNNUJVto3wMvrTFpytCHg9X2gKnlbc/0qJh9SnG42AtV/vFQBbRfq6
zh6BSAre/8f31hD8WNy/+GNMNItscwNUDPz0IvrlEgJ4rjQ5Izkdn5TFNXhV0bMVPQL3+6SYDyLO
Pa6R05Ch6uQJCKoWVgj2qzzzZQex0JDsCCL7GR7mmCdefJNwmJtZK7t9QGslVyfpYtDekXJO/t0A
NjNX3ODpMSH6HZMxvOOz2E8VPy9DWB0mw9pl2Aho9auI5aJufMjytetYdBtI+9kuOpnRRYLO4s1R
KNXkUapglJVPVbjE7ifvM9JRwccK/EPZYyQqEYw/elHLrTB773GxUWLwalpRsJpkrM4lLVVdUKjA
yyMVnMn5dNypU4SrTY4fsbo5gJ9+hG6gf6I1gwfNEIc1TAD1weskNK8DBKopt/S3GIXfDeysDKt2
cq8Mf2phAkoTDOKcEZ+WlIRL0PCw9+hIRd2erf8fDBqTLIkqt3bjAbfqRjz4+UnysGgGRUlr0p3j
QAlwGCGngHUDvO77fe2fBgk+PlUp9nIXgWfk3uB9V3DPwFg2FUQKJzEY9pRqEDui1qAfvRQwlzn2
i6KLSK97UxZYlTzC+sxawBUecDzXSIjgum8YXfrM4Dy9sfakqtfWa9qNHInB0PjvRSwSpjlJTikb
BhJ0cP3RKSFD0vrVeF+gR+7Mw72Cs3vb2y3P2XOI2qT9r/r+zhUtBY/A23Si2nPGEb74XNo1waBD
xe6CObFo02MOC36EJu+Krm4iYahQAXct2nfI2DDqMdZaxUiP7DkjMFvzF+bFvqGEeNwGcIRNNjGd
IDvebuQRFDqLD+HOQzCrg6qmV9H8PiI61nExbKdLJjpHVwhc7ZCmigIsDUBOBGSJDSAlJsgUEed3
xjdOztI23bWLqtSod9q9MxE7OiZfUER6kR1QPLZty9JLGkXieLZJhjTHI4j+cabmuLjMevHzsUQT
H4+dvzO+l/7sCqR5i1q4Sl4+W19dhIGRr71VBn1xE2GYzEeNb2GDoS/1f7a1jqBZtG30Ysg5RdeF
/vEm9i3tza6G0aOvWY/6G70C8SBOowHjUTzVoysm8LCJ+27qt6DwI1jqGw2WFReAk+F/weUTWYVo
058xTISw2/m8LluwOu3e16D7PHDnpyKlo1qnLy/oAwTpk4DKbEa/mPQF9yNUHKToq17G1Um1roqD
MkEEWupwRZhXGeepnpYMvmuM1CCoxRNzLJKPudv1HaIl/Hgtt8fUW3S9OxnNbNoHxqi6z4QqNMhT
RxGMH+Y2FFEeZ6QNoGTDev7NPmiF8eenMNn3cpx9LLdJnwpl4eI5vGHiW4yogiF4uaBLZaBEkN8l
HaEo7lnZsApeHy7A4xJkybilPgTAZVorWGNOustrzRoc0eQo2OwdgDfMHmQuCz9goglWNhXtmyqw
K0NQumJJFRnka8uXHCz6KbNHtyKwaN3IKDOwW9PjbOCsTxIXoA+5GLsuquSb59mBR/7vmq7gpkoJ
3LIRKOXkGXTIoKOjPeAhh5U+OuRnywIrRp6mIYhtIYU7C+tuD+8/6SFoSytLuXnuNmekJjbx4UCn
f+arub3RsbrG4MMBP6PSPeZIe2ZqhNc8Ex+0qzaaQpE1Kc3uAeFQZfOh7kjUsJQcNePAuYZg9EtM
iEBfbufeLGiAML9ExDbumt5R+qATiXnUz6sBn7BAEsdh4iFClb13PrFBV/cZWW3lNYwU0j73oq24
HeuxkD95UR5IlzcVCKJNZuU03lYlxVhVKCoQrQ0Fuf1TqJN5DBosGJvf/WrdVOwe8Q8qMC1pJrq2
H/bcP5bxHzbWSQlvKswHX+B7/DmcFjtXSZUEiXRddCTv9BXMx2/Ol4Yh26jrPc2M8epftzoWKGbd
GH6bs0QzvGkVqFXi9aWgmr5hQJU4J5sgWqbd7RUIKZErtLTwVquwwp+ZyR+h977vcsW/QjHo7KyS
9V1i5o6QA7w1WjgnGF+KFZHA6gcu6cYLIa5b8pTKDu+JsOPor4hyUCsqIBkUadVHPaIXH3thqUx4
XfgQabViR60WJ9WmdyDm1+IjtSWj4UlodujyqUSI3vV6CWGTtMTpXyEcKTNNI1MME4dLJ7/2BVOz
ZN1JfvJ2MweqC97yqH/KL8kvB5i3aezu7/eZjvjuDF+u1d56m3c2mDNn8/YKg6n3Je8afLBhgvLx
8GpMeDHKa9r2k15e8oT9/KCwZ4krUDACukBokIvVO+WsDdPSEkO4nSMQfL/hgsPGaxBBEqE5Pxr2
PagAez2AcBD+toQMalsVJhmShdGcqgB85DijA1QM2OdRY+rKBK6UFd4irYtQNfcrsR9ZsWg3tzXk
cbokV4Ap4fsyf75HQmTiUXFZRD4C8dcm1xAICkSuGdg3O/GqfyDMuskJXcugEtuqqcApXGqLLN6I
IQqASmZnjxjOTLmlm1iFgbL8zY2SEf70j30mnhJnPrf6R3mqGk3PNYorF5TN+zHl1CHZNCtMBhrf
onyhcyEHGw924InIj7cXya8uzCSeUT17cEQVRRvorOgTYlnSVuXHdN3h0+8yk0iQ94lVZa81/J7H
rVCpY8OqoA5MkpBj+9ZjpSZrTgI9pssipcjtH4Jm0+fdfiFt/RqiBYtfU6T7sDf1MD8Sbapj/kAf
5bUgxtmpU+rsRnMbuCHheoqSOi1MF48vSwlDOhlklImloidg0lLCka6xhTySvRFj55Vk26oTdYs2
+18+YEWX24qIdxCzedbdkuc66ZmguvazYSpYHXQZl3Q2EFxYFTCfzf7u9UgcPiVJemlTsi3LVQ4Q
wV4mUGVF+n3RbJ45xgUsZVbzwRWrvViKRJmNT49/gsBlnKrQYRXvxy9LOjq1HDB2SSJkjjRZydYy
B4gcDj0jVKOp250nWVemk1ftFobCT6k52VD5WLnXQzUfYqI+irlAmVbMbCr+BUOIhad1xWJBuuEn
VaS+RFAHoqC0aSqTswZFkyyLgnsaSVStGmkntmaN/jdCnR0BD9LOa2nGlM6JcgpU/6CJXybxFNAX
VqvOwhAvXj658Sn0LktzVp1ekqkuW+WyKEThFtDHY1QgkJzjNDb4ud24indAurN9CaA2BlWRNVpc
OFlxcy+1O44xBZb2/oHEvDU6BLd1pIHmsKCS9F6KfzJgqI6+p8+h2PaRnkmL9PCPK+Eb9ixD90TD
dXqsSBeOMYUv4rMbj6cZ7d1Pqeptrl8PKZeOtuzIQ6oP6E7TWnC9jz1dLcALfeUMszhZwsMgrwZd
sF7FZ9zeozR2A2bngjABvBVVnDtYLC3mzoER5M8e+YaGlJmf4d8Nvgotqvw6AhKicrhz0yivBHgr
HkYjxM1VGyxKyk5yLRw0iIZyB23a9S/WmMld3wBInDg/hX1+hSGFH/Sd7cTJRgUgKnfllLqTwzFa
sOw4yL1QEu7lrsdkI1OCVu0dx8QANkRbd2g6jh35onuu/MqYyMgwUxV5O3DS/qBxGpKQLr1snE4d
0+/DZQVruyp8lKwFoU1cznElLMQ1CHhGrM2tuaFUxADVM1TuPLfUfdwGG3hWu+Xutrx7IiUaoGd/
/KeyWJ+CiuFXPhUKIWa6iGkbKrAg3khTiVTa2YXBQwbOVYg3w716M4wiCgCaGn1Q09w4G/1cewxl
WVcMsbZhTB5RpYR2vZzT81WKUtelCBH7KGoYGEJ1J2tzny2gpsCO2o0pCCwTDaBBodVUX4kTysri
M66Sgt0rmy/w0N++cyfnsuVlNiWtv69u0iVS+kL9AD7xgM0TpHcRuPhBtyefcWgt2D3Y758fbt6N
kPolvKfpf2Hj9p4mRYmLBwU3I5qfifKjx/kY+YGa+YYo3YnskoldXqbuDyXdB5QV4sp4EFUdi3NB
RGOHa6CQjkEKox6WFSP+cgJitJUtmd4vsZuIbyUSjaztlq+RuQ/+GtmLQ8U3J5oh5Q9DF2+yUH1E
Iyz+DCSovPfy51cSGQS58SFy8Ban0tUMvK5bGzQsjegvGbT5lVAWSW8dNIQlNRokbAUQxmBqopIE
AElStuekB0taoGnJRKTK5wp3Rk8NfYuQB4rWIcmwNi5BO8mwRxKxKEPcB0gA5VVQtl4O3pfSUKlB
X1ioS4nrXhSrLw317Bly5+5j/Uw7I2xlfYyC5L2Cnhq8wiHZt9PrmDdup8LXiNtHu5ER2JnlGnnz
sWkmvVsw99xc8AqE/rqLe9tuSl0FIspngmQY2rYOsiWz5gxDJFzukGo18axOi/4l3vsTYnzEWgOt
8RahlGbZCZ6Sphi3mCdILSCyEklpBQ77A9Simzt5C6vrJ9F6ON6fHNFV1ye6wDlTVQFv1gf95XMs
R9H7XbGrpkTR+F9ntQUf4Azq32INyd2rANJWuBKeqOZ/OXZf9xLG2MQ4UlhtWesyf9lD+1y0upUD
ElO8zRpmwxMU1AXW7KIj/zYwc0Y7ghb+3NH6nD7y4YhttM7PFOeLm9I4+LIy7OrxLFqUjBfVXxrK
2fTQQc27ztZYBz3VDPsXzAfMUbZ+R6hdKmqKt1GUaGDPzGFzBSbnlXMebN4MsaQYU2dOds7/1YbW
RPab/is38iSS487n7HfioNjyf9e+sWArpkMr2ygtrHb7L6OuuLjxV6hswwL1YjO1eC8wM/Uc8DrA
xUr87mhuQbDP5luwmbU8CcwrGjwqT3YDkqR/tnhNvqr9fdHifz4SrzD3Jimgrj/9zUHXQ4fciQWF
hQFLJlTQeVcy42qA2XR/860XheV/UHDS8c/Z+EotMxpvfGHSVGxJlNfXVDlP4HRrmVbjSZGmng0U
lNiRYgh0gNPCtCoIO4DoZ0YlVtviXZGXJ7I7ryoy24/yJvMZfwo/vkyvSXupEo98dftb3l32CojP
VgVg4tE8F5WaCZcwQvnXnJ2aiMiymBkJ8Eu96jlpY+QT/6SuEwVyf+vwqGmYcMjC/n9p8Topf8iF
299LDaN/TY637foIv5Tl2tUeYB6SCZC83U3trLcaSx7VuWqcXp24lWrskpGxEaOMbHtgnlGlR3Gq
wyeJeVxTtSY4PUcCkzFrHiWYJYyMksa1chGKgwPcBkCGrJJEtbVrFjXXqtZIwSG89qLzLQcyBjP7
OkkfQpsrwzWDUuOciwUcWh5vw75/jEjU5wxKuDAjfx1L0dFFpUfoYLNezs+sKaU6Q6rtCIDXrgku
VEcnBkrln2eS19kCR9z4IlhqGdMU3bKC0H9Y76XaygcQHF/mspMQPTol+4yDRf4gY3sxhGw1TG33
1VNtHntlyPioYod7GAyWeYaiAZW/UL9oMAsXiqEqrQsBQG8VlUCCjc33N9udCCXgVaiKh3RBvULf
+IsdA+ysnv49uiSmU7vk1iExHhFESTOnvukmGpg+g7uYf4TVCh550dlok7uPpXlQFJUPt1J2msiD
4ZSTeJNDcKp9PlrgXnxcV1Hqp09H+tlBiUNuzjjFWyAMYp3r/YPgu5il0f6Md/3PZ9d9pLakmN0b
sknwpQt5sot9GkBBrLs0zpqSeQHtgWZWWv5IUTmLH5hah/n38o3X8vaL8vTZOZAkG7YPnr/WD+yf
dpt1Kt23yibCjT9DCmftBxH18UxLhO8pWqdflnsFXil3nSBRpbNu8JjVUSJiG71vwX8Vy916zzpN
Phz7Gq6IN+eKjdxaUm+udFJ4X/9tIVN/mmuHnPkhTASPonbeyHICzCkgOqaN3pN5Dx2F5NWdggLc
/VMdngUXSsF+RV6RIoB2PKcWW2ckV7gbWg3ZSbYqPO7BnzyhYGPvtL9Qj40RjA5nGX5PYFF1mdyq
ld09teZpUt2BSXYGBNU+n28DUZAQeHIeOkH0HQ/8rT64TG0ak5ydouVzol7J7wg0PlQWWAmB/jiP
qoUEfDaVyCBR9gziUlNXca6j+sYo25Z19M1MJP3jyOsZPPqQ/hf7LCUFb0ICVJqMqX949N+TCHSc
8mr7qxVZoXNF1wrEXrFBYPp3mpokXljK0ec3iV3+ySFwiK6Nb+Vnez07akY7Yl3XkRMxmCJNV16G
+e2BoXphPDfrnIVCpX9RtYPFuvfglaZLz7gQC3MyE/SX6rNitfhXhuM92mBKnmJzV0ZjKsFAZXtU
YYw+A9t9Y+oAzYjBw7Bmft9lZe0I1GnZ4WJT8umfQLYJezWU4ICaxDRr/G1LATz1fFsMBxyBbfMw
mxpRvbqsQoliszayaDX9H7nSeTh9g8L3au7q9HWeVf6l6zES1jlQ3pQ3gMZCLdpTmy8lPaAwhVU2
zs7+wDQjCahPYzsy5xQkymzMOHifKAA7ABVQsQWroN3yp3Gr7h28sFQ8v/eI157HI7Xbhlm3UNd2
x7Lt+KVO4mBpo+U0YtzNN1lmKE5jfjf4RQnbSMBmZRS2U3bAeFfGZf8/MH6pBvRv5EDTcze57yZj
dZ8lwnpPUAbd544Bgf5EyxEDQKO4UwqLw0pGrHZxWmJ6Ue+0YvBYv9heOLoaA7mFk1O+YL7WbZlb
bMDlj4jKm5torOij08PJwnwuIuhOmFg6VYjNrT4ZDSS4SkyMVhKuSNn+sHJ5a42i32hcBo8s0X9T
AD/BWrU8LdfVJTHucC1MQ295uppvzwMNkVLTCXlr3GlFVl/7z5LvsamoAVsdpClOApEwz00SfaV3
Ljn2EGZc/CH9A4DLim/eM6xMiBTg/KmGeucXK3sN5wwxvsFb4lZbJyCpsKW9TDNhzNshN81bVd2X
B/Kp3B95pWSdSNpKdaMMV/AmtJ02L4SeBoyAareKBMOGaubRSZdvoudT9pFsb1OpRGu07sSM+OaK
Hwg4wWEyJcnl2MGozFeqmKoCnik2cb/mbBFC9TK7L54MKG5q605PTfsMBH9jcCOJsbom4e7bDva7
RvMv2n4PyC3ZYgLFBWFe2BDirr3kWmx25FmTAtOUl0HKLZB3APZuGNcmbQDgTUNR8w9gmlvg8kzf
jOzxriuc6Ar3mFr8BDiIg/7VSlRy1SwQSJtey9FrSmq6qMYgntTwpdcFLMxq0E9VtB92rQkFDkmN
G8rXooriY0lLjv2O3Og645WKZfv7KW0bdxzKXUq9FFNiiIkz0QrEo/QRz/97Upvs4/8s/WvStLYF
p+XU8fK/h2IMcAH/UupWwn9Lk6fzJBUGgosfBhmpdsZbdS4oAZ+eRHOys0RuTip9Zl/x036JBvMJ
JJNVCE/8iOFwJdaPJwa0RqdQ0zfVRZrJS5hOfJxVEc0r7s37eDDaFp5Lx1h8LPmCf5Z7aKu1PRqV
g2cseVRABaKEZm8kk/Zq5C19emca2d5WInP6auwuuTi7VTBQ48f78XrcJCMAl7uvscnws+wU13sY
2vf2YgJPicrLtG+PwzPn6uyhJkf60VH2rzvBAjNOh8e1rmXmJBHoS1+7DwQ5w6Q+o/1gnunlc9bs
v5VVROTF1/RqDuFLsFQ+5EeqeohnEy5gyI46EJWryOZtEwWmQtBjzs5EzbJ3W9u6iqoxFSc+RJxJ
juGEUdfPZLsVoWcMWlzLkcBgwJ+AvlvSQcjFyeZk3hg6toj0Xn2PsqWc0b+crbe8ok91uvbhV3Q1
EcdoGeenM5IuA7Zj7akI2SfkpBW0VBV0kwh8SAe37Zmh6lsPk4yKsSd7Rf6lZAKtvx9rTHzhPsnm
uIOzr6wAAY7fjjf6S4WAuMCyE+d0tzA/mcvXsUPhL76MzAovHsWOKg7yzGhelj0s8ShK72a70MgR
ThuIKHALQRbZ1e+4dSdcpbybG1xHwXu4GOyolqYq51M7fdu6aFYoyza/eWMDGAdWy9MKdHFAIW2h
yM+KLNnccLfW/2LPJuogZAJzHOp8KSB2F9h6v7Cpu4mXrDkKIns14N18UiFYYKresGqDliFF60b4
ZC77Oax9V60rvWjr3KhmMqycq8E9s/Vkp9z0wXa9DeC1cExsNKZ2mxY5xISFUNHmj42F9pDsBmTG
kXQxRUQRwhp5MozBxGP+GjbYB58MSro7pLitLr8D33jaE3SW7FkWrQqu8fWXL1v1zbXwN3lxOoDA
6CAiY3eEdMNhVNENpmAeJJJEkdY5H0MQ2atY52cRYQMJbwsr9IK/g+Zw0hh2+xodN6Ax0E3xVtVw
Chmq8zxDoMFwO95VCvtSySxj0mEDwySKWWi+HZ/g7mBogbIDsZLhX7uECIXMhnHrWINci0ehhwtd
woOk8xR8CB0uHDph9dV+7rBCYEwB6C9fnY5jupR7KjMJZEuCG6k8Q2JSw4lOTtU3NqBG1uEG1p6d
h8wwU48LYyWdELyyrKFQebRitQydOxrEcp4Mn4f0fH/2n8LsPAaTZSRjuL/SM9N5fdokkFmnCU9t
4116UMYw8J0KOQWB6GlwmY0Qf/aRslF3w59Dv1L+2P2qk7UPndijckkMKMMnDNaife5rOg/Oo0hT
vp8Uj+UZ9Os36VFZbyRF9If7wHBQOOTHgVcErd+t84mcKpx/BMyTGJtrsBgNzrSxxLBGMfZiDSBT
sXHtKbjOZ0iV36Jg0LnNqxKofaVqKmbUL2JdhwoozEMtltut+rB/k3q0mQUSssYdtvHFeHKM+BO5
N4y57SA4uUCqQCY2I8+TxJmjAAN4Ab3T8A37cJueSHaAMupCXBOAM0CE4WIDrJba1mlS9jy9bEnz
Kfn7yYFU7WzYIXh7u6F60fxFtlabyOtV1cJIPl25ciKYITjqcaRX49cUSYMsJPudoUJVW+hdl6BP
BSC2FnhcU9kaL+YbruQ2eXCqozlcj8zgnNSV7gyKzCgLBUEAs65xqjucpge2JObopY8Tl0T1VWP3
tZq2z1U0O/ore5zX5UUHdtMJWtnpD5/nDrLqdwhABx8g6D13Ad4TDctZLKnXfre0xd/xQJo9rVwh
HSZwjSJPIWWeP+cigXGh9jgRQjNDkrs8CSAcfzVZRAoliD7jquVfLbxy/jOX3IbBtczYwFS6mJZr
0Ej+I9a7zzAfNxiwjXKPzWX+o7nuF3oiHlTcM+V76yNsiQti4LuTb1JwPnkGJPL5UDKp0ODbXZ69
cOeaV7QvFOwGHktak8ZwcxoK3zhmkLqnrX5QPoazwil71jy4zwYgqTINfqS8yB9pRGO/7p3vdhXn
UoYZOr87WU4xwGyIklZqygQu8pga3gdeKn7TMc/Ys3mNO5frMn0DHuXuNr84kTB81dMvOSrqutu5
Fks0sacsPm6dn/6F2C0OUYiahm13tJwUPyS87pTMRcRhs98Qcb894ZlsxkPDrWU3HqGeDLzehRQ4
pxw7oD73yiQaNAVPAiy60XSXcQcMSoQbELXbqgOb8is/jZMma3Zm6TcAw/Gk6EDMkkMTvl+riXPG
gmWuaEVidv8m3YQ2HiQPbH+A9U3v9t+6Tb9caVsRqbQHBPWok9Ugy7mkY7U+xHowTvkM2uzMt/Io
ssyU1lQVBqceS3YV51lXvUWYhBGGB9aCkaMoZQOnRo0sPluqGcAYF+75Vifx1cmYUnGeYLlluX+f
9z5oYVbz3B0ZZk9WN5P9aP6tm07HCG5e82+2s3r0q/5rDIr8qAciiEASCkJyb/GWkt7JgiDpFTRh
ZrpPHdhoNYOwRdemESpVUQcd4Em9rIrNwk/B32ESov7kRcIZ6NHrQZruY0ddPEjsACrtjclRqniT
lw756oMVr7B3Qw0FGHemHMjSABhAh4Acz5zoAQE/6y+cf9kfHl+VCmUz+IRagsEtijKyQrTfUn9L
kpj+L7nV7bTFT1vHATc25XIvIXXXP45HpIpP1fuTyATWyK+m9EWlMAI2hytjVuJzR92mTpzzGsFd
JCtFBf/JbbSR1HHo/MU4S17sEfYku8zkgajMuekdikS8Ak3g245VeKG3cFdX5d8flXjRhcXGGSTy
aupER8xZurxLn7108c5SkcH+MKOYhd6KTJ16ZXPPBqp35Z1N2FHIIB/0JLi3D+f2qUfTjMraTM1Y
PzqZsf3UuFFGn69d/KMmfyfKVc9t2+c2qP2jRvy+1MAcurX+IHPTvYyPEZtXq/bJCka2mj20gEQd
qt9rDsB8exYuvQtVdUogE8QGU/KRszuXNNq/N9zoTcSBv9Pnk1Yx9gMAwRflOT1+7JPFqQCwZivy
WqxbArogl3i+CuJIlDwRnXDLmM1oGK2WHg0pGwzLTPjUVUONWarRb3tBFfS5U6RcTvzsHXxLEcEE
mUWqtbEqkxBKj4pG7hCRvYlxHXw0+GB80WgPJ0UaSYz+V3uVvOPZ5dVNyNx7T4xDYTOT681YhJjl
mCVsv4mdhPYNjHz1RXTg1QxMFM65w28g6wYWsxxzoVYeC1HrtTSYQmkM6/i1lJ2pXAb/6kzOok6r
U5/Tyv+2mqxTzKCW1qu+sUaZDWgO5wjx7aR+LKoMAcijgTAwexIE0Kvy4VcqHqUQCqDatHJBqYTy
/UGDfWnc2MfUUGag3Q7wRWxTCOvFx3zR9trb6y6KZ2T3GStkpk04XS3rZKvwBscLlIlqOKXzpl3N
kpiZtyL/eL+BVMwXmLz/aKCzScPCz76XESuJXDSO52iJP2N4vboAzEJ0RCR8pxgtmxHzVRbjEOMi
UL4zo/UAZ1AtMBfRgSXC+owQRwfzL7M0gMc41qI5f2XihxSHlhguJ7hRLTphsr2E2KgCf2W88fMs
Mix+fwICH+zUMcnV6iXQUBwto/AYNhJ3R7Um5fDivfaTcJNiZPA6CONo4OIaHWQvaJQVG/+Qvay7
xemGvq4B6czieflwq/cWJWC0dGkEjFnrI9q+cOipQN7/PZQSkIq6t6T7RUEnajOh3/60APr3a6QB
uOYBDXBuH237blKkPpcvZ0BuiMb0JOB639uuc3h0iHMs9iMJ5BI8VNngq180CzfjnL1M2OeGlJHW
X462hyl6CQWvOagHM1MmY6ZP2lw3EG45GcMtaeaMqXMmKGgXallcTgD+yTcUiDfVAO69KXn3xdvR
5b4R5ZssGbrDFg33aRU6txvo2LSigx3cYf4NBQKIobWV8H021QVHWwIW6vjGebHpRc+KFRhWLK/+
HS5Kcmb1l3OtNsx4EYTdnHJhAIvoByzp2IFF3jEaH3StHzI6kZy3uXYQFKqoBUE8EAKg3BiGliP8
563ShYTEMBrFJOsf6/ksiwb6bqxYQdmgxjSCA2s9YPu14KtFOTWuO4bICVAUkOx9x6mrVqS1nbUU
ua7iI8LtyZ/y+++Xu+f6mW7+GFyAY9XxufRrfygP7SKvtSmt4xn/tFv+pqCjF1spf1sivHmKfdVB
0xjfL65D+B5dlmXkuunuiFJSKNKZyp4csf2MjXSpH25nGiBsl0dNu0AkcHQdrs3ntHZ1arVtJ2Od
2dHPcowTojVCwo70eSRt6tCCZEhpwJ9jFqt2rpWTrvS45dw0KBPOWtwCAn9v0BCcyf/p3Dto3bf2
9ihFF4uROOlMq+gXzkJ1ZvwXJsyX3AinM6BCzfzyzxme8N3kX8aZNwpKQ6VYekU+9Jbbhmnn9PzF
32YP1qBU6IK2SbosXT9fqY0mrh6b2N4WYkNBWBC4RRjJaP9v2EzW0/NHeMsi/Z7RWjmKBga7CoVr
nUdHNnKjZecYwXgZL3veWWSn0QMLu/cwF8nOLz7XEdSBWE1mFfKFO8Av88whpEwshsmvAsm4HPxd
w7CudvlQMt+dGr9QL+eNM6VL49v8v6QcsIDyW4qRHiGUg/fs57bMibgT34g+gQJxaCbx2a8xymM8
a90gQuc4XzRXyvXMiyaxoSNYI+gdK+JwdNkXw2mmqp69a2w6D4mweZ0iEltGy6P1zCU/i2o8Roe5
Q6rZ4F/QuSpRI2qTATKK+7yLFENgPacTfbxqeNn4OztFqxljFgcslgZVsh96elcPYsie0bXE8uX7
WFT+3hy8qJFJDm6rNys+SK4fJ3hYEhxOf8wsjpzIsXUdqoo9wNy33bML7djrdBOqHHbRjwXPmaui
RHrniDggJ3xUw36GqtdkV8LYfdd+PLYRvlXWRCjxZoRJjvmBU2w0Gpu1gjNg2cIoHf9AY9tHkOWI
fbCRG4i0q26e8ccmXzYYsxSR2SmTxJ0hnCC2ASmJlQV1cGa7VYXTjzau1k7F2nxOG7AEoFIVAZ4/
GHWndqNd5qn3NVq2VvffdkuWSusC3NphMQqwLIkUT6StZruKl6YOLbbICxUGHdtkiN5Qgi9nDYiB
rek62YZDDO01Q6ySaHlfOul8nCoTA5gNPxQI2l+SjWvIhesk7mOdIBLPXzT3RAEkUaeJYACTsIEi
BIDgDJr678P0EFwOc2Pd+NJWsAh+ZUuIRUK+vonrrNHfvvZmO+tYqS72BsQGTZwO9A+uO74YKJi9
iJ+wzlvLE9krttIK7eHHXqByV7Y4k4js5/klfoTFF+ti0PtaXnK8TOnBAcUmxvWuTZ/u2dQLZlZY
XNu3dZ6GW6O6lf+NEbimciZ1piKPiv/39hEj5y5MH6+5Rqvx6IKqlDgUTfjfqn/UO2j9fm7jw1or
VyoiVHfqs91gxksMoBfWXTZ9mWdcK1ZBBEoHDGzGc6KuhR+zeGdDaMwP/tJCYIKP4fdEPfvPB37h
cWmMhqwb5GzPu4GFZTPGB9VbvLUudybVJlyMJXmxOF8S1WoC0nWvpTWrvgBYU9yPAbBE5N/0PFOM
8kZYjhn5HStoGon0/h8rD3r1u/siAuyGdglYaHEWAK6MCDmNNlvhEobsvYQwCMOj+fWpWJnJsYfo
FUthalhRsqxtSsPzZbiQPZZ5MjAXUlrbwhgbYn6f9M/qxp87BAUEWRebZwO1YwzUf3BuxKR+7EKa
CJJZHEUBTSrr2RadkEKwBqXxMRgnx6gXxPyvyOcNCL++4d/SLpB+QJO1ylrSOW9CbywXK7Det/eI
V63mEzYVwtpaxuDuHGUY2JcHNzKYT2E8Iqo1iqus9fg52mN7e54a76iOKz8+lncMiAW7Lg1LHwg1
0WeZbj8+Ssa4jZ8a/oQw1cL79oIZvZ8XAt7w1p0loD+x+hqDIQTaVcxJZUcYBoCYKzWIvuHGFuM+
l7xfYuCXFpEh5uSJerTsQ0OIi6G7+vSrYcNtdili9ywtX1kdzYaAmvNfb79LYO8qdcgJW5uyxK8T
9sc23NuV8/TmXQPrR/bcgZNkIcwrmia02R1WcU4nRXZ88RQ6u65hN3+/VlgLCPb786DorHi2YG77
k33tN6apSH/cuwdxiE5iLn56TSg7Io4UehkD3qa0XP0EL4Hx4VrTG5eARNO4gyMm5aDR8KZzATNg
RTdxMD8oPH7/Or7vp5GjkphjozpmKP5807wlMwi1JB5uNGUvO0I/LL8ng5K/uAr5ngb7agtptPw6
NMBE2J2qPPdJL1sOHccHDrCETQFDOVQ1+7Coh+rPqS/5hDXKcB8O21EEG47mPt4t9Luo7zGEBms1
OeTXlcHgNNbEFKzgIHSGHAzikA3+lbUp1RAGjgVZPX1wQ7wnJobLImALZ7NM4RoOt3ih+0oOYPgx
lZzBqVPkYtMAPcgnBeQFQaLp6CnPUWwQh88C0vMpEp+kMR+GeFEHgSX/IFNYL7TZSp4gGjATvuru
xIZ9jBhKth7GKUZnzZIcxeHXV6qxqZBz93sZVFIKFAX785P9hJk/Wm/h4Tqt8V76o1sjbxeQP4ta
zrLAo9bVrQHPAUVM7Eq5reL4kHE2RC7GT/l9JDQ2ir3X0m2E+aqYOgNEj3ChSRc+KOMYXsE7wyfS
5WB+o0QatCO/RratDEgKcj9G/0OOW6HRAzxj6670GqakQXrRBxxva7Qx76o0r5qve9RbbQyDRKYK
LQ5VaZZj5KrSfPAPGa9VrpKQyEJ91pbeBchiizkIPXa302zGuP6Cxc8emC32GVAsatWleikYTICM
u24LQG4hSzw6g1rLbYPZC5/WDMZyGRgmJHaTfoMTFx42DcZbVTERqVl7QI4mYOPGb5wSMOuqWqlF
/cccmQr/3hVtyMbIW73lShQ2hVj7micmfVUPboxav/f0sT6royzpUpl0Ll6FE9bsuJszKjPSK5MX
pdk8nebOogUE8BzP9HyBN6TzeZyghklKN29+vC0A0XoEOfr/pO6PRHVayQi5JIv/tsqHUQ2CClwq
xx/8Jn8UtVCiHFof2Sr55Ejz1kgTSaYAEr4wrvCZOycDMupcV6CyaP2X/VVJE6UzjyKyWXzsDSr3
1ujImH/OPsWsJ0KO6x/7CqZAyJxhzrSNdw9JG9jSZN4m8tlXquZsIbJJMdRq8gDz/vi3JP9FGC+u
SXKmwD29oIjchDadb+L3rN6OganGwsNeofrA5Mqd9cmTzynVCFOj+F6vLNqMVRwlQTassQpKpzG6
AIM8nhZE4ywJI0KIBI87oKKjGkZW1OjDKew3rkcyuNEJwX/6tYF2SVcUfqHfJkbqMOiE8BN1mOwe
mOAJ0ftWaYpFriPS5YlMOC9O62eMnaB78RFDRiWLadAWsffK+PBFnVHBUvHsBZNqDwSRa963+Sot
A7fWvdHGQrdwhy5Oy6e+BAe2Mqr2e1GmJeU4A7/Xb6ubG96bbbYooeu+cLqBXZPAa4PX26hvZoiK
W4DjCsFLUZv2Hu6gwRYQTeq6aTzNdhSSmcXfQF6VxjjyX/dcve+xR4rI9vSNOOFUck7wLMlQ48M9
uxFADDEtrdOvDf/AXtOUUMKsy6b9yIsXgCZQEgZRG+DXCWWqQNkeWZs74frSDAsB09wL82UtLNFq
DAEIbOpBSawWmhX81I+Lmf1B1lekgT6JjnWZ28fhE8V54Q8zpIRjpRtEXR7+rTJEFMzTixFmkECs
/gVU5eZvSkJHuvYU1pPytcV1/v29W3kJ6WrhyOEB7RxHUcfmPPgaz+IIFY7jQLDajTXz9ZFf8dfE
VCkv5vRNhHryeMmt6zuIZGjsFCmPmeeKxENIg0wFKlEnTALGXBMsBVng5FSQ9uPQmZQTAxOyFA7f
BboNu1oTp4/MaJzFolzRhO9MI3+Q3VCPOb+KDFKAOnu/VIdXlvx99U+ryimBEdbNgv8BwXlql7Z1
zlf0YSnqZ241mcmE7vOwCXGU1nYQqY7RAYrF760DvVlazQG+tUS9HvCXuzLzehP9odNIUJ8FAMSj
4SoIxicyiE3Z7INOIH1R/+mEVWKrndirrSaEonZvL5gy+NcobnteHc9PuzHm5GVnCpU6S28vxSuK
vpGlH+1Ch+napmzwIk0QjGXSi5JpvGR9BdxqUI37QpMEzfTtln/wIf6JwpHsQbPXHfVqOiFbXw4u
KgXC5gMPspTL7FIfjvw20MY7G/7H1IKNx854afu8OxUGBQZGLvCikNh0Jus/nd38H0rTKiH1P9H5
sdWkxvQKMedcTWkSwKrNwKiU+5oIg3JjIUr5kX0i2dEEQpnlGc3Vl6ecUD28vFUy67ZtHnvn0vcs
BJNwjH5AVWBQTGKEvZCpKOWxOS+w+b9KYce8kjpGhWtoVTNcwYe6O7TGBhTN3n/1ejRPt4VfLtRA
Xof1amweRUZaHsgOAB/6VK/i/XiKJ+gIdbnXZHmfglU+Qr2l8s+N7D/7t0R5s6K+n6psxigzTrjh
RP6CdHHGUYM0Cj28Im/skRu08xNx91d9pwUK2sLc9sJIKUgcWuMCUmOGTF9WN6pDtT4fyU0KYCMX
oPFTOuyLqQbKsG6MltrvYkaRk0ZZD757ueoXir2+mjJVoGtDZtDWENx4XdubYlEKFXb+0hMyKa29
Mt4pvpbVvBcWdOVd56M8PAuYij8cWC7jxwYt2atXxsnIm6FW5E78VA67QPmwt6Ywi9esMcYlZp8X
fJ4o6mD3tlg+D40PcRX3ZLUnuz6dMIvOkhyK5N7VSJfKBeOQWYzPjykUOghHVlMFECGHhFUf1QA0
8whFLLdvg7o43u1USJaMsFuZP8sif5dXM7kw1Kc9mZxffIwdHzX8uj+iqSyLu/T52HJ2tuoEdMPD
56ZByEY4yLIP0W7aLHxuBJp2aRkcEWjGd0YnSHegeyFzaQGPi3b+RqwfBGDUNXLOq6ZKfq5OQi8s
0HS5B9rZkWou9V7301gBQIb9dqqMCIUR9vLr1V/RlnXRwnec+zt8VKPLhnO2xq55dW9ea2iLdgeh
VZXLF1wtuh+WUBM3B5kzcXP9Qa8ZFhynxPIim//vhANaLloXtQpQDvj+Ag46j690dnFtBndoUh+D
zSg/EaevdA3YTLJX15spAvazjNK/9xtzsoepqem8WWcZVHeSEp2k5D2qQb8bSjlMaTlSeOkMWHXT
wHfdEnz5NM04GnIRkIpcYvnYdHGBbRue8SnG3XXcA3nE5bxdBv0HOcDUa5VdhnGp9fvWY2jKzBpm
c0mjAuoO4dOKgbZfVaL1Xi2F2W+9iOc6IkXIL1kdZgGt8qttqDM0GjxZoABEQzTLV4hFGCt9Sm2g
jR3NIBEX7bogU7QKsj3Qiy5nRFW3nBCPPPxkVb/EE6smohNFvz2ffOiJqbtlmoSKFA/QAiNhR4BP
0u7Asz8hCGY6WirVFCwi3WD2m4PQOWQNRa9OBsg8rskAgz+ES8M4dWpNxxcHaAJO8am/nm5uNAPQ
vV1hBLWC+ZVtdVrRVSwlcyd5F4+dR1DteZqgj+81QuZLdVW9tkvOcCHvOZastbj/UI2WXM5nZoGb
AVFy6Hh2zo9MwW8qyqGX+AtfDipJjoamcT7yEkgm1w/7E3uDHtIa6VRBn54ClYXFA2RB6ksAazS0
ZW/qBRPvVfYt1UOqXM2QR27pacwyMa9m00sTheXx9PVjtR8uTWOkmUKLNKWdqVBfXZ5TkMPP1SCt
S1mUVnzFD2Chbc9I12qFJVF1wMzbO0fYUMBhP8nTS5sjxhddIxLTafof1b2A65l4rxLYi9pi6BVH
9biLP4U8Z9kqlLZRrMRn502CeZtXxYp5nxRg7oltKIaEmv8OAZG0UptRRR1tyZFXi+qOSM63SWNB
01j+2s3XKByXu8JXLWNo4QLNlL5OZSbWl9NR4zc3IQMIQgrRjAcIT+RY/4gHeFgIt4BRZBk/+Lj2
xf+VzFqtAQaohiMnfxyKYvGU+BxNUfH3+b+cemFMweB98eaDg9o17mk6f8kKpSxpRKFJgMpDAG+a
jxJjkQjZI2VpEUM3f8KdGCebbNBeDgdszNTLzVUk67YVpZWV7AF7Ib6BwAUEi5Ke0h6yeAn5i1LR
CfYyic3hiaijCWTOx6eq0Ra7q2TvCquajuTcIoSbsUiyv+NLanNgCibzH7lqyEYbqJY8kAkprdRV
8JbtRHT40R2JhH2e0JDjezNfcAmbghWWcRcZVJLey4ZmQSjWhPlsOlf45rM+gSfqUeATFZpqregz
CdxcLc/oev31N0QdhqcJ3uWscItjeG45A5CZ2V78+HsNAmv+4VGNQ72ETKBDdePk0rDmI30FZOmx
yMKYrPeoXJ077gyfR51AFkHC8XIHtvt5fVgx/N/cWqpko61wEFnM3N/pD1fEQH2errdA7ZqbVWeB
sARS30kiqa1sQQqt5h5wv+UFbLwVGDsXWPHAC1aI6SyVA4vFBMuMOXBqBoyhnHuSzMotajSzKyR3
qUVaVpYNUVLGmKx4XC9fiCVg24UtuWL4bxn+3b2ur61AQbS14JJw0TIrLSl0YHY3PMscM/Xx/mjd
RmD1PribUQAXQL+/KPGfX/I4OWIo/bA+UrcdjFLBN7DBxeVms5ykih6pCOt1UKxaufvUuGv7mooU
KUy/8C3nhw5ru8KD9+m5pkdp5JopwayUGukbKV67fryL2xRxuY3TA/BMhN9HM6qIErUt2aRq+YCq
9uBjLtP5byMl5bCnRJvJxVvnMTEc7ysd0zidf2gZI9Du7MMB/adXJgDotrTIrNSRxJ7NG+nSp60X
QM0dQ0PQPYKMQX2h7hEfC61DgXHO77/hwKOakQqP/IHLn6DjDS0nwAsAheeWdryjFnufczxMxMfY
cVenB97ZXzT2s2nIhTqN/9j+Nb6yYG+HpdhRkDOddsJoIW9VEBquFvBjEzA32YHkifWSS3+47nlg
yDNP7J4XDuMLAchKadrEDVN8g/BtEZyMi+BCB5k59jxdLGhFY5DjQ+eYObvq8kWKrpqOFnGSlKHH
YF1PEI6gD5u7ijVLgbF7V8INY79jrGX+j0b0ZoAdIG6qGKwN4drWrnIdK1CvYmw1WlsFFplK7cy5
jvE69p1cMVx0EVfjaszp+CudZyrgj34olWfJV23aGO86fWg3cvLent7vNBnQo+Q6gYlMJ0X+2cA8
9x3XbdVzuajqHcEvk2QI/Z7Kd7bFtIJsffojxyKwEmoFT/R6a4LUWjCaZ7Up11vYJgDLaMSiG/LM
92RY789C/+RlxTQ1By5E0/9jncIcMQ4grkfH1s6PUursm13uUNmfHsvR6Ny48FhnCT5WwNknKr5+
yJxUNnYQg5zPBdIEHmjoK7GTceyZjH1NbcScqhV/ngAmY4LjkIQfTHaVsZZQMc6vvC3vl9XGw012
bzyKEDmdRXWY1rCRt8QO6WfPDDhxhWCxeOc5OMKf92AdRSSAOXULxyCO9Wf6bzucFbU/Cl/YYqhG
lPipKtJq68VpCXWFY/TlJpREdePzI8RsNXAmW1NcUENCQ5u7oAXfoiN16J1zRT0iqCvNAwbEYXDX
++OCWfuZ3zPyVQ3HJ6GHRKjiLmsTc1gEUE2xycSqzs7pZVg3K8VaTNP2SSm0Oxv2JEyaklMVBPgm
hrPch3v6gA5QBueTPhbOObcxGNtsZlJuKavusbNbc4JWY+pixcS+ipRvLuNYgHkKvTZJ+yCKC96N
rt8mrtGchy+HV75EpRBK1EUGGCNzVtMC7UBI9lVbQoA+gy8v2xAYEG1ARJ7kfjj+fcRKUO9kLeRY
bQQY6pL51fKyjSPSG4jPbYbAKJhLTWlCDqi7f2tOyruTEd5r+xXuKdq2xe/WhxH1VfKpwOO1WNsB
hXk+rEPzJZRiGBbFa10xHzNk+XGXDpk4FnsATUWWhKj7EnX0IHLbaMCGW0IAb0mX6vknfTZgdYt0
NrBN0z0b/6vE2+sKUAGPUyz2MmhGW8vSejq9epRMKkABIQHigEbfreua1CKAPS6GABj0Kye2876d
zDm2Y2DlnVjLT8B0YptztF5sO/p4bnYSTYfXqoYZ3LIXpMSjWCFhqaDCHAhIUtdcDNN41zUvzou+
GXs1ownFja37dMaBIAA6IAao2S85m0Km1OCx8HKlMNIWh97o1C+p3FXtwK2/eozrSOeHxQB/Bxps
OJ8G5lRdnIX699+XutZ0LTcBars9ooBxItlOvATr3GTxyUx4hN6stPm+raKbkrK7fBU5ysAQ8xMH
RK6zIsdESSE2Q1xti49hGNlT65Nb4CnAQQl6pOcleiVL9o0o6Lyj+y9Q56d/hwXzZ2034v9VTvqm
ffM5Js5OQdQO3tZuOqeLpYFgm9F8f7ZChfl7nIXV4pGE0Q9+K1VHMmUqkY/HHXCWdADf5Mr2L3f3
gwgqY3b4xhQrB0y7+uoxC5kej2455qgnBFWfS0bf3WQ8JLrejP06++pDY5jL4nzp6BM0vfwbTgqa
O2FA8qHObYBdU1qoo9WCcpFoY1JZuUTe/vfwTaLvTfZCcTg3sl3qZKsECa0tZf6/DCL7Z3QAhfSS
LCB0s2j31o588vwyyLxiVfRL9++sT7HF0GkGxVg8SjNaq0Fli20i5D2cUnlz9mSpbT5oYvbFQbSa
f9E6+cxumX77kG9sZ77TPelNbGIRwiIX8rtAwgeefZer+rVlcKMvFD35AsW2bAGaXFUYGIh1CBw5
QgajuG6lWhkBsiUiT45Z90SVJI+92LCMmmouXef/1rVoJdZxIRG9ZYlH1eW4ZMO1tioq5bVQccsj
2a4jUwa9bFqr6eTAPiYYDNBakRkwBa2NaOn1AxykEeleOINyG7FAw0LFWp7yf9K0gXyY+vgaOx5a
mVtsN0MR/jiH2m1PRtLUr5Uok6ThseEz2ERdiaNueuFrJ2M1jMjBBp/DKDIAUhuzq31kgza7tqyZ
TImw52ip8exRg88knpSMGB55PJWPJoq8GWJpSglpIQ/a+lspA17YPwWFqE8tXlukUE2A0QidsQws
1mLQeTeOyJildJIhzzyOMqJRGcdRCeGpn/jPqd24SHzWr6WO1jLLil8tM4vnelqMz5JvOn8bvvGn
Jtj0ZBzUGLikHXBxhb0jXbgS4x67Ei2MHvxLDjtOH4ax+gHG2YHuCMmrcF3c4bWCboNTTutRe1b+
ikUcD50EzXyXqlbwxdSRcGhA42JpZVsdptCMPXZAaySxY/x+6R6DlaRFOIzR/gTT4o+eUaou82Ca
u6SgFst4yWf1tNOaRsqexi1mARLPg2MFoIKqNFWA23hjAQ1dlrobOoasqylpbFKlG0BG3bbbZGo1
ja8T1I6lJvZrruo12KXTFrAZ47gz36AITP0qYvSuxh9aYpEeBd+r5L7iHFHbk5DAHbFAg4yxvjnm
9ZzvmWxHCxuUdmN6CCY7tmXT2BByJ7A2XXfPfEZFkhbGCLei2apoCaPN0NKOG56tUUJFgjozmxdg
zidYsBXcMIedvvkGRgwICoppmYpQ7NyYdPMXou4baKvrqYnOOBAf5TCFVe/iPPdA30yCoM3ncFTH
BRqa/PHVHBpOc+o3LRpRoIRFh2hWG6NKez70zVZgn7/eE8qvesblHT3EZ9rw9uZnFzHK61M3vxx9
Wz+SjcdpufZWTElyp/aSjA/SUdBkfQqP7k6fx3lsmFxrCgOUAaC0DUTT4YGhoggZZqvA6ku7H6ns
Z3krlrWg2O5Rfn3xoLZ60XTO7EfJLQFBiS4kNdyBlpxDP70aDSmCJe6DpA8eYN5iFlZkhiXBFhTv
qrpb2EXySDqZHRtR7mbx5Mf3yHQFESuRah+U8VrcoifyFdoVLM7CUui6KM7+3HpVKQrWGenT2l51
E/7Ly6l3emkxU45GzTbEhP891SDkRVkSJunpKKuFXj60OrkaBfHHrfjau9nj9kA6WRU68kcldMGg
48i1txTy53FPtP/3vCOmTMUEeZOqs4KE2ja2vtReCLHiFhfCFqePTTrpHMwP1LvZPW9LMvtqCpj2
33E/2qjCjXSNhSAJZ1Bz5JzwaT6o9RfO1JVZkEB2CCm7+nyMhupSyP3PYw696NLB+lLBP8Id864x
hWzheeOM+pRAYOfQmZb95PV9s4C3UjN4pW1qThwuXFbM9w/yGo3/q5SsdIZGRAHDfp8mEwGyxk+r
Fz9BI0qBcUfjA1zZDQyaZlAAR4o69aC2LxD05hv/NTvddOA0EPFO+Bqh3piGxwjKTycr0bVurE5p
lJnZZ+DJ4fdDCXk8iz7IYQvJWoPMn6y9Qm2KdpKj01Oew/eXEUt6a0olns6azg4fXZH5OZ9cO+3q
FFNCCl4RyXetQ6DuX+bfDm1I1US6Fo0EApTUbWWb9pRjudoW+S0cJ6ugTWL8sKK9kVe75/CwyAv8
eYU9KdbPAFuzhnspgfE6gRJSApq2vQ8uZQPDDSozrXoKvJE6O8j/8JFAB4GTTEYw6dZW/QpyebtW
yD68Eh0tYFUhw8vhdqDfEi/q6NjdOk60+uf5H/6j3eXLltOfSQEI0PCoZrUSUY+ghGuxpw6QDB1G
zb7vIWp8eyaBplhZN7eWTV2Ede2SiHwgQzgJ1txe8GdNW9gmvkQCVzVbmHKY7gt+lfpo9T6FlB1n
7XhidfOvfD9t53N43/4EU3kQSxhbtC8QaF1CaojAHRUsPgyghDYeh0eHIj2q55k2QEPxVxbDs8VH
CxAxOPyA3RKZShSVs1jj3cg7BPZ9OeD21inb+nDwrKpC7/1s/rUlC5vevW0o/151hs1nlQEOFVFu
aqWhcb6cWIIbELO61FqiYYaMlamJItbIZCWPpWYhtqYbfsABKKgTZr38pUFR3/sJ5kaU9QO5AarE
ujG0Y98bNtTIas4VIAQLOePtBFORw5Rw2ygwa6rnJXsHJNDVbh9WQNdEDF0Q8+YOigG5D3M+eteN
B5dNCMkfs/UvHDWmzW70zeXd3s5J1+1ZJTB5ghdrQaouMXNM6WqqBGw+SjtD/J/c7+0hLPd3ebNp
zYescNVqRKwiJpH70XSBDOVslcUcNFXvxGq/Uw1sRARbZiBFwLEvIQP+BlGbxv3EoAout1kW7nBK
TTL/1NlPLYmk58S+25iKNtb7DpDM7bXRzmRUphuKyQkphMktHhYarICwKAa5/hImFZezI8LkWcKd
BJ++sd6WjK649ZwTNG6zCb/lCDCTzSKoUyLTHudTfE28gIVKnsgV7uQ2p13caWMDxDpjQPba9J7r
OJez7isCHyyS+8+n5TOB8j8Pnx5SwN2uPZbVmTg7K+XP18llRH+mFP23qpLXPiJxM7txFt9j0hfO
VNbiKtMCgfUrCQi/zMMM1B2yuXtJ8G/fX9o/2DZrY+WdlwO81MA+M1RkEoRbe/o8Rp1Nr4ShTj3u
Lzw2apnlKA4YDmuLiW2GWVzpXchZ9BFAXVJ7ry9Ggy4HHPTcvhuOROu4gMayVGFvPxKSjjxIfaJg
KLKJN4agi4lAsmEPwVkarWhTjt4PK+oYlOXxQf2IlfSzwNQfRmcI1gBhzwhqzib3SA9THnSfFHoV
M4VYsawWyEUcKxM7rN4T+ALSXhDNzYDqO+TseWGYbSYHdNuJlkK06g8XqHeY8QqUoyGsB+v3aQln
EO6/nXyc7B/XMHvLIhClIguyeDIWMQlAhFrEzKEZpWv7yHB2lmLsbF/J8wd2dAVRU1w4+O4ifxEG
yXeu4edPReBwr2QUHF7GAtL5NbcgUOlVWjuU9yLFhR6x0ctjzHix3JkvUX+LOYKsnEdz94m1zPxE
SkGX7Q70o7omRnKSyJJSIL/EpQNg5EGVfs6akrRHRUEnfvXYgSGMAGOW+h9NKeWiQUFO3PGFRPRW
aFIMQzbjer5//Xc8bLEN+21rws24bnoa8Ngt3C8rFBVw8hc1oztjyPkDfZxff1jSwLrYNH3zIzzw
ZSImS9QjvbqQb4+3lF9QQ5X2eVbZjdjTbytVC/fsCXunVfNHn/AoSd/5NLtjU/yehZXBs+NJGbSX
9L6UQ3iJzQhmUSN8MbxF5g5nnurB4BzdlZxM8RX2R/A+G69vn3cVOcFtwGcvwwk8AOl4a0UecLQ7
Fff9n5A4TkeKIXAKNJamL8zJIhpdEVzZRO6tyuEol8wmkrQvM4hrVbPAD4t6Ms+Os5zB9iMcbQ+i
UfM8l5TMse6VHyeeQc3MZnd2dwASECjKiCMPFfUt/TWv8BlaVhRVQzzblS2AMfZiFsl+bm8PLNVT
TcIruBSnFSgYgHZartlCqBVfOV+OBnd3c0o2x+9s5mWB9EEv8C3mbN2CdpH7o0+zp4ajzq9v6448
/EzwQX5gI4wsXPTWIMOs54JyH6U3rEMTEh9otmlzIqZmVltSiK1n0u6Hm0DZ+UyIcT4sscMV2Ec8
jyVPkGaDUw+1UJD2I2WMG75gRJSbTnkIpXOFpmt4BMA4ZpdvdmLTgRuye+86i76GgEzpM4ff5fey
+GoI39DVPpgfus2gu+9M31MnLy+dvZ8NfMNFCEhikKtodeFHQ5FuNjs6YwypIh6vr7NtbvHTMwh2
wBS3wMmwtHno8dt4jUuRLYfT1fmX6euEZ8uY/4e/ylbYfpaKZnE8BCQxOGnnspiwBbTZM6+id64C
qADHGMNUsmP392c9dhM+195M6T/pjiuI+aEYIGo/phb8Re0sfhoSy1w3ygvYa5VxNyb5AhLLIaK8
KRCmrjC4JKUk2m3ZdjBTKD0LtpnnKzWWdwcIWmUH14+LfGR73JRKMnAn1Jznou2cf1DCYrLq3wdy
B9aiuLgSvREFQAAQ3Yu8ziLdvUQd0UQhzQslNsJUVUD8+7Y0Ah2v58umKKRwLfCmbBdq/pzBURuf
qnQwcMlqjyolxDDhsWf/hyr48hOOtaIMAPIHt5LF6XYfaLbsD3Ft11PEwX9Qvptv/KwQxMo7rq6T
0g0YdcIiukscjg+L1zJ4xcmfKgD4K2eQL+3aqTrLbvVyQR95hJPF0CszwoNZNN7px1tVMaf667TV
NvG94Gc5qUUQsDaiUoT6zbxw8o4i3ikq7RtJZGL/DCOP0i2DDTRLRouLhQKyyygcocnofVnVOOtd
OzrQXw+CeRYZUdQO7vbGyu0N+1M9jOr40ZplnF2niUL0AvCiK017x4Hn1DZweUtGeVhZ2Jtan6Pa
TQxg1hmlqQx8e245wqbbdGmPTC2CFil/cFhIXaUU7Z/TWcRJ318KIaJogkZE/5CNlolN2i/Rk7R1
LpP76SUqbaRvTHinnxbiL9IEBQXyBXgKZuJPHAFV1k/OzmIjzyik4LW0oKPzd1dbh+vSLjC/eInc
CP2lg9oVfosd+D7w+7FFv9J4N098geREYlwqaLigFZ5ViQiwyCJ2J+KQeXwXpvd54u9GswBZ1Xx/
HRZ5zBf/wjYrs+bPc0DS4n7ViDR2ctuXj6tPB/eTCo6zCSmZdaEQti5UCeHnwqx3CnqtaC77Jfeg
iG0qgX/LJv9OvaeOYvW/t0WEnCpLNH/f0CTkwemQXPg0MV6W6qibFvpRUk69B2KwQjQbygATTSq8
A+KWpHhxjVZJeRpZPbU05TWYG60XdeW7zSU3UHHRqFRIu6LNVeBTPIg/zCcV0pUajDQTQ8bdCEET
hmMuNOIKkYdr8ghP2dJPKWiLvyHBCf1br3YxQO3YoGpPcifwOwf0V33nqqjwHFVqyGjfsrWIeHwr
27Ed2E+Ug79/uq5I3XO7d0KF1Z6R6UnQq480n2RmBSiyTIEQ5pTv1eVHuvHdYZgGvFmVS1K/saZ0
glNcVfdquknC4TALgEiSlsO3ZeNAOnhUUluY5XBe72qR63nREAcfZC7b/2gB2wc4JxWbSZYshrt/
dUno+JdYg4XFVQV6kIA+VsbgmA1c3hL/+WeqncT0ysVwmeMUUqrDb2Wd5dL4riIB7+Vfkf6PCfo8
loR01CS5RRHZuVQimrjEOcqGi9yTTTHvhxX8rA5Jp5Thl6hoiFWyrnHU+krre4nCXYoA01qP+kkI
ITyO+u056L4rw0tLqgxHmcGKf1iYHWbIwHqgGVGXaw/LwTTEVINiKOFbkoWGz0vVGYc1MZEDWGZG
5eQCIyV0lmWyGgaiPx8LzYai+wRDWIQmb8Xybu/jbFLAUHvsNmk55wuD1sSmC50lP3QB9oc21139
WGutphzU9S+DpOnvJA9HyDI4dyZIqtESZYn24+ykkAIoZiULiv3f60emUvP5WAhc1EqJQ0+972ki
JnBspvzR4FZ6iMjAJobkPsyIy7lejHI5zOSZRYss+yAijRjRWX1FCy65RY/vxmWH4ztvwfoc8JV1
aHuh0ByMgJC8fLvFzSQOSV5hWm24SFdfkE3PoCn06XklihH6pWZ5qBbGIYTZZ8ZJq8zp9n0L7ynB
o8NlC7lgk3SBmlEyp5HSubt9vyQXnj6/8uLoJ5klxrB0UeZtRmpHpbFfCK1lCqlMVYeFeYfmjbn9
1RXfGDBqPhuLHbhrwSZFl/JyWOr2Eee4ptxWI722Ekhg3GVu9pjtuhbDl39eF4Kl91p3BwjqkOA1
+/1/kkOLIWyq1XRbjkRyf59XvfwpQYeT0qLkLvmIxxPrVhYQIPsXwCaT7iDCuUk3TRALoUNkIQCp
Q75RyzGL8wT223gC6hOWYPKSAvuL73xNUu0KqlhH/CXqAz577+c0zOgji/p/JzUGRQM+mPL4dXeg
kRGIeUWnAnT9CwadIIBWthz4Cl304CfLzXba2u2IQ3g36sw96ZkUTiz+sEJdxLkaPUxYhymv1XwB
SbK6p6yp0wzh5RbzRJg/BMa2Xu3J+bPEW7qYyvVTeiOcA07D8Wd9vrVIPgQ9b2O8WSx4dMQVOtN2
RcnGl4AsUs6Lp0ZTI6n2QozuSq2Q1BqGQ4RJUXJWVDUcnqLfyEaQXAcAtal6IcSV4QQKobnIb76t
iUUyi0vWDsjOZh03KIwLdYKww85IEnZe8SsNOcPpJyYrxBjqEsdpY2wuEsyT6L7GnEv1ktZANk7q
7TL5X/eLA1vow1Jfm6TqG/kzqHJuueyUzhtxsNf1JwjT9YYitu4rWwpwu1VpqDba7QY8OuqoOMPm
SZeWA0aRSk5jx12+4iLTJmUXmfDXUUVsP0SglGhnnxfBKRJcpoJmcTA0uYkJWI6kf/xV9Jw9T5jE
cCW8ECwM5hjmQ/i1jHmsxYsiTtxCCND5is5jLi/M5vUibgDgRmXJrS8AP2L9/lgW9YZ1Hug3WitJ
KEEll2lt4oQvGJzgeKWqPzsBQnUNpgP4O6OZ1z7wYq1fT6iPYSz3I8zQFUtYDVLcL9Ur9DnfdJP8
tnvhbNdW7rMCj2iFapA8DfFJmhka32L23A8S6O7txm+tW7eYWr/y8JcyQsejADNN7SeZ7tYsgUG5
liFxzqKDAOJR6f6OHEAyqHj2QHGMqIq11f6HEL9Y9sqx50J7wT0EwUlD4WlDLiJ2TPpBbvlvnE8F
acVnPib59EQGDUyffBb7RCnkxppvSkkvxJj7YD0gzWifhTZgl/TEuSJMCj5+oY9j3Ioe4QIq/j8L
jQX+JvN3VhCodaZ/YTI84JiBTRbEhOt7Y7O9gXllxpAPOATvPs8D5LgeJRFulx2z7zBLG3kGViYt
wCVtMLo/5Tn9BWw7zyC8WN3r72VOz1f08XNLRZQNQNHWBddyYZLzDuZ7P4HwsNvcw8Lv93xJ2vSV
M12w9GNeT/NAh4w/VvuaqGEb9pw5TKHanImVl4ByPcE3Wu1j8wcSivBR+88cRX76NJ5qJCmvjlfG
sQYJgUBVqQK7OHVu2xciBIhvfkrqhm4iy+KRIO4JgCOcAMJ713y3It9zjMw2fNNkS4nAzafN0yyj
LvPlPs7lzOJ+ffFM4vdK+/zbxi5djFdGzincN50CGxfeHzEzUHPdtm7tuyQvCCvLVy6exGQqxolb
g/vAetGSmRYrMKQSHZm5PCu1cC6FbxuQrefqAmH7roISdsgg7vINPE/K7BaaLtfVoPAJjS8TWA9v
Cc810lxEZ608qxSMUP5uBjErz+b03ZAF44FkPELS4XKRh24Qs2Y/MW68phO5jECtL68cEZ+BYCql
UoDlc7djou6TsH8r5/AuHDSt/P89LkEP0fcZV6KoO6Y/DIkuzzweK+SDMDP2cc7l3dNRaXblmEDj
++uDwWbVJAhIiwT6IbiWgOCqot3VNxczGqXaf7e+saeGRIZxjnMbJ7rZge/7Gwxi6AxQa4dSauVm
zswKeeYjJGxGKeUwZPYdyiHYy7sofrDtPBmYktiS/ikoYtOhAPasOHpFX6pwJrvMRL1/ZEt0iqQN
9yro3e+XUCxstWrympCiQ015dqNoPAbw5gQ/2uW+Tj9tlNq8kmEjgbwMCRk5t1JjOn7Sps6cwGwx
vwjC1FFOd3Yi3uoy7NrB3kcLDUsB85seeYjvxWi14/yRpD6bMw1V35ZqBO0z06gjgmB6Lqm8+q54
xPe5lAWQefiZ5T5R0aoal0f5QfO7KRZ0W7e2xOImLCYbX4JeBO8gURO5CH5jVQfEgfzwoxXnpQwe
5gxAHhNZ6/dc1/1X0Us3emIHQ61XYYBr3EvQIbfBsP/foE0wFLjKhnLCUSU6cdifF5K/aV/jBRZq
jHP6w3U3HGBoI5ldfSFW58npUT5BjtTVwp2E7CR6G6eO1FDXFR/p7QJ45+/taG/wug55/T3/AR27
u53zJF/2LlQtUzO/ir8RDhKMzR7wjY0qW/zezQFskOOuO0HuLlEAolog8MSgouOGby1LpEQkNkwQ
7OeBUE9cEIQTY7Gv0rYuSic0NUtAfmyBQyemwj7BWc+YS2vKgo7Tq1xhd1EKTIPBOCJxNtTRiqC5
Z4GbF13nhIQRy/0o71cV3d/nOlw9QLrIKL8HMEikm0dCoDM7GevPQRsSblE357shHz3A3c/vU7fx
QOUXYTxPrVKFBahl3i5YZiFVZgu3T3T032oArcEzC3sQNPD+RyE7hP45z8+XIhwbnz5Yc5J1ZvKN
cTUH7pQOn505FAbHfqmr0C4TTJ5OvOnC32PqOZC09M3vQg1kj1cpTZIatx8tcVB9CMlB7DSOo1F9
BGTNst3MWSfou5YBqg2gzUIN3RiMKYdYcUCYnR9h1zHxQEbvlhTH6siBHaddOtzgZktVw3OWswpL
h0TcZhArnQv5yEhIsXocas/MTQWH4vqGvhJB+B5IWOcZ722WTwDpvBZslHP5ffcV+6tazJSa42MB
W2LqsMRwabuP78HqP/3zNG+wPe39rUen6r1Q6X+pcaptF0fGO6kHkxSiEBhW/kHCRiqWnIJU4Ouh
Rs5sZz1xoroxoU354BnxkSb0+v4jGYWbiE1/KdbHgwfaXvQTaEVBxfFxL7Mmad0MNHcKs4QpSoBD
8ZieS5l1+q5oEH4BWTtNAYjLpzopC/Z5UWEPdb+dJfKlScVgZUOMzYYV7u80ZBTpAh67dfl6rA0Z
bCHGbOaUFAj774IGMQKopFQG6Y2WAtMdBOeS6QrA0BhMKVggEpis/TiPCCmuzxURlaHDJeweM5YM
/xUjH4ZkmZEUdwxbqXU6diddXfmy5jxnA8zhQZo+HNj3WH3UkHV4DLA43Pofkhha6TvWv7hK7wuT
8dYsT2zByoZuujaZpkGriavmAdxVax2VMSyZ3M2tW0MAw038kvRBTBAgMDRovwWjQ2diURh2FOhR
0/Zog8wHSI32v7z3Ti1hq8p7kvFa9+AAXwjETYmBY9qIWprX1nrCM63zwX2snkprD2TmuRe6xkYQ
sVgdzDrhUweXHvUNTafHWr+HcKp0g5qlAQyLnlE5wSNQb6gMrochUu1OggKidnQzd0tHod0ct4WY
t8yxhZs4K5vBSyWEonqCwuT0IjBtlUuO+tOpHtw8mV2Sz1Fh8gtmWqfDh6EMNDdMBp/z/iaKZFzO
zATRDLf2iQ4Z0bm6CmxIFfkEe6zVX0FBEkI2egGNmMTiWHPz4RNtg6DpvR5cB3sANC+0X9cfuOVq
c5FxVT0SYMSET4RFmv/jdNMh7ziIGzRDRsPRiFkuZZ7lbSGTmH/Tafaw1KuQIP6Wagv+DnjjTehy
Pih+CQqHFrew6Y3MVUV8jwrIjNOxenEZUuLqY8VHKOqqxCu3X1iZ/jAjcMZUb+stUDFfhUjdiJOp
xbBDDneFzehY0rCXj/UwrJ6QeCULmcnQ55TbYr98BqsS54WLjTtRXhxbHZVM3goYhJ0z0Bgsp8AB
62yCHu4O3qASHnjYT+phIEgeyu/QWHprlvIfWQx29kwJ56ean+p7Kjol74/KZi5h9KB8dQ1Ta06r
2RDnXFrl+ezE+MNNhr5gswGQ/ZMGiYUiKO/1f8jHb7fCkBKBzzRsp/2WZoY01BazlXP3CP1RVvgh
FlBJ88mPalSsu+ZTo2kRpRVkRd9aymy1B+dUiC6C6XX2loM1Xp+PSmBHJzf2+x8uGFBebqyZm+xz
z533XPyCDJ8tGFtBBpbeAvqYtDyixGn/G6scDkbCqJhjhPAitKCee9UJ3nxfRGZPVjw0r8tqj1zX
5JG4BFH8b06+jEf4TYzKnla1Nd2KgIog1XgNaPmxuwzoscij7t7kY2QSE+5ADFYnxrCh0unukLzA
vqjiOFsQmSWbnDI5Im4RMYervCX5Ob+MoLQZkyIqWfnmYyuvksJwpeYfNSXK0FYbFIXAN95OVpGJ
kiT7q0UPLO+AN1vhq4YZe/AM5qBpUQXsxhkt7j/LxSH64LfcdEX0hMG3jSl7a3kYO7J6yNjKnF+m
QWnbNquUNSmHAqYXDydnf7b7oF4AyTM+wy7YZA0plZ8ORFo+/8mZVtx9GBtg0jcV8YDg9ggxHJCr
+jJegE6Gcvo4hNZuv7F/1lIsiwtgYrhLJFPSyyHrcoBVsyIv4N2KNPuB44nRY8pNRzJdNfsrSuxE
ZLHbseskoENai5Eld4OQ8elD45nAylHAO1Vj/FVLOTMq0BUAnxYSrcxYv3gZXXxVE0NwOWj+FMZ9
6cIf0E5J6tgEmZ+nEyv7JmM/lphY+VShoeLUojcrbphM7PsscCnkDmSHMAIRUCaxRtKupvFNDAOD
ddPTUBSVKOGtelNjdY+EXvbiXdPCuNZsyDbCUnKjZQB7nBV3EOiim2SIak7adzqVBBgyg5rpFy5N
4eREi6PUl+fQ7V6ZMgitBdFxs3PHV6E/FP/4iCexvIYdG8MjpCAdWCoJWPxyKYQoRhuLU18dyiGI
ZE6rnl5ki74rYBr3hwHj9skoT9o9XHNV3yQIGw6eZrn15l2ZhNbRvpptF77vs+7Rta4f1bXsN6w9
5dEZGlV4WA6Vd0QnVkaGXntoQOV3c+BVm6W1Vc8x+gc9EzwUZ2JJkVyHRCp3Fx2siSlqTrRcbHWa
S5vqd9/2DwSTs6yod2aW0lRKnM4N9Py2kPdRWLx9kRQS7GidqbOZzJTAhoHeh2TPmdZbVQV/ID4N
z0+m8c2sB1zmRsblipPNeQIgOz9KFr2KD5OZvE5PrF3uaQfe4E/KwdbD01sToDjnZt6kc2MwHo1Q
8Ux8OeWRUWX+xKKiXWDiPvCZkWI7GsKLEV568wwReVqOuUEfY6UMMh7SR/i95BVkbwqK5gAtKraM
K0h2Xs4QyO4YO95f9hX1U6vzreAkN+r+ssJNMIyIufNMoZLOU9MpLs6CYCiGz3MwVZctLnm/5L85
6WbiWOgqWa9EbhXZapV57qUeGaTS4ORyFytDrgXov+Kjc1eAGegX0W2pQ+oULCZ0aLSXPygf6WkU
hYcxjQzD1uGJpZZ4ndP+RKC0MOYrq753h+Oq6yNQOb5oM8mK68fxM+7ekOB2X+K9OXwKFwhwBSgy
Ib12cYAtUPcxtLO8eKp9LW8sPJeUstXY2sy9ZWRkh59Hj3m9Ul7FC4Jf/Qa/EG8HKHfpF4j603mu
XedcWyMVrX49cymea6R//wpFOWz7z5uoP5R+pAp7RcLrVIroAselsSDAWhbwphcKGl/HQK/b0tVL
rtHQ6IxQbl/P6Gg+oJ0c1VjmV+2qwLMNb7V2USOIHO8IpACrD+B/sB0c2PMuZQ1T5zc35JlCRGxp
MNl+FsCo+9hIQUZrgKGeZKyhS6uw/Q4GpjYv/LbqXbmOBcnP3I2dDJHn5TEgIsjsy8DoxcGs1adx
eeRtNFQgK/xZuuxglOAEx2U/7EyqZc55jF7laKqsN6dpNDS8DfXagjeKL7X2l1kxC1wdy44Ch+eS
D+mzYFvZIEg4GP604fIhIKKh8uVmdURrOqdcnk7rfcPEScC3L+bzTltlaCWz8eT8ro06VgA3AFrT
Fs2cAsGXcyVmmLHY1rGpwLDHNFe+ogd1LBXFyFr0nCTymYqlkR+lEIWxdGp9usD+LBT4qC4vNIKP
J4ixwVFPijRDtF3GqrHK7AlIfsHviOg2UCwhECMR2CEXqq4fOrO43Mefen4a4CsZ12hTHOtO6dyO
64WBq7iZZg4gVkxw2XyiSIDeNlVqF0VZagxb4hhHwXXJSQpPGVbjgc0TcNdb0reNXO57yJlCKiMh
gf1FHYtZd9JiMoqE18HMTptfUDsF4B/NZhWenDwy/nmq2JNUtx8RZCG8GIpgPTtzwKL+NyVxQ5Na
yoM6J/KzHIjrscZWJccD+NV+KAbOw/fJB6R0WHe0gKHc8tVe5HxIJncI74ZIBXXsz2TxOhFvjv/B
956bgbHYCG2MAktlWYL5JS+y6atBp4aWI05wQK1N1ENmfdAbg+l4CQvjtXHsOnkFS9qlGMK82qxf
2TJNFuRc8W3Ch98O/aJc3Fdchn/FTFSqcFNtOJVt3NPjeIwYOl2loTh+jQvMKppMU8FIql5CnBSt
iT1qOaAjnQctcYEiFDV66/+Q5Q7iDBU7VHaxhODOZOOJKhVw1tJksK3yBFMaJqypbYvIAxI15al+
r5sgEkZYwZDsLi617fV45RfjqlOevz49oZBdPinNayrnMJWEXCgxNMmuE8CyjAuqjqq2pahVKTIM
wgSAZOhNGGHdn3vKF3wT5hkuZSDfX/MEcSwXYQIcCbpLZ5Oe1Zs3WD0lcycg1dmDC7EizpxI5RpN
HNm/za/kzkKvnD7C/ci7L+GNL8ulBST6bgvNoe/fEfkqza0AqWAb6if8/LfFkIBPWTiAV0WU8lPG
GcibTizBWx26SJ9geaBAyc/VcANrltFJ29joFEaNkp92QeC1en1u+sMmppMWzHIcxiTPOZTJKNaW
9MSjPNBAhWH5pHBU6UcWzdv1dGvqeMjLxuaT3POuiALMolh3fbvvaRqxBI6QnpJzj8YmkBpjeJZX
68HXp0CF4bytOrTCyvWk/iWzlu2cxYThIW8Vo5ZHPBObBZdAkEkF5Hc3kjByz3PEHtpGD4sl0An2
hDmQfbb3xhknH7TbEHy1PYmztIPhd77vaXKyTgOJiqok36wWU5TDDqB/FiY+uQ8mLCzrIHHOn9m1
plShSGgPQq6la+SBKrzVXMSTheUCxZdKPfj4Jw9R0PzaT9Q/qcHgCukQu7/Zt199OuAGXRLtEIvG
jB1MTHdqjMWN+NlDuFco/Q8LBHChIj94bYABi01YK7dqRF9rW4JpTByYrCSsTKT5BnBj/dweKuQ+
NC4k27uEwowMw0GJUqpAg7QM15XzK/lGOLq3s3WoNvoovXB8vV/aBMu6DsZJluNMbqoAVd2NLwge
dHTMKzIseax1YJzDLGPe7Di1yI6nnZqYZw3WlP6mQNiy+UvJ1TZgItuAoP0kich6OIZgdRS1u9fc
2I4Msr4fHRYM6ATJlGVk6o7okowFQ5EicHZef4mLZu6oH0QpY/384qd3N8ylfQGmg6Ej37Qj+Wzj
jfkAh3j+rhKRWjm0+MaEy+GStR3Gk7KBT53H+OGfWfz4XQBDFy1dXU15kNMNdG5Ztbptp/TGmyrS
7WI7b6/yRsw0PxwibjnGa3Xs1gRG4PoCZOqn1QAolg4HOSzN6q/+dHA2IQb+pCEl6SIqa5NNS+Cf
CTPY4+pZwrdIByRqkdx35p/+ISRFBknxZYdEEqI1l63CV4VYxLeNtw3yYazMXdKuMJpEpCwJ7gpV
somNl8d/RgnvP+bdRJVmXR7+e+ajy4LFVJFEsP8ZTLkwFE357yP0Fsb4aSub9c90aopcqVq/P8kK
criygMaVca2fofdGaFYrdAMlqUEfZzDQydj26ctWLEgSSuKr9QMrZOE+14MvusjrIUVh0HH909fH
EV9qFF935rECGEKabg/UATsCDg9N1u+v2g6PAauSul7IN0EEkKrRe2Y2k6EqJJ74rL7q4og2yQG5
ZTpvSFJ3DZuF3eJffXqSLfDh0jGyjhAE0mIOi4II0JoSzZyXY6JQmKfPly6biKAp0FMIBaYsS6fl
LWmYgL0hnsehL8hJlcAmjBm+x12wgySBfVD5zwZa1/kAWDcElpqQD4AHwVFvf1zo/j7V/Vehr7hD
zDXz5E8H7PWHSLTqhHvLr/Adi7nZVrieMePX741QhJbeCChndUo2Bc1+wTtDcvNbpQXbDAZycye7
z57+D9p1gYFwLN8DMb40iEYa0gvtZ5t5zTqPAgxVpVD8+DhYv4xrQfKj9o39FZMfVRKMHq0dwSGO
YuyGmjTanDvlHL3fvb8wWvT6gNUKUOGqryiOt2HauFhcFGpaaOgi4E9SzsSw+JHvsigbfJcE0xdJ
5cV3xyR4hSCphznCr8G28TxroSLw3JaA08bQ1V7agF3jHQk2RWHA0XT/2pEyGfU5s02pllxncqym
whu1EjdFcPs44LihPoI7cgYKS1SrUCrj6769gDejftLixFI5tDAYWiMbegFRQd/dHHJH+AQ27gvV
DS+S8n6tzQatNyF4skfJtSwqKVRGqyM0NewSVmtGTnJ030En64PHkGlWaf8LDteqvEpMQVLvuVVl
t9JqlmEoZDf8wIFfY+24/CIX2D3kW8328H9O5dmNccXU1FcE7gJ5PN5WmYMQpowpzJoDPfCQJEDH
VNuTq0uAgCmN6eoJAbVSXfaH3OF8m7EnDfCyFWOfRqJ80yNARDGl+mXGMAOSjBvlDjquKLfXnjY7
dnAjOoDDEsXIysVXh1jOTUGLbWZTqaOE7jO6nfQ0tRnw6EjyYIScarazXQBLiKyfa+aKTEA/eTcO
H13gF2zonvUDnwy/f5BdNbzjiSPdOHDh5mka4UuhJF+OsSkhLYdrr9nGmBSkPzE962hwjgJ0J+TK
tDPkIV3BQcPqoBtUvoctoi6Sk9Eq9JtwTgFOQksPnaiay9NM7DX9j8yaSIapz16Ka+fvOp6RyvXe
BoB/jBu5xQoG/cin5dyS3tRt+DibsG+sC6zq4ztOMPQ5qu7kTc1h56gD7tt1zkMf6bUxv3tLCgv7
JHC0QBAFhIhUFtQ/JDphSalovN/sfFCHv1G+XAhAIlh+rYFEjW83+ZON1igZheV3S4/5n/SmGJI9
v0HHalITBG5QbjtgHyugOkmQNRi8BJ1/0dZu1zJklngiPFiyZCqUUbZY7zHURTqWagK2tKqrkepR
0GXeJQktCvRurfWI/4Fy9OUX+zSntfgrY7wbH1CTNbuIcGFzMALEiZj+Mh9HAkrQzJe3XNxDQjOU
2oxDDasbMSiIy0RGMYqzRoabU/irO3rNbXkR4WqYprkmG6jcvt6k8yPv57yb+SRx8Djkq0MH66B5
E4L3Qxp7l1xFjR6xRSd93MmYt/VW4lCRjhnTnv7UrwPsVePxwNyuOCm9aFaiA9yAAn6XmvhEHFbT
7HmSGOKw+tVFZhqQpCVNE+WpLsP7gq5DMfArXcx9YUM7RdnN/s8MrTebDu1RqZZ7NS1mXFXnDLVi
d1TBNpX0A0EzUAwOSopdooOrh1YOMING82UDjVRh4/7/hpZvAWkJfkigfj9vhxFdUkBtyQLY2Fm3
32F2XaYdu/uSI2GyzbLVi42i+L0TXvl9Iyt8bJGwCWDkXAcNHdf57jiNBWeQWGMOC5jpNwU+Ruid
bp0a1HqqZA2UjZ7S7LVHgPiytI+XsyqFrUnO/a4EmtVbGxtHGvFO8kAVw445qntbExm1s0Ak4ncP
xDPlUVXiAS8uzhp9Sqk/JliBxgG+ZFC+MiL+eUpG2PKiy96YuwkPOFEbhe3b0fkawJGkKRAudJF5
FPfwRuTWnaxbjpjf6KEszM9nzx35jgnU+XZOSPdG3ncysYcID6nHTXnhoN0VlKp2x+eEQUmilMZ7
/Ji1trKVE64wWuQ9XfcOJ12eRcvwn3azHrw9yf4kdIX9aHzQvJ8O5Ar5LGLrazu4rSD3BxYK7pyL
5hE8VcK3UsCB+76kWOr50zVfy4Jx2oKOwtl0iZ6cijzdWkQnlYyR+FnFDLL4XZDqySSrwvEGzmhQ
7WmkaSx7Nh1qxSf0L7x7Z3wx0ExHGjGmulNKDcvpsPYWe6irkg/NmSH9kcc/4voRMpgJPvn3HPcB
24SbLFK7VG8VI1fEMLLExKGS1U8J3j8+ZiF8js2+/DaPx8MauYoYtOHTqd9Dj2tYBtS9cReo2/An
4hlv98UysjCvmJ93h+DntgbIPqU1WzHVs3G0nOK95B32yFVMv/P2NUuycnET5ithnXFvcDZOAdEe
jRASnKDS7OQZrbDAz6zB6Qv4YoRMUTx5NlBqyhMu0WgMDUIn8mhhqSibvzyqh7X7EA66e8qvdpRI
K5WlAWml81dc/021C/KIgPphLbWblWVBiBQGT68E+RfnqV0Q5lUW7wWhafOHwqZEpli/4htikMrf
e5vef98+nu1Mb8cV1Ry5KvJ73dW++yAxNyYO9WWER2E42hL6gmKoUB+jUrd75W3EwN2KGt6oxJMc
OcmPjKz8c8bNMJvVN4fJrYgcwty+JgXDxmomZPkIlikWk+LBWhSkb9QHvTX/lWEl1DU7ZRUMt9gV
gg+oUEMh3yKmUTJef1v2Mmg7SLbcnJgzD8pBN6KJClwwOwqYDa1F2aTWb9YsryZU+CWCxmCBmAbU
cc2XRiXEucvpOw3QMlHVMAyTg0XDjWDEF3jG9tZquazXsvidsCSNbsXq+N9cRj0kaVCbeNsDPDmG
4rpwKMbFp2XF8d3kC7uF0uRx0QJ9Yy0aK0mKqm4vlny7LltYzxKU9GbmOiKXPlV0dx2Asz12kqgT
8IsxFEObhVGfnCOmcgPZ4fp5SdgjV82oOG6ZfCgL+E1wvWZV4Q7drtAg2vz12gc7KtY1l2EuUHY3
ukTgVlWDn7prXwXkF50TvK4c/D6ad1nk/RlUfF/yBtZm74MB1G4sK20givY74LnI/pohyWFdcFVC
YwIa4s2Ubdyg44SyMn1nwgzuo0NfOlhNkGcuYR8ajRGknyPLUhVT49WxaxdGt342qUXmARk1ebWc
E2SBF6BH5vR+KfcnE5sRqRwlNSR0LsT7Zek/py5mpOMPvXCyLLlMXuFFbj4lX9UBKXXhLj0HDe0o
YLu9W7OOdk7nELkfBuhsVqgGGRR7BGnPHLBDknY4HgsEX6cDGuyoWgHpeWbVk48kFIORPApofrMc
a5DS0N/vD1g/31uQV1tmUgJtFU7DIJxxAFji2iXVjA/KlEUqh2u5cqp1q/tcv683pLolRkkicptf
uuXNoTQhGiRojZXSsfjjuklibTSJK+l2mfkIc6Th2RBCGzXMp9hlnIkOS8jaHYlZ7faJIqY7sDM8
sMVcWpJhitFyKHnKlLjmVqgw8u8KznacON/tSqOizaYk+SozvGhHvcxwagxifU5SAhJUxadt5Uw2
IVSpFs+R+OwWNzqyqhHqr0FIZH0qvDaW4TXLtqGqefMXC2XuIbH6Oa+ekylHvFRLZ/J2uJ54gmjV
L9uKgtSYbnK8rYWtG0a6QKehLHEnTN8YScdI+R2FWyxa1aX0hQrI3c0X/4rAVETD9HmpidQeyJe2
jWbuHoaLBDeVCpHDZmtEPHkv0bL4ERnBOzWrHoasIhEd22rQkqEgKqGSTQBHHgDe1pi64wG0oF7p
Ol5ZTIcdzB/j2CCy8S7Yqg6divzXkPxr9AStTbxejUn4Ngyw4Xn0gVJt8Viqd4B+hvKMJgIBQVhV
uHlNzrL3Dq8Gtzt3BOTLZMPLpZsH+SG6rtFLZ0Y2yPTvGLjm4qQPzcC/h6qYU3uWazhm6rUA8D3P
TxL0hbT1Ek30xLjaM60r1n72WjvQI7Ar71M2B75rbSnuCYDCA2eq6vJMbdt9yeBFMbxsTtRM3MC1
PpluhSUrIUpibS6TS5ubLVzMKB09FV0+/u15csT1dVzlr7MdD18IlfvmYEuOSjaX/tX0GFhGyGc8
BAwI9yuxBaDJffoHTU/ZcVc1tCifBKrQ+cnH8SOBSRbpT1thYsv8bwtxB2vyWRxK+SuxYIB1rrFV
TBMBj309qKcdpiuCTFRylVgXAbG/gf/I9EfFxlo5nKMQ6KxhJRQFNRCAIXvgfzTK493LjW1Qx3se
fvDWy5mrcuuKvTrLAA+YuX1jE0SSMElFT6WiUffo2Zk/Dv/cut3FsGAWDC/sO9ZQo2D7xN6jPYTs
ClkX8GllVYBpgxT+2v1YpaZyUTg7oLDXTyDNTjRjGkRkB1uSm9xVcQWMMTMnbBdFizqqD+uGKE14
kLx0EiQvlpedXFr8c8pCN6mkvCXZbg1uoXfY5/7vBWq4qAsYP30IBSjvFDczzxG7LUAfzIzGKAEM
ei4LHn8M7i8Y9kUVm39grBVyNWIrl5jxv5gm2QxAkDyCgBWPwFurXvuBTF5QAJXfmqtvISuCUdAk
zfOxgkJTEaskbaPUxRthQKhJKbUVssqCTetTgUL0cymz687eUbjbBe7lf/GE66Q1F+bNs5vA31gf
YTnR6zH3+CiKcjrio6nFtTsQufYP7Yl9Eraixp7mrnx29MDUyZZ1tVKPrRdRsev+IC904VKbFwYa
VvZMSXDrQajnWF0f46ta9HZMoATP243vsqDm/fCj8QLsAv/HMNV9r8R3ULAapnAjIBmRQaBJn2Nh
FCnSuFXm4s6YHAj52JtIiV2w7M0PA5JJr4YjFaisCG4jdP9sSGVuMxk6JV4OQZM1WcGauJsW9JQP
zLQKBr02sCbc3+vU5qBO2LnuyJCtf/4uPP/2RSFowHX/PHdIQnPaJ9uEgXwgEk9XULjEHgcHreuA
P535daz7xMybe6pbJfgsH1tJgU611hGdoALrwOw8EskoineaHIUzCpO/QWvKHzez1B3EmEKBqv+O
TqOYJNXHf6/ZaXBYMqCMNpGusO19CIjB66/vMG8SPM2VQz4Pf8hg/INKy5gqLoGGk10rJUimPQZ1
q//0geTve7E39avLs2QMMtDlIHcJYIf6Xg0klsuyl8oMEEI+GEzodDbfw7cGIGEAqhWrBkr5t8iS
tIuEWY5ccIjpIhtH0nD8TUISWqAxNa8tOxAiTz1kx8wz8xFe36yBC90ewxbsYFebAycw++hAJRzi
L5rpumWqLLYdzLIWEZxGFZZE3+PoADFxu+LLFSV+bVWEyH9ZU6f1iCtY4RSXuAF7E62bPKhTlab4
j6HMx7nSgIoFuNbxoYMRh4GDAsawXc/fn3U3HrD8L4zdKw6Np4yEW7LQLy9Olz4llPmFAYH1C8Mm
+9DTnvKPgZqASuDjHoWw+j3jyAtw0+SzlApRDrpmV+89sbqK1PqKC0W60H0XSVH2bAw1f0zovZPi
JoItZd0JY8shVC1gGilD6yTbey544CGg/cDJBY8JniUEbJ7g95u23+sX8OCbpATr7bGVS43Ph0ql
axqHsgkOHIqpX0jgDiLJz4q4qngZGl25PL18GKcp4Y73NXmJwTZG+3Gp/E8L+/C7hbxZROxTV3oD
4RsL5AhzTS609O0BLKYj43KrfhcUHFIdu2OUHnVfyCwL1RUS0IXXwT3bmt14tpYA/PXMa1Xfjub7
FPpICWQ1uCuDNxhWkHejA8I0sdwMc0yqYQX8xe8hfPd57bxpJlTf5Q5Z0P4bt7NJBLGaIf25v6uH
RW/q9B5phERp51XRl8RhMl5qinh4U/6PohabwGoH3el684bTX32BuLWslVMbXPDHTtu8rK9aEP8r
Z7zhoSf7UKbvqWXxYn7/7LEo3H8FZAso9KmbOzzs4nHiHosv24IPCGqzI4I22S6nU1j6Jlfb4Nk+
c29k2yPzUYs2T1c9vEQoolgmp7xZeCyBgpGZbO41uaIT5L3KFxRIx3ON+2mmNBvuuE85w0B0byX2
2XV2K2IvKAII/IcPDUpgNnaodE3fkwTQD6c24K6qMhVbRRfqraicJLTAKgLgZETaNeON7b/T4N0O
v0DL5pusMdOr75nMTT+oEWN/ixbsusO+Jav56Ddv7saghQEV6yy1Jmm6zvDdyWRppOxTjXhfR6ds
Y8qJtErU6Oh3YbbXzJ7gFSfybqv+5Do0rYheba9PFHDNhBv6i639OUA/kaD3h6jeNoBFXTrDZ8mt
WqHHdth6jLQNqmEV4BCA86aUio3pU/Kw/k98+YOufAUi+neIqpOctKcAtUGIeJwt/kx+RsPHu0dS
J9A5diRCfWGLUu5ulYFqX7KDvR+c/Fd/9W6wX/gUKccg/tEqor6HYM98Ol3Gtqu57/OPHPYjsUVt
4S0BEoPkkBoHNrikeiCXeG7lSnUSTEAD2u5sBK25K1r6AXA6yY/g/YFlLEudmd6cQiOIUJ08Lxa/
LiODdY+fVv9fQkByR77PjcupRwAWgn5eJL8WU7fTA/NvR8XrZbhdfXwDodlGM9yiYbi2sZu1M8/k
MPwLoG0yKwLc5ZeYtxu+gvQa4P5LZgAZLF82XPqIQ0CcQcvztmiNgCOiHl5OeCDJp1+9dEgi5lKn
0UWKeyFoPN/WDoUH3OGvw3MOdxEar/T6B7m3Sb5hUUfZIq+c5lKLdU6RbzpLCH3mmiWKVP/DM7M6
5OTGQMyruMArlH2uQKAJD+rYsPYABOz10NYRpdMQ2MITCYpW2PpkKRfVo2qiytXBDiRod52FK8VT
h6gvyv8RtlIpgSllqH8zfrwSW3kVTShaqM6Z07R1S4Wb8gKbXNic4kQ6dA3U2P41H8T3kc5iJYqJ
VLU+2BwYE8IY1OQ6OmsUgTCw5oMgIdLA5zyywxmHSiEG7dNRjxfd6S6jATGffQhnsrEMNjX6k4lq
7KjRdMTeQhxlfSmWqaoUvA73AUx2ea5WyVThqfLG/QDR+pzlVfl7Y5oPoREEHSKEWb2ISOsAHgo2
U3fPtALe1k7Gje75U+eFK0POMEPvLh3bo6A0ZD6DsAiiLnLB98unhQhkzH/88C9l0dqdLFMyj0HF
J50RpGDlRikXNRye/8DrHSRaYh2JMzXfNmzg2Oa1GaBm6fREBPwVlFXFa6jXR9gH/j2ZA3s5DhSd
hZ8xYl6lXot7T9cGDSsqfLHrCgMZKeMtU/MsL+uJfrTuzLz+j56l1vKlAz9mycmucKEv7vyLIYIT
DUiSqCDLiDGf9DQFm0WUAy77vKGhJWLGYKxzvreYCkvjwtaTJSf0kAZKywvbx2ebuzgQbVemX9sX
lWBULStX35KDd6TSyBmLgetNpTv1vx4kqw91+aTF0eQ6Zv1GhJScWiMCDp+N57DUNUgwQpPP0f+s
hYXIknyONJZHpq7L+FGaM1xAXNeIV8T83vucXWuPsAql02XR1+bMeXZeBWc8gPQbZwkS6RHIUfX5
0FgKLTO+PK9PPzChfOUjtsvfvEsfhZCKL/AqqUPsHfawRd5bBAOK2KyqHxqEnZ+HY/O1MN32rlsu
g4Ji96XEsqOO/O4t71K6t4uX/k0fJ6hg8LYfAontdsKigHpZKlE6liFWBCBSDqoaY6fEaR75mjGh
NehibaG7Uq1xWN2X/Ru5MIm41ynPFc8+9N3A8QHGOy2bwjcJCnlrE5MihVrX3BXeGopqKJomNFl3
w4mm8Iymijz3F4qEX5xiz7YYtJvJPBMoXk1oeyGha0buDHoc0QBNDUAUGwvj9tT74rZ1bzTvlAIO
/KFtue08XwS0CHrc9dvA9ii/6MDkih9yTcGZM9wlKrT5fefdxnCzgnjtk27Gfr1iWi7XHIbjRCF1
6W/p546knre2TFIU3bV4bV+NjoeD0oL4L6s3jhpLB4DeNqq66GLGb1yw7qEfYYi8XTVhCIuvv6X4
/PbUTma7Zq3S5R49zP6TIggFcj5p10isFypAQ6VY2xn32QerbSoDztZxa9mCn91WKf/54vc1UdrE
oJE+wNu1wql8Z7gGQPqoLpAN3xsBOFZlzuF6fd/8cIELFJDsD5LWV/mrUlLWyU3u4GHxrvBZzbQi
L4d5PUv+flVc75rHAYlk6kIgYywcyyTKSkeBv/8CGfEI/mxeHhSmJEHelqWmtYgxslo9WHHMHz1U
2ndL3sb8pV7s4kXfde1Z3y5oE9ARjQ18XjRfEGvjoRgkKMcs4Jq0YbqQPmiwqjalse4oqsUr1NDE
gUMugg7PoE48XELLw4+BTjAmy+ErTVjam0C4yA42TguXy08ky0ThgCJJSnY9kpKDk7C0+q53qRiW
Ms/uiPCQmncGkJ3ZOpl96OSY44uAq6EMOVc3ubec1vWBeYdiU3gXvWbA1zvRNHioejlmElwJsqRX
czLDGYl3PMAHRJbDmKRncBuUxhMbrjilGRCwCnuHpzwvoFOmTZyPLncbyrHstB/bVQXDY6VLDQd2
cbAZpaEoRAaguxmp1U1BmKh/ArXDL2J5+DmHpk/G51Q+cvPCquewyQj6Sg3gjvLvOFP6wAVCEWhM
vQX9H7q/5UPW5kn+mVmNZurlrgy19XGCV+ZjIycEVw+fKgrZVDz1lS6vhDaBJhNKZBGsXHKfG1oQ
TVoxDrFBXS/iQSBEizfoTZgCX0rpeMhhk2aYjIgEBNv1rAqgqHer+IHjVxGlXleFyx1RlZpm71gH
nJigeke2xfjf59UEAa63oqqvm/L48g09dX5yyaKAa1LUS9KzYZfQieStS1Qiz0014KpjTZ8FL2WK
0fpoSIK8KrjLGmy3WAvanmdUuqn+MJBX+BMWwzMytsU/9yUQQQ1nlt6/y557PKR5gm5aBmXV6+gA
ZL8+6cmYo649aTxhF0q2O5WlMRFWU+Zo1kpTrNVQ8JMDLy/jeGr7XQX/BtPr+5ehr8gH1syY2XU3
wtKBwH1p31TPo+dhswcBqgc3CXRqkIEfPGPAWJQQh2s6/Bxwb8K6c/L0zUXxYJECKm4Eh/UnyiG9
SbDBdYVqrPk695A8TMPReokqHUVYFsJ/JFH2HOSExVa+ZdgxYfV6+iMZxK/cqhyz/GgchekY2HL9
Cy2Bk4cZogGdz8T7XRy1DDlofRvsnsG+fpEAh4I5KwzjXJmRYpXNGRbCryvt0LUh1EzghV+xCm9X
HzAXr1GlDwFRQY1zQ/LNt29gQxKxqxS0v1MEoM9Qg6DqzGQ/udcsmnb3lWBaK3LdWc+M8OIOeZQJ
6Mqx9G88IAOUoFQiUARnQcFv9vmPBIcbNr/GyB8CXgFdevCrbe2mGE58sQ4yQ0EWyLYa/HsMGr44
P97Tb0dTJdbrG+6om9ityWxVzgkZb+Ba4aCj5SoyTnnUOJj+pd2LrjthEERMHAdWe8WAmF+2xwC+
QkqnVS+8ZI5lLLCdL9y673EoqXLdxVuoQC+i14Gqb6j3Kg7XC+kDZoxWN+gamYR080onpYdkkqWp
nm/ctoZKulmGRHyXZWJe3ApLBPvCSCfzPCeb5aIcXQWjr+wrQVkj5eJbLeD1P7f6grktRLLzADAF
WbBPyRXQl9wvMJTwDxWcnXAUJ+hFFjvbMfhclhrsSYkQLVueVGp63c8isz7VavDcmkLziEGHaN0H
7CC4z5U3bG0aAl9OOS7j5gP1IpXFwZsKTKjuUYonwE7RDv9vD1CtMjjiFoMR22OOJN1k0+Jf7vbN
olReEY2SGfIpGhBaVLkB1mEV7YwHlssAhARGECc5jQdBb6Gn9iQK7h6cp54Oh06wtTzOszLnesfo
sP0/Ag43vQcST/yuNHM6Mtj5XmLum/628unL4OTJr8OwV+BAEDDbTiSAeVzJ1bdNvUmr+keKEKmL
K4TnPVX1evvDEg+VIRN4iOu4yPcJQAMLJo4QotxHIUsoN86hW2dEHd4pzouYN0bvVaBmTJOM38gT
RwKlI1FgOsSbVoWC4lwTK8fOlDyWAy3kmFoQK5X1Je5KqBH94W6UyGkkeWFIrB1XOQY3Uhc76Nzk
6LKLQ7kptLEnxBc8v0/Yzs5WVL+FTbMhjlsBpSnLUHRf1nZGvZ9lRsRUyQUSMSlC4xlbZMXjkzz6
OzBkHI5dCRPGDhjQQaiki4B7xALxgHVTNl+0q7NfgeLoqnF0stn/LacJv9/U6CSvoa32wR97dlql
14wfTlYBnJBTVrlPPFWI2ZU3upxF0xbj7BFm3aJ114/Py0P4JaSICw+YFLsJldCApZLCAcRdWDIp
Ki7uEH8XDjXJjjSs3egvzeDuJKXso3XcXzClmfCSyaYTbambS25ZYJXPJZL+PQBKSysMPAIzfaXX
wxsuI0HNkLEsKtM6FMIxj/3PtpklAIrQfvyIaY7oO46duaGX+ZKzzThYLqKeDcSGsnSvykAR17uM
yzIC4+fTaMrYizN6LSrA4aB2zzrv9NeMgGY7I58rEmCnykZpkFmf4ifqyG5TACjXjTJHQMcP3+7J
CMU6mlZZFQmYiknOqPE4BfxmEGP+s35ErJaxGfHGqoTeR5SEvPiOkW30xa6VAKAXXEFkPTZ0dkmE
ba1rH8pWdnT+Yjs99+xZSJqD766sZG6I3UOJzhfxsiw+vSwC3+ND2tvjak78h2mk1bHdvS4qXmsS
t+mxGo5Bfjg5MLFGYwjqLmbTIxB/XtwxikAPrmsuUZw4RwFQKycWCKulMAj1Lgt7vat+IyAhEbWx
nbCnhLf6ZdnA8eo5+kzs7pFaxBnKVJ7/JfqrGWZsvawFVHfgzzFC0dUh8IoIdxbivrALY6iNGwUV
v0mFBdQpIgq4Z4Geo8Prba5SlddbxJUl4h3jcRMXLGfVcS6RgxoUjDt4viPTkm7b7h1Xw1lbIRJY
ZjEc/UtRwi3hqhJUpSPBlZ4HFsvwjqGVhIEtvZYj/4HAmp0t6mApG7VhK98mt+q+7dlN05/cdBj9
KRE3nRqIPQ5mORbVNMjRJe2hscGCXUDHKG5NNPRj5dP0irZXFaXX8c7Vnl2iXA1sXLSG0KFvpOUb
jSlTMc5xFFa4SXqPG6QStPlokCylpHaJAD/14I7IAiRXYDIqu+H4dcaJsg+gyZWLexYwPXOexLNL
NM4pyBqAndBhVf/2Sklt7mxrLRUXhhH/lBwf0bDTGVVBRMNL3W2q+myzzmRdO9nG6Kp0+79apSWo
0cfxQO9PIzqVdZVi7YHabl++ttiD+SXVtsK5zwovzu5lfiVCR9b5dv8PnFOZ91mgXMCLzBCwCieO
Gg1AqfDwkZ5Ru0W8H3XBAHV/E7E+CNYC1CUbkDFYRefVRSCqxJ63WnEqq+5uThCR7RacFmFCmyCw
aQZFPQdFkWVhQkMIRRvzr0kXHYpEAFF3EphbT40GhakB7b/z/MDB8FLZl4aWTO4nyn1mE1Ybfx9E
HBv6PEGgMZcsWkGOSvETpJh3LZfaTqNM+27VuGPx9Bjs/fPrCsJOtCsGwLaBD+zS6x7y4nCme0Jo
RhE2iQxHGF/a57mKfcY6reoqZi/U7LiM4mnCSKLjLnfy8X+cT2c2QFh+icfv9gprp86S+lfm95cl
9WPSbJIMq1jC6xkgAHJudpppRviLy9+uHRZPRRz1s/0Ph9zY638NPvwKuxy+0wclzAZA1O0fdhzT
Cj7EzWh6fjkxZ+8cYaLrl292Bg9h7YvVgbTG/rHI6jd2VNNhbHVNc4vAvHv4TUJ8QpbewqkgCGgv
RunlcPSOS8QdCAymt3fT7CIB3fTJQDc9x0qOcFqgyAUNi4ce0QTIZqnFEv0K33sdPb4+vgxKyrfR
jO1kqXYgUM0gJvZjzRIzS0KLlb9BBIlvE0fM0rarbJTEF5qf82ab6c9g4t8Pc+1Y0cAXwdOT6WZg
FaBr52Q0LWdLJvi2w1xlwmgYA3ITpTi7ujQ8FK9xk0dZ4r9tOhlLLTuQFy26wjlfoUlYqxUTl3cO
l0aTebXH60xwTbfOvR0J/kdSMQ8Z29u9NMxSDr2+u3USj2ros+lz0rmvDk38v0AWgefWMP9py4Ig
K9PdR9zVFXuCgwTFtXMmuft3M6coiUIqsrRSHZRWxIGbQieGLFFKOigilg7G6Nn9uAilrNwabZ6M
VlR0fVq6FqyeMn1lPXEzcbTuwPb/Eyport78z/Xiu8pm10iqei1Z7Qob/c8fZTt/b74a8eNtulB5
HpBKIkNjVixC4q6pBOIRQgCmPqUFh28vjy5ftGYhAwB0slrX+GBOh0jhGUugk39eHI97GOyUMJP3
Fd7oDjh25N4CwM4lQHZwHzwnfoe8nHTrM08kQvYbLU6P61YzylltlNm3353lP91Ty61crFCsGdiW
UkFLqT2FeAhr/sb3kti6toWSf0VhR1EePJ6axLiBP550oo69JTIdv597UK4zrgWGutox69CUnVZm
e8sNmWtNjYm6/YsT3YyRWEwdD2C2FF55Tu5Lct/z3j7Utk2GU/p0wMR71jczZzESTZP2jIUYza7F
I4XFojp+phWu01bCbyfoX6Dk4+TXvsx42MUtaIeSbSbt2ZxQMooBn+dvRKlAqXQrWm5n4YP+BLTG
Hp5XpPUX73YtGvNjis++DMgnmNqFFbxY6Mz2VqS3FrTbHXvFLA1eXXA9xo0Olq1BQIDrgireQ3GT
Pwpwb+4zhFHGqBMDuAvrHmtau2ACLX4nxDRkPwUn43I/j7Cn6JD+keh2p4STzPsgpeOc81JRswiu
Gb0ELSOjN+TKSEkmQhv2Hiu6x7qf2dPO+CXQiGvNdijJJNF39nK//vbSo9pKB23QShMzX6bMsnUP
VZJW91VFEDu3BKhOwA1NRE8EmjDIvgbH4idDbNWjP6zdK6odtKwJUqNO8Sz1lF03HLMn5UUk6yqa
pNHu5IoJxF5V8lf3qfMvg/rTcAGgFqCZJpoXMFKoDjK5cfSPWhjV3z7sR/gdGS7Z5OJ58gOi6ca8
Kv+av7szC/k0fSmhegZUGRdQD2LSabIgiFYA8C/vB1yogtOBbwXhDUHbfslHHRzT9jweijNrHN6y
8ceqE4NWusMhU/qt4Cj2GfrV+noAk2hQ6hlsMJN+oC9XY+D8K24ZWJ4C1lpkRUoFOzwK9Bn4Dtwu
okg78RXuco0qY6f0ntwzWn3h+YRm/0zhiPBrxhJCkbj+3ywwaFm1C4HHDiIy74RTpjj9f+of2pYW
58Gkq/mzomD1nVcX+c6/JU639b8M8uQeU54N/cLKdovcFCCzY02CgcQbx0U2oQ74RTyXOeaV+M5t
VsOsgkeH8K8v8sb+W3cNyjhUHIE2jTIv/b7APZg0rBeG3kI4c1HLhYkFexEcZejJpZYDhwMzHqck
a5RS5ZD8cJmO4F0y+/Cc2+APFyug0F22SZcQP9z8EiqNDLp00IJyvOagMvcWHU2LrvGy77FFxAhN
rdCdVp5lIN47dD/DeVwlP2AajmgNH3etcJl1tIyr4zb2l3FDFI3RuU6Wh+bTX7jzTsdyS3cssJJ1
GGO1vtqjvMJ6+iRCUqQBj+p7vny86Prpn5K71E4uUsZzdmqzw9kz1DGxfVc+7b5esuY+fOURoaeJ
BT2meh9VpWgwIJdo2+vP4uKjjfE3UrvBgV51eCAI0VQFG4ZpwmOU8PDMtnmjyoSycd6Ic2H/NypL
8SQvklAaf3z+/FFQn0b5Vjx6Mc067F4XpCs7C23b85STF3Axv0DmGjSHo/kCOszGhRoQzecGO2EW
94Du89D335w1UkRdDcdHalOosw6a0wJfcue7ZkAKHUdhOJkSisCAE8rA0nJCv1c6qymfihm+QGpS
nKgr8CIDKPVUWMZSdRRmfA1TrDxtU40On+Z2a08lGqHu/2Qx72UL+WcjBlwbNIB8kq2iDV3Ezozq
qAFWRwAxNxMqsO4EcyNrUIk4yiqy0VjPHUPrU5DzGue7JeJubTUKONn5EnaRaULjiaaB/id9IQyb
2mXY97SBWcw4zh/O32we4IiSMZzvI0uHzX7CkmbgzWtpl+S5gkaeC/2D7vg1oMCH4XRkWtEU4qv6
OGZFC/jsQH7tQ6gyBOd8UONhcC5Np4N/tpvshil3iKizhrD8isBdYgtFYjyyH/vanAPMLSzQW8Eb
2aD0sYKevTMggYeEz6h7NEj+lF9zkp+koMbWFVX2XLCfG0k1471sqZtUn6bXAH+19za0J+9DKpPe
4ai9uaz73prfdH4J5hXiItHnJgvDvBuQj6b3AEF1aTs61lXHYZDN4GW+TRS86k3BwNmmn00FFBHH
D+yFYhuqOe87jfeLdaaLtdYsMR/fXT584KxUbQzQwNAM4OUG2b9+Z+Nmj5M3TQiWkspNSIneoy9y
SqGEWbAxzmWKCccKJTp5Ww1zDfDIT8RdAnbr6k2sQQkQkpNzmwnxgHoswKjY2erE9CLHB5yV0rG8
0ALu0H5bvxHRIkGcQMf3IS1W4AJ46G1d45wsn1u3lMscHjR09e/C2+K6pYIHZK8VM6ofr/t4wspx
l0U0NJ6yKU9w0ZK739P9sEPhb9pzVuOr+NKGagQuddx80P3ImrEUfhC3c3XtzWb2VBR+W9MhyaSs
W9tFn5TN5yO8RSRSa3GeWw+ssVzEJR1zIqI65bxiQpk13yyET/YGR0xB13JdH/nEjhTllQfpKlIR
ZQdfWpXK1h2z/7Oh+zddXrN2FewgxeUCdFBslCasitJ691SZdQczQUMb5ZKdY63+z3f+dwK+8kw1
O8fcsFMDmTcQsdxvMOUB9T1yoarefnaTWMki0Wik1GMaEvqjVyXjaFkVybnJPxvxh5gkGH+mBM75
bVGUpA2qse90KGXpIbT/mqz+fJtKxX3s0jPV6ZI2QKrDjKLusvAh8glyMZ/3iNezJSXcSb/9Ig4c
+5fNEnBK75kjtcIZeIwL4YqejJliOjPkbymEyDbqqInasmM6uoNiCdlpemOFY7S7WdINlWV5hx0A
VEWo8acSdpesSrGNlkfkFCISPx9PwtZw3/MhXd8b/4OjlKAUTKW/aY8mesYpRBICU4JHBQo++ffI
tipjy6JR8UHsyJw0xm18/LPoQpS3q4SlKjeXWW4dVTvraMakH+dM1RK0ANXdjY5yBRLn1y+2OhxV
ZxZQxdFvCD/bpKp5DfZfIeO7Klolml9fNmCz4KWt6DRfi6/WfC88D+TexGNP3FDm491LOynEY+aH
nl4ULyKvOicoTF0usN0iFXbAspMju9S3JzpbH+cnIhvhrngdVUMRKD8LC6EXeUIbGPs1AbYg7j0T
We+GSlI8mv0PBuWM5fLNvCSyk0k+JOg5ZIndSLwQrpqsITj1v5f9fyv/YbUsfw+219TQVKeHvsWT
8Qja7YGlmln/PvKHLt0jakjxGbkAmBlrS0Li25d22jzLoGRKT3JnjhcrxavqoHTkPfrMDFDr1cGH
IcHlRZJGrLz5BOekxMyMKCGeJJmfu6+9GvxqiC0KC3+8Ir1EIy5Y0LIYKp91l5staOcsT5aSBI42
oKUXs8uIUAXZB7qypxOF2X0xJ+nr9lrB6xEAkoJZCH3+lPVEt/huYZ6LdY2PqCr6Jj7ZLFuozPLF
hzA07SWaFzLqEB3zMVL4G043y2p0mJcaJKZduRTbOSAp9mB2/A1IwjaZoKXPsIYAJrc4z+VSrPY5
xnPr9O+/4uf2APJQQjv74+LpzdzygEPztiEzBVGNl6AwfBPEXnIo9OOthHAhraSo8VbChlkfnT+z
Md4PT9k61kfXnnYpw+2kEqpbO8ngNIurRdvlaGCuHWtDvBqdNrmP06RgCKIIP11gn4cdSaEMbyuh
4VpswpYYXipPmDLJw70D9EYLEweA5v4bh9LuN56pgpDD8nIdaOQaAPIuX441U0SMY6SNcXdnE2rM
Gud23/i4f/FItUyUCSj9ki1fCzzgRhXEjjx8a7zCicxYXfuKGluJVeyZR3fKYB6XHSpu0d+GrHRf
z81v+LYvoO0D09JTA79mNMDuYIl+pEVF7zq/MBr4AAnyp9nqFYXBMZkgPjebZVJNOmpdDVTcPxyr
35AeUxBdgMs8fiTsKNa4besK+C+nfNfS29RKvzDm6qi/cDxSCXKI0BAvkAXU/27osb4Nv4MOSiRG
rpz6sZqPFTPgQDOvC46lDVQAEXsJDrjmYahKtOrEZl3HS3Wat0ZSBG/DGesT3LLj8iqLMLyTbCkQ
G/ZrJkWFV/pqI9MRukgA0Ex3vzNC6AFKfgcusZu5ozMP7rASdHap/DrpN6JIyetJIZvrQbbWrdpN
vIXmbILIzKxnydSkj+tsvxMgDT/ec9V9DEQ6/lmd7hxTv+7F8wsu2Z8NqPzSyW+m5h4IxzUohox1
/b6d1RjsWSi3DUbT7YLiqYglL9Py136f2hmZja75XRJxzrbHmcyUxqi7qFbJFhInflcThvx0wYmv
Z9gdVVGJyV6/zOcUK5pxwAqOuScD83V7V7FBH3FXmTDYjldRPaOIsygXemZSg3p+AgaXz5JFuWP5
+dZLyShkYsOvp65OZxFqAl3/EVXbnoYVJlC7IhT1F0QPim9TIYvnYFCEmKt0Z8RRmNkTdrujNztO
DmQ4HSNaoT8fSuHTTQcqOqeVbUEP42vYj4kk254DCujLN42rdDOAgfLCYAbZwqpNAKWaZNJtNG61
xZMq2ahRKEmvaosHn4oQ8zndoq7eD0awSWHqL6iq8bIZq85qBU5dxh+DEV24u2SQ0avx88URjup1
6lN0Nq4p55tEnCe3husOI6ASs2RRaQdHZNj0RO2irYsi3e+FYkB7IUbBq06Fd720RTr8ST+gWPhT
4Z0qERjO2oL/XF7vDEeCZvBjopCWxn84Fl5WAPBpjmCTTIFmxC7TtI/RFxX9Had8fBzBSc+jDsEk
oL5796bFOOSJEVxEsg58R2EMyIv9GZvPCCMp5dwDw/hJogGvxsnopxS2VvYHm8LugQDT3oocduvN
YWDWRYqQ2GQWPrlWcUW2pAM5TiJILvAokZwKQQ99o/PDQHArb7xHQWDt139uom0y/eRqZ65mQXtV
TcLyoK3u/rJqgdTIydrqVCjZwn1pPDzH5RFtDHKjulJ0boOlKjHlCwVjwprmEJQ2hLXyBtNrzbfK
eltQpq0rzYYJYihgAlva0Iy0sk91k9N/+4ypQxN1i7Qxcd+YnN6JGCa48OYcEenjhRUNrkidAUTf
aaFwkWnuufW5xIuZlrLmWOx5iG5eA2w+TkWtNwEnQSuGw6IgTWwFNWENeWdHOMIpRiJ9Pm0Z3IT6
9ySqIMecw8U5Ezy7SFsgtEAkiqMLZXcScckGdWHfRKFfwnQAjPdPGEUzXD08oTfXM2UJNRdiHD3x
AAPKCEieZ0NmC9IqtSF0P8xEMXXQWSdJA4qaqTU6aLqPFc4B9++0l0PHUy34FlxQeRjnopU8qD2q
62aDqCSt1wes+ZqvKvaRL4LUFqv0PYLWljzFOb6xk2+hVgTBYpX18bcn8UvQsAmvSPjCeDyA6KQU
iyhi0Z7/mmw1iFER6lzHC1UsxCKpTqOZjwS/5M/CiPUT219l62kCGyn2F/aQ96RD0W/QvJYJYXzl
V/XfvzCNIjxwZDQNJLmOQjqJb/wOtKXihuyhZtA+gJovMlMB7O5wZNeh+j4o9zvVqbtNoJNMm0LF
cW6EUp3KuuSwPQ0QKcjKfm0kiGcD9rV4ix4BPsNwDR7aj5YdqLcbDjSIWULE3zdAMEWEA+vzbZq9
x9lCudi7Xh3fSGmLJZlOG4cP3TH+IUbnbFDojv0Vd/jv5gCUsWhGDVaDL3wE7PjO4ldhTQlJ6hQ/
iSWdupP2ieJ+4Ri3umDAQWR/tRuqtHHgvFapOJ8+Wau8Tq97WopAUcM9g6Qihb+8tmGnc9+Avs7m
XG6q/rEq6vWq9oC6J9qhUQhaXpNXJAgXX4WqTMlTDMkixWah6iTkHIzo3HvuKIISecEfrkLEpytd
tS1GBHxg8wJfFkxoqqngDUAY7MLrqGSMfzSJ24wYm/toxP9ApbUnO9hfacPcDOk0Qj68XYwny1p/
MTDJ/sOBd9u8o2AWCEJwcw9OiOPe34vvsGz/uq9RTY6eNwDxKSTNuwCjj5fAmJ3J62tiKvwUYk1Z
RCZTKz0jsZSUCxeTIAtaGkfEneFz7z/cfUyi4jz6QND8AIri7jlOElp13R+1XA/CDV4gC2XX76Vs
kXwur9TkD8OW/1xEHkmA4WpQtJ1BUIbt0ocA6Ulq73Is08mW6M8FPkmJeWS2a7fKbybfNvip3QD2
WHO90LKCGafr/u1u+XwwFulkiaZLQD0RbIArk2R5gCLsDmytCv+OJzZ6lQ+2VRdNXRCJibwFGXhb
pvWjjgk9APpI0hjsI0iSnJSUiM9rLz3J+4BSJTNb0IEyZ/PHH6HPu9WFwCmjaCQ0tpQeZ7t4tZwX
ANxv6H3SBkabtgYnk4NHFLGrvUW6QhzH59PRK5AYyIS7hKKy1+ZnXeD5scEtoclFW5kSN7BoncMr
KRkz7mtETvxRQSA89Ji8Ycl7kZsp5mDwlTwwGTNkgLBFBd9hB2wYv1MEfReGJe/r6uhMNzNGqucA
u9Ib5zqTdO+23ZB9MpP7pXLY/kh3Ht0ZVpojNR6KSRbNOdzZO81E10Eh5ASsoYebohz6RNjlrzxT
MbrJ2t7cKa3lJvOCUVoHnCTcODovSAvZcFOnbvWpVDMDFtJaxOEJImLoQcNGx1J3Gqg56cCFQGWF
G/Okjpum+o2MaAhhWctH3v1JkMaarKF7f4wDNIIRjvk3XkFQacuyIzlA1Czm6n6RTIhzmUxhGIKn
yLLOrGd0e/bVhwQOuc8QTGIVK6AMUDfCsmIKYfjDwDZgHcdEjPC59Y4PgvFvSqH8mlA7Zzv1rPL3
ZXr02m9FHJSRyyFeWu8STEotDbs+9aiqxz+Sd8ryre2wdWu8VX5fnFESI6bSrMaQNkkwyMx8f4Dm
3MtCNe+RHZ8KoCj1ZPBOKPsZlkLyND/G9DHzfJP7v2xrJd6U5i+O6ay8BqQ5Dj5J9JiGbBGlanon
uWPWp24K1sqjw6GUv5aPltF4i5DkC1+8Dcuows5TXtTvpnA0GlIzAUUrvm9itk4Gm9Oid0MqJhn1
ATEbNXrMZtqLTJALqo9NFpL1HvGp/RUmobzq33EQWc7ULPuOnzP0+einhDk4/X92vipyBhigL1hj
gLaLVn2kOJozdGiaI0vAeN5VsawzMEeDaeWyTSyVjicDA0RBBPqAZgpa04Zl2RBkQlOlNUr7WSHp
stBBnq2x7bmFy2hZ8JeLqZocS1Yiq5lwOosj7lGslmxjCpl9GT33ARa+vFngR2IAoCct0lTYCUCz
d3NPan++xGV7c0O/D8EYIhfjvm4BZwHhvMxEpmYkY8nZD2QhJPPsEwQiS+H5kfIgawErPMy6Q1mY
bNq3EQhn0INy2M9MuTXgYWNaP61nh/OvA2Vu04gFr0/FJ/Cdi5oqip2UMmWp4WKZ2TZ++iTVjD5D
fwRfHPZruoEkZWCefQB+GFmthwsAi+ZuZu36emtqdwKX/xJu3e7AcwkPxav+MRP9xT4Pf63jVfUz
xP5EbjqQ0B3h1UjP5qivjg99tApk9BdXi3LN/uUcB7RcUjg1SUu2YOiaLP4+zQhYG/ROTB3VnYwA
nNc5lh48T+D2Dwr+TnPXqNLnPSGUKy250LvWyKEhZVUHSxVNLFXDvSW0kRNHHTiee+ZDdwhwNky9
dHUNFbFUh/cYooUNhVX80Gtsi/+4azv7Qf5NpNPdBmCTdfp4AZ0hauV0lOPvf+prMmmwEOJ5D8Nl
3kByFdSyYpTy0oIadlEPdNOzCzPLEHD0eUOzmLfFYROcpGptYKu58ohkD7tHc2wE0aCBy4PFmCa+
Fubhl2BTXwfR3krtC7oVAgk2CxyWdOO2Hv5iVKUSdzOZxyIF12Ur9LouAKvC0DA5zaxg1mjIlo7g
b+PdS0XHrluRUp/PL2fSdyRwgnmQYgra/i4zkIcPWY6HkttzMoO2MuTbDVJSoXYyC8gcCOoIDfNN
3PC4Vj4kcyqfNOjvWaG90sv5RknX1OyjHEqL0YcD5NWSMmvZ+l+zHb3te3Zbo2dmQHhpbGZlWA/O
ctadRnDGVG7WIxh3pDl7OdiZHNXIAFIgWt4pRb0pimVM3w5S5ridydYQVlY+bBsmK9tuGOoM3RXT
5bMjbBy/QP4TLATP0acu0+ywZtJfionKVdn5lAIgjL5zL4w8OSKnHX8SKXT8039TVNU+ZMyzoz5g
8M0+ia0bAPNo/u4wYH1xI4Q7UQaE7qrsJTb+2dscdBtp8wqvYMOPyXvgaUvI2PlAtbC3IOle8cQF
KSYuDSBi1T262iVmr+8a+tAya4EeGAaxzTodec1kKqz6sPTswhBU1RxNU9fZkNjNHNkqMyVZTuOs
r0yYIOp2oEtUK974hHYK1q8CznoQAniiqNXpDEIqV1mm2n4V3aYJlb09Rkf2jVgKYkB54WqjgYEA
KETtx2G4rTTzBwbLUQo9Tm+xorkdE+SfsZMTV3qbxDOwFkcqjCdbrMGahSG5plwLCE83WOrAcHsP
J4VKXluE+hNwwBbikgWUiqGgaa/SdIHLmJPYxzvNpJ4pg/nMxg1ou/1ffnORXTwyzyHgIK8GJmst
5LcuGeOb9VuMejJ5NQyuaO42BxqdFSFq2cIhM/IDGNEn7gXBtDTdTWinNlqt6T3iFugIIeoEBRPF
PzrR6amUt8ATj3fEmCUXVmtGfJGGg+j2+Ye0yG7gm/Jloc1wgufT90Hmf4V7ailELfbz8a+BIGW0
dGHOuGNaG8d56pUa9lVMED3h3A4gJ+z9e+58QrHueSjLUzyYgGpYeLT3D3ubYdh0Ep8Yw1m7U4LZ
VNaMrltKcj4J9BHL+FoBdA9W2s1HB2UN4QAbonpkXw4LmZjpWuhbXFCEoH5dWlZtfNLD+H9TygWI
IUTezZtgKTiEVQdGpRG63jDUSPVIdnl9wvDOU8vzlqgV/sQe8k0rZc1tvT2jauB7Q1lqp3G/Ci9y
fuUhyusnpYOM2Hy0aEYMrXrM7Z/utUPP1oqP4XK0AQeN257HCeciWJBxzYH16AzbjQZ4jwqndjhP
itRf/GNbL4dfTVTovFKc3rrfY9QMyEQuGSJgW4wiFBbSNeIAW3fs+MvfY0wM1DitovvjZbGNWOXZ
c134qByg9yA3cdZ3i87YY5c4sWkZluB8NTiiIPwPe/UiD2w2G6iWSa5jK7yEbFikZcKAZLVVEPXu
tNUVQjscxEFdzRfMR+OTRT3jhZRLbI+hx4mnvOyQwNO7YqifbpNrHBdiPHLadi0xxZo+Zdtq7N7q
hQVj9zbN/X3pOU3hMEW3usu0kxhGf31BdQK2jdlPEGfKWmlBIqV+sn3V+wq+DV8B9NFH1HJhKTyh
hVq09mJQjrrR31RX74WN2opzpwH3On9HzzmG7RHCW8aDYnY0Vba7KPuZ+EbV7RMOiGRg7VIgXmQg
bR9kScmO6hr3keiUQfQF/5SKwSFCA96kHxMjLBnGBdU2mGIlmT49yuE130viXojud5UeCoo7fXR+
NIt8zuRy9AEc5JlwsAzV53Oj7P+VJvcPP92FLnaEMA7gr+9BtgUUCcAv0Cc2q2qPV2tkDcEat/PD
e2ZUMKQSGAYOYyPRrmhGA13/QYYIxwsaJ80C/3FUykjEry0cp1RpbXccWVkRXjeC7xp7VHbZlNaA
MUF6x1wEOoYok6Do4uMMXGpfIqJZtJfjydtiQU29GWfsQVeLRXacBhkf5XX4/Ync5fnqJuju5AlK
CCSQC+9vp2rycuM5mirJOSQyyugyTCCTeBfAhlOcI3lBh8tiPbfVCLXpKHhn+gH1ln9xxGVF6GAJ
pxZYvvrlM4SOyAx08zqT4d+VYm2IOJWXuLAxiuobgucIUdauRsWsjIfEwr04Y7THUgGuZnKc5MQQ
jC2z6VWGQpXdFEvLKNmyxpUR29JCXeb8H8VLOEgA7qbsWCLA90jcR/v9x1A1cnbkHXI2fSumhNBq
JH+IMCF4QYfbYcuzT56t4/mQntjozVTkZAv5OBUoT/6XrcwUhRSNXLJOaqlSeL0YY2yBkaS+jtlN
mMFiYa0usCZu0EPXFHy2+gum5iSReVf3iMGsYnVhU8iltKEqNH1DLYgUM0i+LPUh/G6651k+GE68
c5yvyOiGBb/yYncx5ROIcxqtjCZs0lJUnKU9YL3dnRF8+W3SzM7ynF6WUk1m4/qKDToqrh8r6oZz
1DxWr6WqqPYGhrPqfatXdomqFsy8kZP68dRYX9kj443kKd9VEmND+NCqziX3ROSNwDmtPnndL1ut
/BKjqewwVfTC18N+9OEo1wDKeTBs742M1lYliglHNLRBN2YfXbyqt4RAuId4Fw7Y2xF8G7VGzFu7
OLcboISVBESjWX9KieDFP0vDf7KZcUB84PYH3PDwhY6fIz/92qoz3UR/EJT7Jd2+0LoAsn9hQF+V
Xl+hn9Rs+yLsakEoDJBIjf4mUXiM4izNqKQUR92wwAdkP1ENjOzxQs058FdtUQy03nX9JJ4DUi1F
PYq8Si1qWs3QlJfyKQ+lrwzLgsxr4i8KNlLn0o4n/Mg0KR+nF39y/IrLkwH0KSjbDibbxVyFzPcJ
RzsysXiBWXLH13ZvLtxi776Wtlz2AUKa51w9wW1f+rbzbidQSL93yRX9OdMSg6GARtMcIKMW5RBE
sjowJu5FOcJs5PWV+uHcV6zHaRtyCfZ1bIWq4LTNvoCbTwUBfU38WSZV6z0FOCgnBLiy8ZrYNSWr
NyTkXQXQO8v5CPBQVmjmYWMr/cVagmcNa/+7JoVHEZUY5BISErQK7pm01GsSbecJ9EVd8PF/8cLF
AUCQBf8oO/z5QnITFKf0JqL/ciMhjjqWq9qJSsY4+Ia6OdmQw0c4jgpLOk8psbKKj/C5FbqFGdl1
syt4RKimzmVCYiukOpW0H8SgEhuymGNhleXlwQPWC9IScIP8d2aEmliHImuQqxY8AZgz8L9cDPPM
Ej6DJ7xuMc0bGLjVKXLzMMbZA71cHauenGPY18wWWpiIYTFSEXaL1Y0agVBaUhUvN+8TNfonb3hn
bO3ucPjLc9GfrYcybWKjcGueQRho8AhzAaxX2pr3iSR9FBizvgqe9EUkTSIk4eEdDgpf9wVlXVW6
I5ohxcggtYKLD/H84rIZow2p1lQpeIuepyLOiRb9ItvcEq/X25Bpgo+3TJ8rOGv+zGpSIW+3n06L
T5RdV4Ti40H3PKr5m7x4Qq4AUr6VOllt/yaIp2Jl2JidXP1tZBir3UI8xFUA09qCVGCUrIdEvFLA
tMpkfEciP3RTOk36Jpd0sPgjRmEtCtfuTAR6QU/lwgHwDVn2oTxLh/Uci+YnJ99R5JCspaLp7GCK
4DmGlIyuiMW2k6e+M4hXb7LSWVc/VTmMU4Xeroqdb+7PyyB19CuwuwxwUjP84yiDCf8IYM+vPNFK
uE4tgOwI4cIoDVcf3iOUcPfiBLx/sP65bMZxpy0EAAN4+47WrYlikm4fwT0Umz/D+RiFiS/Qg3Fw
Hhq9tjdGRsuS++/hvwQ5Mg28YvDmA9Z78N/vdyxvM41W5gX8dHVJ3VB0Rgdypw8mkB5Mj3ctoGPU
wAMvgL+HoBKHy+MG40d+0JMwDAPoGuLpbOi9N8UTGvGC8GaVuXdOg5KfTymE5pEeekcRBhpbdQmm
GCf3tplHH88ttr0GVx0Kp+Wn9aAkCBqZ055KW6AUsBvIz5Ul+lM/GaNB6ziPuHNpQgnanEkEuktk
s+puGzGozd2zyhdhUac8cbXOT+vfJKW0KoXOFDtqHU41F93tfeO79mQq/ml+ZvSW1QCOVBMKZCSj
DFsJuam01L1+9lIFkI/Kv3hJrg8cfQCwJxNjl0SWyGpk0akxccq6mrl1f0SGxCYOxVuqisN6fmVb
9kJIxCeG61MojPQfejilhdfvXHy45o338QY+sH5f+umJEeC316aymtQSNxJvFRBFLr5lxjE3Zw8u
KUbDDdlTHix7Xbw63JaAyvRLjxQNUCyV0ZBPm5RFPKW9hEiDH8d8T8gw612fOO/bVsRHMXL/tyaU
LQnX4dTOi1k/SZ08s1J64L270BUCgx2iZi4OFhCvszQCLSVstdZinGDyJWhFtuXqy9TNyHqIwLmN
ZVjIVwi+g0MzeN7kEwrWwenN0357CwlVTBv6JCmh0GWI0A7xKmZLADiqqt+8mL1On21HvyCEoiDK
EJi/x0yFd0JH1ybMvmoI3B/KXB/VIBT2W3pm1eCG3pazaLq6xk0gJk7Y2SZd01JJfS3OBckKYf1p
9IxdP2PhaNAYjSiH+dwod1gBzr5aap4w5nbtTm9jRav6mlAm/0wtMIoUUgAx01T2ROR+8yK8hhVk
rk/NIXe1GLBxcmA7cqWaxFfZeRsDHuB5uiK2YJROgQAV1mWi1E3lm1ocfGEwwrSvL3//fAZ8bqSY
+k+0zzEMBdx9VkWcjzRUlrBND41Ad9tp+XydOEOrhe2RZg/69uWismVIUbjZWwRHBvFguGkBvXcv
SBSovjwwDfzzXbVP8vKQF6Q17jbD4HF6BCXStKamyXX+1iMwbw7w9HUN0jfRyPRgtkvDoM6m2Pac
R4w6DstQm9zb0ta7SQDfyvjvvA+7NRnkQAlDN/H4ihThL/sQXCiEfBDbWpOlVi5fzsPiJGhM4DhY
hqAlg0MBUwJZIzYMx6JYo00S6kfbZWcokginjIzawMNueu2FdLHnLo8/nYSeP9cH/6VovgveyRpj
vKFnWubQvg146V9sDjLieBV7jdI/SR1VXC+kxVT+qEGtlHCQ7lQ6ImYAQvoQs3Ek/cixYCCZjxCT
KdHjUE+nGy1C7Lf4tt22tzSKtkOrVS3JRGP53NaKvf7U9Fy4mQma52+V5TMb12rYSEAjlddxAnAa
TTJzfuEfcOHyJPy0m39lP9ja26LpeICbtSk3PBl4vpCe2LcPBldWonlSb0rQVeJAMixK3Bflb8cu
NlINEfaeNm3WoP/OlP/h8wO7FMOIMvZelJoXDxBk0GeLRlVu7WsGDZbtffI/TPKxhA9V4tzemww4
toNWRbVsBUMM2vXdbZckdyBrl7qAPWPmbHsErQj+kdABskurivnfHDmNtN8nsUZvWbF4lkAvZD9O
3CTDorLD9IKAENUc5+gE5ErtkhlgmPSHC/WaONcPfCd0tfEdUqrrXsrRUQYkdMpAzdWEvjBDHR9d
OPDE8WoTXXMK0ltH6li8CZ7dFsn1F4xsHtERuzDbxNgBWngcp+rPnRQNpm4x9lCR3sq3B6BpG8tR
J7GP1I2Y80LtiY7IV1WEYa6MaOmXR6a5Px3mhr9iJNwzJe3yUZv0jkKhlFflHBJfASxUE+5Uhw0q
AeTlYL37tUsaFmIHMVML89QHsZouP0IIdUkwpdum5RxdoHkhpCL5qKGN90OIMb6HuDKmw0e2NwOO
zlZqsGAQLuI4UcGCWSyjeFKn9NQ+nlygg4wX8qtyjultIT6J1XjoPUQ/NkYSdWQjuM/pDVsjZYyC
gRl2P0io9yWMF8cm8F14W0Qau3x2hlR/hs70y77nshNvj0nj2KlP0JRdHPUyvSn/Xpiuh74KRX+V
j2xVXGVCshG1xQ/cRnt1Xo0TGGe6sYcnBmI2VkjynNi4zL8jqmlqLpdTRmfKaj1OchdYNAuNrVg2
EfqjTCTDzGM2Nkq9QsiG8H2HeEYwgcoia+0ogakCVgezPcPKKlZZuWnOL/UvAU66VdYABeQPzi4t
sPGiQ1dQiGRR2J2becmiWzMPDVIRRA0piq7FaeDJzp01HulTFxDiW4nmKO54vZW9TEqFcDo1DAlh
g22d83zKd3OjX90vgnqtDSY3RBuWJMh8HYuxBsJuiFQWX2ru6A+H4bHMb+DSLeuuuYOR0tcS8jct
E+GKDrmPYyunKJrvNAFOvFow9f8i5CFAokH5mBCACn4Pr3LDPfNqlvMhf+9UXiuerMNMuFw2oB27
0hfCmBmBdsIQGEOaJMCnKtvKXcrHJIN6gECv5frgQOagWmJoMHy78K5SC9iVUweAvESKAjp15q2W
lq+z23oC1ZZohOchJy+waFwoHBMrEwGHOcoTeEuz0O2CDCJGRVmFD91OlJnQFj0vYfhsaVaQ62Yp
LMWHB1JfmC3NgmxlIkchaH2sM/gIFs1DMc9b2F9r8ru8Pltzt7aKZOdQ6WK57/0F+52n+t/+9rSQ
u2m5/IDm3a4tGrJE67W1F6b63hcmaNkx3cWlvzntRBlXhc1leUPqBB6RBCOJ30XshnjtFKRNpemP
GY6n918kICdMC5dLCUpuPWzXwa86X1bbom9L5uXpbPfkN+nOWJx/pkchFwVTKzDmPW1bris2zoPP
d25Ax7g2YzCsLfyzUmA+1VBXj6G3qQXVP7Kjt+Ou9VxWg/b7wA40paNvkGK7O3V3ZD23jA5NaqEU
ed4Cc577+F+1oJlkXxcOeaPg8rJiY+zCfZN/DZNVuXo2dxkJd1XlYr4evT0i+2o0wArFawsB9IEJ
wl2FYUB1nxFg02hiCbyvx+Ab9jbHhuBtH52zL6LrGeCakuc4zHDhZ+AMwx8yVvW+b7WEE2w10zNC
Rk1NfRO2C9mhcPXEYS7aykzEWEcZv1HchdSd1ofTIBDA65bFxvlUcRNU0++FUjng/tnXiyAzjw57
ShBHsUr0FsQsLHGwncGf/0g5fB5F3tZL5ZUekpeQ+Ut+WqX7c9S+iAKBV+F+wbxNTrWpFlmvYOpx
f/YS8YK2VnIoLXNlHiCaKB/3nKI+RALi9MP6ADNxsMMhgWnzmVygseJ2nBf15upnbu7pwa9QbbXh
bekC5QdhFRayvxFfvMAonkmzZ2qWh9QoC1C+BHj5Bp3kt4ULhB8aJ8j5HUrp5VXX90HokRWijMqE
02U4XDjYwfmk3i1nbDGnjut+CD5H8bJKDiGL6euliF5GxgygkrukVrVxLhyYhbqXTi6gZYs0pBZ/
8AA0M+nHxSLM8YzGvlXofXyqN7NJzDzYwe7BFNpWhqWJInUAv3GdKtlXfi50R5uihqL4t1a6zA6U
hBZwOXbgxmmLLk3caC2n3Lf75VCPpmHib3jNwSyV/xtwKhADPLi35pvUPQ093iIB43zghmMnn/9M
nF/WXQp4BFHv7zgal4sBIVELYonTXV7O29mnqmlDodmwDSl0Ytr1a6shInfN7hase/NxqCuVyREd
KyinLx3gS+/70BG3trfilYcyke5XCWrjn41QFV0NZORPWO4Fbl8jhWz7rq4qo6N+oD1s7lYNTESx
YPMtzoXNItz/52BhLV9Rt3RyUx8IhajxrBriyZIh0EanxosrR9YEZ/PgFlstW9vF5UeGSzTeAIv8
3Fiw3eIqoZWhlDhpdCxTElyGLShXTYKMscozeNtex2qx5DUMi3QMEbFS9hNLp+ixrdjkQU5Ph4uV
//3umUvqvGn2Q5vR0ivzhkzUI/28fOZu4ZBdqaMoDZlioquaOkkYwYHD7wONhRQ1Mb8Mi0D5zg74
1dLVNOzfOv0Ay160TwaKKweNkjk30/GGRNohu7n37fP8XEtd5RQLGBjsAMxj9keYMboTQTSq67F0
eBXTCMZucOMm4HsjUhqw1oFfUy2tjUO5PTi2rKzOuKDowKlJe+GnbTS6so2sAmOIeFHB5LH8IiLS
awKUMp3XphBTlxo4FVOXUc1yQBEFWrn2V9FA9x7OuxHdBWWJA46m9bHkMNq6WcUHza4M+eOzx/M2
ZOh6LfbnGgCK6H3TYV7Asv+313YOy4jVpe+PRvyrk9XivryMqpbXVQT3OjbqJPIVu3qjfhuOH73q
smPioRLikYHLaqjY/tsvwtNVJTO3leaZ1dBQ8hDYRdf7gFC8KgrmUlLR4N7x43CDnvxfcUthkwHv
t/9msH1SYt4B9arGSoKP8XxU+mBYwtYhajP6eCwKXn4RiVxjUPtmrURSsTQiV0ERbp/i4IISlufK
bVwVsJGWwBVBVMeRMjdlMg+BCt0sAyBepZE0HcREZo0RohZqZ+TjwlWRosvuCGkmxLtPmb+xF5la
2CNau5/EMO8Kn10lLIkYeiA3G4OBCZl/oJZp4F1G546YGfJQi5k6tIhmyG38VH3o1JBChpZPhbJj
nJTQsw9kmpGcbM4jS4i8FoyJ/foovAP0MG4P3cpb41qz6jy1Hkk/rF1quvOEyTrKKVAfuyEbU4VL
s4KHXQ1s/piREO9zqtA/5Jeo8+Yr5qMlpHewLTqHc1xA/TZRBBpKlrLyvAya1y53dlJGO8+W/qzf
H9xvA5djhESZShdJ0ugajA/g98VwSUUkB5rhg5GRkSWPyS69Uiwaslc+M8KLJb1W1HBjdc8Iejft
2m5X0hSvJg1OMZUfJp1mVLw0sFp9c73O9GMWBguVPelIn/dcG11sbEWIZPjNP/OtuqMWsIeByh8p
si3WgzsIZE/I62PtYQiIi184AEL2LH1WtFmvnhY+tdVUi6v8ZgdEDN+n9+paU2yA1VIHAQc/hBUJ
BcfVdbSGkRxPrSGozyu3i2VZ3h98ehMctsoYWTs5QXx+EZawRrVj8NhZ5FWd8uUW1qEsp4xfTAnX
Ij1zRbOhD6qa27ERkp1k6suNef15ASGp+/9mo9/xaRayHg+WeNpYRsHvfsrl6FCmntPTPUcVhUvU
lFgCDGZzO8ak18hjIQxEh/nWPyuxYdScuY+RceqE4KpdYXqYLa7DjfrIsF2IBzczQs+kZ8Jf0cSk
0s9I7B+6gYoqqbQwz45fWYlIgWRDY+cBmZQTynboArKN/I72yQcP1t0GiXRXMnWQxw9HPuUFPmV6
GsZUiPyWtO35BYYflZm5DfaSUm+rqWYZDkezQec/+SMLNiN2mxwaBVyPxaaXQU1Rat+EPQUYyvJk
vmbLB3mQxab+Wm0ne7VPAecKbthywJSKDZXiFCrz9FdqpWH5ykS762qgqwqX0ovLdLisjhRMT6Xa
6TeVSi5wvbgl3HV1U4L+COJVzY2jMO0POOsYRn+zhtBV7fxeQiaFKWbQtyhKqkHHo//KA0I39Ge7
3/2v1WqBuSJbJ0EEevsWDe1pYH6j2K22YDaMDxDw8IQ/nGTXG5ULTxtBu7B9DFRtYIqV70h7Ejtk
FVp1yu1O78k1pSSR2BE5tBIFkjH0olDONyf65ZlbMwUwz48azPNCzGTxqIf4d91Ek7othSyR20pT
oNJIPU/xY6B5pOCWNhajQzgj8bafsNBMEkKtIyhRklcZKKeNMFj3FhhQvOKI+xsAR5h2EBWr+bgR
czJ/FIDG8KwU0H/wsFfNSY9Jog5TopZLEbnrdhUA41O5cqXImLmrikjnTzS3w77spu4fe+dvk4kY
MfJngCU7s8fkVhCSb+Qhr7J1bJRukAAgt5YK1fF9qC7q5vNFywUUZnRNcLeFGgLxaVmNL+gjhqb2
NHrSGFk+JNl/XhztcQaei6/p3cLy5wkd5XY+qP7gT6yG09DwL3u93Z6VRrvhEo5iZyEqTQziznzj
QECbpNCSU6Nqp5V713GRk0ieH+iP/yCOH7OiRLGPtvRY94eoCh70rdPYBM9Wth4KTMNPsU7p5zTZ
EDjJTZJYL+Duyq+eDLeTwwuhFO+xF5rUBax3g4IZAYOu+6nH3RlcBzdsM8F2kpKWI+0HJmyHAfNz
PcWQobhMpQfOaHY9frn7N/jRLQ2GdyM/Gyb5wUrGwUOAWjhN2309Dd4Nbdn+4nLil4IDqH5hhK08
CWvZbg4QK6BP+IJL1J4FWFkVOHvsK4hNVju7do/iegFCE7q5OJJInr9e+s/vHl2GF4SFKOgvBdrf
oM4wG+uo01X5ArQJbCvzarLRqZYZrO/QEw13+XsfcAisCbJEOF86kDO4mbUpUOi93Zr/Xb5vZyhA
cVfNH9L7/cHC/rkQn4Tga1oh+XtK/wnP0uYVfKQNNec+i3o2+S8zKdEB/+kg45eApMhNLr//pCum
O8d33Ljc1V1Qsa2qo0qB3Ndrz9KujU8biLgqsohVLrPVrF1Z8nUZElNDJyROd0NYbNnl7ourkws5
wqklkgX08IzdLLPRkLdulegbuwc+Nsiu2mLOiypXf26JXpMo5OfaytgbQ/j6YHsioh38HWZTp9Ed
IbQs9plVGTB1mEgIlz2DKO9rTgtNE/48LfKtBoe+/Y9TBVE3Dji5/TlpQpVfbW1+DzsyPE6XuYuj
rRRLBJ+KBIjgjtTPCIns4R2kq02J4WGCp9VpIkggAMI5EIPCJ75sTqaPJwn/zsFhux8ynytnnCyu
wZoSaVbzIO0pCbxdLyLPQS+tz0iIcOeDPzbizxPqt9+mIVZln/nVvb7Dw4TeWxLYzO5n6by75Ido
XI5n1sVU9kmWbZy0vgbCt8hLue8fI6LE8YsAe8Tavqb9Imosj2EocJZNH+0Ewm7VYW9VYzn2f+hE
Wfa1Ogtigx6p02LEnt59n6FzmBNo+7j2LljzJ5yZYZB9HMdnJ4ybB8J/W8iRuI5DGwSTM/yfINnC
PFuFyLci1xEvDPO6U/gSHdpKu2lBRkj8DiW8rKspBbKg5zsF/J41O9RDSb7d9yreeHGhTyEBELoG
evO43A45nVRlqqv5/UOYb4zZx6R2aQ1/dRK1JboUHW6VM7PxP/ByP/4qKUsdFxvdvcYnaET/QR+G
5pn9e6LOUq8xPfZy8YOz2ZLIZynn+XWYRFUIVEYjN5Upa61liK2wmd5QhARMdwznXb/CMHkdXMRU
czc0ezsMNaoJ+jJ3YHlD6cBSEu1oZo08fw9HSJQH54uICaJeSp96LTjVwqw3YFsDFO66qtoyDP+M
mEkU2denfj0FtU+Fq5ruwc96JeUtHJnDROsiUY93sOLSR9iccLHynJ07fMbdPFBhrry6WmjNNgDh
cmYMK0ZUU+p0E8SyL3dlMwtMHQaDavdzzzFzr+CfIFY7qVb7JoomZzZlTAt03GQ4oZF8Pc5epa/B
w7uzbp5Q/55kMOEgIQXHGWf4OahzDGp9oPeDA2zuiiiLRS1JVc0N6mxfGlCGYqmboziStFJ7twat
K2dMGoIB7aASWVI5qsN0ka8/yOOkjGTZnOemIhKgjInHsVQpP0KDAk6rjVUeZze9ZPcWSgpZuGKM
4+nFHE0HXSt7/9nChOOPLOf5Sd7Rf3EaqRIsJ8QZxymGzKePb7creNbsAQgokZVZuub4Ffzjaxl9
Nf0E9ts+lH9k3wH3BUghG5zhadv10WWemCC5e9+R4Mz77Pm+e9IDknAcprZypDEdQV3QQYF2xt2Z
Eltjv1mUFPKkLJPSVB1Id8P/4bJXHJBtNeiJHJO3Iq2OoOQQyzjMe00anD9a0YpGe40zN4pbXaB2
dNCh2hRlq/u0fdNREZIGByfhJyiBmBh1RJudqu/UY49/kHFN1IcVi8d1Jzkow06/WhgCcLsu0qDp
6qwlv3paW4J26epUC8iM2mRopfNnxTzViBgvJr9y5Ye7DtIKUjgYO5P6eUQi34vbzPbwNYbpbgFn
0EDrKTQhDf0qf+VQaRan5uqIOeqXukTVM0h4RyxOdVA5cvrwg6P4/piwS2tXZEJ2l9PhorzzNCZc
8IgFttmesCf3vcqysvYmCraly+aDonYr08XV8NDeP0EFnS1x/s5IQcxOI1xnESxf5GeBhOVhPydh
Ws2hnBUGDXH4HYLDpPzPb+QVhQCeBLsCiybyZqPv9XMobfUCCUA38oo9H1443eyVHEIYCjSFQ2JX
1GyhhPm1ywvtjbHDyPwICqVBprE9ryB5QzzBdeNvZNv7lcj7TdpRshNaccoTKBhQ3Auh0ajWUWK9
DGMrCAFv98xFlo3Qsh971Gb2CuvagrN4ndbm5JopxRQk1qhKX8sImskuuxocrtZdEX4NtAdu7NaK
BWS5IyT795gRxFUh/zZuQn9OvfPA0X9qkEyYsthO/rDIQ3BdlVbsKqq7g6Et6KKKdEWkdzsAMMfn
nLIWx3gGLgjoYY5vQgWGJd7TTn5gbt3zImMDkvchuELsXYSue7rFIunPvBoHU9AjG3EwXreUAqXu
z+yncsarAJzC8Qbyt0OkcTCeVCJf/KNzL6Zwh6MBzcjLdXBPSBesdd3Urc7h6U6T1ZCm2KK9ULxW
L7T4rZQQ62LOkKEVVUmApMiJy4SyqHhuLe1itJvuvVY3TiwjGOSkEp2uTB+EGapOXhf4rhhB5iKu
Im/F5HDaAVOIdTSj8j9bcfs+SGg/dw0uwO/LdyMNKHsdUGyeSjt3NSAbKgPN3SouVoAtiBJulxT4
/3qZIcZ2bETBot4sm4nJEbMyF3TigpYmTzyrXn4ueNJ1ECQnVp+x+spzJvYNfeBXKU9lOQJb2QxH
VPdURuwIWsxrJy00c7KlniWMMeUtLKny9Tsqq19BcRq+ni7MOH4F4G9Lh9dGrfI/kPwgtPFF0isA
uB5NqMdrUJkpMT6cin01U01iHQhGB5x3AOYY6xvLFK231FiQhRKHQpyDjTP6VD3OgDYsALGsk4MR
D8dYjABdePMrn0PrqkdH7tUJ8qXlKfqA86s9N662uyXuyWdiK3/Kx7cATHbevYhru8wF1x0zo2kk
rxQ2/Ef/9hdHZUa8Jy5j6GdhyzHqUFjomNnXSei9f/Op9604nLvme7aOw8D6rrnwSTl1sAyc6BH5
Tx/NsbeyKP/KnsaovubxH1RoAlLetGRoNsu6BpOAkhKicChXdHLZMKQbB12wEz/KTupIPiq5nqnp
UO+aHDDJfBN0ukdTSK/B7/Wqnch1vFEuz17dBMJR3brP4ewHxbMpLxnw4L9PSAuDOSuCYGGZT0ME
mp87BeLMja9T3S0+ZHRuS/BR/FqNjNQmgxQULoVnX+fA5+XLn8RCWLsZqMSnbXN1X4JB4SkS/XmC
jbCXwi5A4qDwzVKU2yHelZI6f05+AfUrzzK0G6LMtp47V63KBIPwcE2gVUNSQfXv8+J4RSHyVRJZ
bjbG8D4UL5kZJZyWqmo6ErRkpeGvwNsmrEjYYf1UtmgUT9QtrThPJuKVIZ0IiVyECZrvhp1aN7EL
4kpMkBLjgfGAx99KYYMP3Slzj5C12A7s28+6ZqUl057Ra9l7IHDu0IFIMSB+1stAO52qCibrkQJu
p2+8xAurI07Db7uiWfOA/3mdfjwbvjk9Ckaw7x3lJ7RKytipP5nUu/T3o1UGWaU/uoBI/etSh32W
XPiFjBXf+b2+hFcvACPx5ZWTmZPBOuJu0Bpf76IjewTZguUAitv/tV1BFtWel7oeHHwJgsmCS5ub
6TuR3BNuQwDZb/ryXjw6+a2GDHcZos3K49lmU5sAXHg3QfTSI67OtrduLS7XqGbUegR8QzvoWU5/
DhoKCPGDSL4E+JWIWIOkNNET987lbIgYIMrQkDHl9130LSR8kxg7JyF90PBbQHS8c3ThbwX6ZYZ0
AnsIt2so69ZuxrjOvIp7A9A4UUKK2whi+9fEhzgtRGVVpqTNT5eg4ldUS+fsxGfL7DCA1P0DAfi9
Y6w4XQyJ1FiUA930QzQynAwEWJWrYqIjwj64bZWiLaPUTZlqQPKDTqcuRR5Jz3hd22xhwd8HR7wh
cZwL+COhHy1nrPRRWNaL57SSzb4j4tJi6Reh73yft+/gqCitUmHXKU2pjg6Jg6rPqEuVYJEt+MGz
WWgW6BY90JOJiP/Jyq3pM+iHe67gx/sZwk/ItB13vsc2ZktGJ2V708xCpAo8fjJul/O30v1r2u15
W/jCI7iqvgMShugvRBSS0+nKbxSNJwMozqpmJXV9WT9yH/xh3ZQHn2WUGPboAUG9zhIihTbHLuze
KJE34/rQnIDgVAjGPYSMQcWqsMZ4AvvaX5xkp4epeoRV1qyjcNnZly9mlE8vp87wBJWGJ8L+Wogq
swbiTgdUCDRoOr8EMArMyclfu2//T6ktK6xMVSJMthMeEii1OdDQTsb1vmaw7twSckcA2FVbpXBE
m/ROA8MqaMl4skAue0cHGzNcfFceS6lRwACoEb4LIxltdXrYg4JHHaHTmEP7uGobB5W3G4D9WwmK
BIqMnvDzfFlE1NSD4eVxXIdJ5aLDAenoUUj/QIwVpMBDDuEB4H7pNIkCEzoCFBwaFtt6AG8sC/3h
UOdqTuOrGQQcjYs4nzpCW/gPdihcKzS5zp3S6hJWs9ftoCKSeErklhdKWX8SL/OKGOd8NtxpOUzp
qZ46bl8K6T4svRbFDkJBfgwRGxjnvYkH97bWGPXTUsv0dnTOaSokgd9wRek4fpW9vqct9a8EYSIs
KBwW66MmDniXc4uFY+ciahvDD0GYHiJxlRI5Lq4LyvglTff73p2qvTUrmY39u1kl07TDfvKWyRBp
kvTEUEoyDrVJxhJnMHwpQIBRt3HnjkyxtYVqEtuuuV9pCiXLSrwdGMqglCUMKe/CKgQ6V3Hrn9Xf
ZBdv0gMbECq9PujQ2Usr0VF6zfUsATt2BulDzRXD3GxUX+NICwF0URAOwkdVhaEUhybLHwNoPRZD
tB9JR9hHXeNGCWJ0hTlVCqUfy1dLQlR06hZqRu9AOO7UztNxYjJkwnCVBfKW5OlTDOhSnvGwN1sZ
68Mf1L0fJ6hJ8lO5gMKa6BAY9HbSF8d6m2b9dV2c8uHds7a2LHyACvQoiSkZlitlXrLWkyLJy8Rl
FloSRLAMGPFU/cAC8pW4vdZjHXt4gCbYm2f5EI5+zNwDKyYJSd9H7YlP7YwxbAkkXXpxefXUzFTw
CKuXWHLitcLlrzpMP6WCELpFmoB5tFezuUwjMwCccBwg8IglyXryYymrRPwV5tOzvsb4PvJ8Qqjw
y04/tKx2akIcXF52YDeKeXE5+CdVgvoCGNpepEhmIFd509r0oItMIpFxqjZ/EEoH8OZzPKvqqPQ+
jgYzKU3NKPL5vQchadKfAGDafOXRUuw0bBUQeTK+suwOzXZkSezYxEgilmaee6YolizwyBxQb6xt
eh0xnwfANcrseWpB5eIv1Whu80qwslJCIhPwvvhNn+viux4RaViI4TilQj7tD0A0yI1eavU0KTsy
Gh7kYEsQSc11eRzgCR+PvGkVwqzaX8RhtOXUxp38v48CMVXHQHzCe1I/YQeHii/OwWyA0ga+MCzA
TqYdcy3Hh+BPpXk4PYeOuIBkF+83W2q/wWs86MaCwc0ECzKJo4Q5MpmpTqHJaxQaVyWET6c0i+Lt
WsXAddX3y9BmgH/XwGQ1d93OA9LAzB9K2PWMTYJglSAtZvr9pLcVvrbtlz7eLCsjXKYvqm1ZroCW
YMl7esWngFCpxQGVZGVL+CK+64aaIPmaOjPUUYqSKz71E5gplggXDe//0LMO25UeN5Kv0WjJtNOo
+GMDajhx5DhICi0v0VJcrQvcwk6mr+oetMZDtGKzvRp3YEUHHj36WwnhASrOpDuvxq2MOYbm7ZWl
mD2PWNWVHz2Z1bBBwhi6EjrZynuEdYbloOiV11udpzb4iXUKTLsB8xtqXBJrBVLzd2Kw/2+5XOOw
ny2bcD72/oozy+r16ps1l4sROC9/I8d40PJyaJdvFasLNyphxySSDufRWFCP658CiDCLAW8+ow/K
emeduUnmbcF+Yzbc/f/MzUkEu7FJFsYhe78C0sTXMChodNaZBMJAn58N0Xq0GluH/XmqMQc7MEy2
F+4rQIWgX0Xk7OOVwMx+bg6zQN80t9Ajv45RdTPa2PQI7J10cHIJ9ydGFlB20sIR5CVBOFiYMu8v
/llQeRkoTVEEEQEDlICN4OToGamQ6MYHSfCTMj2mKMQmC/GSpRb6M6bUndnI/hIfw905fOU9zHGX
wSNQpZ+GFhJF2ENfaeDHUY5yEI2XlatLSxScV+imVakoJFjLJ2ifRtOIlb7HdBy48Yt6LpUcmCvw
71JxP9jG4bg69mcDZKKAD578qbKLJdJOCSB07TnwttMX7PGM04xKRVAE0shUpPZx20HHTQxuJ2AF
CSC4pkuXbngWpnvNGOUedxmKCZay4vGPI3ybzNuUUSxhTp07LQwc6N5ERQLxPEIlg+L8sWArHXqi
otImT/Du+1kdNJBjywVGNDz4TKHNmfqPRlz4+Y921/W/re/M6Gb+5FHLC/tcbT8+uzZm0JzKZSux
xgb3BwTB/A3ZCMJb3pSvM54OEJ+PCXZehBMB+/m4ra9sOMXRADaJc+rXDXh1nEiDkBR5ciHMyWo5
xTmuP5rKe92e2wtznrvfd92JJCR1+B7NfO7V7j9fbNmfcWP9vMC4B+/vjNx5uujrMT3yW1bleUZR
6OAFtt410WG+xqjVpFxe32e0g4wwReQLkunbdnbcj2Tm3brZGy7V+7p96DvEUIo2TbmmYk9kuBPu
6dgrJOtIaIxKZI/j0lMUWdh8K7EXQ3MGGw7uq0/L8Aot2jWB+U+xOisRqNf1xvDNzSowntn9+7Nb
UU2nVhgRGK9KbDmmMhpusEvQLSEZ+OkXX9jT1qhYHTvIlo8fBVXxPV59+gnUhdGbjGTEIs6NiWun
tssPF+1u3YmVq5oKAEY0ujST8T5DO5he2UDi6DwVZiIDM3ixDY/YX9z08qJiniYKDG4NHMUfvrP2
uAm7t9juetpbt9TC4aFPqoQE+w8sSBTPssspFu0TKvWqGCvVUrkiBRP3Hc2yLyiLXJlA273gaRIT
qt8vDdhJqU+ny6z4pjGLPPW0i3+MbRY/MUTbpHUJno8l6QiI7LgxM8iK0RFqcZH3WzdtImOJUfka
wkRqKJex1QAv1dbb3AclQPxHiUerONkCBZgUiagBIZ/LuOEWfppyUyp9f3y+nwNlTGmqA3eUYaw9
THu+mjmIYAqUsNqkrL3Zl4AC0ZtqllsXhzW5FL+fLuVPAacUN0CU/i0j6AriAcyzBNg1TtU8pIIp
pA48AIr1zbgMDfuI2HVPVoNRqsh//eoVV/hJOYjtcqi3W94UxGsezNpuHflQQySWNcD4RYVYN6rs
iN21941GlI6T0ylEbqF7m2WqThSPlvTdXZsbAR02S9IgVPE92yyCCoVi/6/qZA8jE60L53UyCy0t
radK7P1nxOwwfjdoyMPSJSg/B3xDn3Z4x77hQE8tnncXwYN1GuGWKGoVmaWm+RJIYTAeLkEgL7Z/
RleY9KQKzPaDrP1mMbBbtgLuLD8Ox9dW9ViHhRdiLri6UW1MpELU0Fkiu95yQyuKKMITRaWNI7UE
z7oKuFaGv77oj6ktTF8yAJtc4T8DFMYzKv2TgeMYV9IM2/ef7jMAx0L1gE/HqRBLmei/O5ORhm0x
6tb1kpXm5oVWZJP76LXheB5UPv+ae5WmLOpsoKNeoXV2gMfAsMtx6SOP0bQewc+W+e1XyMQmk6Nf
PT0uu30au6e9HSrKYR3bC0tHlflQkuYvDCjfQWKadCCEzeU4/+kGy/SBQFHTWsdo8LlETEHUcU+0
8+/0bTeNh/I4uEdmIMmrntVbzq1ROhFUENNG6LhRkTdgtLH9ciYB7cAaHzyGxbEu12J5ypitu05G
NKfqmuV/b8+P9FKl2XAFsvFCHmn+aAYGMOqFNr/BwATIQJx3rMAMCXvjt5jRdLy3MunShoGENXt2
ue1pG1NwGne7Hy4+ijlkWUpiuKMdn5bJyoTNncK1sNq1uLkE8v1RmBsiF1KJdfJsM+R/vg9fw1oY
Gcy0NkqZSeMXq2LMa53oqGUDvHL+sGiiL8jjZ6WuLl/E7060CzWTQnazl+AN4Qm1Pi4VMSw0U4R/
J/WiymZdiAcyAxqijC08FyAPZOog/4ZXhcC5HoC7TA+Hl//BSCJfmxrr5ponaYISMkrcuJbxdEnr
VOdM1I0qzTXoTaF4NvtTl44l9Ko3R9M+PUFPC33yKfQnEjNLIY32rnjphEVXywI2WjqzKNmtK0/D
P9o1Tp1+Xik6LbyB7vjTfrXrjCZBWJJPOEur9ef2kcy4UT/niQdbGopoTE7+6hYkxNFMNfLXE2/2
TAZFgqjKpnsBoyGfM5RDTqppXFJbewjSyByw9GqTf+X6z0Byehjiv64QxIcVACOKOyd0U8ciKCoO
Dj1Aza7LR2QkD0y+yFPjpfGobABcYzkwXZufJxZ4IwYqJPXyYXGm5w6dO+V91HPjLN1O2VeFe3M7
dO4NTz0mNKaROxq53mo05r9AqMYjlz5AsfdAYxMdhkmoB9lfLJhv8xBkEqTh5ZfqvUUL6S6ciL6r
o+k13LvNvy2DVqBSVwxsHRTguQyU4adkwpEJ15mb0BFsio32AZh6kEw++9M+/cPZe4FOwHBzWl/G
Uz+7sLcXtJRGQRZw6GMSetc2miR9e7scchEHvK6YseE0hnBSjp9EoWXw+ghfF0admb3hd0l+V/Uw
QUX0nJNcinMcDcQkqRCa/2clzjqK+muKTxnE21RX0jXhUUU+ZF2VBcXrjAqEhJEFnpggbZboTxdx
O32EVSNfB4eS0zTo3ZIQrd/FUO79PpQZXWessac/Mm7QrW9m2ca9Dzetv8NiVwJjMwNmM4R8qX1g
VIzc9O8TuU46LTykbPiMSIS0+k5kwv+t9pD7bpRClaZnwv3w85qxPoEu8oRM8U8btOedZQPFNNrS
m5pd3bi95XrjbpDsp/5RKHaKBt3v+P7bqla7IoeCj0Q/dhbljs5an6F0iW+Q5B812lP+EHJaOeFF
9oOm2tVHrFwrmnzmV38TgkDUbZLQNQ2wWwdi4PlQWJdjL9+GrGyX192R5bA5GF8xF8iyRn7bBFIQ
GjeVF3vNC+3/kkyRUdW8jDaQzayHJlSkVdU8U3CTECEluIDAfbu6ZHs0DhkfIbxm3LXNu5asmtsT
THTHh7s/iUB8guhjkfSTIpnxaVBe2LCpWbACfbkkSyMgt7Nm2+b4YSXr0IhQiYzoaPLjXYM/oAjE
83n3NZCddJixVShA+/VelKM8yyxjES275XNmXrpcT96Zoob/BT3NcacKnGU3M45y4/ZvMOgRC3Lb
LVsimG9SPeCati3Bb3DElHx0E6C727JIViA0KIRVMqRcHoq5iARM5g2llp4QMIU/EpSWhvInC/jr
tITIF9/qysT0FxL2GJBTKlXACCK5XzYoI7Gszobb/veBJvZ07NkcMRCeWmu6oqOwlVwKG7t5SItW
2aV7v6WASiKSQWEvdTk6B7KcTR6/b6DswvND1m3wglQ2MUnxIwGY8MySyN7xrtx5cAf2m2UadjFO
e8ckSnXCBTFOgrXihTI3DdfcG9hKuIfEejp5HFVI+pkYZtfSGAwqrGetC1+QxAusmA5C3QyJ3JrP
EW6tYCTEQv+OTm3NuQd2QWYoT6O9VMRsyjqqmiWO+LZ9VAb7x6nmRyrvYqKAveUmNflTJYBkE8IF
TjYoU57VbgWnBrbxrImOyUd1jBwEYR/QWjImvMlknV6UlkJ43QtsuKIHjasjP5Q2e8LoF/98NIof
e7abh2LzrloP3XpQvMGCsEyTdaQMTVvbIIk366h2b/fFucJdN1vBvVe8td00Rq7SD9fr43pq7U39
bLCT1G+FUJBxByCeFsDd2IOav1gSDYfLsbo1lkv/6JB6cYs1gK5oI5i83yHroAfPbe+DmO2+qZgv
oE9ql49R3XQ2IAmGxz1yA4AVF3x6xvk6gk6SZ6Ww/06W7bxNqmeUrJDt1ry6g5slpeysy9Q13P/F
Lu7pfefhe6S+ni7PFmeyhLanuoyMk/18B0bdN8HMS+G2fD9nWqecU6LFJD61EMHUMbdp8YdcVZxq
Og7QJmik5zoi1mHuX2RAkEd8hq2xEXc43cr7tMXMNlXXkHCj7K7bR9vFVoJTpcx5AwRZz4/EaovR
dHqepsh4V1Hjx9yar0eAIONUXkZ34RF9XhrxbSOGK3xs6mHUTh6QT/YJ2bT18BP3cwpeQ64Ggd/u
KezfWF/RLcdH46Hm/upE/OLdySsKNkskeapt1v1J/AMDWF244gzD1mvst7N/RMjAtywcHntpP164
uTw7PiSwUwUbXS+tItbtjUB/8LXOEIsLX5tVzEqIuqzny7yh0/JtDrqaCf9NHoODVcaq9oaD/mu7
atY1OIRCB95xWvf1jk2T/aZhZ2/k6pGOQoF5/0FGw/b6Re0ORHhAiARQD/DRD7134wltTEQMDHzv
acONkymXmP7wu3O1ejbSmf/py3n2fq7gTsi0D++vxZXtrtUFb8Qary3JsSDVRUkA1XDnN+ltpHA6
kkr94pZIIMH+490vN3HcRteKxE2eC+H7yYwZk865+EkxQwob7gaMDE5awag3C5nCJGZAziC2c1uv
dJxviznX7WoP0CVlXGLzTaz01V4eZP05U6x3vBeJRzExGyQUiti99X76cpWJwyRFbEt72fwbn/jp
JAnXjZqS4s2ocKxwuKbYOEaqXVEZ7ayIeNjABgLAxJH5Ld3mcJKtDYSw+9ncEMlPHeYLlgbdFZhU
f4+064vne7inPVtQqXWpXCLjGmn5OZndysrw/m2XnFi+DTbriO3eU3RBCUGmw9iHlP6ohCzbrDKx
XhHw1lwKVKbI4vKbi/GU0tIonBmEcENewEnmR4hrICxXZEGhEy1XD+B8ioQYpaITaWzPojeeq73n
0iO6Xsql8NiuNn80OzAVwr3EhJVbDZsRGI+V5ZBsSswE+H2Gq3vEFOgLwBVFxIjke5CbxJ4YK4bs
DYpdqFjjNvc+ilTzWYDJGuK/JqNOIw7XaHAba1kWoxxdr9xHL1fTQihdB0LyWEpaYRwQbl56/ky7
THGm4XOp/aWiOYnohrqBONphBQhO4Las3Fp5/H7uqVOoCu1Oe1r1mrHpHsIj3cCRh2dXM7drUGL+
GCn1bVFPlISmSfmw9jbekh8g/xmrQMvKKo5EB+7mjAXqZ64rnLyFh/SrheVEXQbW9V5dBvlwUSQ5
L/xmKsitgZQGXuIVLaT8JsYHkDKkc9s/Oo32BYN4CoXEK6nEt0OQ2yWVSneW3U8j74+PzcCvKDvT
aDnIYFU7znhxbT59MIqp5MyG9vjFFJjv/2d+HRPdGf9aHGMBAz4fI/r3AHrlTH6LYR6i5CZAu/tz
z6VUCAFL4ExgJg9q0zrxXvhn0szWceYieC9EWguqmmzvmJGFGtkn0WTxGOLiv4hJwpVXgq2c+7El
GyB7049BfTOHQPrrqMfhNn+nIXEfuFBKwbozyPiM22i3a3G/jj/w/OL18xBlAa99gP244i4e8YkO
SaGSGclGLKlI31fvBFqFUKPpfLx1a/Bya00WVYbJKSSTDWvVLkuwfA7IiqKO/Vyz8WswmftiZyUJ
JyztnTbIp0tllkj4h/GR1FvwDX56jGTEkGk/VF5mdOPu9+rQA0mo+Pap8WYe/OKB8wXd5QRoU1iL
NB0yRcez3MGmi9rMEyc5De4Qn4u7n0LMU/F0eINVQQA381cUVAU6nw4lYjgFkH4loUzYZ+SdAp0t
Xn8/fikw3fH/rbmIpOr9hTRjp/MuqoPEq5n8J8XFjHQ9fODSmfYt+HobAZbuEugBnlH8fj9++3eW
4Y/BGko43mZ410SMWwNFg8N5xeAY53+KH9nSgCxcNLurW1I4LXaD/9OwPS1/53DfzI+Dpb4khFn7
v9SxFY9MRqBm/pOcM3OjLBIJ6XbcAs70bpoqfUF39gQPj/UUwS81MqAAIV+68Jl+Enm8n3pBnIzx
MQPHZtBYJzwzlEqWX8ceLS3Ue7PjdZcRPLIeknFqoClcVYdI1m7mBEI6/gjGWiu94Jw42Y6lJxVd
ONQcEMMqOdfoWLhaNnATecrD0hkv0dGtK4rBxaOA13OmGmbgJ1QHFSXdSZ46qzOlj4f1HqRDkTz8
7sDxHhacocY/6/P+LIVv3R/BQndb9dyiOAvk7b7epVYBGrIy/hjvwKcKfvrnkRdq9PpVr4qVJJsA
RgUii5QAwGAz/1vqWKYic3bUDTKeA5rMqlM9h7BTfQLxOBGibujx2Xr8SnA2a5wad2GlDiZMzuW5
6NQajb2EU3HFSH7p33hz1rkeiTHlc7Ozhy1zTBHqPY8x2wI8MvsYy0Q75ZLOvthz2ya/EsZ4ZQA7
+Q8FY+0c9y3RW4B4nmQ5clQt+bfTnSF3+MuIreRTLz03lPAthvtO+c36F3zafYm1K3Z9Ve+oSsG4
UGQ4lgX8TEO1CjoVxkqd3Wd49Uy4aV3X31l+xzVbbgvX3RKDSCEZobHutOAawNZOrJkVPTmrYWuO
b41lDftgH7SwzLa1+zj2ebGMMjEncKCdtATZBCHfFlwMDmIMNv/jUyvMEjtK6fTKzyEBwGF1qH3g
n0RVwjpMjycgiTH6SkP6Zgzf/+DzWRw6cjCMJoQ/RCAHvQVYCJLf0DlavuS3yrojPJEnKUDOsxaG
Fc2v1F1JMo/6lpfBWeTZMKCBmeWNmqOpKWjqJke96SyxzOQ58vPuH0TNCB8WlMr03UxyJpDZXn24
XRGMGSwpEfAOEM/jEdpdnlHyqSiuIy7CS2D0jrfwnM5LA0WdGlIFmPNEpvJvBu3B5tsorkMZuNst
tM49UE18Lwo72rO2Sg/krzoYaFOQpwb24yOjPYNiGBSu+/cBaDLUCjsy4YrkKPPE7JeQqYG0kTsu
uRL1EXDZTgH4bjFCmebhGXgZtRg9ZHIQ8nK0jns1iLOqBfhsVmo2VUhlYnYL7M8w6L1jAmMkLxm7
mbbh+mlHI57n9X522MMq0UiZJhjIfsbUwiD8L7ANpOPBiyZ2/t/S+n8yIY/Ytm9EeRJKY2NBxESv
YLotm267xv720hqeLlR/pkgfMcWp9OZ0NoCy7CNfNMxXDYUKDZLfa3nvCGdcv1Cf8Rztr85KRFWT
WSg4HkKzmuMR+V6QxsvBkFb5oWjBVWdfBBQPvYXeBhFrM1/A6AC9NZ7E1LXkB+VkKRS9V9FWwV8h
EaH0sjNBtm78Kh30o3NS1F4TgGWO27FB/P1jcXx8h8KaU8pWDhERL+o9PIB+Jd4sKlfR57pTTJW2
4ApTbtCZmsMq4MEG1YTdUZpGC2Mw92LrB3MUn0+FbCBOw/RxyGuW3zIej4Q4l98DutLa+t3+9TbL
igsZQOhPK4ZvnMs2opLNWbmP7+qsPHVOEAfBJPLF5tObCqGsXPjO3Csfut+7RuQAD2NCKbcA5o1w
wqgGi+4Gg1BYPQlHDj640YehVE6haPTs0C5WTFJauqqtP/c7qbOTr0oAgWmwf4DFJCQc0oaTtBZF
+2cNG73Uzn428kNxYJYpNrtmuKD8cinCdId3pBkZvdmXHUSd/b+74pz+PzclCrMuvUyr6XSbheWq
+fDtYIMwK+bOuu0aIQHMDF62kuVLsjaQQO3SwfX2hRne06DbJN/6R4oCvtPX2zFTzdKmE+So2fCc
kvJF0Xf+POpSCBRy+2OlaB40oIONI7X5+0rba6D3V6WSsjM3Kx8AkKVqrFm5fIbKXTHLK6zfAtDg
zyq0WNNZYFjE+GmDP82D3iedWIJ6O0mjRqrp2PCdbi2A84X+ioO2vkFmBFIBZUH6rk0oxaFPl2vo
EJJKq5cN60HkKNF4rKwICIGQWaaaD4cjUSZd6rZ46HEUdNJD+m7yP1L1kEQH6RhnIxc8PLnrVkoO
XI19+XdMHXDqlSI7j2tWHWlnCAQLeOCIfD2/GnU9i9+11WxhGkyuX43AhBkGv69LiRH++ROYtpFC
BZQ46zmhpXp/ig/Ou5WRmKuXJotB9Uqi6Avo7V+dtB1/sZBAvu4gZl7xmd07f/2D07mOrQaFW8r2
zlHb8OAMp6bENWbKBfTQ2ruxn3Hl8nPQpDVGa8jNSwv/CF9v6KmAZdW2evqUY7d4ibPY0DWY6kL+
bYwBVJghB4/VQbfy9AJb1O6I66tRL+mWYFZvqi4iiRFdj6KhQKgXwI3mLpLb1duv4pSJZYwTkfkj
wOkwJRQkSNMMKeoVt2LqP+FwNOcuDdWYa7UniEDBFXQAMaCEq6RqnJ4qsSCSgxrZaIJnoEdD5o9s
fUg2I1KD44qiLfT9YruOpwUE3FXbGSmMUx6OmOWtp9YdXrOlUZmN0IDCRRkJFdT75Ae31UTQOXXn
Aq2NMOhTN6qIs5z7uQuSbhyB/vGKHRUqNy+Sb3Cq5oO7fPOt2wTSs9FDguYvMLeyG8zcO0S1quMU
HSwelHDmT/9/h6FkxWKgRz6rzr3Y+YB4OXhQXuI4crVWWB5/GYvXqceDUc+cnMKimnnAEjKfr/1d
mIki3tMm5E7LkgHIIOaU7hsW7rfRW54Wgqs8skzmCOFEPddSlcHiEIQgq5/BF3TJPSEineUiA6B+
V/dwubOHtLQSnV11QyLXjqLM5bAMgPN3Cq9hammwllDu9Pay5LeM0TNh2gcAcTo4Vxg3ftVe2ZfJ
URyJojX7D8bja9PSxwW19Cfh2bDT1aov3Y9fZg3MW6uDrn640rHW4v+DpJW0u+BU4qkPcdSWVhyR
9YbZxjhi6GzWK5doa9lRcHkF3sxfX1N0qo1Qnc0ltafzeLGbPGHAPs7eP3lPvHUm5H00ls5ZOvkB
PvcE6DKJS07m00LYhPuSCdtjSVPuLw/6lRzuwak0hcbmezYyueYnuopHCHllo+A3wgx4zaE8NJ49
crmiQJEh+QgIIZEcsGkxMUdc4+U46/uBLCyIn7mnnwanYcgsHpCScN1pMJjew1FdYX67RzXRToGr
4ly9Brg1DGWOq7JdE8nWzfvMQhsFLDRV1sHTZPMy2VTl7I5B6y7hZvV+PnY0m/m4NvFvvQ1oqS2k
pgpfC/EkqUfw6kYKWhwXR33Vegj7PfpArZZhDxKaSWsh4aISFQvCZdoZhtcVFMGOGec57wu3wq7D
Z4SBIFyEIeuf4S1euR+qCojVq23yBe/DEdnA14VRMX+ZMWOUIUIu5r9xxGhXvTdImVJcjOe4/rYe
7XVCmmPK/8yo/4WNZ1GI7Jc7UAXjzyPptOqWujg+D9/k3JESqbQJujXDQ4bHBldizO1roKC87K2Y
NUvGNNTqQDHUcT2QuuLhAiKHnuXoQZrY2MhICwWA1Kh5sC9mdS1CPEdOhwUvXVaWeMvwKZeMwHhg
PPUPJtuEFHm5K3Yrx6/Q/5FfZ7UwVZsYmB0EykbohaAt0FW26ZXrwR9xwNpEwW8e3FnsLz8FtaQ+
/zZQp+JmmqLlcIoSCVKBwe+X6Lu07k3jAaFYJtENAN08I3kA1w/X1+BLl0tElvWsIR7YY2Zzb1x5
nzEnZ1M3blZZX8beTTfXdrKpN7EbXcFq09n2xV/7C5ge2s45hbqdRqCCeF2kkQYKqks3BOwQCGXV
qf1GdtcXstlwx0I742MqUfzcc7bCXrDMxsEx7inZaMpTgZ0lpd+gd/aDNn0IyW43kGNVXCFsUAAU
pcIDlfHs67J2q1VWjiHUz7YJngI3jGF2cnCE+L7fdhtoHuK+VOkXQL019ADgDcYRjPvmi2du9AOK
sRTIAwpzPUGsA8ofX6Ml4OmBeBoPuP+SipPvIF+2JOCmEk8MsyElmqvnqO/sdC1inoOik39E+y1G
N0JeWVVBInfJ/pqtXcF1QAyAGkbhKzAUx+blEIeZdCaRyYymJN56KH5UvlYfYoPJWyGOF6sClaRR
/WnD2jXKW+Q/tDqWXELcj/s+RydXn/KuDdxDPlDXeULHKH2WqQlM1qMrFyqicm13hDoi8Ovsod+a
iN509DXupE93uwwbEMI8j/wkqK7Mx3ebcOz9CDE7RBHey5luD6kCh3S1XUfE68U/PEz+9xMIoiug
q0tkfYs5HHtMOSLoerwSUHYKRT+PRNxF2dLHoHwvS8mYv/tqkxyH2o0Az+lZreG5N8BDZ1RF0Vx2
qhGtVJ6QrXp6Dowx+uyY9jx6Cqtytwo3wybayc1rQJuyq4qbi3Waekme5DY8i05P1K8A5gmyQiyv
VD8NLbjuvdXR9RTsxLzbQ3qhnwbMShiPLOTQmKY0DlUwo8u/hzsIvUmLsRnDwwB0QYbr/yJTOxst
O9RZegQAPZt3A6fvOPPcq9vPjrrKtcAmuJReJ+wrTuaiyHBgQG9y6ovTWW4oWA3+TrnTkD9bklsr
sw2gWY3Tpezsse/f800p/UfnjxOd4dIcA9EAE2CY+wilLqdJp7sJlL8UAg1U6gLvA/vmgPEnN3NQ
bVKXEo9MqC8pVSC2AA/AfUcpPAzT8WMi5nc3qY1jrd0SGBBHYN91n7A3oyZVu7lLW5+9a2ure/Zq
TRtNw3YBUbgwNbFYATRctkizFNro99rjw1vKdanU53+X2ifjrC3cG/50P6p2ss2Z59JLotofpY+D
WMHjcq3n6Qs7G6wFMSRNybnIDpHd+YUiTG3nGB7EYwIqCqu2IK5VHjZvKQC2yJSVSw8fnmqVQE5R
hB+ZOICwVpB2gQnlVz9jkEsljrO+pW6I7EiG5nkAYhPRgODyo0L/iMg98AeBDw7hNcCoKuScNntQ
rHEbVUTw4FfhkGKS8YTOQEACjsEnaOcCVo3hPZXbfBsvVB92o7thNhRx9q3K7kjz05PaKquWMzXV
3le7uqd5I2inejx23rMQBHOyFwfZ1KA5FcURuiRqZxlFd+RzW3KEujvq/oPeWW0t9eElv0zOuCbd
2/VLaR4ViKoT+SyPxRzJSglWX8tvpTwpCTqQu2QrO56sR1iWX6pvyLp16r2jUn+2DzfAba04vLv/
G+W6jZf5tp9USLAb5CvTEp/Od7GMMMUxYHNQvCSRcFGJh2XgVubtRFPvQlUUnNU683liL2a9CrEK
t+HzxhYQoBJAzrF9Ns2a8Q3mVxE8wJPxidxZn5Ly8b3dRvV0iIqE4Uv/d6CeKeHmBdjnpJnVoRmu
tuau9hmFVrCVCVh1o85Qo5h67ZYYoru9P8NO+4vahdCoQ5wfqIFPQDQAbqlv8AIXJuvlLSYkaXir
Qg6GbERF4AzWz0bIYku5gS5IJ+5zbEQC7BcMngkSpX9HoJE8ooJ/DMX7tM1xWvbzmhss/6728xqq
O6HC3U7HhVLlJRzcr7s2zPBPilCeK3uWCE3SaRtUNEQmpHvJPYawx0Ot6IDhBQDZ2dFC+ljCN9O+
bIqpEZaoKCcGUnTOkAhwhShv247zWia4h/bFRmya3w770ymac+iFF4bUjOAZGtLY8AImQHbhQBKS
CWpqid0Ptg6F7c9j3jr2QoCa/YZM9NxVQFq2tdoYZa7VO2a+JIdQlqzmEbfwFqY/AyZLJ/QLUAvI
1s7bA/8/USko7Sx1Mv1ggIQXvnQh6+C4lUEomCVHtkTFjbVo/25vXeGJd8xhboWUk/kuhs2kazXd
LMMJhgg9nUEcswkDET+WmZuqW+xuw+rKRdDVKximmm2abltzBMs4SXEcyJODqZBp1yTQ2I12bS/0
l3L3uXyExAXBMFd45q4Ns//isJBNac3r8h9VLVEzJV0DxH/3RbT4J4sa/S+E0gAKTdskmCFdmiD1
xA07z1gPCnfoQ+GfuibCnynpyQIR9Ts5ww9qdgz9gVmVQdsQeux43CoSbVzZ+AKZA+tEuC2fLvtP
zMUib8fwjDr1DUMSubtz+DxpVLWSd6TVgVaTt5C+4TzYydjgr9voZ2y0WyUukL3mnPJ26Blb/FHv
NPFd5BxA4JKm9dZoUa+bDSGdwXyoHuXOG5dTkdhl2r7LFgwgriGG8tvjHmLrd2MY7pvW6l0YHpo0
HfiyrpSyboVn7+wbeMGTYHJmthPBn+FT9NwGcp56hSAD7EGOMF9T+9VqakgVbPt1nFiG07S6a4Ip
4RUtFSuO6J6nuL7/ZMviGpBtnzbCt2Ijiu7vmJ0dZ6o7fiG8QDU9e7jP6YzN1r63T/PgBgjlJyd8
uxs3kyyZzpvwDIf4lSvG/jmfeE6Gy7V/D2VHk6uRzBJyigG8bTCpGTW6E9xZj8jVqwf8A6lO+Bwo
RF01gF/ctz0sHp5jsON7FrxVPLKQZH36otwpykVFVirvQaPT0GunjIjZ+huMsrcu1Wyy8ibEfMw+
g87IMxf6qhUEgAjBkD1TEzG7qd/GwxeP0mTz6x7XuudqQiTFGvCKHhkuGaApnoWh743xKsKyEG3X
wO848Rmpaq7SVafuhKMrzMhhvkmuVjJGbRysgMLLQYLiLF3UcIKnAT3A2NqQUELtxJkojEVmLQPc
962/fMtJ4bjoii1vEm0Jq70iFSRSyKxXdejwpLEL4m+UYIVnu2d5bsXb1BBO9mQvuUMvultCaidS
sJVzbNIi1RDj2wymD+xGo02cBzjpyfDw024l71m5b/EC+7eQe7u1QgvmqwKEGnbcC4wdeErKQyhe
pB3sjHbRExzbmT7KAj3X3wFPmm9hX+Sz24kP50PmzPH9xNDaSQadjUBvNXQ1NGk3SsRFW7XC0cmn
DubL3SUYXp3TeB287P74zMzJ/61smUs9Conre80WyPMELpXnVxfow3fZE4PR2HOLscNmXEQqpFq9
ccb+nmyZ7lh6SafkH/LCEqZ7oOftXTrfAo+RYh5nArVhc0QwKorwoFWS1cfgzMMnikFdbXGeMfS1
E+mUYLlKTMW2hmnMWmvqvjH+crr6lNX5cPtgFf9r2Q7IOgp9VtGFO72VqnDL8nSx4rF07lX+fjNp
dK0Jp23LeihzsEbSYHEhB19X84tT89LmfcZQzDlA6mdkvwp6RAQsdRH4je7YrFFyLFPsUwhElUM4
OCaMjgIEhnqtKygXiE2zIbF5pV6PCEpkJ9bjpWEWOHHF3WcAUqjI47ZRX/1dbAj/Z8KKx/YgKg67
/4UBRxUuq+HoNPOvF2AHPA0V0Qo4RKZ9TDQyRUzdQS9ULN+Dq69Q5ZqLfUiQE0TQRj+2fK0XHFay
oMpNoIEFyDgrKjQUqRX142/aRAj9uvNsf8Jew5h9cMb3Jl4dG9q311+V5muNjLetKlg9UojyU7Q2
GCIFHkgq8HJn/qRvPBKSd4taLpx3UhzoGUiZuCVu2yXDRc/5bV8CMqsCOcgMVoAwsvCDwtiuebMQ
QGI508LwJcPpPZXOgH3vEWdMFBM1BnV47IYV/OXWgdXhQ0QvFWsKImN0tL18/Mv7AG3D1Ev8qRBz
OZR0LEjnZfpCfj0yM+aoaIQ3mD3ew6dCfIucXJW7eXx7FIiNFjRzVYW+3zI8/EpFc3o937aeXdiG
dAI2P4JUBQQfuceIxi+6ricHBXZWcq5Qg7x/FwVWD3cIK2s+QOH8ND0mFNQ1JcmyhDlXce+T6cHQ
JSzRfX7sOcWlx1ra9Ftwj+VSWF8rwO8M0Js0saHiJMs60N0WBIQc62XLtLO+LKZUy8KrDXIe62gF
SzA0bu7rqU/q5bwnphPe37HGNnoDZvdBWsDCmQH+ppzvp2rVdNQwQQMMcTdjERW74WrP8EGv1j+U
xThpLEleEnG27S3OYv+dFKA1oOEhtbjh4QpbqitsQXUDnwW2jxq+xef9OGaEFFnbtOIxoQDHA7jd
d7FhwxfSH6zIoETagcZc9kobM/KAC+pD0ntz19t0athjhKwFI1MCM5OCK8pJyg5BTi/izG3PaP1k
3oy1NS1B+USQIS40Z4VxxLMDC/+mHYKhqNdtRpJPkEJ61MJwgefZuEKXu3BxgeorKD13JZAWXiBq
GwUQQJgk/vxn1q/DOiPBEHkiQbcgmr9TIOhF56BrFiA3Hc4uXONbMqNa6e1+vWwAfsYzxK1ocdxN
McBC1QGwbNKLcJBAqAzXtwA+b3O8j1Dpmd7uwf81eTHO/pYchfayklcnabIUhM55oZVHGbwsFbHG
9d/jeWYPWyLDzeoSojXZud1DkXOeg9F1yreIhicBYKQqlYinbARQ9Ux8rEW/dKSiN8oAMXVWgb6M
mQ/NxzRQRKJO3z2JlUs+5TmZVxIz8n9HTDeG/B0PE2CkSSExDogqcBI2oTKtWvMd/A7AfjJCDDII
TWuG55mN2+w5zI+u/YazpjMetCp2dM5bXkZmsC/RMpR5JDD0h6msQIyuDBDrk/SsGL6awi28KxEl
WAXpxqT9ME04U8l+iwlgN/OmJhG/cOvjZF/dOEt68nsYz/kpalQCi0wytKYTbOvN9MUIJf/BxF4c
yN3pxNaH2unTGSAeXQpHgmvMHkms7enWlvAIG4ydFtp6SFHlOTxH/ULxHqJHLkn2RLLs7HnGIK9m
4SsiChtifFAi4sNkPO2vU6gQgdtkmLtGSPZf1xu1/lSZz7NkRhbzNxMlOXywJV7f9of3vrLItBFV
b9jH0R0rcax+/aAmI5gBdgyTquX7ZfQZhahoNlsJ7uEbZp/nU2p0m92rRPd0tZ3V4psBpEAzuh0t
kR02zGSUzXwsBqyRVfUsPIS2A+Cx8fYoNw2B7Q5XLwjc6s7vlrbm9Z1VBr0/ErSfY0w71n2sSJ6K
veomeyjlksD7Rn7ELJ5iSiAPB8pZPRa0nvrh0R3WWsCmJFwfsW3O06Kbs4luK2uf3yL/DXGQzqId
VfseqoPD5ZAaADK/k9j/PGqNWGWYsjlaPjafMctSlul65xEceab7JiWTBXG/Q/fs9yVQ/28vV7a/
CvDUkJ36O26MCM2De1JI97RaByGbsm4qsaz9veoXRUlmpubAadES6ObfCobQye1sRhf242d86H3m
dDWPLFTb/3v4Un/ty8SHIL4Oqt2znyYmO6C8VjbB/Gp/ce3Wk3ijhdMIkho/4xmx9klkYVeGA7fZ
pRw58LTrk7lmLMrm4IeZ7kd8sS6R5JBtJYWweP8yHuLXnDZ0+wV/HCvJKJ9r/EAFGy+gQ/Ws5vbj
AG9GRr+ouduyV6bXksIUbdaLy/TsSvZLiFfkmey8h+beGvRdB4WXcHu/AXbdrM6zED464Gpuad34
NW/3hPfU4ftAJ0W8t8IHbkuI3kS6I7G/GUnXl0LeizJbUbi5wW3AEMrQgR4HE79vATfoOk6fZhZL
QEdZi8D0f1/chzRJ1+sQQLA84QgJvM0tY9R1H1rADA853qD4lCicFYWbmD35VfvOl3CkFVXTpdPd
BCjoxtAF9cgj6tr1Nc6bsrT61KSafIFr45777OikWSA4cLJT4i0yIIRZDZes18qLCIFk9IJMJjqk
T/pKr4xX56m/kIcfRUNL4z3exgzylmCUpUL6JSccMoVLxrkaNrVgsP1yQ8FDmFyVuUCuNZnrVEnn
h3NUR0E9jIEb6SSM0re98OQ3x2mKy9kM06uLX7tw7J4dVa5T1qMfRJvGe/QfwynWJsIiD25C4cf0
puXUSedfDsmLqDR6QhigGBGGsHqUjXjbr/TfWnDaPnSkydV+JkPGB8p1CD9gjFm6Cf+xCZcxT9bS
dyR1lJwdM70JQpTOryd5tgqcEfysMSwWGhA0ZD5aq+e/AjXJJsRLDKx/GrpeHkqlAEi3RbLZczVd
X3wPQXAUNhr49Dm9eHcub2DZrzOpjoGY2KvAKKHKA9hdPP7a1BwQA/+GbE5mzgweyVrUnB4i+Qra
vLSHnZGDGuLYRD2ZkZrM073aYH+ROgw4KvC77ZWRQKohbQb+fN30U/eV4d1gPqUocpWJ8WgLrd+A
cfSgFwEjREVrI1g92aGs4SLW6xRTEkJ4/RnPI5LxV6JDjEQuMbUBXjQkU/4FD34wSbtgS0fZuHEg
tfzNZo++cQ34iWXuCXOU3H0MwyqIoHL3N0iz0VNCgfJLkPcEVTVaUZI8yf1siEdcVLtCbxlBgoHm
w4vlJ7guolA1cz3qs0YFDbNKchGedtfiUhg5EFIoepy1kRZG//6LUpKqkqK+6gstGcPkdK0cLmrh
TsHxk0ra+hA8/pCgjd0HSrtwJrKGAPI9hOD4UFxB4Mdrs/Qqfb3YxFAI3KvaJsLunF5ec6l32Zsv
przppKR753GcponnML8nqv45Dwi1fapnT0uqHNKYY2IIXU9B3ANAz8wPwg3GGwQo5luXWPXHhkmD
rjMFoo3kPrHQ+PIdpv96RyNBsyU3eWZiKqz20UVk6wOZDzyZXrwbTSL5FYNyZeHboVpzV+S4IbPM
rqxu5910r0C4hEbGe0vetbsd0u3F8ps+zTcsQAaRGib0WG5GavICBsYJrQ50BhNWjGUqqaspUeQj
wCOxKfPKAhreNQN41SYTYzSYUl8oVYwkXxZ/IpBREAo+YOOHilYFpPk3LHRL1X18D9cnkPBrrOLr
06sMB5RXp+kKg/suDkC0jNxCt7WK0YIrWXjwOvVDU1Mhopx1sGLaEEvE8js8Ggnn2dvkun30cLQ6
+JZKI0fYCc6bNv0ThnSd+rTCaJCycFHJPUk8NucfqrHKh91Wznwx/meGZRzjbeyQf1it81QG+eHA
75qA/9vzMpDKiWihCNekTOIyeUJXtwDQAgBPqKJNN+l5lvzS3FFXda6AjvQX7UVK6SlkDWbNwDlZ
pXVDeO28TE+AdjoR0QBBIj6tEsjv7UIsig5oclLKLMGWOwBhZGUHePGYOWq7g4BIC+iUzx3qSPFA
g8D3jUPrKJdxdYoFlDRjTEBQ0909cnTCqJDSj4grImMApjs8POCmB8V/Ylx8gECxz6v3rEOoc+vP
fFhONYcAMSAygv6WcECbBej/WtShwkp8gdvenaCoT1quYsFFdYPTcDzGpUt/bO6Cd/uQlaeyYj4K
uXKtrIZddHYX8iwpw+WHhO7Pap8Eh/6OaCju5yuyZ4x1mmWbWPThiPXMgjkbXIPu4m+jaCYZn08U
YPQE8dQNkqzGdzf6M6MzlYQHJ3byhRjULNofAhKJgNuomQW57RGJbtv650ppM1gW65FesyGTqTV2
tda05aLPMAJMmrX2+A7mrmnfrPuY+f0T6K2WDL8uRbMTuDSP0q1caeDT5O+5jzhWXsuTO7pVvX5q
S8+nJamRo7NrZvvEVaBEiKjJG0AIiA/gAa0fZMUH9eU7sUHT8hhaYYBBn5z0aZUoeR7cbqdRonQF
KHfQV7P7HoV2bzq5jiEEZwbSkSQvWhCBX54+vBnKrkZg0XgcZXPAk2Pi2QxZz87wGODVWjs/qq6J
rysLnPqsU4JA7Tpfwy5A2/vaU1EueOYiFedYpz+C2egqiqhwzOvb6biMMhWwqU/gW7p7cmqTcNyr
WDKiflWWEE4ghW64+5rKKrxwvKBgNmpB8/GU6Ymcqi4cxqkH7095Eg2SgCnig4lSrPGWldX+7kCk
7e/Z2qlFHt/nNKi5fAAR3KUiHkfpSBOu9b1FGb56mRDHMWpsRwDa6BYawXmTJmHgiiBT2OYCtRRw
0jab6Qcj+H5Fsq5wb5lQ119LVYdrr1Ubugy2I8ele/fgxYfyTqljDwW9eJOG0wuxjOUWkGmejbYI
kSPmVMTA54q7URiHWtZTM4QmulDsEU0utFNpczLhgvW5wWsgwD1E9qo5/+pH7GY38fD0fs+yIqtM
zhd8huPh8VAbYkYnsMEMYyUelMgYRi6rrLktisWX7m8V5lhkAHebkbRPQDH9dJ7ZuFy6nf2msCnz
oP4OKpWMzY+QwvDzWpKSQJZrrOUboLCob+rAcHlxM7DnTjmBshAwhOm9ZsAQm3fPiW/4DYE0KwvN
b9lWAs3zN9tQI+Q+UWI4LYk2IewfwX/+eQ2UCg1U8Qz5XBSS+RQzpa1DS2k38BtoOaev02QLa2ag
i0ImFdimoeqlAS511WLtb+GjT/wj+yqjSKzi0JVBFc4AWwy0aaDDsEDLsbMeUstkiaImCjLI2+My
qwc4h8OWROMHKMqorF7Iossjneyaf/hBG47neRIgY+E2Jf0uVHS4XATUEzbFzm8T/8Z2JSihVh6s
SahbhaCIcH8o866Z7W4q+3x/bo4LO0Mqo4HhuX2LbZpDsy8Uhlckhq2RaGo4mXlj1h15RsTuYzWT
zhq9tvkdjuSu4h0wgOOTDR3oowjDpk8Rm6SeoXZ3fYOMB94+6AjBAyYRSq2Ut1/jOrYtf2N4mb3z
ajoSyAkMXYHajSX7hNtHS7fV3nljZW70FVXRxuLWARCfpjEdbPl/vzwR0v3Vs8W78KxMcqV5Umo1
wGjBXR0JBXA7V1o5kd47ZD/wK1MLxjlPmRhTQYLw6M6EMU35xVVw7UVw4PyPtYHC8zsESqg0hrxe
o6OVTQSBmV5NSavZ0d4BErbC1C9NLW1kU7rIIxHXt8rPs6srs7aoRSSr+Bw3vSbKsG9t98eeyhvZ
C7AvPKmpDtBU2/HvpTI1Vy0YX52yrQgXX15T6TAwEdzeSEtB5bDK2ZjrEeZSKlzJ3s99d8DdaHzs
YyDunbuOEjwErmCebgEZ5PlMPJ50spJIkOGzHvxP+NrVq/WQSARQODZIS/yFO4Fy8jujMLNR9IXF
UtLbt77B5yMSKOWRyWwmJqH6DDSBi5JWs0KUrhF3iYR6AYGVfsorYrdvy0jorOPzo+sEwl30EH2z
m5oS+WNxUDYJOS/xRHrvSfEB5SlCJVXCqOmsv4d6pbrEhAFerHLATeHkQ6nrijhBr6A6aClIf8ch
ROFoyb1zvrclalv2PVING7rLPZMuhJB9gS2n0APAlOMx+W5tb5HYp4lMx6v+4QJlBAMHQ0kUzVKy
2GV/bG3E4W2k4fDDXhi6sElHVdtc1gN0qMVGcJgxXyPt7kIDPGRkcB3yUQLOE2Yu7uDO7/0Ds/Zr
HLrChpB+17+b7oRIhB5d4ESbzNc+RIMbNdRXfgRtC42Op2m7xK8mDHG2aH7ncB+lLiIt/FvmgoIU
MX0f91z/OyJnhNjc6Gq5BKxzBYSZwNKaP1f+EVEEcyJQRNSrH2wzTZsjrKIdR7zU17w+RnqRvS5C
Ppk3BIu4Tm0LoUOq/CtneqiaUgZRH1eLUUl9pU8guBIv1j/XEmRAAI6R5RG19oS7zWtK1u0TKG9f
cVEFPspzEhgoCw0owpGG5Kpy1jJYlOaXbcsf3wuDNjPS8OJOVXi7/jxVbtItvnBLt/SOY26sFnB+
lPfUHAYtChQTW33wpuSqp5V6Q2T9WEmB1j9rDo6pt1ZF9AgcB+iw02Y9iob0gm8rjwdLPfJUPdPd
xAoAeEQ0giKjQjBoyLuvoWDw5MuPKIP/dqyI0oVysEnySWLzWQv9gIyNb2jcNf91gUYEWR0OeMcp
9Q0VqoU3JU3kgwKbDPs5dFBxEGIZT/JRCNzpj/4IQgFykLlDO4bRb7nXfnhhque1YX3QsxDbHX+x
b0Ep7xMA2XWBkQEOTIh4cDigXv/09ly0LlNQmxof2FTvMIow6TbF6ZfM9YNdSwQ+vQFYfrNesMUz
WEw5F1epG6a7aC01yS1lMYvrhWNt93irWfhUlS0G7d8fsLqk5fhx7KQDYrfuXM0Ac7HQqWLTdfss
GPPuHl+vtCMbLDuEjhnaO4LdSN8E0d6OaK9iVulS+z/11vwWNHMkIxvdMBbfxXLBbz0CW2Da7DuF
9Axmi6ykYUfAXIKARL9YVKdPr8m5ufoB7b6f/4fos2Ehz3iVgYZnv2BpsEfWLyiRQ/6HCjXD2hwz
61lEfApZP/Cr+hBEIzUMf9OwsdZ8o0qarTXQHVUpCTkqNZYPrYb8y5Aqx61+Vw07Q5+9Sl8MYv/j
yxQJnae5RRJKIIxQSnULWqLhWUjM+ltwUNFy2NRyBf7sIATXpWu9OMabcPyQYoc59jK/pTrLmqd4
bDHO4FD4o9Kd+K+gONOFg3B8O0S12YDw8S16ARIXDdKHwX611rrlyEsQl5//kXQ4/oReNahiC4Gf
Y1tYTDpiCN9O5P+kvrq14IURdy+toPOsK7o0q4NQI6B0AczUKNXJ+lccp2HhWhk53SiFGiZvy0SU
Dt0zuHmKMXk4Qn40/13rISDeJU57mpswjTR+x7XLf07F3735rd3FnfSTEmCeniyGgmhdrIyfR87U
Gvf2ikkpZhGkQl2IyOWHymzP1MWnywFsbP6P0EMP+zGsk8XZOfcNdNP6lKqNnvNvs6v5q2dgKIMa
XY6NB/HW+7KFY/vbEKsG2V+CHMxplHQGd3NjswT/OxyatJangKFdipxvEry09q936+4kYQI/zM6x
Qv+guUYEOBIQ0MJzH5KaWcbSw2wtEtELNO163G/Hm5ocsM2EFshJigMOJ6NEQUQDEw+G9OBwLWS3
n/Cah64pYjzZcI13gX2FjdKaJFGI30lbIciANjmdLGyuOdd3Vq3tvqLNE41Q1WSnTlY4LjHYyXLF
lWeUlMfM0IMVZCZK2ba+Red1AJ0lvtyO0tPepM22N/pxBn9q7darDS7Mt632xHtW5en5DcXnPCVA
tggYH07iEWHkfwFeisvFt1XyV4qTA0HDY/HoDcokQL9LjHueFn/YJXGUJA51Q5jxWHovqmSb/0Ds
+UfibmMH5S+paOoYKYgltMFWMnTmOcY4u9NljYi4R84h4sFwWkX9eZI4tJds/ABWGvPolZ0K/yxA
nH6SuzLzgoe+bdvMvJ0RZtChdxnsDRNqsG3djB9/Nv7oFhrOgMQLCPuTnbLNngm8R08GYVuNkKpI
Y/5SrpSBJ/gOPYuCsARbh0uDB3WSr23sFh22s5b0KhmDJEYeMWuIdn6R5s5kp2Yl+WM1Gqt+sKCO
aa8YH8qc1lkFEGdLsZoGcMkoAqt7NIzi/ffTdYsiC7qaZwS9ejYwTYFEdxSz0wgBPNH8Fli+jRng
PPPap9SYz+rOXi97JhxJ4saAR7fsTGhPq938GxaaTBeXGaqSYjsL3LkQBpruBkBVkq+ARqC21/jO
gUKYsOROVMs1hg8TUJZv+XaSA3LR58ZZqCYE7wXB5pDj7WUKnoBD3LxCIoIJGpuD4EDni1B6qAez
zb35aOV25mLK8nSwx0taiK4af4LSfaAsekl51D72iMG8iRf0RwWU6g93Cj8lvx1r2MPlQ93X4Av9
6+HS8SSpm6QyLVNoIXGiaCzGY5ONR3ezEkV5CWDIdcgXps0mjLnx/kBDd0IrNA/2s47AMUXuFRnL
QdnI8kuE39fbQQ7SlslKnAY/UUhuUgH9rxeM8r/b9IvvVBkP5zFUsV2mw060I9mEFePQ1qxaLh/i
S2184FME/kwB+2UUcoKpa6r14rrfz0ae7NiIzXrPSmPnXOdq85ZOhWaMHerJUKsackb7ZIXQWjjX
Cx5FwvKTfX6Iwp0UdKN5ihEgodrDIFq8BZ5kcEsMpUqT0F8BZ2Ck6uy0AZMvDuKvChwA8+sTpUjn
OszSlrOEQv4jOqIOjaL5AfwYhkIoJzkyKOoRS0sN0czbRcJ75AOIjcrbBxHuDJWTbS2HrwW7n3ji
/8+oZuURa4AmnI1zRBK4YwlEsvJ04zWN3DNGoEInHNTBYzA0Wg+/3z3aAr5MbVR3heWNIH3XDwVn
jZNlfTADt68NCW0kO8wy0vnR3ZaQPiWVeCXjqSQHkvjbNVPBfVuOnzcXM4NinSfykxZ9HIXxnPoO
HkGeylBa2Mq8xYW3MnEM+W450GNQkNQ9n2p6SAWGatyz6BWergGmFzq+gN4cPqWLO21UFO2Cqsb6
ouLzwa4VDq80r7C4Xn1mYqj/pw2eMNAT/y6kvBj0zo7Qi4O+zgAWr51u/2P70Ku2brvEfMr9GXna
IDBtKI7uD5TeyR93hCOaGp6JecYFxWLjN5NLmsoVtWQBYqrY378HHcRSmnTPYEBvmVcOHywZpVrI
qaUsLo4aWfHbmDBNFXgA9hXgSTneaT7Kq32juw3sFIOX0+J31Jp5q8G3SF9t1I1/WqGaFkgPfo7C
TyXKoVquLOYl3/aSt5LemAr7yvf0kyxWEDrSrnlJKowSoji+oNLPPy67wIUghnSIVwQFku+5ZRaw
BuvFmXHqYa5drBJOpcmKZ4MwmPZijlAfflaue9cmOoWQjmPfB8dcpVQSOZZKptcAON5apsEr9mpX
1bYZdZoP4wlFnzepcV62EOEI/hRSCdigDe8M/jNxrppxh7sccxv47t1UBZsP3jBbnrCf4MHTQlMQ
yB6gSPpK4YvF1++N+8mNIRC2ECKqnZUqeu6dSEENs9c0OhDlEwJGidgy4cmrpTJ1P135l/LUFsyU
yshP9QoIou1Xbl+rNsavI5MT/aV7ZLMeMvf+jWK20L7FGAQ9bn/ljyyr8w3k4VJJuotAdA99A1JC
jrcpCohkAN3rFluckRn2PiTCchNe/9vO9NRJWgLLlFrrT53cRX4tg18huK0cOcw+kmc7bJP9EMx7
ZhbPqFaopyAanlLkvAdOGkfvv0D0iLq3x46nRytev/qcyby3MWbLgh1/xvw1yl1dnwfHBfIwRLih
3UUUSYc3EDu3NT3eg2Ate61rSKQHb/e5RobGH3qDVgc77ylAMsAOeLywHj/mggD0BMFc3+9ktnQS
d46VEVSlFWsK1K5igRPiVslpzvkHJfcCATP+FqBLi4t5cvmCk0EovuiUAV/KI2jMfDiiz9/uuwKY
vVCaUKf2kr9nmB5QwcfhKZkT9delgnqQwtjwYcX62sFVtvAsZTjaeJQ/9RYE4xKQICzFiYvQbRRy
WEzTbNEbRJ483G2eQHFs1bDhlFNuTEz1WUXJV8COVIVJJSisKqspptZBcSFB3yiR73uyku1dylnO
IjFq9t55HD2kcmx9PzYNcTAUC8GHHFmUVSkuVUBKYpwynSXmd1UlWCsjwRXt65XSAfWoWQBbQGLJ
QWloTfpQLNWbrSlLywMtfx4knX2jf5vgY0W8OIsvGNJNAntY/nZPJhPD6c8AFk0JeoyE9vg5oLdz
oTNy+IBu+TTqgrFv7vm+pcEtsO8jaFNJrkIGT4VuT78/aIFWe9YxeMFpZCyGXrGas6OUUM6egxmX
Xx75yq/eWLjnhVXLG8ajYhoXPLNAgrDOc3u7w+1fxUjETPu2d2jKq4yULGw5g6Ir5lAeB6shZpKY
Xu42ffgvf0VZYuIuWuoqgS4lqM4mdeBi1drK7KdipRTDnz8t5DJa72EhQUugWtaErr61HSFsfEab
eslcbX7d2JRyZ1llQg2jk4CtQf5SN+M/FulEmD4gPfmpQPndB5w5gsm6Xx07/AyCme7Aohty8ZEB
edA8z1j26lyuP/UrUwLKZ0fW83VIgL6FVRZXwtouHrHMIBUlZhQOWznrbXagnGGd5bmMp5tdwQgZ
jrB0QzxPTOYQjDv3Edt0kvZMga93oZYll1js1M5rebpmKO8kBoqhOflDYpgBPOrBaNqzyb5TiKOb
Xq3QNiHWo4Yar2bkw4MM56VNWXbhIRI7DtjXtJGKjdzz6kInNLIdEj/PoOFsZ2gmc+WVEyuh96m4
CyVQSzNJXaxPwPx+1CXiyWydOAQjbcC48bKzRb+MocHvnVmj5RqbGQ8a4aTcefNb/LRWFBiZcx+l
oqr8e63PFMu8G3LVbrHIYLxNSJPqQmup/eQzpKq+JJ+hMe8LuK434wvg9MJE/klKE0jkx2n/aw44
j4yBwMhYhSw6a+Dflt0ENQamq8sDxCqxBfazeYb/YcBih930GIT/umF7b/XUd9znR1gwOsFpIvOE
HaL9mGnlqDAYGqWPjMk0i3eluABpQSFF8G1fWwzIC8E8cnCPAAO1HUoAhAKeTmV1Z3dfBYKRF6qZ
Mlmwq0p7vivOGTFf7TayTUAH5choYmO2Wr3KzN8XbMhXZaqYRCYtJDPuCe6L5js7zBWdHhFvjHCx
wFRxI77JbcCe36tVpuMDSnnVweoCKmR1j07L88dLmhNyJhxRo9xRn60GcjR3NB78lNkRyeUQcPOC
YOUaYss+SBQJbu99+lL5Ih65EPx78ybA5Tn+YneOk1ydrIDrVPUfLgawvWrWWI1YBZpLbc1psINY
Q3DqOYsSih9cBXb0rzClR7cJnnGO6YgBFS7+eeaJbPGPaRWq0M4+Sca7WjBkKgTSrI/w2SOYpub9
Ar5sHMo3wsPotLfXi9Hl51RQEeFfxbgNfsZmEPWng0ggF+zBam2iobuNCHiQS+loxMz/PgG1r4bf
aGyavhrXIsLi2y857AvlKJ6szRH+LscEy4qmHMvzPlCN5ad3GSmD1ujqZjkKLJ0wVU4aRK66w3WN
qrmUIufhK8VQyk1V4YhClIvFh0pVySx5GGDrDCekrYSHWYHqzO7+ayZaktpVF1OZ2CWHsvo8CQg/
ew3Bkmmsr1kYhFH2svoOhBO/fJ+jq/wayhuLXlIsRQVXtRYQ3E0qAmyOSfTdyoNpgzDJOHcsiN3l
MZ6voGLJ+/S5Lq2ikgTQLLJKR2pFccEA50A9swAFpS7cjRgErovH+fdM8UOB2MUhinRImTGjBaBg
Y46F+sJ1q/QsYoNhsgIn+S2Zbk7pw4rFEEPzX5QVtYvm6svegj4hmiX05Y9xwZOByEJkibUqdgWd
VHB1UZpt8PKJFwvX7Kj8Tq/6t4CplzqKr5WI8+CgZqtesXJVMjWFhr/dd6xTCPSnXNhLIf0zYo6L
fz12e4aORfttLXuC217v+XChsSC9Sz1F9lU0R2xibzrM1E16bQyHrafypWKqrc0EHkxv4Qa6WTr0
fVc3vcgBUzxT30c9kXfA6HqjB+OGLTXLWoGjXAEWwcioDwgzZN4yCk8u28HxoNAzJRQNQc8PB4EE
xplaPm4YNSXm9pgo7BPD6NzDwnajv0mE57aRbvCAeRSaWtlvQyBrDSaMPHXW7b/xYZPVbpkhYn26
/LYX95h4+59ndOi+ifb1TNBcXSXhkrG/SptXKXdjeKAGC1B6SjvPeAKva5S0lye112lOKYQ7595k
E929jjq1Iq6TWHVdOueDsTxdja9JwNWDcABsSpYQ5WudRvfoJGhQXePhyspP+yMdlEzQeehkApmz
/3ATdxq0AgUnjfv2m8KOHfWodZFZwJUJfvnOkZ5T8pSSwWagWkdplceRIEYS0eL5+U6k8E8LsA9h
g6LZdQilticzBmf1+Ui3VBKM8job+dQFWYGCEbKQ4V7Fp1MivcXJIMCQnyB6XMQD7gghSW0eYcUl
jQQtIeKzaxe80Hn0rNW0CtxqiTISKakFF4IIZwfyePVlDASf6zEoAsCNqDO1qLenfvYMk4RL52jM
GDRQVR7efNPKjdUNOdcFg5qHydaZ1UVzErHXeHpKgc1ChQY9MZ49eZeyIlQaC5qFfLq9LIJopD8f
GU3jDSCN9wdOnqWfrJv2xjyuLkt/M0/EdKAhvK5fc4bmzEO55+gBqbF7uM7drCCR9goOMuzMj43o
czEF/M5nOwUT6us4EptPT48yn0FxvO0nQNJFEkIj96fEiYn9nVWEUD1ABQeWuN2nAQPx09KFL2Tl
IFaMsiTeFOTdQS8wIigr52edC8bjZpgAr9aqiOT0Syb9bpjuOO8XgPcLyuNr6BFeXX4CJjK/q/83
pdYO0EucWtB8l7/C7/Tw5yxrL+oLsiwsPm7hFTvwRbgHZpBQBz2GTfoF3qfhMz1Vrqpu3aW/LMRs
mDm2zHRhmCCyfkgc3EY3fVcxw1TerxMJa0Lbe+MZBda8vz2xa7bFPCC0BQvoGldXP+1kYWi9ys82
8EmY+JKT6cuZfuuHk88pGIEYcMNT8UCPpR3PJ+p2+QP1jv1eC9cGOUZOX6aDi9mDkEQk7JM44eEl
D/q2dgvkKfqk6NIoXjRHtKfa0tK7UdkYGYIoqPZSObuSgbT24VIUkHMXP9dCpVaTMedJgKR+3GeA
EB/SD2SROd9OnVPBguv+DsaTKsjV+IPUmR6I1vtSk64G1mxaaQ/JE52X7TgQTIzYAf+bSh1K/c7s
51ZEi1/XmLGYwCUcISx1U1tD3QoBjH51x3Hq9Le16xQ7zzYtOEkrPBPjNfeMS8YyORVbndA803TZ
zsiffCwE95FexFFHjlgQsDCbjY4RztTlFpvhFow0I97ltYu0yn1/q5wA21/3JrCkWqHAsUSSL3XM
rJdbXshJ8SV6gHtEsIYqan9kd1kKIWBEK8/iHzL8/3pnQWl0J9G+ds15FeCRM6o2bC2nocmj+bce
CxpLxnvUWElIDeH1kGup39tYb85ZJjO0u9P5X9dHMrhtxldcqyoB2bsnAcq7gAAX/fJvBCw2kymd
H6hIG66oJEvNBunlIgG66NMuIhiW4OokZNEWO/UW84hqL4ZUEtl76R8io/6PYPpffBzvRE0G44w9
ocTmfopIEzZvr8gYUk3qQB6nQ892B7+LQHsuAry9b6/8ZtJsXnpOXUwbF3AM3wX0SpljikXSBhpI
FQbBzwnJrt9AlrrEuqji0hkv7io4FZDGGpVuR3P0ckcF0tGHLeqabW+AwqBbmp6akVRkpELMXDMz
OmgZ9uqPDiNIu6mykQ2RHCRR1qTl6uTXcF5jfO/FV4hSfg8sil1Opz4/U71rEKiEbVlrg4BhG4zj
yueGEqYSzPsBIHPUe53fiHlcGk6ih7yvLya7mp7amJTb4BHuroRivwvr73C9+aiz+CUCAmemHhuh
U1ts1WqDB7MViJfdC+e523RMJqOiINEttKAtMouB58EPBf9mgdObL7grquCw6v7lcvjooIMOcEtT
t7fYlcByzCJLkbLFnXdBsko4FPO0hEhUdvXG5HdS2gj2b+HAR8ejoeiki4mabgOhODkGfXuu+WCA
1mcBvEInPSc/9ZUJjYBUG82QU21QZjXwlEsNz6WJFvcRh/KvbRV8Fw2g1UCHcf9A4BgKGhq7hx/U
0c/PEuR1x2uSdpNyrMSA/XhIc0h/MbAYcps6xpFVxCVfqXUxWy/OjWYrzzF2rc9sx7L4tdibvnfO
+C4XSc2miN30JD5YEmCykRzZcsemsRYr2jageZqjdLf6BmvZ7tltbt2vIaJ3kmEAn3WvXbWwRiuk
u2xRXKmBLJE7mFKeq1UCCESw/owRjvMiNAqHVFSyBjepvbWKNUHBMhlVflb0xY7ib6i1xh8Id6tB
xbODjYzW1lQfoKuR+DfG9XTNNvVBD0cgmT84A+ucJtAsccsPM3QMuLAitnBgASxX0Sjbyx4WfpFA
Ygqv4dMAFT3vAwQGqfAv4pDvw1w7TVZ20XhTHkpN2fzc7H1A8ZqNfD6hNLjrmsdmytzao/R0sow9
itUy8C2MsC7qjHR5hm3uuE856b0Df9H4AdkqbIUrq+59xydi/w5ltQ4lUIkFVIRCTQKC6fWjYZQp
9JC0UkgY+r0DqjClsPjOtS/OWdTMh87xSZsBK/oL8cCRQRF+vvkl6s8XwmIJn9q0FZm98kVQuJDz
IJwTlHLQWRvy2V7McwVR0OOHztsjIOf+der1S4//TgCeObb5fghcB6F+A/V5OyfuIkbkLg7lu978
BKpBHgWGz1k3yj8XxBcn6JF8WTdtfwHIXzZ/MDQHhRYiWW77UuuNeshmB0bXL0NiaeSdrHc2TCBU
M9tBPRlCVeDNMe5ft4K2mEKn9UOvW/WKOL0WIJZDr3xdg65MlAQAUjCtPEa+UtdAs3iHyB4SjDbu
l+8qKv0xyoQJbheXRkVVoL0l04Dx2nkNk9lmlxCkadoTSyZD3a9im1o9sUeiFYisnqVDw65tbgnX
okXFvIRj7Mg6LS22z9o47tVdlo2meatdn70M7vAZJkaH7BW1RqaupLTX5QKwO3Vk8en+qYLsWRVj
o5xrcWyEZ7SXSFDFyLc/WMnNsrYktIiv+A9a0XjDxhiIcAXxqlH+RerhxyJlkhMEuuI+g1FdZCF1
S2A+ZVqiFCD6IMci2GPhtbfmz9ajlt9B4b523BOF/ZbUmiq3uHRzco/XTL1YH35Sf7OaEPSRkUgH
OmVgabSToO9aqgWRtmwAHJEgt3NolVnBgR5AoP5l9d2kogSMEpAhSFFbn1WmftE87p7zZhGihyoC
MT88jOT3s5+8UWwRfl06iizDsRdeHP+OF4UPYbjEAxAqFjQZ1kmCRG7Ql/IbC8KXpCz/pGEnT7C0
XJjsYD4CLs7V4H67l5i1124c15CVhJeQTQdCeMNEmuGdJy1WHJOX9pPDVGt/BNqyYjwbt4MH8P7G
ZQetaUity5wZTS0kx435nk0reycjarwQSvFgCznaKSLOwDnyO5V2W7wPfVVPUIRC4V094sfl0Fjh
yfpi6KOTBPmSrCiKrGU+a5oOFpa+4qircrVVf1QBZy08RWsNNX3JX3vohqrB3NWKvyfcsXzkOTNh
7D0GbtWws+Qp1xDwojzAO0/G5SAW4j4Ls9AknVJGw7DznXer+WzXwd0/9ngNJEkti4UxulPAnOs5
4R/BK5IEBUbs882WDNMGb/uV5mJ5oZUs2amZOTJCzVhRSl/zbpfHFERGIclOnKA9XRUlfkFSKO+4
1HjBKWB+Yb/txwdieo62oR1VqrpyeLOaxwsK5fEsiq60Dib5DTsBP+vNR1Ji6sAzK42RCYLDjOd2
Vy8nGvFOJiWAv4tpp83jI8xpQ7j2Cg2ALS9ybsOSJRF0hid1Zl1Y6yaaJKlT8HPblctTjwOegzaR
qePsdqAz4m2bVLb/xxsDOU9ficFeyBAanqxYTDB5e5D0McGrYYn8xM9/ZOK93+zHdseOl5cUVb7x
S6ftW3cD6+cT60JKwg9+T8Vx7ccU0lHAJWPdwj5FQtCU4fc4360ADiZEMBB3+fseaMa81z005JcN
3aRvL3nRtMoaHsoHh66+4kfLa72XQBqIoCrv/AtHbLlbSh/C0vyJyI2IiP/GCNj46XXRd2+Jy5mM
GhUr2SUqagdFW0GtmzcZ952ltm5mnRWEMYqnRy/Yd/KD7nKp4j2SDYbsOujsm9L3XlZRONSmhoth
DNvjTnP7ykYTu29BVHVrhmtjLKsjjNgTcnl21r3CmZHTVoP3BbPHXMbgSNcbhTp4Ck17vMvfrRgN
zLjj0Fhv/zkPtIfV5r2WGhyWRwzDZXwvs5mam7g0Ox0yC8yOP/aGlH8k9D+G/6+7ifP5QSKSkdx7
ZDyZSP5kW/Z8Tntp++u+JgASWsjHF5CrHZZpDc6D4TLvSPp77hZrnZtXkgH9H4gSZ3viEOLVxXPD
7OVDUBTN5/s1q1lgCZRcMZnvuCB6DKQLyTIh1N2lNPR8KuDsZH1hLn+xOJwCJbnghbLYVW5fcb7Q
v6f/qh7Lr6NaFPLh/KaLUN3buM17pe4V6pKJRKhXYPkz6PT0blqybbM1RtYPykmMQG5oU7jrAwic
gtKo4CLQlP+OmGYVDy5D2c8PiT3x4kcMfhWswzYdhkfC+OM84VYju0FuxIp9Sk3PQuscl9MzZ/RR
MmA5dMzu1SvK3HLjrYFVHLfc4LPPsMAYpwEj3tIj5g5wn5UmkORpguzfLKxcEf6xWOEf2HPg6j5z
j3OtZmvGKxY6b1v0jny2YIAHSuguZpAdTSg9WGfeCIP2PPHoR/9pckGLIj/6rbHuha2gfMm5drS3
v5Sd4Fdl+km+Rz1Sd+kyZHhgrDMc7TevmG+NDNQwp/xpx7EDIoR4k/dVHHnC7rhg0nWEPrCDtMTj
pssT0Js+tB+vuPDGTlobsA/8yXQ/ZjfdS7TwPE9/OBrZFF1MNmpJa6tTSVELKxa/gyratqOeaYGW
LKQ/6oVrkOgq/RV8PFN8iMuoiZV0//C1ovkvAuiv3vdxxPcGVOf9Ez0Sa7OVy0ALP06wZ1G27/Nq
DspIVkjZxdY1MhpjJs0/gKtdRt9l/5AyN+rwYbYD2znn+vRbWQ1dV0pSGq4Qrbvpx+a8Xn3Ovjpo
Fi6vWr6yx+qfzKTQiNoGFb72UH3py+DHr2Z8fZhMatiPNDeZIcbjxcCu1LapkrHL0qBee4sF5BY/
YiC+0kY6buHFygF9g3j6dlGzRNo7RgKLaJe0nctajHNHKUm2EHfmuwJxkPuUbgR5FP3WSK1rEUxv
JRcxGMl3P6EVuOTIYbD9oHupeluvoqdM+8fj1Y+EG7DnKxEc9uouaaUFujOp/7rUFMX9RQqWj0om
VliqbYBTXj3RoqGoe+nlQ+1JEjmqYK0U6t321f7vRIrK1lUX90ZM9bjjxY6w9TqxLdHWI6ClYVqh
rO7fFU7wRAr0+ikZ2QmFD2JufAf73TQUJystRVrDTTSB2FMCn4F0tOePnhVsrHFkfcLYPGhwdSXO
i8K38xZ4h7T6trmPVSXb+k6Q+Dp+Jz+6rkRcQCdUgtMz4vg5e/D6ET3kfkW4BTQoV9JHqgOga0PN
ESjHKFVX0DwZB7TxTe1wisTNsa/bOmO4NBSaD1z2pz4Pv7K3XKRV0z5WN66lpLK1FbPDJZxlZhqx
zN37CtI+ieae1mfrraA0o1/CUTyTstgVJgVPmm1l3vk5vB0TkBovS2tm+43OY5hDWtJ0n9zsRkPv
pjys8xREjnuCXBtmREnbXEIMQ+oIZaYv3kJwJ6NfEYJRojWSamMfaCzxaLyY4KoD1z1awDlm/FdO
s8O0erVN52zPywM9M9z6IvmY0dwRmrifspj7GMUYv515m0Ze2IntBe9fz9ttCyq/UQSNdxmSWLaL
rZoe+DZ8jYgwWWrC+/gZg7WNqipGthlHxdmi01cg7eZmtkn4ZaSqaO30HnJfJ0djstW/WdITsh87
goCZBJB9y/T9g8HXM4cnMQI3T4Nx5Ic2h2fEA65P33ZQZXbJz6VMkPg+SiLayJlVaJlAu+EK9WhH
PIFWupu1Hy9Ap2CeZQxzLYsNkUgwgrO2bRAaglKXPnnONP/4xycSUB6nAlzHwtpSgH5ZXCRtL3v5
IMxXg9zZ1EClegps71QuEg7ghVjwT2gdV3U6BIh2uWtBP4tvQMDkJ8wUbpJDKpX8Dc6OhmVMcj/+
fYvc33c7+W8QCUytW/pG/SjvsswtzJJTmHS2ILXhOon9M7jFFfgs+yA4U24KJPCufmbbne6eyHGs
hkgZZL5bt//SsdHW/JjEE1T5cVGRwB0yffUdrL9aU01KI++Cc2p+LXg9bknQyTKa5l+afRlI+zCU
yKk1dByH+OBVGW8xI5GgGVq2/vTuQFoWeMKWyrKnA1KfPzH1bCf3ZZQiri3sID1stso+5rXKNSIE
9mkbtWNY68ym+5yF3CqMhcgOWZFHs649N5941fP5EdwQnC6qF7uhHyCwUu8UUCr4DKVrNz9RROOm
PIh5sHTMsi4ITW2zX2+jh+n6mGrg9WZWqpF6a8oi7FLjfDR7n1Y5hyDDnUS6YT08vE63q4K3HHMC
DEvFjub3YkcMgptYkUFxjckx8YEy19bS6M19GZ/RsXM6dkLlcIrP4sAEkkFKVXgmdcj5nw/vHpQT
wjTHKvSewIXakgmxiLVn4H5QoyNJYgko2S9vik9EiUTro2DWisqLGZJMC+8ENWuJjaGD9Eg0bKUW
qPPx4no2U5pwalRSdupfDDxAtiBiIfK3FbUa002P9Iemc/Q5tHPt6WwKUf+FqEwu+5YcB/fsz0pt
wTLI+Qm/rYQO4UeN5GLZk/npUS/aizt/dy5Xah3tVVS//K7KN4gtBwPl/OctUupR/N+HU6MRHY23
XIrf8FzJfmw6n9264Hm5wyrqohV28nZJ24mJAaF6OeGJiZwoyCE828vpMDNAt0xcyU2Wt6uvbFis
JWrGaGSmE+1zZQuVsjotRFRB8wE1Yh7NAGfqthvSNtiUpMqPur0NGCM/n0l0I2JRIU5LLdWCciv5
B6zINYdpOWP6PhJkR8/XsrrXGmACZwt5BNSvq65hMK+P5lDq06fdJHtd3FI4WUJZmVdIQ4GcvJsA
tBl9TiWZr7AIWZWAe2cA37bJaWyu2D4CCb7kNMUGIs1C/+UpMZ18u8umcwcbkFoFc1MNwaOZAfJB
+fX7gRktYcnQkzGVAqHo1Dk4PtWHxLjVHrwrdi21lc2WJiGyUpFYr/v/l3jvvqmjq2U5hn5bcdU8
CGJfNDK4K3SH/IAd8Euz5TlnK7ZRIONgJmk0i0cj0yggyEHlip6zuU4fPFebb5BiymiGx+rp+yim
SH4GIW5EXe96eu803RUd7Qwl53YFIpbHbAABSYHfLs7INuDYzuKqt5LdNhWXSwXeZduzp+xEBYIu
QRhC48iBSFI4lDHuuOqWShEDtpyWyJ+W/4wEmpN+7vQ4COS6Wp9SC8Kw4hTW2VSPjgs0JpD1o93q
xGzf7bt5iL84+hTtJDoaEegoxduWi5cJKJiJ7tc2WRPTrHXwhRCX2x9wbc05efVy1aS0L5gJ9xD8
Lu106aRwtOxRpxiU/Qnmh9SfL63INsinZjC9Bd4h8h/LVqON7E4RmRA9oS4PBDBtayI5KlxQBbVV
La0ylpXOFfHeU9IGQSkgk0BUjk+XKe1Iw4X1W8dnWComvRMN4qw0Huv/4Ln7g7WLIGJea7zXuNwS
xevFlF7EwYM5HdraNub7sKdc2fKHjTpozSs/gqML+8DCNYXS5sknyJcYo7eBrcCLIxjxNnWKbskW
KeKY6//BvHS7EPwRqpMVwAIzlXjbKPRcrtdJIvTZLvuWLayb/aepAaQRfuwvQiWMXh3uoj8no+X5
xFvJJ4geq4Mz25uFk4otWHX0pov6N+an+XjuQ4C4OEtI4GNt2jkrOx25N7eFQvQ2vyymMay41PZl
L9QfJMNi906pdw1xaYY8jWKgHb3mN+hCvImL69zIv1OAi7e8jvZ5gQr7N1UcZTPh370o1MRbmcZw
pdEFdmZklBfveGCkX+4Qpwp3EuCPPSM1bRG+YwBK7Ld1dR/j8ahfTCjB2Tx/BgSPz0wyaC59YvNX
QmJk5mwxx70Dw64LEyP9/d2I7Cfs2g4As7WxMenYJ1wPqW/ghLsXoOOm8n1WeuoXyZD8gKvzcZV9
BlZVDWdj2hU5otnNJnK5dg2L8172A4rlEI4uaRO7VFZyrlI21shz3A8dDkCTLOtnxw2oD+ykAcWZ
iG92ewQKnjCsNPoRMZgQWCCz2GvbUSDiHafrm5hGzCA9pjndzWvxHyOGZoHW7BntRvT4g7lZbJNN
Tt+RLDUg8Tdx2uFxbgn4FlaBDV2JVm5V5BRlgpORE2FYvN0WdwdCEm81LAIM0tmTgIeW/j+7xNFS
AfDV1oDS8VLx8hH7QHJraV8y2YO0UpfVy2cFcvIJQcHCbUb6LawsWPbtU71nNWSerHLnSJvOCn9P
i4ei62PyjpJSDgrEr7+Lq+VtoHugSyEsv/j3yv1k9+faux//XV9KBl+aCyzZ3NKbFwnKwCL/JyYt
x9fn6wjGFdHcmC0NxyBG3hf/iNT27IpK4IkmPCg7BDootV6v3L8TtGDWWOKteFMiRRefa9OOVi0F
NbPR8RjAlPvWvVmk0/Ovsd2NgVshFVA91QV++RkVy1Uvgp7RiWfF/wnFMJX1jBc/aVY3Cj7dMGnL
5mdSPvLKjDhZoEgRKHUhMGIsFFnpKUg4ujg1Q1XDRx+NiXnWvUlA+o4xU2kdtBZ6AFZxFwIPdfMn
zuhTA3euMJJO8Ywt38AmVCAlflZ5wBxghrYpZBn18FhjpK6EUBWvw+S95XnXx5OQ64gpI903w0Iq
SFwlsxuJfnbY5zGw7e8qVlNiD+0HDk4HNMOSjYCjRuPfbc3mvHG3HVWuM9YbiczHsiDEFqMJ+7hH
x9WVKPQ66VEfzt5zXR7xjIVA0WRte2zKOBSDWyz0VPNCArbKU2EOqLdVKoNXpfrbjjmhHfn9q8JI
IZhfh/3zh1X2/KsLsXK5XPMWqstkhSPrNX1GBPITuvcByfkacf11L52siD7aJ610ChPHYDzkmMNr
mpccV2Qi9PKjriYXogyeNTnqo9n3TsM9oly8kQFOmXWNHJhicXRA5NEudzRfLy2iiYiUTmm8H0Q8
DOGb461uNZi1gSFGP7mf6Th4W26O0/iHWnQqIrgBU7pRPkAtpNL7ezyi/nL8by+0hiHpNdPHB6k+
PdekvKQdbuS9gYKarDFe9DV+mPCEhBXsAcJx8hIxoPVznnUTEQVebAPXcdnFWGQUr3HfNjJrIb/N
FqO8SbzwtIUdCuTDX+k/PDBOu6giQPN4i/5f0bgd8l/vWhBt2Ejl8Kb+4nFY6+tUSVp6AUSF3Qh7
7egpqAsCvk3Ob+eSIp+iQjM6Rn82YgosQayOGnI6lnp0C88qW2xucmZomJizcQtcr7U5T/sjmrl+
ff1Z8/6ZIYbsuVQWLgFjXeegykV9HGGC8U3bfHvYRApRzUtKBm25CBhIKJ/W3JEJ1W4aiH4Tpn0o
CF9gHVv7YRcminuwazh8r8u2FHxRre1f+v9gVsgq0DsT99gmzm+2wxKsK3KSp6Hr05cvrrGbT4oc
sDzZe4B69YsHC6WB1tsD/6/pOJgleuGDPgK8KT7N3bx2qk0NiFEQ8xwcm/2gAuY5jr/1nZnRYQwn
QZi0Q2CGMQw64DrjRltQFBYm4paisembZZGOKTEzVVTyomFBAxduPHXlbbZYCjwl2/Hzl6mpZ8Kg
UU7EItg3iTMFDYKH/WrSoXTwZ75AdQ0XlEl3Nzs8sq5c8h/paSr/vYq+r/jTmIOzKRu+KdH9nPNj
65N1SXmNZgu4/Qv/EDqbr0COrS0i0DDggjV7Wbqm1c3GGkPwupXbd6giKy0kXBW2W5GXP3kK3GNR
kemmSba+4pDMD/cOav87iiniTf8PzWlwwbL4hgiDdFuS6xCxIGE8mJODodnKu35M4/gKg6gJnYvd
uAVwqEzqwShkSWNSaM9AWlwHaM3cwUNv0tvToFeCh1mX+QvAgTCgIKw+EwHZZEu0yWuzQ8Rf5wsV
nzEYawHiE1Q1x9UkwQ+WgK8DXf5MGe7PBBWaSL95lB8jQA+cnhbJLVuI+OTVjxSWwT88jT9cNNXr
WA63XZwMiqKwtyI+V5HnkNUJovxEsQDwRGp2UrJCmgPfXdHOc9MVXIj29ttqSQ2r446byMHsx93M
97biQcJ6xarOR6QVmUY2jaINxcW4VcWDjVZyloleNoYHVRghJb4nyxjBncexRNcPN2loUprym+z9
cP5XQZK2eIJXSxy5OYJWKexIjP8VVRhBdCoh+FWFQFYLWYYmL155/ApC+Q/MzxuY9RG3YAEP8bTl
fiAYX2zJSZam3GTt3oihEFtHw7Z5dW1lFuYhhrzki/I7PHADoJSV/R7Y/zAxWN2F9wS7UGtwzqtf
Lu+c2tz/vJKQS1DR1UJcXsAQwy+GHK1o3G537CZse1UNuZ9UKK7FIA0BwCrW7L60GmOdmsj+nenl
Znia4mgIY++7UyqVie2xvzuZFb0JW8JZMXydkR57iYnhNJ4iJ0gavA3MCAL3Cc8BPdJffp86nqaz
MpM4+VlDe8SijqWPEjPBSi7wbU+rh84re61AuZad0ssDXQxmYCoj+aIvYM0yk7f78f6Hon7KNR5D
6qQNAQJLVLPrtzpnkCPe1NtbVRugzqM2L2zt6Fmddl4ftr2pi1WJ2GXgjSskCERfiGfOwkt1Wkfr
00T61Vvr/qu5HEkPa99TFsdEa/6CFH+OZwhLjnHVIRXk9LzPkwUCOxi/1qiw5YYyG6/oLPt6nNC+
V+mCt2+arPBJVaY7cdbt4gl2vKxaOYZpr4xuFFiMPEL0hVnyArVjzGN8Gp4cGmOZGLAY1bfHi6hU
dRoPKTnccofO2qr7/+bprLvAJe1XHR1L5+MZ6JblInJUUaS8q8Ar4kMKJ22I897v7lejMIkNCeJF
KVcDAlOy7eSs5ywmS+oywhpJ0Kqey0Q9gtBrvuhlHoY314mnjcp+Hh3BWepa7PcLLw85gHPOZARK
YiPRGz4iuF4wuso3FaXFxaTOa4uAKl6EyUDH2nf/Tq3IYPfFByC7RWk/vkuu1q1vfWwygUghrJtL
VLldfS45YRd4+oTkrutYKiC8K0fONLcAYrpjyILY1s1SZsUi1KsWfQAal5oSDLZnkphhimCKrcE+
y4AEIOn/wGkJawNHHmU24r0II3mDzTUJNEavzWruJNQbmlEozLZsgyV8I0KRfrwaguMe/9GMSjSG
Dcb5jIZf+BEqU6JWTyh1zX6Np0ASfcU3Ag1kbx0eSUjQxywu+4v0MLMJV+izp0Ekih+Z1Jipdrq5
dU/5vzszaQH3ApcjJoTdtSGxTOhSw5wEMY9R1Pm/7hxNULlDDBtmtAXKHhHOJ3bSc6nesb1ioRYK
Iv1sfiUilmzdMBtwrtjJyK6/D7/gsGlo8VUYJwoy0LJG2Hsx3oazURxfVsLo03v0IuXCAjqbYQjS
cSCg3XCSv5vF8UQDukYulb2j9c/YBkupNCeEdOLSmw78BrA57HEJXRRVbdsGECA+zfFZ4Yb9yvID
qj0j1crg4hf+4lw5Ontc8LOU/NQsyKQZheC+qLZNpbVnmu0PLT5ew04/wBOxcbFEgvmJ6Uwo1F7Q
U2oaqIHzTSx8ENPkdmeb7+a+6h8/6E5XumnMuNJv8SzcUxkydeBKjSSe2+fABUZkXS01WU0vyPAD
7TsckdR1vrUfUtK0Ai59eO/hY1tPmAX6U9J9/7hh36OVre2NrBtyu8wcINgE5IVSXdtV8Hfkd7mh
94+tBLL5nBm8qTexrd66xPUWFlWejLZk5mzCiaOsieF/kqF31kAVjO5FrXYrd/m9MHmVffgAWm0S
XvdV87ZUmhILTM3ERPQWeJY5kym54vPFVaUIr55dzksRlWRLbyzyarslO9eyuWDX9LDdBSu67HSX
tEXMwieXggd54dcc5bzR3LSvKwnPuk9vOj+9+nmvNQwOvx65f3bnOfZZB3pgIwm3scTFf7k4nRQS
unMd7wP9SrfEPOczQieQ0CoLV3SRUVzsedqLoedUjpcYf80Rra+xUiXjwhfutZCv/46rV+vBa6Vl
Uqs7pxHFp7Rjv0jR15K/POYV3nxfd15/REaysw/x76Q7BJDN+j4rzxgkRpcEJjT/1SiuZhZA3etH
NyaI5Gdcx7AHtc3IJ0ZR/8L82UTsITIuKdekSKKvc5/ZYaRYRQbKKiW440xSjr/0Vz5brAFECU7B
1MypjjF8bH0KlSSo7+//C7cHuhHjWtHpx+4XNF6JxhwHFkTivz+6VqJVgnDnl+iIM9j1V5p4ieyQ
Ywhs+cLt6mXUGfNyIf4VBKu82I/Ym5m3VdiFoV8o/SpGUrc1CRaMI7ovYUeAqs+CuquLc+joDfHA
3YjT4VTn/ynop6S58sRuH0un88CvjwGYwGkbm+0v4x1VBTUyg4hWJJDE2Si7lMdG2yJ7eWBs3Ld0
n3AAs4NvPamdnxHzX7bFw3zrGI4XVLrGz4uFFhqbz8WhBaWNglotT1W4mwJCtEaAPX+7iR2r6ABO
69dXM8SXIIGMIAY7QGpS88xc7wrrkgfSMj64aUxHWWon0mJk+Q/OzM63Ql8Xm20jy1oXHBEIBhFq
ZuY+7EshdAtUBNZuFhSiWa0nzaUEi9zzWWHk6XP4CQ9+nqZXqHvc0WCIrQ2ABI1ukryuppR2J/5B
i5iZ9o4gZiBSYIvuKYENFs9Wx781dQoy/qog9lZKlr5IAaHnUkNzm9Sx2cQGCXRNa7McyXNEya27
aIaQImXgJZoHkwH7LO7g+CFUn3NYUbPcaylRX2bSqeKn8Lcf/SI4tWtaB8GWDQ+tmEp+gU4XbVSI
ZVM1EkDbkEJY9VnoBye1NIw3grN1j/i1J3xFiQOBqsazP2XYcNzSnGu8FZdGcleG5htRGTrWQM3Q
lmg0BM/X8zjb4aKqm7IdvEBUlAvhR0nOUe0MnAbpT3PxaQI6gGinc7KgAuH5OyWihXFambHax6y1
iGaLTkFYb5xJ0e1leHKENfc8oop6iIiLKfVEYS71NDZYrcYg3q/thweURJ2RptjKD1OSC4eAKwEA
IvQOHAu7QA6RXZWmq0Ek7jUP6XQ0SfM8LSuiYb93VWQhOIMPGtLmRhq8cAUNDhd5Xp6fq6F6qqqV
MryywDFC2Cnh2DOyfxy7d7rdmUQ5SJtfsUkef88+wZhxCACm3PTLRRqCJh50G6tVIwNgeXYNryn+
v7P/4Dm6YxFGASNAX9AoClkpc2wjhtCfrb3oPO7z8n8EBFbrdEjHHR83Nb8IkdM9+InJUikj7Z6l
pgpP9bOKBc0+yGLcDYy8xLuLSPaZ1K2niQIkbC2SOTwCw7xDKEuMtaDBT5Hwy/Bafze4LH+vqFhQ
msE6mJ6tyjMubPmI12Kyo6GzSGSZrpnDgfSOBbH8z5gAxnD12H+HZAbMkNqOMArwNdgsZB0ZjzoD
iciTFSYOApfwCoF3TbZvIygtiMgKIFpV0o597i5PNJneFttCGVm/u6Ia/nk8fi4oud3lC3UmLFof
ac3Dkr8Q5f4y0yFbInkrJAt+oRceYmTEVtjQ2vJepq6/aFS2kWtnwAjzn4EbsA1b+N3rLNWYBsHz
uS2qiAqgdbNgq0M0KR7S5OywwpMROKabATA7E7wU5J3Dlm0j95ILx4lwEpOWum1ACaliyzixciNT
lOnnrLzqC/S1UoRMbmbSCm9RlZ4j8kvCL2Rc3snk6wAesW9uy3gElhZDjo+rPnsEie3wkYdRuUlI
igL9eUaM9FPoZSRRhY7mv+f8l1k5zb/NXkf7/HbY8rMuHjr+uXr6Fpa70us5Whbpbs7PX/ViwPyX
ZwoyxNQIZ+jreY8vNMJiHdeqfxC87D1m5HrXhU535CRFJVzE17cWf0x8H/wxF6k6KOo4eDdRylfm
gkFN/xPAADju83tvmC3/jsKiKUdXKfSVOSumH0b/n23FLpdSR7nIw0fJU0nM8cpxMsitt/Xl66Tn
CzOPQLwm5o0QogE3cAyUvVtewc1rmu2kLs3yeaa1pDL0j5mB6dFbauwBQBoFvTnEQzMevW2J+8ss
Q4p49uOpKUFQbODoh8g71FAWEVJ83roBZJmMEBt3ieorYG+0ks+XlY8bw50+Zsqg0r+BsVzWoCAd
Aa9v2i2MsSEnjFLYYi7dcmU5VQbYN0wvwcljRKt9C6/4thQ3L4MhOAd8wxt2R5VQOH+7nnL/QBq4
Pl6hCEX9C3DWPGtoBp25YWWiW5DjJHImMJ/Nk5ZGyFC//WZ2lfUnAS1Mm7sCgg6jgUqnrpgcMlsW
acq3VtyIVtrxgsbumwozsTkuXwkWy9T16oK4nZ5/rLYFt1SnX8W9n08NVGl1yG8yHySM+ct1Aq5f
VNMY5DM+Oz5PGZxOaogzdprEKJ8D3rYi6HfUQlxNTblKm/HXaf+VCzD36IEUU8cC1vWMlslMAn7T
rwAgoNTcjV36oTyQAmuL232N9zGpRQ8bpq6WlLN3hIf/LsuNjKk1Oh6n/J+PTF5Kzjw679Ls1sZq
Ij7D+RJ9eoPBD5zCmt8NYFEYxS+tlEvZQRbDtcfMPg+XzQGsxVekx5UPDwji4t1GhJTPoYfEh9zA
GwzbVwOklCwg9I4myd/3GZF6eIgSxgFB+odv2QRdrUe3UVrBp8HDXfHMIhluyw5Ag9BXslRS6XND
WSiJ/Z4EsnoA7sOBq2pOxXFxQuuEsadRQw7+5CmrvvqiikG5Aog9zEUZ+/a/xnTl189hFzImnJwt
QuzpwOC6IsL19xDCQjI5arj5evXqebbpLv1n9fjz4sE4Hreb6OPbMRkAAKjkmiFtSiH7JfuOVPn5
i41iWCWtUnOvVodNnnUxOmyP5rGijvp32pXv8pd0KNsYNoyGuBA8leps/9V3a6lSnOj6y2m8L5v3
4N/g5rMsserXfxnCZe+o0Q0rPsHy+JtGmtRhDcuEtDjUuhlgFLnJ/sYFpD6QdEnXU0mESnpVa61L
1NvBRhXq/6dcqvijCfQ1SerITUxOeyTs8kwEFE57SED9G1esAKvGQL3UTH9UZyRnp9ufcAyPrYJh
Q+cLN+zLxbkzDAYDfgc5UMRrTYQxGpdEvUUOui3Q8PtdUaPsufxvxEr4eqXYPXBtQkZX0v0c4fnD
8FzzzV1cPM/t/jm6Y0pv1cwFAs6sbOWOG4hLhpB2CT0YNJ9FvDL/dpb5+FvNY9Hs04+qi55dcvXy
rchz5vD1fbwc1v3o9FVCjgPzs8gMNJN8/d3nd3tIrydCTFfTxUWqBSAqwKfEsp0AEMnt0jFbolFw
XuS6qm8PXyFr0ef5roMFVRTzct276EizpnPwkXn85u+Fy5RtLuiNgDpKGYL9T0foPumZvFH0oCvk
IUhIQjbToGhWT9oo+Uh5Ww7m6ObBC+6tQ3PlqjgjtS/qYripwhF3X1S/pjXkdCTIltI90Um8HlCy
Shdj4xuSm6sxm1J1BZpFzzuj9XzS5VSxxn8wzN1bAPb/7m+Q1ZBZ2mRz9St4HgAHKG7RdqhN8y04
C1zRYMMCVohgNZFAUYmk6w2nIh9nrfqMBHFDVbmrKktyJO83s05VIsN3B7022c8AWcwvlsSV6igR
JbgQgbvEQFhqhBSGQAMJ1f1hC/iPKuO5VFRuj0IF3ML3zVlWSdEqZMp6YAIu04MfgPoUL89KcAtv
8A6AGq4dTdEbFNqAc4jugVoUvVjhbP3LcrQEdQVoTLHUyibDrwBFM7ELSTMG2P2ZvHVd+YXqlXXh
vZAmTTaj6GEsiIIFE7VFOk5WlL+TFrFjeVc1RCr9li6aPFWwrxE/89pQi5styGlJxKN6YycNQtAY
R7elV0BFEfUSAvQn5lGvQ4e8bTyrA19MO0Z5J8stFEfbSqyi0dy3EUeHMjQSkWRSUnUP80QmvBBq
dOG7ju7ap9K8ywA+gWoAXk7I/0aKGM6iYgsHqROuDKUtGwUPVXAHIGPxu4AlF4Zj7I3WpIdwKTH1
oyC36XSYDZd0Gk7vcMm7vWTCKeIwYECkIho3/sbeSZli3alwrz6W4739Yp2jZYebUDizBlAMsHNv
rbvTVF2ogQ9xJ+TRl+fkfGF7zt7lAog3oJUOaoRY5DdzjPp0CerF4b6UHYc4HBj8D19FgeKNkaJO
sDJlVxzMBf7veIn9kNz4P8vEVf4APmKCReIkfQpFK6W3m4pxjKOj15BjuZIBIO7pc9eaKlLglJtv
TCui7YxwxfrT7C5JQuywKTw6ESJDFUrxB6E0kkRhU5V6xRNl7PeI4B4GnSYX+3XcBLhuokS9HMv5
3d8mh3ncQt/c/bw5AYLDVldh6CUGOfRyKHJxtUcfPd+PARGajMHIR5B+UPG+bkXTPQeYgnZYims9
7MDkQSyx2iX9fE33oMjffLqqy8AQOfPRgPeiI4nsDH6IiJ+RC3lhmUSa72gA5w1d/A8gVNfjKjCG
y8zZtnKmzOMLyxvvSr//GuxM8xsh6o7pzouqpfwia8ir7WAFDkJOjiRiNSH7lve2+YFBem8UqVxS
Gpt7zW6h12wr4exTrSqLIkNTaYXcBTRCtjRsgUrRTlMKJVPlVvYZO3gwpklsmdMoBTGrKkoHyH6R
J+pIuXmfjy4s4aEK7BF5Q4shLyel4HmgMTJLyWXo1RS/JtjmIitJ5a8+U1d74XMMEdf1AnPp//xh
aQOCerkYIA8NNlQy8u9FcOs83WU5kH/9OAxe8tw1G9SIlgdmeZ/0jc3BqalXfHGwS+tirNB7GyAF
4da+zQe4vdlC9VbREv3KRz6trnA+p8mSM9Txoq2bOssnCTXJxr6uoyfjvprTvQcr2UaX7g8uhLxQ
wHOZM/jVn0Mmbsl7QBPrZrFxGOETOgU1e7AEUk4cSKxL5IzF5EXcd32OJkiRNLQLrCAqP4FVLk1B
Bq7rvxyrjqtY4LXmv3fLc4rZvnxDm2ZVln7rLzxQUPzaso8iqL4NUUN9NVXNhzzctE4izCAKqfnt
uTUBdttCFVyIe13GxZsGqk7Xkbe00Sf1k49gjWdIfiTmA1b0rLYQWQcyGpj+o3Lj5levjj6084yb
qLR8nMpYLMtMUT+nXttodw+S6dPI9qpAc0UVfRcK576Qujd114TgAxIOsosOGw20e31vVvPlYU5V
X+fiIkSh1jmfPEj7bVwm0y9f9MwAZJjMlI/pzpbULbmEelhrpS0UzQFv8/ruIrR1cqE6RZgMkCqZ
lMXO7vJzz3p4iwEutNAZ80Iz1B0NmCHenNAau5IXtk3P97BDetrNPDRcfkhzefdFIMAedhu1wgR6
jQ2V5/PWWv0i9WLZagHoNwo/I+B4eyEsQ8JqonGvvW6/EMtHcqAUwxvMZP2cgiUkgbH5vBFt2bGn
hWS9j/sIubNHVV336ceDSYdk9Ns4wUdrwM98d18vZ++EjkuPBh1GtH1hOV8WLSUuMZ+tgDCMo/tK
hBvSOkESGdPZG0CVV0KebkOsvBxRJyqqqIWTWafBVKvM++DzTmggLsL9NM9+9JCLo5pyU1AtDMwL
tiS1eKtpk5UPQloQL9h3Ij6j3f5zaUESccOq3r3f8zzSTjYxSY3qaqhm9h5nK6RmUkQIFvUKQ2uj
s9mZ7bJv0sUgYgS/kKOsSWRypZU2SBV717KKHjxnr6VhFVNG5+eIFlE5XybIIPkwFy26McVsi2i7
8LAht7jkonZQ70f4aivBZMR8IGk86UR1qttT0sLeVCUCwIAsZm64zO+HJvdze8buRmahEBLOU6nD
OMZz3qB9xDM+ebowc2cjCDeqMEvS5AD6X1gYGID+VXxPoT2x2T7xK6sg2Y9dyGdZvuAbLnEGx3M9
CHVXEzSBV6shHGUF2nj6xpwOpRS4vDhFqdx26SLZ0B6lWCBhS8orSsogEhCnZchbfaMS+tnAknOZ
q+s1Y4ZZ7GgB9cBUzX62Y1I4pHIGDzgIbJLuTp9msMD9KpgJPNFla+6Er3ZvPD7QiNV8KOP8nPiS
7OzakD6bN0fe+uZ4eYXEqqIAi7mWMfewcAszCqnhDVtB9x35+BNQSEojThWwql8pP0t3zOJRz2eP
BxpMSUd6MkJAu16Yag7JLJxbZVm5U/r0tLTpcZP4xsESEpNirtltPEYdwKIctFP4VkyF84M0b5/j
P4jd2IHI+cJjMP73tUi7uPn7GoEJsZUsTGZ8u003wtFsZ+XzOxycB9r9N/N1GRqMbRclRmLVrhT7
DXq58+2tfWmJqAMdejgodsXAuZ+u7KqyZcHw8XIhHawYW/b9Bj9xYIykOMp7p+xXD7OYz/W8pGfG
+K7UTUOsQvfXkQ3xonqLeK79tCSqTw6sV2eQx7IsqdzuiFzJ93Dr3q190BWWYrpxIvH7pbZK8Ynk
3Q4hz9bUzEA/XkiI+AYIzz2pR8yCToP9CYiLQxVHC9arODK1/jI5/ckEs7w+tQNWHOuHKbwGjtAN
+rw1Pm9ORCqptfyyXZWR4SXStR7m3udrDWINVYtabyhKBnFkVkzhaEqZ4ePVMW7eOnfs+nOIyxBY
FIwOTF6MPxlzZNsIZk0KEL6DgnqWvkmi9Js3ucOi/qOPZA3sUiweKYIOg9+UcuyHAJ+J2uAfItqV
4Ug/zqka1jZEzPyYGsciaJ9Tig6/lmR00FqSYufHRvJsZzO/m0F29p6MzUWIaC0UWsJ41QBZrBOC
r6Ebi2RjW+IiiUrACFhA/V4L1O8at++1n/JL3+iemMKW0TmAHiZQYPrtyu2goXCvP2iADUyOYjqb
UlvqzxGAR5VgVr3dSY26naaBhd5X9dgXmu+Bl2juolkXpve4C/KW+aj80xUIT8g0qH7aZ/UsELMc
Jd1w4jtGkw3mJmiVS+jok7AL4Zttc3snuU59mRd/l5fqgogMyhrNs22Dazg/YKyOiQbov6zJVM9k
ZHXw869EX3nvFEaPvL1PFM3Gv6kaXB6ckIRrIyxYggoOLJA5qclSwp16n3qUKVBj2mtla9uR/9B4
Y36O/fyHJINxk1qAw/rH3epawKJbrw+OBfFpzOlbV/Dsq8biwidWOyc79VMjmgwfxivTnLH+CoT0
lxO5E61NVQtRgiZertWrZqekhiHdnoqVMlaxMJo/jPD77nVlI7je/mYfd4eDopFuCA/NEgdX2RDq
R3OyWSpgBR7BMIB7Z3ZBpFEr/HMTlmn2Khgf3DZ4cjzz0XWbuUQfjAVbvGJWm6qOE4XBbjtk9XIY
0YP5bGQ6yS7awNL1++7UPWwIq5nyTfdc+wLrqPxSRgn5GFVDrFtlmqf7WDWuu2XJqPHOrm3xGYvM
aklxfmq7ivH8Fl996IBa0BH326O4aEAtkGIrC2PifBMx/VdOGMqv76oK53/08HofvlalVhbT5XHO
VIXQX1Pt7mFNnvooOu90LOknz8QNBie7S131OCm10G5dc0mGTs0AAnXDLv7mwWjDdbvZuOeZXjq1
QWsbxn3ssfoOMtBq2bKezjZ6jqGIzBIlPoSPlyGt60LMjboinhDiwnz5VyWgGKBNrHtINdxpTOLZ
x1XATzeT+gxBlpZiodYPZ7P6aDs9o/kAnxzczw4JLKnoJrhUc+K1/5+CbfLKVwRjYSD30I1kUrs6
PbH8AXAMGhWOnOtllmysSGWY1y6XQ45U9szash1htV8w2DHtxDBWyCjwc523Dn3Puj88NcDMCwK8
bGxHoa9ORkwzOBY6dK9x/LFnHiKqA5I2NbclNqaM20aqxSngS1sCfGVuJNyyBjD0LFoh1SiqQAQx
5zhswzfwH8x+G+B1J2UOJe/EXSQVoiN0TG+FXB+kj7dL5QSvuRK5BA2W8EclkeKm4r0kJ+NLyRNS
rdsZQ6UtTQM2346xRkeyR+DuCaGmBJM1IdNfmfFeh3KV2eGPQUl334ZqqTQzIYscRs1r/eqRO4DU
FJ9dlhNlLgMdLl2sHdMuZjk7xEdG3iwiO8sW5kX5Wcqib3wl0MfbiqWabLzI2qJlN8j6RdcJcyP7
B2wIyeX0k+Ws5KRbLkRSu1RFJrYVyr2fnnoQf9ctDoOUaLZYvQmpo7MMGAa2ydAlhJOKeX641/2/
M89lsKi9x+TGeGdpbj2kv2dVWayx3Nv0XctK0zGT5b2525ZbzcjimvSddeymOCLhSOdV3cVglbtN
UogzLu3fitX+39LeLfPU8yAMVX+8FTXZRcdXgEXq1qGaznRq35n9tUvJ3/MiF9oBneWsAhK9tcpg
RdcArYxGyj01RwEuhmulMgZRdsp+ttPHorQHtnbVxtYH7P86rCNANiUzAqv31pOnw+rKAQdgDdDE
JoIvj1xfKrPCEN99IsoGWK1fCcl6iOkLqOYZga5wftwh2fFUbYHHipFX3GJIfrazr/K9mxpHi24C
F+RD28VYk9ffzjcoi10mPs/SOy4JJxdUyqb2BLzCceHdC3qmIXBOCTHBGHZHDsii9HxHZKTRyUV9
Dz/PFpqCKZBU0ZCojLe177iycBVdgrLINtf2SeSk4FTvEC9+UoSH7blYnT6/ZnjzIVWRR/2KzFXh
j83Sv0hUz/eeCcj5Amms2KK3QFFBZsJovo7IIEyR+ufauqVhIPq2QN4mYCQ59jJTirenyezmUgdP
FqvVMlxv52t/LlOOmqqwapqpYYA8rkF/UExepiSEPIXcGfRhL3SpwJSgWlOmLjL7hkdeBw1rwCZz
UUalLEb/oY9KQHwXelTKT4zZ7MTZEIoFYkt+tjie8bEWRWbWRVSRKJESyUzPghTVNggus5dfU1Fh
kgoD8KHJSgJ0UrURJlDBZ6eGH7Xxx8b504W9UoWzKUjJug6VoCDh3uKBXRYvBtUsrYW3Na6l3BQk
8HWZYe3uKwPR0q3kgjRndjCDt9PF95udosgkIKsWbFS1iv/0lSZ5esAsiZHDzh1rmMFdbkGv0hux
Kg+QFpbpSkqUrGEsbIRCsUQwCASK6M2ChMEOa8rolL8Y57qabKSG4LmTCi8aH9y8jde4nfqkjMow
wKw3NHeC28DhluXFrbCIpsSRCVCHPmmL2A/lluNq8lUQDtuOUEkBr8/1ZSmcmfX/VbavRqyICnwf
xPE82O0j+b0yJPCBrLuTlY+HGJfTJaFX3xcLEwUf7hcwHuUlDGVFOehd8xbtZlsfVz1IMXr+EaR1
NSztWZyRRLm50rvmmJkmgLZ1vimk+JQ2xtHVFnT6+nUvwUwAGc80X5JuqaYpjl70dgLtBpfCsVTJ
SgiHiaLpYTb6280YHlbbEEZcwcL33Nj+Wc+O/zEblLyJ/YLKj7xRkXT+zHG2lmPpyWfGTupQ1d7P
F3lAPf21Aks97yAlZ+HtGj907XYf0idKknofgqEQYd9SbMX2ySh40mfPx3bUpUy4cSl8ayWSULgf
Mblir2Wh0Ml0GKAB8SWdSrXSWgW3gz62dfcCwBx24RF7YSK15oZRBD5O2R066kAWVA+c7W31nJ0c
6Zzrsdw55Zjzayor8MbNMhdxXjikHPm1On/ix2akjJr+3fYPNPQ3lShGbCPkT/lMJHldH0R24Y4Q
mzlPxVZqrF9VhWlSch43kLj6eBkNWJOYvqeYlX12obK+YGfbx01cLtYgQAO1QJDhfwCPkHfvp1ZK
p4X033Vzo/lBZkJYiuz4iymMQFNE17mZ8VuVL/V1A29FjQsxSCeA9n+aZat5yMKwn3fMO1up3EMY
9ChNPUx9nTbYQkkZdZkLW5gcSxaPRI1brincOD1/aYcqZmHwwQV+Wrzqw+mvOt0QVh99tfnHe1J9
zxt7WEV6cxN184b3SDI0EGS4CYmX+v38/4PCw7T0DvV4eAhjPaB9F2/p1FrzuZcUNcWjEB+fESWx
tlVx6IA6mlZx8GN8sUbZmSO0dyERANgbGdMwUuEcldF/2QvBJftOFrIPMpW+Ol8n1bMAv8oZ9s6b
MylNje1geSHKEP4/4VIHPHuB7hNymSP4p6Ehk9ESHTVbIVipDc+hfby5eHC71PqvX31XQMfmMg0p
rC+iIQUVAN4G2JHFzXiTmAliYYHjsEBKYVhlZwQHpUeKZGSqgVlxv1GAm3hoYc/0LheGjw1cdszA
/d6hwMI6JbO98SfPVOw7rs9+qRIUhqG2XQIxOaukV01VQboWU9t1NrOBsjL+Td4Lpepq9XpKBE90
RvQgzhQbV1nyn3uPFUSUhn65Oa8L1TdgUFX2IZVEWLC0s31hc9wW1t8pe3dQN8vxfp8LH7N+ceD9
xl/BUSUojjwL/jvmrIUshhQFJpDUCRm4uu1PlZSxyX5dPX1xn532MQkXBEi0b1iV8A4Qa8Psrr/L
hqNwR1qAjQNbpn4Q3MG0pTyM85Ia2rYNnT+CNI/KI49QxjdMFkY/L4MagjWGcbXx2iKVr/4npXJR
tBGupNMYbaCxvjHPuhIlxuh6c0F8l4Z6OtZFMezCh9f+kMdnodDpozZIU1ugDBLSZMj/Q+Tr8Ywe
RRjzj3WaX80rx5zgXE/7MfAYrijE40tIXKXh4cDsBipri7wBzHN6KHKqBiBGLr4LpHJWwBgCKfoR
Ntu3CbTHJpFfDXMj38MNILkbbjHzfaTwM06RyWQZNa3h4tUC5e8clPhkqLOR8pCuPaBDx2r8MAJa
7XJ4dROAOAI0TRKO1SQvCZloZaDC04gv15H3JW5KaPHAl+fQd+QFM+R9RgFTZ3aB/t2yTws1UuEF
bVTJMjjOiiaysNfLyxvlyoS/PVn19YFOTdMc1vPLw8SJ8TqNBew+NRcZO16oNNaDt90iqT61xGn+
YyYYGad9iQsUkVI4T3uJn/XSNuphwHJfa7RBhBmjAIT7N+z7WYGkIbQyFLUvbqw+hz5I3yH1VaND
ity2+wtxZbsvubLP1RhbMynvNI/ZuNjleUOOYDlUFojW9kDroY2WdeQESZIlgoPOOlVsw6ElFXsz
KicjZZHHPZxRyoBMLfiiMdYVaKBxrizuIRQ2El3l/uu/HLWV9UOHrvHjqkam0lSG0rkyH7qRYjKp
/D+dxcEseZpGNhiM/DcP8QDhcvgoBFC/Vz/5ZmgmEcLMK+IzqIgIlxibvs9xa21xHmbQDcu580oh
QEC1AlhetiXPzK0jRT8fr2rSYcAhRW7DZi8W0yTzxrGmAa2ldj8HMyjHHq9mu+AJEoRD41qN5CNG
wbqBkVJic3dfpBaFiL7IhnpFYtpSC+TdTr165497gupMoeri91rZ10p8vPnYWxxaKs6SgyONC+/Z
VCEM2TPPmTtAkkKW9H/Xu92A4zikrRmCjmKFnkK3vLppyvNlJOQUlstTftp9YQNtTjtX/EmEr1Du
/ftrmONLOGn/59m583/UXkPV0T8ViCut5kwdnSKRjG3mxxNP4YI5QBwwKAmExZ3MRRk/pgw+db/j
p+ytR6SyKZrnWz+6Z2423WLJB4y7d7NbBT9J8gXH8KchvYLHR6WZ697GtjEzTFPjn5NEm9QbUxMt
aXPK8QXRMZEkVn6wEIjOySc7Gb31kPZdJRVPoRpeSU0UFhX5oiERy46/R3u53Zl6hoMWoNo5f3ff
60fPQCUVlbr8PEVNlpznjX+v9UCThjZDmfE5DVyOOsPjitu1Td7rNWM3ZhFFVrr+vDpC3OZZAcih
S3oKZSaCDp5HtnXAxy/CD14TtHuLrXkmXiDjlMXqWvL+mq/nelio691yZij8BgrOtU3sNB/9jdmN
o2cjW82Ikkfhz5KD/EKtpmdg5zBl2wCMuQ/oKbTvEvS2O3f1gBbe1aeuVbJRBVdY1v0FdhRaDSKa
GBF+dP2xtaTzEm+lhanOYRpAPVC3zmnKK+SpF7BG702RVrvG+LPpRrfP7cD5bq9gyWYTPR/MNfDQ
iM3vIF0beOanA3iOvCKz3XMEjQ5wktZ/mzyHSzGaUBGJi1f7jJBnED3n04fO/Pq3msqFeFF21Gn+
Ldcm+A2qWx2QDeg/lUddEAC5o/EwjTi8Lqwp2EX81xpJc2Q51i0kwMT2LMoPmdP3qup/yT74wo4R
ReY2HMaPVVSpAuk/TGsEkG8cyawJQVXBjfY+CrMVZjop3FRePtjBlOjCQtpWFhmfb2td+WiN4eHk
mIytago5f2DltnXxv46yBBzL+LKxKyYIeV6GAUh/W5TX85OO9Z1Bq/d5y+lWZuDdWpgPXeBavQ1+
nkhk9so3JINSTE/1zp7CM5uWN3hmkJFJur7Rb3BrQfzhfutgDoCNItXHYjxhyWCao56ETxi/fqpG
hLVKRMFcPFwE9qqQgaxve0fmnEbfOBHaZLr+VminkAPA44/R9aOSPiy4XnFvdMNiyXPlOG28xXtA
u/qT9rCWwT8o/iy+yJv9k3Aqvap6Tq/idVy01NJiuV4ANmtywNneyjPasiqQKpU+o6e1RXeiAMPv
Fcujght5FFuyIFdy0BbbEqHjLcWZrZaeEr1UKB5ERZXST1j/yVql1QNdDb+xUwtIA/HZ8PwgnB9/
EPjSe7osiIEybQpo3Tm4ZcKp8fJj2UG6tXvWs0XJ1ObpdmjCl3OqIq0G4QwDAsZid8ob9znfD6tZ
rPktL6j5uE6bKqEp1G+g1RH8yFch2ILgXBkw953jyk4l9ppyVlDtDvpDUWDPPPY9MLycJZmqWiKw
TZM3hVk2hwY9AxBxA5epa1HRPFqyYE4gf4BgAq7pXyyUfowX+JZfonjNcVwZPKh8Org9Op3Z943n
8fMRtMHHxc8RQGnINefcLXACqkngKdvfVUiz1nf4+tr17Dgtp9zySH/BBh2BRQC9pbIuufDOPDM+
YrEsKBWjjUFU31zX6o4nE3JoJRGBnvyUd1ppUNkA/PeU56Sa+izB/nv76/R7iYkPyEwdwAM7Bryo
brlLYGxek9avFPs1s89m2jmF/YopEAbZt7iGdT8PimtyMQzGuZGtIfNetDWCNE9VxMh74eML8Smm
ecldkZnPw4v0a9ZTNn7bZhrauMtgVBfTChbzXCq7nOHD8Ft/xCgHS078N8kLNTYaWHTBQsEy3txa
NIBj0lyE45xu0sM6QVhXC1CngY36Xkg3OhTMYCdnoopGBxJNmRwUC//11b5kJHNvHcbhCkLp19M9
i0nM8Zq+NZTM1Kr/p1WVveItj+3jYRVvJ+NHOv0SjX4nUV1XWX3eRLGOwNDjbPeFFtBkRyZ8yhJN
L7rRjo9QXgWihYBnmI3etjVNSXBs02MGVZf40sgqmXmzI9tSwGgOsWRRBQh78IF5E7KhzBeDdbRI
b9aTY/W7ASdxGrpYiHf4hWuUkGjkq64sm/SqdaheICDpwB8tgAXIw2KWzFNNvOqT6nxDMqN5uO68
uftJqM2YKiAZlhQDHAq5q9aF+FBHHA03MOkH9l6BUH9rZtRR+v+32VBqOq1nF1BGVO0lq5cZpqNW
wNYgSh04HmCfU/hRPSDgRAZgrpJo/Q/KFagoPLs/VWAccbIBgPr7XIVp+iTJv+ppxN4NzF+W+x2C
VSUzBg+43qsDNB8OQk3wZgISv3HtB3tj7N5u8XeYV3swhuS1IAHSGZPes1xQ9RD5rp1DSYs1op/V
DvDUk7hIp1apZ6WzZaiai1AXeYUuNzUunxMgvQwMuhOiC7FbzD/vcqLXekXV7qiUWIvI7/EErXHC
qUHHJ+m7GG0ynqTBkHdw0WiQKO/TJYcZM7azDkU6AdAt9mCpR3ovut15L/OOH5l0z9IwhQfubdHb
5SKPY8CBSQpo1LhySwKCBN9FxCpnDMDnLmad6L6kMPhIEw+6RjRkjtIJiBdrtiKo8J+aLF3SqgAu
51/XY1Po277esdUKgl7Ai5+AsiNvXfOp22aS1+DrFDFGiocOQfBNfIFEpa+RdJpuZI63PYKZ2/tH
mrA1sRT0uXYS6+nyYOGYTdSbE9HHhh7FcTSRodVUma/3I5cDor47uClXlQBeDRk/1dEPv+RPurIX
eHUmP0GlGm0aVyXsjceEu54JlcSrsR3zmWriWN6Rj+MrXat1dwnBk5S11zFOnlFGvloDaM72/KxN
A2ssStOqQyrQ9/05IGq32CoF5ihXewX3wzMP/nV9QNnW6MJgVPv6Oavzws7WjtlNJp6OoTUmvz1W
5piWoeWn3BZk76L4SP6uL3QY3bOnzytwfamo2Xky78c55pdbwAduWOFokKoMUx2HLl70lEcIU/Hh
sYXSFLOFmbNua46eGvvGCkQb78Wfw0AWAbnb6nLCCa8OFE+nOyL0J7WDa1e7OqAjJwiNOyhvvtHQ
ZA8nfOjx1sCOltyYTxFXs+APZ3AMb+Sb7FRUSHilbN//zVdcZVUrYqbexWDOWViIqUS8nWDhV+Jt
MXGSLAnZxKqcTXv1KWx/O4xCG1cTn2DsFAo9pr3Evf/AFf89UTIJpnT3zFBxzDCL4CVd/XnTicR+
Hd856cXBu5CNNqvUzddk97G+PghBsIuG58s31/v6eN79zxG+8r2QY0TxhuZCn1dorVP2NEVPmyEA
JjM7vju1zC4Q/0UUrdIhiYx3CO1DDnumK6K0cFRAxZMr1BwQrsyRw7kgoRYSHBJsvAqL1ncROTWa
mqDx6QaK0iyU4iVSTGjEtlV+3+IKsjoEY3WI4ZVl0T0WLHd6/4Bkz0ixKkolHCIq1UP7MKlI+Gf4
4HfFDzjYM0/q9GQRkQRW0NQMyoiWVC004BkNXz1c9f0IbKVsg3+gJ5ZQNH8eaGeu3XXaEDoCnA/z
hRuuQwKrnyCKwaoWjFBjvb1nt/aSVkmfV6KDYJIB32rmWnm2ZKEPNuFglkW6dIXDXaTYIT2Dthf0
YndQN2CghollodrhBEfTACwlCQoG25f3MXk2gNNBpP58h1IKEG4farp0rTZz6ZtrpoQPsuTbxDUf
aFV/cC07JXKwuzjffhZemK2M+FlysAsvpVBuE3PpaQ/MnKqzubaY6GBc/E4DfWCLTTPhgUiWLEEf
OAgHMz7xe9KddBFnUjRgXM1DcxmpSooXmmNoxzMvx6CbMEJy/nEd/J4bPNbHyduscDFFYCVWzLiZ
pV+BVfkoPvJzpEKvFdP/F1etNy7myJ8p5ftz6j4wWrLQd1gZoR5+O/fqMIGCFpseQjVAa24AUiJq
bD1iWQS6B7Ame0BPDwF4LWSukyXY3Wmvt7VMqbiqX27iBwVD7RD+OdC68buIzYht9VTsfpDUgLAU
7pb678MdfsblfGay5VRhUCK6QUiHxABl68eGS90oZfxlO61bFwU5WJ/rI8AcKRUq0FUD6UzH0FJj
qWp58x2RDMo297txnm8NFU9SDqhnnkQEM9seYYIbh456Gw+zZ88JEjNdlenaN1kZuHz5RyNKnsUS
m4b94BfmdCncp9PwDj8H6k74dDinjyyPRAkrqq6EYYYTePqsCdjIBglczJMfy3P7IuP2tMV8F6WB
SG8BH7Sag+l8DrJk1yqAlBIuXCRZ+MM4lzpfErgsifBB1vXmRgOiayFMQcXfNDm02J/pnW1Xr38L
B1HwcAbWMqk3V2L5VxrpIE78xcx9F9/fjSYkKS9+Y9Pxwf5S/mGw+EA6EoQnTyluGc1m1JY7I+qN
cFSZlYu4x99iWQrucOuOTrQLCE4sJNjFB+A7NQf+CYG/VYcZ86DDe6DB8HPlpMEHkstrI2UQXljz
o//vydHkb3/+RyCUERpOuJzs5LqeXau3p4KQP7EjvT6jbVOWCEjqypjZ2Y+BxZklj7EUogKSuuLl
F6uHfR0Ys7qmeYGQv3ZEB3ioFucwSySDt122wTucV0IZCBjNgl7K5y9+B/j885IW7lZeERpVlHsv
RdUytkRGfttdITen8vP18PjO3MPc1TOZLdq+I4f5mCve2leP8S1KDzgkXoD258INuoDeFN+ZpE9P
prc4OCB4rp5CninP7g5yMFIjusa4aalWpVo+uFCQTp1VEoAvuN3CgeMBSjjHeiIy4EdEFWS290b5
mJdisRC91HyGuaJGAUbd/j2al+uw0k5zR98+6L2SGAYKczxa3IVG1sLaRWcF09wPBwtc8h2stjgG
4iSAuxdjs1xirZEEZ1FakXOL1ItwwG6gCHQl104fWQT36PWORXgaMAv/cjJdpu1hTIVYPWdWkLbO
pbnR/STgI8NjH6aix8Z0UFweb8VAIwBzfz1v56hVoyS0lkujNAJVYFammbPMONRlUn72B9vwK9Cl
TH+BvmJfXPVoo9C/+PsSl+ws6lGn41hzicn/vJneAAlS4S1/+fI4QOhpiKp9KFQfrXn9bw//fkYq
tIHhgNt/FiumoSNkWQVegJluBwItnaOzGGIdVTxfWJ0ak5Zsu2BsYqHoqlLFTI+KJYcUaOK9T0x8
CSTz7RWgqqFQ4pKeHQkz5hcVW5LvuCAbolOfq/qGC/66CL9w2AteE1NA5/S5kDGEZKw1TX5O+uCO
wetzElkt5+YXpLzK4q4v+M3YBRCZoR3MtFkmE1gLDc2ja/UmXB4giQUC+O7W2xrKWjc6XfbY2wmM
tDAAKaxd8nmHVX8lcRbudsjTlc5unaKJ+vhsb9pGtM7NlgivIXVXja+0MqwkPABxP9q8sp852ilN
RPkR+9vUWOeBccd+bDlKRx1v/gDc5rWp0w3cb6LljWngCZ9wgiD8iUDe0S/KLEcqd1zxDCgf3JN1
3XlKt3KymqKgR4/EhVbacy2R1KhAa+Cdi/TatCHZ9/m6WxJunw9GspO4V16M3RmhwyxjADXC0wPw
O7oG9WEAxRgZ7vRmEqeVpiHBJjdwLQ42hl9RnNPvtJ1F7LDqg1B7tqcvOkl3s2d+5bakr2+AFkR3
fm/2O0UsmnCzlkVCvMcN0cV/tk933/qVq3vCrOLIAonvoRx5z1jmqwtaVb2/pw+2pGFmqLCDj9KQ
JxU8+Xm9FzqN3eGbU4aBECffVkicvdE7WJ82xmloRYkXunE/NMkBwjVGXZucktFJVGaFMmWDWRWV
cs+AjvAVPqnbIugDHa+QmUqd9yhc6Qx28RS26zqOuGalczmAOj/Dd7dW6Y01Hb8PM4vlkh3ZOKmZ
tNLZV6xhZHrbJ76E1dKELM+Y0H2FKti7wOEVPI3zS7JnejzKP8ZdF6fc56U5Qivd/CRZQZKu8rQ7
Y4X8D7SqHFvJMlUr/OpR1+epUV0vd771uUyRY3sedNI5M5OwxufBXEwTz3TNy1RS+y/E8bXRuL7u
m0ivIc+ptzNbovF//m6NAq6iSJnAePfSPiR0/A+BaVsmAFXUCf/qol+Rs/XbM8EXGQw0QS89LEIm
i+j+kNdBTGuQS5nDav79lLyoFv6l7H4zyWx5FB6rTecIR3aLYNv37GdheqtpSDzlmpTXhYMtsktH
Pne56yBXHhglUGnEyp1AkbMRuSsu5tmz2pfNELDeOQDAkC8FiFBsUpJ96Aeh4OgvHg8Y7n+Q2uRP
XNSN2G66lENLTkf7jgBjU4Yhyi2NyfQ+O3xpUA+rivbMFJh73libQ6beEPHqITF7cf+RS2jeO82c
UPdbam9TAk8YjHbV5SNxj+ULSRaPGHiUfV0eTn2VK99Ez3NYfPaX2qMdUQOQK/nGcx3S+hApiEO9
w48TEzpi9e3oSuZsN76Om78nCl3tJemeQ0ZXOCHdilAATgZ4foN8LKmRgOwCDol0G3W417SCPVXL
TT81L5TmSlNl6u+hL59HtVN2P296jwKbbNUq5uZVfHMihb2T7kQX/m4PMUSC9fr3zNUzMuem+H3Y
Tew0Or54naUaUDRE3RE7zGpF3BraPkwfWwQtUOgdhxJrvVGH92xxTybDr4l5D+loGFXJShtjPBnf
0l+Gf/2XQAoOz9r6REAUtw1qi/dHoLEGi+ZLNtu2/sl6bfgZIOtS+ZrRWaaVhRzRtR1ECkkmabRS
k9xloaWYTgNHCB48K+GW7eCATYHiGLBY2E6rEfs8bDEvXaOFBJ0xKm6TF+AfbZvwWQWlJXCTHp0n
4JfnKIypnz4j19BhAtTJYGZyyUhAt2HxY8poVLkStmYPq4NA5IGcrJ64ZPXEvQI66dF+gjGG0L/J
cbz3uPRxqMpfAxkyDWoXoTNGh84oXWIfTccXdCHGFn4eG8t2l4xI/B8jmWdgIdcrcxgna4rL3K0S
X6VUoDex6M7yOiKfInSTpct6RUm5E0AHxNUnde+q1p0iGdNri1Pa7FKkgICTiVmNjkLeK7MBeNJb
8LML8eZnT2aEK/gBqzeIhpQOCkr3W+UJ8BeKdO/OUsJ9grW+SBA8eFwt0XpkdH4AvnlHDp+aMQvC
ECQ41PBq4bC7kd5MA9IYMAme84O1ictRK4wtrCaZzLOIkaD8HbXQCxz1Wbv26vIPPkEpwMbZ8rRx
bsFUTIWRUxmFcHQO4bo0kaTjtXagluS+Tu9q32Hgj4c8Qw1Sk5GFoACsPSxoK6w+8ia+jl3dwQbM
sRAYelDBJGViJQFuQs5vf+bI+5Wv/j1SDH+eKKr13iUz/AEEosv8E6PW5obXgit3HFNzhILMoqCm
H1TKpNRoeNhk3NSFspqida10v4ARB1o8dp8acc9JfP3uPspCXYfLwboCOrfd0lIUBwIySiXBhD8o
45i166HW3dRldfo2ZOBzKO1ZZoNj+0aJkafavB7hyNmeSLGbHWSp0mJoTplIFbjvAd/rwm74RjGV
jBKPEj7fMSTSPRCga8w/p6g1+bURbMPhsKLXH2Fwy3QfSTr12N4gKjxo7I8ewtaMKwPUVhL+fIG0
5STManI/dj5q3qaSxuayXrJNWj4wpoDwEa/vVOVJGmW/yi97/riI9q3TMCA1++Gx/VdipOKB4fB3
JjKub+jam1npw6bEW4tUEUqIQh2xL0btqJxZn5jj3mVn5F1spGbCdPqQoMQj32c+KTZ2yaE2oRjJ
2hs9Zd4/a3YxW0GR+evfFBCzXcE7IVVI7HFHICVGO9XVehc5tbPerrlx0HFHCwxwR+QFP1o02pmb
73prSOCeK929Zt8wjZe2VqI3RkvewP69mNnsadmDn//NwWQvEEqqKBYSYEiTrthY+SDnhd5164hp
HzhRSh9r4j0JDWObRjIs6FCZxSJMh/I/NV/bmXLrO1oacSD81N20PuxXBbQIdszFJ3K9HnXLUQzF
Y6Ye3FAVDv64Spff6FHr0jdscu3OWY2bVBNtR4cNeYvNc0+423+5OKr/2rhxpN5XBkgyBP1SkM9/
UqkVgjl4kt2HQ1j+JzfbPCXgz+MVI/UXfjvPK0CaTfWxLeZaTw/5VRLoQBg8O2tdt6I4mmlwkYpU
eTqs4H8w/78tghohmmWE6kUGRWnSfHWXaBNENI5g5s0RAC0GEZw/uKqpvMLGgIs9MGCSVBDGmVVb
EDtA4pNbZgJSTLcSKBChE0XyaId52bGvT+gLfGUK8udIFbGmjTMqd8ux7fHWW+nKgV67WecZ0AHd
SJGcEozJNHTKFpDwlA9ekhgywqeNqrEUW6qwB4jPC+9WFHlv/2Twf/It/J6wCw2nMjlvtv+J9A48
dkxhdOlpo28TK4+W2d2pq7IZKrkxPHI2hNX0sFgOAUbEf55C8+Z6loxHq+ljfHAawVDtA8J3TWxY
qXqd5fE3xafZaNKTUqQ5Kti73I2HXJ59nyv3JEzO5EBiMEP4qyPt1tnrhNoV9lWPmzCK+qsxOkEW
FkiSDWQg5MM34pR7+pOkURL0yvyvx+QXf1bKvgVPu5HRW4XXDbBIe8arooIj7KL/YMwyV7jxs9YD
zcYbGe3iZgZBpPoZQemCluK/5Qzdiswi1kt2Ez5qYeoPvS2nA2bJnNCZYJ2JjhN2q0/zjKgKLbmX
RJ+gl40a7zLo7hpNTT/0qzED62+htth1VCD9PDxaZCeWcL435EzOmSJaoP0gr6Zjfln4w/zaUqY+
BzxrSm6Ls0t2Hyy25yWsxMvw24EHI6vSSQa/oFRE/fbVF7vXnmyoedtEtvYkv3ubR6RA60HBhMB9
Vb1VgoO+X0nbuOVfalUqXVjdejxYlReXTKw6oAJc14JyFDKyoaMcNHx2fzauorI1thvPr1/wNq6m
G6LovFo2dr9TfHrYipmPI0tcufa4XRQ5GJZYtijv+nCjImuuGoEXo8gkmx7gaK4Io+L5sXpsb/N4
rh663dVGREh6I3QbiVEXxM0bYoSFdXoMCiGWdlHHLzzr6xqsqUpuAMfIgjr6VpjQ7ceAErNPUG8K
fx2O+5CtDSMya9PEHRdwvkAdOwjEnd6ItiHpsBu9+Q2OkUchQiEP84NFMZz52G2Ontx5L+rvoBZx
QGRd0GAKAExVOZsqJ93MpxcwuS3zAUc1q3mXNyk7Dd8D7o2shwul+NLb7IzX/RqtBXlQTwUKEgPd
YlPe4UKiEbssIGu8Nurz9WzCHVn9u47CwJl7ryv7EHHYfnpYUogRbz9EVxqKRbYakzAbFU6rdAv+
PdzKy10COO9bbIcsvZNQLHKbzDJSP5i8BEVmB22fXqBqAhjqUqtEMKnpHGgvD2ygVXwdZ7wxAeXg
bLC87b0lW6JBO9vUvoqWAu5z9qfgM3xzmUrJuXPpsFb6h/OwPlhFhPvYDzq3EHwWUDqnaJeahcBs
oyOMaegCh/+NOpQjhl363VTqlJMVq+QSBZOittC5gwgNA/WT2cNAPy0Esh4w6V7mfN7S3WiKcnsT
E7QetwVNlC4o2B1uF/AAaRG1aIl+fiPfZ0WDjVvsysCikazCzjNGSVoC0XMwF/mWBjBicoswg3f2
AdLBpPiVlAG52KaMtSrHGjQsJ0kTRkORdbnR+RodToAJDJke2mKMZZYmNho034z/BHOkGaNRi4Jp
VkEZjmWTjOQShC1i7vYQL6FUIl9MZsT9VCTXAg4TUW5ievN1R1WTMy/rKa/XPRvv2SWWQ7tSJEoQ
H7Kj1lPsh+rm36GKjC7SpPMDUgAi4aeZB/n0hWbdDdTOZI4RuP1LahJQgddBDIGwUpTKFnf/jZBL
hili1mbjeItbsYKR6u11Q2ibsQut2KU5kMl9DkXrJqKjzn0aIYMNMfms3fRJKQKjSyQR0BFhgWy6
pG8yY+dMQ4rx8I1WNRLdtvn9aRRueXIam2EF9yfkcLjkszNkgdf/owpSyQr8MMiQNETJ1pQyNWxP
HtJ5nxrUKWlWhykybWZFK/Servhhxh/9Q3NltbowyYWZtjQGM+PZ50TEk5exHbtFcJmTdBkhM4Kp
tD0BcCX+2Nh7WZSK4Xt0Znxu22NcitcH3FWr1aAKDVV9VjoBXZFmQ7KdHDFX4O9ZzKToglV9ig3E
zGWfrI+oF/8Hua9QCJnYTlFhy7g+VzWNgASLDsIm9GjvMU2yzNSJ9ujaBnwPmnuEZzllTjj0SKlh
hzb58iGM8PMeCxXlsF/C5oEkqpqcTVoKMbNl8GHFdpTblYAYTOzipFJbl2ZWoyXGmmLN4KFoWLiy
8nO0klMwrG+2qwfrvz6Yal+BqKRN2qz6Vtbaxcf1yWQU+WOygdi0GOUijPqU3zrCzfo4WFHlOpwI
bdorvXKb2I6RGpr2q3nI+uGo/Pet9+o5qesp5STwj2S02Yh8SJcmo4CHta0JFb8fobx6I0HWFGQN
t2PQmdBa+fc9X293Yg1E+lNgvIB9dIrT41K+1pUR+Z8ByQDblYMaehhJmGlCTNYpLfDtc+hyYVDI
pbXOqE7RuP9/m13pLjobQiYX5UiiEvJz3NH0lUHr8BX2DkryVWs44UcwA26dnvBKSyNHQLuy+1gS
7BxHbw2ffunh7bLBppXWgtg8Uwgoud5CVdoJ4Pq5aqbtuPHlCZpKpSt4m+6kgbjtqx3c1Fv3f/OY
nbA0TqJqPtevheb4KmLuweoK3Kjb+MRkOd9IzD/4JFTRYfBkoKgIOHFPkWNA82jGannkaLS9Og51
JHrqqiYU7BVEPL7bwJzDYyVaulzs/pW/1T2CWGnBYrZJiHmngnLPXT1akZCJr+tok21FtoR+nNrd
1xzFS4NJfj2T214e5BnGjP7qUgpDctPNUaY7Mj9yMZs0sIYS0xOvyUGbN8MwKgjYSxMpDwfue3Tb
PIACzg4GmJbN5eiTys9BRqkXN3UI8i1PpgsbkxjAHSL8OMqgTrrS5d9n4b4G97p2CuN6kAr03tCH
wOGNfU1ioP1g8D8G+5ex4GfKahW3cZR2PUzRJYs1+MvU11aBM/w3yDNlZB+V4bbJIfNJZoFod+Yr
QlpF+kkrjo3ukviJsDUxsWaspxsINUXzNx6Gi2GE7asiUNYey+vdm01GZf8DQLZ6GU0eZvR/7/nO
Pjg3FLxQNwqOr+tS/JsPpFySlN4OHiMT7vc/5Jl69vK0502jY/zYdN8SFY0QB2/3utzYisZqzwG+
3PwCRQ+gOvVsxka8pqmOAOaCnZid/yeCddMw0EexdRhQ/ymn8fkLSKmVprN7TjSUvNIOANUfoRpM
Xa2C81tHBMswukszVcpJkhJ+LzH8fWrX4jI/XH6E5TXrJOSj6Vncqh6OjDWcB1+r38pJbrx1QvyZ
ONdswv5P9ktBvqX6J4zGPIcbR0Bjc9myriH472SsUVwSudbVyglqOhC6eLWyo7MBOY3x/g1RaZNH
0+73RupzyWiUnWPwr2PM7/T38UNjNAs4FhJhUlinUI9gok0YGroCJKdPFh8wzlop7E+Wjdcodq6o
NkDcq7yIjdMXEAl9eGpMIF1qzS7tf3n1ZAj7IJcoWvcxios1VmEJ0xEp4vY+bEONQi+1ZhK9ChI2
3uurgIwImE6ubicpOwVPaVRwE3VQidAEI627SBzXGpW/t0C6eNlrilKfk3G8g6mn+dJ4SlN3iy3q
2wDXQ0ra+NOo/UbVgcPajo3ObJVDlVEL9o45pafLMEqTn3m/A4r227MYGqALFu1uJXsDMOVnFhLq
2CNqQFWgdnKk+PtA12DHq6ci/z9REYCoXy1DIE346w/AkE7CBKFd48I6A15K4RdHcL8GbEg+lgCB
P+YwdykSuNQf1lEwljyd6ZcYPijZluj7moHTNfGGzLpGGKrX9x1IWHzKRlLhrWHXb+meOn3cz/kT
0YjnJU5nrUQuao34mIryiVfEF7Si3n3JRoBeS4z8kpl9F9Y8diEApAgUFsZ7+bg/Lhz7WFeYUDtN
QHzbhCDwtD+QLDU2vEfJAonKtHt4B0Uup5oLc4GmGhnt2d/g8abIl/KFuPPZfFOMKePoejgtblL3
tRkZYJOazh3QQGdg5VpnbFkucDRWg22EzKi+x6OZXezn3kM6f5Q+ntoCj0QihpWUmb7h0sno5LKt
XGAgiT/S+4ObyqViimALrMPzNbxF1Ivr9l68a5qFOzzBEsEnZtr3Mx9sZJ8+k7T9KJ1W3Zc6Ifcb
+JVzSbNNLGTOZvgQJPB/0mw6d2bR/084ZCuPZB+FCp6cDsfO7Y5dNZoyCy2+MMUF92mh9btsri5f
5OFT82N5hm1VFZE3ULiVZDqduu29zOR9LA6MQuEhLpXHhr9B/KhI1EtQgRLVh4wlD+VRU5RaRIHJ
fdN5JpoBd8GfgbSR1b0HyN3CccAc0T90n9Dvhn7vBi7PxtJ0vOsWTbgVMldeB6huPVGE50kIKNQc
6hzt0r6HFj5fyg8PBEUAxMW/Aw64TlmnMSsoU2HmCqRng9Xqw/tWqlgiRl0dFHM4yPxtheEdLFb9
R+EkKwUzN/Hx/OI92Vkp2BynPte1IYalhidntq9tma3wqJiboann0nP8TTsdDnhx74aTDPljPx4M
qxw/Of9RDSWGxzOuIBBf8SewJi4PQKHfKrBEdd0ZD2FGbm/kLdu/brPBw0L4YNbK4v9Z1Bl60oZY
qsIpoUdKAVtoc5wD6dbZlAt8903bSi8f5yhF4hQ073SJVeMLzdSQhi8pGTJ6kUPwxgJpdk+H61CJ
O1/6qsZpLzN7jMPOwuh1kqcTSP76R99yu3QubUJivqjH9zeWDy5NxMJZ5763UK5uzEgmNj8GFvpg
E6s2Fvra8i375iyd3zT+X4KAdC4nSL0WliQG6++i29gw9qIaClz2OQ0liWoxiHkszG5VV4gJOfro
b2aCNrBow0oAhkv7qSC5/xLL6nxq2jFEH4K8LGK8N3DMsA63BSy3sb2gu5rO1hHgtYgAIQ3fKIm1
YS7p8XEatuLdqK3LHByFAJY4WF9cGJ+5WHyomMpGei+1wklDwgsW+JNcIQ51AenldL1M6KnTot9/
+cTYoTQDLqxe306FHRUDoDvM0yeQM7KOal8Xif84lJPWDaxeqxot+y/BJeqdhyTWPi36ULVeUy4e
F45dLDj/IKN+Idwt+reE/DknZ3G4AaBEn9rGTCPpesnPo9w7zNQGngHWHcnnZyjnYmT0MS3sgt65
p+BwpKysrDMgXIYKk1AI4aVbm3XQMzkspjBl3c2sh2daxIoaKXirskLVv7u1IjfqjE5ifMBzqeqg
DmKIDyHrPgtFVP0Cyr0Slw4CH4ubM5qvCldRPSP0ZPMF19tihIA11Dknx8IU0Im7IXgk+QtFS3fB
Uws1jGTCqiJ+bVa81IO2I2gSWmv4QMfWp40N+VpuTH7ajks4zG41XUyCVrNST3S4k7d4iOc7eP7l
sKDVWo1sF55fniSSCVhsQ4XDRDH0SLWF9m0F9Jh4urzyoFw53Zm+gkujDQCz7eZxxGKAJ93+w09v
t5lXE9UNj6UL8DXhBX/R5wSenoHqYFM4Qyo0Q/EvgyHRBSQnip8M8R0J0UNhIiScS8pIQ1cWnCTb
ETyDL0cwkh5c17GKMR3y8h/Q9+m7twF2RLHNtqxNOUmoY4/ZjZe7GDIajLRpo9rNjRnZOzXn985g
wWbIIto9SBWy+TU3vMzx4Z42cOLaOE6QpXvt0+JuqeuK19UijTh4F7Khgs/aC/2mtJ0Gx9uqKgkm
MLMe78Gm4Bfs1/SFf6HQJgbbVzmHboAetthuECWKtGspytBk5WsJDwkgXl3o91865bgXAfhprkCc
2BEgdDFoXG/AzH5O94GJWdNyQ66MzJvNoLp7gn3W4zv9L8IqtbnLNbWuJZrXe5fpbkwxzOPqqNQp
si48aPKg0NAT6laXl8f5lnxEnN8B589uCNLqT/k76Z8yEZ1RXHJk5xbPqTnzNDgc2nrS6e2ScMpx
1rVvWIQKe8WAdv7NT369dSY1a4ZcpWOJ1wjrFOuqt/pvFcy3OaABd66gEbE0xFDBFNpEkdG/nVa1
qypLR7e07Ms17jJ4sO8+3pYUCcuT49wfSsTcBaVHef3vmQMtl2uMEj/MSIEhkNLuehJH2l7aCH0U
ZmVNfQ2NIg5fEh58v1JaeFaMrNDX2ETI/qoyzCjIvl4w+L/VdHodcGe/tpvsITC0uFJ5mkF2qf87
droUG9vCNWW1K10JSCOYAMQR7vjE7mBD0wA864BHZGyuCwnjtXySAvIl9SYOADfmayjhU9sJALSc
Krfs0XBe/buhiyZYItQTmav0faBnxmgpV26FzQw0Bp+5+bNMdwhNHXtJV+q3TnqjU6jI4cX/d8d4
VF6N1kruaUF0aLEegt21XGnnrsXUJsV9k9lcwowIiQdJoJLqkGuYqSSprJynopJBPO3kLw94zQH7
+vanFWSmwqBbbBBzjIHtc119fyKIv+bqHPeuJyYea4hf8sr4hBzWggblrf5apGfdNfGX9bIVW89D
sc2rZm9ZwHKDYEKtF7tJtlND3S+aR9XPsGlV07mbgkE/z47Z+7+6U9SgJUtcV0mskkWbLFIzd7Bc
TTORAIMFicLNmJ7Jogp7D6C4gnRpwuyRMtAanDGiVFbKu2hoQV/R8czQ32txpY3uTAWdkEvfmRut
NtPW6Uvkdf9ga4g1ubBwInq8qOx1CMOjSRAhST5n4fJauTDTZ12ibXSDsezpEOrSGi6opUn33jy/
HSkLECo6e5ufGtkpGMXD5EP0Kd8Ea1seUXIltE7v6rKlFPv1hbHjuBi3oiuT6HvYmkvkOHJ2ePB1
tNucoLVszZtHzNTaOS+0KG1x/rioY/mqkwYiibtfqKrJxtSj5KdKHIk5GSB7MIL/RMBWNELeMQad
nD4alCHxoiclsyV+Uf9BVWzLrPsP+W1SbT2Ex9Vy0fTaA5QSsb2xeHOcN35OWxoZ/0xM0Ldj/OU4
pggbAj6GtdX53/B7r/dPExmOxUPihnJDBh1/M85rL7c5t+cvcrKnXpaNEVIQjuqy87ms494oUsD3
u1Mji+idssIFEj+85prCQtzJBm7++9g2xKMAm1agqD52cm9uqpX7Awl36zXVUdcWnJjmHhhQ/GgZ
LTAcGutR1xau2maXf77mThBq6JhB9+/2SvKcGy4GfdqCEitFAAp09ur4P8d0n1L2zzo/brtgcg84
cWX/MZsYOoY2+ERSGdIOLBlkxWoHvtCiKpW+EsCy3G3Tm6pvYLqD49QKm0DXRJCZfVQtE/fh2Yii
fYKtuySbW43g0K2gXZ1pYSJ0OHX88dxtY3yfPhTyR9PkMMJBIbXr0srHVFNJfevUXghRw8WVLwLH
sLpYrnueCuLug3tcktWeknzfS4X5Fe5zGsPCohqnRcPo9Vk04qCWU7AvuUxXvO5RlTj2uQjdiAPb
jc2oWdMtWXWtVntrFX+c0pcKiQddm96fkCVYELb41m4l3hoqql+xAsvFvtSIs5SlmP33ChzhsS7N
1BUz3NocApP6P/MoJ/ydCaybsp0/od1404qLL7cuH0MkAqSVOsWKl5k3DxIdTX+bIPDzwY5QiwpL
EXecUDIWEB+ahcnfSQQnBCEPudRZl4VuxB11Bisz7+rbLrM8TxpeV/MaCg5DqF0y6qu4vHI3sZ4l
qqg/3QALa4pILJfNlBixYs+8P87ZDm9WcbD/89yeCITyKexsWlYLRgX665MvgZMIgKboYzkaHEsZ
5cLIvSeZI+Jr/6O9kPR6LNhn7zenYxIZDCTh6kOCjZmVO0i2Js0z9VPpRHIIh8IdBdgEPPrp0rqM
NNzkczPgxJI1e8eM8rdNNeR5r2MyNwmxMTwBxT2pj3VzPnzAzUFpojsfuHWCOnhEBKCkKgkG6xv5
zCzA45IDG36eCca9glMZ2WKxaIZok8Jb6KLrv7kIEFsqw+OH8hkrTT7HIunVVsNgb88Bafuxp1fa
SdykcPLxq26UH8KJGzZlQ9iCQX40GBzLfwAc754xM2U4vHaXZLTATVu9jY8GtZ8OEVYZ4key9kWi
TRQaQ7pC+oSS9Un6T09GbjYkQN/m2PyBpyeFFrBuKrQN6uE7LdY2hhR5lnNzmUtwpOq3pgoq6AF7
jsowlOAjv4617F9IkAnUg0hLe/QCg5Qo4N8GwCmDD9ncT3KlpcaplXDbAvmrHqk9iB5Pdpu4yNRY
phdhmQOvIM4W1Gl2AkEDIZOso/2sMU4cvrFoPw/+jUYF9fyTVyu5KbhYMMB2fX0LKML8azHgd8bF
6ZTVxNZ+e/lgIQLVNPsVUAgoCjMMSNhbvBA69smxZynAn5mD0/CK+3f4sooWTizJjhGhBxQlHB7T
ZhzgZC/vN7I/Z0XmWLhjNlzjrE+srQAFHcwvdcUaxpDRmLkk4uWdTmrpYyB5LNPw6u4D/0tfvjJM
22jy49z3RjAWCfTWSJhFpFomOLaKXnU9+osGrZP/DCka7yFbfF9izaGhujMmNwH1rU7VdFDzYn/r
bFrKRzjjG+sK+UixiEx496s3e6Rjm/ewNLUvwoRVAZJMsQf85wJOKs7SYIQmVkmw+zuCkieBvfbI
nUmdh+MgcY4Cn1JC6y3rmfZJnz1dg+/SgD8Np0rZw50vWH6CPSuYdSmUBX4lwrp3PXlAW82JNGC6
w04AepoV6DHc2+Lk2GcsAt+YphWj8T3C80ah63KbM7kbV+82lU9aEUNVaeBozez0EfvWxkrQLNDK
hzPUxjBW2MmjOLmZFz6XLT0PD6WKL5yTiKh+DnuRVmr+U7Zei82RRAln3GumJ8AZddpr4rL+7OAg
Cd1bg8kPdYt9pRyzD1G1bH/jU2LwJXKXRNS12YnmLwxFisQ4jd8DMjXzixNMWL3qP2b9kN593WZK
/LYt7L6QkAucZcQTuJjfXyAk8HWXz9Z6uRzD5rRFudS+QgSsSk0vkAFDtwEDnLmCENBVuxKDZ8a1
9Q89Q8Oksmi6wmnP0nPB6Dz3hDry7Z4BGtyZQMo5dck6JzWAri6SvoNVgXnf49kRgDcOTpoSGebo
nLrAyBQNAaYJ43iWqYtsVNWXWgrE6vGrO/35r2BcalK+jml4oB6cyXx7R6YxnljwA2Br/PS+E1TH
vWOpTbunEJ55CDk98CHpQbn4jBTMyaYy6+vVCq9fuwtpU9qHr7KyYKNQK3XR9zPxfJSPHo0UqRWe
LsnV2uUXFlEwCN+PZ8eOgA/Mc1mB2b/ZDQSwpyghTZBn5l/uIgWOml+nAQWZE9NinWNx9d6Gg/oV
SUluNFfgsGfviQjydvryf2Z98UWSgo9tWlavy9sY/GusYVWbeN/C/PEkryssyRj6pEuVpHuaUZ5p
Ky4PWmR2eOE/BnchJDTkejQ2+80rRfT+AcncRd2WUfMDdMos5nQBwyxvJ3mnkEoD42BqNm6t61Rx
FRru8W4T7679S6X2saaZP4TDo6eiY3ALKebaI9miBewYF5Ey6sahg8yIUTNDW+jrJxL7N/+LFVOm
GXk8j8LjsuUwA9B1jdctsLcYbSeyMV6xOwXxkEhB/AFEUVvmEzcjL1ziO4BOKN3eGqcsIhbl3fjE
/b8OhPID7Be4Qo3KwIU8VZaFRPlpv7T/V3PNDvAPxpoQTSY4Nf54kWMbz0d0LsF8vHbNv1rz8dKl
WjoyERwgi/CJ5YKypM5mRJmqkHGpN0YrTHdRS5C5zJWiBHRZv3SWKOqqQUVv9QygOgPJ3/pn1e6n
CBIY2TiFSJw0NrEAlV5Yw93xR3ZBvnh1+NeWPJTXwR6ER4cXKnMZtmk1CESiYgESHrYd3yr7OcWI
RsIqfZp6F6r364wA4LVBmPUYuHOD8Hs6xAjmTsIxgPcQbgcP1tnqwXKtZDVC+GuDzph59aRx5p75
HLG3JNsgF9dedbvTUw4llVLeytP+RTCDPhUfwvqpu6FB7L5rpoDJ8QXnJqJmGwcC3oHPxXlYCetx
GbXn5tXKBCgUo5d4pQRFLPHv4BYAFz+S39o2FRabCX9t5mnr3KNbL4LTS/PIPFqj//IzKb+A9eHr
Q5uK5+w2RypqfNbUVWqZgFHeKVCaRiTfIY6d/mxjYDwwvB8Zx2q8R6Z4H8M+BGzWvIysXiQTfMeC
psIL1b77n1ZnSyXFb7tfEDL8F1/J1LhzL7J3jruQGki3GxkibrT30146wb7hcpC0CaD3FK8gZ8Hf
9niwqwpsHUyjJe9D9q00H/Wzgb04KwyJRBDByMgPxfHzJ0Q4hr38Ey78We6lf4Qog4IOwmST0FY5
ZWyrLadVLsfWv+K4UDadYAsBy2K8lIlCFdVyTJhTHPn1TgMf1Jd5a0ZiKuA3bHz6H7xnOzQC2pqJ
muQHHJuqUXz5IghDonA0Mp6DxNyOt41dTYn5/dFN/PhQv1Oltt+C53H+GDCIg7DW0vlSTCw+pR5F
skKNPmLwsqwtDBtXEBeTj4ExjHcWqXIMk3/ob3mpvLtJc1itzmTvwp2uxZElWtjPZWxkDfA2bT20
2hDLsE2tg4MLI9ndX6j6nfHBYYPlc52EeUjebrpjY4npeHN5dNrQkXnlt7+gPQcBAiRP4+yFGVto
JEeuoqTQ8o6rlZ84UEDz/BwXkNfxjcngb/WSovQt+TQjxrEipOZW2ugrepGL9HYoQZmYeOijcWj7
xJSUSjhQKisZzsg2al6c0hzVT7pjDss9kbsHVF86S4UiJ4GJtepae1yvyQ/iix7+9uj1NhMKmMb4
tAVGgYZKMjKEjuWHtpSCa0WpT7xV7n8fj6KXCDbyiVdGaWJWdmtpGFytqi72rwAByIrKgr71PPIL
qIWUqrhSgclEv6x6ceQzEZdTcRYwawuTLYoeVYsHTpgHftRX24RiNc2J2Yl9N0PP+QihCyhuTgGP
oMCs6pa3vjNoQBqqc8gavuh+2fTlkGAOWeP+qydtLWUcZEdYxNTdJKDjKpRNrHTmi7P6Qh4YbyU0
WSC9FuWHvs0d0oSo8j3VL9P6JMDuktDzVWSrgxlVtJJ32XFcAvaG2mzYvQj6BCIspBQNHA95203r
egqHDKR2ZOj9+BsyFiJ/7v61KjC42agoGhB10cbTQPtEGrXfkPaeg5QoSENE44z2MH7IGuoToXtZ
ER68VNiq955JQu1767ddiVt9wHp7EgZwmxvmXH0kob7Zw41wtP1/Yn0q5V0fchOql8bCfsAHaTfh
gLltQSq81jJhxA68swxN/NMjpftM87ZjZ7DFPWyXTltVYxVX3Rv7Hpw44F7CInmWzGnCnUl7p+7f
XqY0Tz6MkkwJMDmNL3C1ooF2/1VlIuyYdsDEHqGYG8vgzUg4I1d5akaxMqxUjEHNdjWDInUnQeC2
wkZW1Re3nSkIHe7l7U4dbnmnJceyMHWWmkzdJ1zcmzzlTx5p/1aX9D5D0zfZ6cRZ2zq4TINCalBI
EgNFYeMjjfD8cZQrPf1BU5ZkLJiDAjM4DYQX4xfZjAbrfi4AARZQKXt1MLd6PXteRcpp2G8hGlhV
Pw408LJ3GOt74aeVRgbyAUwKsbyX9V68vx7xEi4xt6N8hX8OZnlBnOjO6nllA74Ta0yQNstmTJtb
W5Czc9hNaus4H+S2a1EGNeHV5Ip3O8rNv50Y2RTbZr2mavi5OU18WhnGm66cBvueKp7dN4umAeI6
z6a/K09apuUki49wMwDAKt91xE/6OYuNNvJCilE4eX3cDhYsPRc/o/4ICNgbnPeWaX15JyqknsqE
I5jviWBvdG8qvP2CVNxrgWp58D4rrW9r5JriUH9CaY2Ow2bizQeqDLc47W4tRjiAstPf5tNRDZcO
ZxrF0mxmyfSjhy28DTz2XgasNeYName2O7xBneQ8MLjbonPOrSGKwD/v1gidQ+dDeYiTKJ09LlFH
IIM+YVgS4onBxfFnkQoXsSWo6EEKRHgAP+XGTkcGcQhWRYhG7gKmwATK3XQJYzCjHZmkQQdgzskO
NAscN7Vgwutynqf1ZKa78ZblFU1DEb1ECzoPBfOvYATqeAXPE9qBfBRFvBbfj+qld3uYPsk1ypYS
ObNXL3/zVfmxO+fDDaiHr/CC7zC2f8QvGowrYL2LZMmVj7o9REJSh14bDprPtWIcraIPXs3ac76m
KiFfgTPlkwPEXR6L3XAme96ULbyUo0lLchcUscqD8CScDFK1+nKti7cT+QsUdJs/bwt9OOs4yosK
1cT4XQ+GYtOEtZfNfRmkl7OYv15zttupZinFaFmxbLTRBO24BsheYhdkRNlWL+NCY8SPpvLO53ah
yzSfVuJMdR6l9NTOgovCdZ2tw/JW7QMoCmz3tMZu52/qwce1XKQCrTZdf/B6oq5Xj+U50v3dT1/b
JMPsULXXGIqK2UXwL27Bub2DzAxQ0qd/fWiJVRhVEkXJqf1yBqrBV8J1eizhliBec0WlJGD4ANdB
Fa4QeBlCMo+szG29EQWxgWDZ1XbZfXvWNLaXhVcnF6navAA8Yg5eSDYIqdHvqPgZJ7H6pigZXMq3
gY1bjjU4wJwFB81UGbyJFhisrpnNA3qYGj5I5Xv1vr9DQvpu+Kd3YEx+anh3JCmD61N07AISzzyJ
dOxYV2RO2mrjSO6BMebL8V9Rb0H2kr3JOC3QXOKcPTq7kyyKGIR/2mZeZxZX5ftvm4LUaFhvzl/H
RrmcUFP6ueYcBhUSYFdUlpkeOS47QJCHflE9uBvbnepJhqNImedR7ky7BuADlpjIH93OesxvpIZf
4Ejcf+PhkFTty2WHoGP/Rdvf0yfFAIISfdGAhFcqluy998QAaHHtYDYhab4+2TezLoPSXIRMHSJy
KbEG615t0YEaHk7ooADcGTDw0aXLGQVUbVg988OYTXwZfebh6AUUxMq0bghL4sZ97N2mkuCqCo7X
MmwhhuA/2z6NhN16XYr5d/xRiFzHQ/tpusKPrfgnqYHsc7MNwAneX3VuEplKcYeyVPtRhbT5y8Hz
EqEtFwFhdpvQo12IEYwvd5GeWza+V4oVHw8m3zvxiN7zeSR68RQNqMc6tDJ7psi1Uv8SBTRNlkCy
GQ8gaLyBL+Y/sYpH5mwqHnX5q9q/jSfFGGPg1q1bmC9sSYZIvp/GA6wF+iCofjfTH26IVLWS6/1a
MMdBwFNj09pj/LXVq3X0ut1w3BtsV4T+o/Hd4D+zlG6sESPzMUq7rCV2I3pWzxTzZ35dTlLIz3CJ
1zLaR7t2SMB2aetJE9F7H2JMVI+XZ9BtdpLVTMQs+cTiVWjC8VBvFpUMi0VEdwK6oGhY5mob0CF5
6y0M2cJIqmMfInipYqBM+3OyeVAffeIqlqol/grGZneU3jqR6UaaLxMpws8ashq0eJDseVWZ25HV
ct1HVzc2try2s0JzC6XAcyRiz4CSE8QYmhfBZdyxuTI6Py5j3Z4KmNemrkUjUUWzhblC7cnNa/PM
Jq7drB4KxQdgcHIx0mxYVHSDnC4laMeKXD8gQM8J2XNZAA3WXZXHnPYsEYRDOdoqwl60xOGLjRxV
hVM+VQRpzw0GBbm5VKJk2/LmNa3usYoBzuYDF9cOBMBqaOD5RGh5aQs51ecM743/mkdjdpTQ5VkT
ZED3vQPUQqho56mtMAqmb38ViC3boEAOrNQuAgGc/4WdPm4ctdvr9z+B4lRMxC0llF7sB438RZIj
iURDJDsOMT3qtG34eQg/P4s/p0b618rdu2R+Xe9zhSGPpxnvLzq2qJ1VKKT19yDfDHWFuKWILE2X
ly5tDzh3Uf/boSeWG8WBq7emUiAZvkvJRv02x3JYa0HdCwj9hdlAwQG6mJSM4PyV7TViFzeSYhN7
M/otVXu0NwX3Wd7FchhyP0/yTGGteyw8IFVMseRsUsGSutHJV7mDwgFQkLhXYXvALUx/nmq/9Kov
qeYLQOcPUNNnyM4W4/dt1WpkHv/0EItqPAMaWFE4m4O1C/1cUV4Nt6AzjbrJwqRu9jNX/HI0k/4z
XtPdpbRwDQ+Nynz+Qsm5Kv4EJZXZS7VVM7VFgkPuwo+iMepydSzVP5RoR2Zr9b8JHhMMFF3oFEJi
QFchS1Spq3J18Z01lL/jTDtJvlNZaeTE8s131t6cWJfj+7Y2Onspjke4Brj3tfXksVUIW1XeD1s1
DwpmMHc959Ju/9B8klvpIJp/t+kEi1OjPicIpHSF31giCXIrqjQsnm1K8UjdullK/ApQyWpvTW66
0Kfd3GAFPYX66ojvKwqKLu/CcVajE0WpOFEEm3S6ueoWugmZg1wJFx8brkdW3HRV/J6+AYr0vKIR
TkK36aMwrxHKDxiNUNrw+ktHd9+9SQTSTyYxxq9sl+UGljp+5aKte5q3Qvc02/URZ/b5YuF14qUb
Dz9g9qryHhm9c4HvUmwWOEh473MCO4hbaVKGrF/1Xq+YKI3U1G52UbMIDqVgKwdl3MI6e2SGwLLw
bQgbjWF0BlzVAjEDVZ2qZ3dUQfpqurWkRP/fdevIS0uJc3m6Ut7G84/m/C0/OLaOGW3MU7sHQWu6
XanCfHXoTBAbe7iZnrC6nBML9l/uBpqsw69u+zt5XafFZHV1g5nstv0WhgYAOrhw7sThpx4EzgjA
msw9IBjVyFCR5b6kBrMJOgKnD2n+Znnz039L/cy0o0RPPurTkwIKhcD756PogcxwG0H/Nf0m2ITz
LHk4oqpgtkG7IwvyKQn9CqhfCZkye6D5VwXkjfpwSsMSo/4xamzmnJcNETFHNAWRdZt5wQyI87ze
idEGBsqgtrVkEuC6+8IQkRlsxRx+L1nl91DIIqP+XJs1VvBMzaVaq19EH+Zr1eFwxHEQWL0BrsId
kJdLlWVgSkKi14NE5LgWyxgJtc7Z7gI5yIAGE5jbRFoouMkaGdgwYNEg8S7cpoWUZHbBc3shR78V
4JCGsKGrQb4vD+anE36hCPbeJgTn19yECqU1b4r4cESXp/pn38K9VX8wKFNWhLIjn2qUZC9eQB+P
y/ZSgIeVnavKkvN9CaIrtK7Yxj4iUk/Nmjs3V/FLXqmGCMWpYEclFnKo64Z/X6RI4Pyyl4rdgFK3
YarG4xSfqiH1tyfd/oTBG8DMRLnEAZuCQw898S2dmY0xG2Duj8OW05FgM8chp5mxpOIfvCpGqu9O
5l+XdqSXH0yScj9jXGmfmLTDisLRLwbI2bBHi0ka5zGLxJsUnZ4b5+C8ESVaVC2TmcDb2e34F4WM
jK1CbKuawfZEfJzxJ7gYdZT0/CmYY/AH8ebnUCON/EcrJExjR57tJ/vNzs88xDNoU88EdQBgvCaR
Bldt7a//KhMlOaT8y6aeDmGkzKqtZT3rDJmTeI6Uf7KzcQnzMNAyXb5aAYTlZO+EC2clnZsAYmrL
t3zFm+SKf/Y+kBZi0aNfvW+oWSdreD9xB2t/rLqwtVaLBmHaiJPJ5YQkOeyByE+8DE9dkUlpJgzu
XMUP/jf1evSN7ehT8h3kutx1xvT444JZ8WpF1ynCUfxKCZyxdrJSHiE4hSQhvpdDtayXDh5wxxXH
Rvms7Mdn475xrr2/gJHHD2RvAc1Dogz14w2TpSnstzySNVPEEUnYbatQcTA7gJehpIt66pmzaPjM
t8F8MbNaBRF1wIs4e76Hyou/6/0WWKn1l9+6DrOdyvFk1/LPpzSoIlxpJZ3EiQKekmuFsbDbsJx6
/bIk7XQ8g2WJmIanSiY7rNhC2jnV9j6IoYX6LsiM8PEEgiZ1kUHlYtG8WyVMPPNqVVaUAjgX1t/a
WwWgwi271MTe1A78Vk69/YM51qGZxvqLkqnJWc6IJ715Ue+bwJdIUBqJuAg1w+AeDhbqhx3TjSCO
cRzjQPctwAD7YpxH45uGOgRggrX1Xxntsj1H05zFNpFgXZVdAithm6tJu8VwNG6SnMULocG/Gcwq
WNn3W+VTx4SPPEc+ZKColbXC5/KJa9Vd4fDwe/QzgiB+1KaDV25nVTzP27TbNBaDKikmhB4BB70E
sPLTOL2JglEiXNpKXd2HmlYBC5iXYQ1hq/vl/RiLxZ3qR6IR7seRfdwHe46DPp71gI6sQeDSXho2
W9qJXC2ikGoqcwm8sVCM96zbzuo0epuncdLkWUfF+12pcBITXgONGFR3oS06pfw7Qp8tMlefIX9x
CFeBcbWXiqlViv4q+tC73DMgKlG6f9Yu3o85ccc9mcNNp5ahKBEZGKvmHQeUJD6rT/205oHnv6Lr
7wY4bfRRipRtUH8hm9suOfPu9kTCUPRu14x8bd1av+5YomTBF7S6vx8iSGMneStzvPPLweNcR3pM
wOOJMI5oX0jpvEMXTpSCb2ubj6Zm5KPgP/9V7/Hth++aeOGrizNvgwBi9cqzpsinLopg08G7IoRh
Zx8eLqL+PEbY4X01vV7v6csTlt1RzotLs950I39EmLllqxNiM5wRiIg3lkmbUDh4CBblnvdx0I/h
xBnu4lyMtUfD7ybLJmR8N/4zl409e48ypbj+uWGhRxnyopSSf/DHcHb9H1bEcxRnZTZzHxQ9NcM6
tjhauPSauaMRvoaWrIWABOiJ/9v5HQprEDiqkupbv4Zz3rgWVgEKuxVky/+ZnoeIn/8jdMpJwGOE
meTdZtZYnnzxu0dpbPStCNhKQpi5Y4zDMQybcxbDKmGkCMWCTGEfjHSJEfr82mdyZsYsHkYAlBZg
n6EE7eLmmn1tXj343ZkX4Dppak9JKu0wSMCFkVippar43Zwt+zg1VidDD54jEZzyMNNyrkyhIv26
aUMvv6iXij6a9/rnpvXoOnRGWwRRcKhlDZi7EUwjBbcjBoUPArp7TFhrw3UHkmK6vN/I+d4JsaP5
9JQLkjC/Zbi5fWcbuzmaANXRg16C59I9c2E9I9+txNo8sH3C1ZgsPixtHsXK8o0y//eSqID8cuSK
b3R3ySRd0fN4qiXR4m63g0O+g5uoThCLO87vvwWilkQ4Uk2ytjNFlbIpVwNGs2JSNlts8/oa0Sik
rJy/9aQ231LUJfouqYgrjnZaB2qjLlKgP9KQDjlOZ7oJop0F8RMxwtIxPDpkpp+8ovu2hjX+J8iu
GJaWWI76R/3hEE09iCQYRZI3+FRfUjBQ7XtoAOM16RjWwQBUjuDY3QU6x+Cvpo9aumJqh8oCqgU3
Ff03Mh9iHpCCRMEiSWBiGrE4nfeyHbzJcuGUIJbwDDfA9GGNAcJexflTen1Te2Pl9eQHTiTp88XC
32gOTH4oscTDBvd8XTmwFU+4Lq692/8Oo1PmH5BGlxeBGHBzTH675qyuMH+2152dmsBupogJRYHx
NcOmpjgASO2/5kd9/yG/JBnJZgpEyFuLd5uQ4upm7N8fsAHn2sDAxNewydCcVeEbDsPLT3hSg7m3
wn/UfE0EUAHRAZSyM6IH2CO7r+XPHrL7XTmLP3bSr1orHs0lxKhoxn/XW83t/t2HxlRz36/Yecu9
Z5aUpWiizyV3gnKco/2f7udXqOGRAW4wCXwl+5kteGVfa73kmcFlfOm/qHTIDjnOQLBk8iIVhvdO
bJjkCXxDuh7tduIDh85Efuns2rbXid6T8ohxdWEHwglayblhwmnJZe3cDk36O9huvXIH8lA3ySS3
hdQhCfs0THYkmsqjb69J3hnzTm0uMvlOQ73PdlxfdS0iJ0u6/jZ+5Wb+l8GXXOCDgPkHbkVCWM8G
mVUuwyMRii5+vOawX/b7KUb5S6HMeiMnPgcQJXKfRE/rhT1HiPIj28sYEJeqWtH0VRd6ADFdXwPq
wMCuGexfdUnwKemfbPccPJ1gAGT+LsA6LezemNW6fy39sgpomk4f8jwWzgQmGlyidO/aHYEnFKY7
DUUilVL4KkLFDgcHnWiul9nVN2wkTQEMsmScwzj2x5Y+4V4yX58rZvlQNq1MGeTU3QK0FU0Cx1pH
DD3L1t9wp6UTWGI5FuLQ+T2DernsglGHDRC5OhGkyEh30njONQ0DvdsPDWciIsxPq1DbPd4FChzF
nDKyQkKe+J9fcIrdEJkqW93LX6917s84eBjQ3ZlVdwDejiooTHa8ejA/h43H6GVmNR4B0etHGOV6
4iNN1PscBtdMEcTTDj6Z29czeHrs2E7wsFURxNidiOLJyNQkKgbHTRIjgomlMau7c5L9zZQBqN5W
5WtL85n2d1Fz8SoX7IzIYdnLAUjS/SJ7k15e2pNIgBafEFv4bZcW12TcnKlcl9bLYTj/vhNHBFPk
u7cEhSF03ZPmvB7xCbFctB03BoUfedfZ07UMydkfInupVUJhAzk8iLVJcVWKPIUsPmmysxO6BiER
RbI7xCRDBTx0aHjaVudy2jrU1ik43RiiMbh7MBoKhONrEQ6CWARCixt/1eoJM39DD3QTrUNG6j3t
OmslBuTtCBP5xbMvBJgw1ECAjagzvoWkg+dyy3fbMxdjXTwjBJ8Qhil8s29YjAd69T1CxudSXEwv
ZJi+KHQlL+SOwYdAlb4too1Qu/GG2dCApml4EBlAUktUb20jkfSVHNlVZjIbcjqeMBxf9SeZMh98
67M8jXDlICugfPBw9r07PyENhTKj1ORz0vpmRDAlo/QQkLDpCvLciKKaFSqvGGPypDZegndEA3nq
uQhrtKD0gAvFXSq8ZCRteV1qg2pcUpJNmP50zh8Ud/oiBgHJc0l3Yhd97brasDdW/FqBuABjr7/j
OAZjDC0dzDRBGVL9v/UAIPLf9fdIK+VZRijWHViD8xKMC87RvuP2lNN+V40fu91aUgTwU/GYcFHh
w8rgZx9J8TZJTO4b3xqcDaHCoVMdVa1Ji8O0wgrE4dx8I56Y6tgIyj9VHsOZVSo1ga2cZFSskZQq
4xuWtdCeORsHtnHYcSZYGvc2vWWIhj7Z0+LeZY1DEwJTwLEr/N5Q2WsxzUIlN7f7sHJ2rio7lfTR
DQRdw4Ff31Ifg+olaGXtvDVpP46qIdCPLoM2fBWzrFY+8ufGPhsScnJTdTIXotA7OQiapFW7aHUt
ZYEAVQT4a8RdXt/i+Ntv9G/yTRLbuKNibBe23X3X2pjGgMUMDU3xOOiPjb/J8hlXRlh9ZRHmx4pz
rWXneH52wEX+Jb0z6NAL+XeGEQoS2Z7TxZr2l8QPMoTJ+Fzg2Al/VxkS9HL2++O+WOye6IJYyYaM
Z94VZvwx1SgLz3KO77lchESgCbVDNEVTZKywI8aGGChGCsgSVPUyJI5aAWYpOHY5Osb9ZLEQmYkm
tKYBpjZA88kfBqmaURhR6Aze77sX8Q7wz67dMje719ALJrijiJYu6KhX9ndzqkHRHfF1IEd3Hbfv
Ikh9LEsAhhfiaeRr89Mrtx9dOhr6U6Q4qHHZsIoueR/nr8ipPHa6T3RI7J2bJWp08q4oq+GRozpd
HHij1wJ4qTh7Bz7AYI7MX2w23u7C6vPpP36gR54vEMmYiflGhtDsk/FOey8p0VvKqgzpXtiIADs2
MkUKNj0N/54bPgUiFFDPkpNQxgdSDgfZnfxScFZRIk3iv8IXHfInUgAQpKCw3mvZDsuaZizsZikh
//cPAxRPQ4Rqy+9DlTc4evuzascoymp81dWvIDMDl0CJQ0QPXF0nV1O8hKT9Deol8dtDoER5hYqA
2n4c5tEB7O/jVzWJ8nKcsbP68D10h9ttSUq7n6Xhs6bj6oPCdNjF8msha3s7NKiO5FE/S5k5okvd
byQ78228hw5JE5WPBHezph5TgAm1pfqKchybeNR9n10k9iSQzX9nqBM2Py2txdrKGFEZhkSCEl55
TlKGND7fPRD8ach4vCzjcEBusLkiQHE4XzS+LGQQsrmOO9MzubEScZfn5BLGPpqX9rX63aXb8CSR
NZBpyKFwXUugpZHada9DSmbw6uzVLBHscJAH873Vg7h9FKXVB3vP2ySjoq9UvBxPQ5eubJeVKJhP
MAxG8q9V14vNHKh7UhXFxDOindcR25Jc/YUAzP5iHPqOXYeMG9BPow3mSJ+fMAPLldFUVuXG0iIi
EsT6woJb4+Co5aY+od6/Bv0FQWA536Q7dcnjF0RzWjsjLAcaIVrfp3woimvZYB9G2sAgi86XS7d0
PWlbe57iiA40sDyt2/d3gcAa0bR9IoL4cEM/ujIh996/FHkRbBWnQa46WmoFZiCjmr64tHDmXFPH
8CbbPmV5bkM+mIe9Cs4S29N+7q5KGswL4BkjUeq32SKyFcbwIw1Jtmo9FCOzFRfLsOizs3IEEBO6
u9HtaUaCvwm/K35LwubCCDnXIo9QymQ7JFDlC+DIJ4X8NkYrPti4fM8cy2ypBQQPL9mFJ9oX7Jyy
XG9n17i8W6D8mr2MDaWJyTi8qtpSrA4+jLQSUBJEUfMwJjMBhCyBIfCazv5MFay2XZndQph4X4pP
KgxRJH7IuEnr+fNodmpBfS229LL+QHUVkOUgDfA/q3k6N6/I+h3ntHn7X+lLzPqaj5Oz/a41VsK9
ft9cdAdIxD6i+TLb1LZWa2pCcPkGar1SDK694mYWR4sRudsXb5+YUSD47mIExQpt/moxx4u0Xlbo
NbYuxOkhA9K6B6ZqJSA4ARqa+UgPmFDzt9fhK0YlhmjmEXdh/IxUlCyfM4Bq9e87yj36X0MQuCc9
bOvgICs4dSgMlbd0Qv+HfNS1HPHDqGBzusOb169gg3liaktlwZiyGIRROMqZdvwA4UneS7k1CEAJ
KuEz5MCJ+xHwvAuySGWcL/x9nAc/K8fbuTGsHgng0BnTEztofQQXjfy8aQ0xm8v2xKg5pVgwP4V5
zhIasfYs9wDOMdGO/g28d3NFlCHx4vzCourqQUrcxXdGv2sv0IMLxSz0EHl6aOvR67stVM4P0K9S
ri7Azk/z1A1u6ZHmvs7cBYIQ6SdpHoGnX4YYBjLLw9IN4rSPemc8ayMCOgIft+juvGqgD19ve4no
klAx/+7IzOiM1HA1poSEN/38zEdD00z213gptkImX6cBCks3Iib5l9hx9B3Nw8sMpmqVVC5JKI0C
03wM9mCnknKJmkCo0IK2P1OoQqvv1l9JKp+UjuCEz0veROatqvDVJN+8CvBEabuH0Sy7PlSEeucb
+4TtIRyoxGjDdP2D9c7qv4pvybDE8mX9xtN+7BDMbnKLtmLXYEHKKclCuCg5bAVMvjX4XKgT2LNp
4xgik0PZExyGnBEUL3LKBWNKMIz8d+Rt5BZ9ZngW6g5IY9B8eLeSL6whuPKQ1aDY6JAIXg3bmvM4
LvINms02gHE6FHjsEQR8oQp3NP6c15fZY7BVQfpYbZIDxzXbtdsA4VTrwNf/H+EOg6Iml/YMAgvk
bd0/w6e0Ig/my8bIjgZ3gUQQ3iAnuOtKuMmse1ROGGfFOMtZcfRb+yk7UzJTmCLcyG81FEPbPLd2
faopcR+A9qcCWji5KKVmw7Et/iNPyLw3Shm2LkAbt+Fx9IG0ezkyE9/MPgVgM6jfUOOcnx1MdWqM
GpqTPGkBR0+U9wsKthUfPR29opxQAktrgcRVJ6kV63WcgMLs4AdknyZI7qkarY4mEfnOk3gnY3UZ
lSaxnF6TWj6hX/9zHnthRpTZcPbbcLsI4504jNLBwHyBQluUJs12LbrPPstp/X0OQrAXFrvnfAhx
I/8sFGdyfAu6xeMzHdWTe0iHwQQ1af+olbbg8QyE0/MvMluA0TmW+VKl6oeofDVlx0XLiSdEzBQO
0QCkK9rxcyZfsSb3SBH7WV0kdFPcHij1PbLyOpVPd69PzGndgaaZi2mBInN7WfwrlLXksPKRylrF
uaz7HjjbIjKZAISlZawE9g8udzjId0c4gzr/vW35EJaY0UEulC47fQLskeodRPY2WVF/63SqA3Cr
3BObGI0RROYVwb4lJGj93eKg8CXGSgtW5oF6pw24XMmXdmKsslFW1aboMbp4Ktr2CkpHyU0tRnUE
lPMyn+LU/Pjlvt2v6w4kUeMQ8sF/6rrR0mwkn+t+gmQ4aVOCY0AJFP58pKrmniQHoOo5RdSEi3cu
EKPiIfwN9qmVBAkTkb94qmhTps1ggIiKJZTR9kb/gyWri+9XI5xG+KkwHoojDXNNEy7MnPOodyxA
sYeItwrVAMZwQYKajyO9fHx39j4PNpWtrvSWblGp/DeRGYaezzko6cuh8qlr6SWZWVUT5MyUFxhU
Vo1UWNFqrbIuNDz9GRCC7UPDBshwvvLFQBVax/xRpj7/GAiFThjOWtdXV5dYuHycIx0kWW+KK2R0
R1xtMhD95EWoEYjuZaGzFVFUN0B0X2y11Cwkp3MBpzkZu4YL2eMoQuky6BdvRKYfh95vZGNXMXyi
TVt6C8R4smRt8HL/A57vmjyjxuMsXq9IQhr4ZXJb8SZv68zpw0nh3DkddnBWCq8XWCPDhmp3msSL
vbhZQL6DmXR595giKugTzXfz568Xn2r43ABywRKW9p1DmfNjT54InKvo936ITwVWCagZZY6yRXCZ
JmBls8hq6p0ujIgUNfsp9R+mWEvmhKPObxaLHDeeNPyZz8i3WbwG1NG+FxP35xw2bsW5uJuoU8Op
GXG8CDC2QvR6f1RSdymyi3ptYupeUS87VjiyZ3IEAX2D/QFcDSuVXkyCgBs9BUoX2YNkWiF3fdg1
06KCEyt6/UCO9efpEInAUdZySCVZo0zPvVM/a0aK9ws7UG/Bi2rr9DO399FIiBUvFT0A48gNZHLI
ZZF2B1cxhOIFxK1oMWWyL+/X/OvN2cAqFQgkmPvbXdguxJinMga3JrlZuTKyI1vyBjZ5JoVRxQR0
RNCdtc8OOlNYnxXzaBhhip9BX3cf/rDuun0CC6SVtbHaoXlPg/JwdlkAPTX/wxBhDSI1B9bGpbky
W1CAeJRW8MGRJYOR28VG471gZoWmtVPZ7Kz70nnhCw0ZRH9zAurky5+Lo5gihQG/ep6w2XhyIYrO
oML+/6gisKzX7Y4ePU3MS2wMl284ixR0n1BQK8NYb0en5/Qo59NVgEBgCSClA/tVYkDdPZxjA63w
CIpIIoYtwtVTkFmA6LdNPrclhggZ3T/KoMDDJvSXGu5mRsRL4v5H8Gu+9B/TJeTAMti3xVv2APP+
tkNjFyMYhjVreBO3qViPk6dacmzEr4ONtHfe+VsnV5ZZ9KhXxvlAj5xAdbEtsg0QQYlFY1EpMLmB
fYGdX850EMlss6RBzHox/riI2YNNF1QhvSoTtUSp2Qfptyhv0xyFWOPHPmLuAxe+LAmfzzBUXhH4
gu0t4ea74yGNuh26r5+HqnlSnbJobP81WY1Bt6j+8C7te8c8VNPrHB4+nJHLVfbvCHR/UqBhkJKb
iC0rVxVs4joUUxoDMQlZtD62Vxjk8i1WZZ/XOIhR0YuTD9TReUUG18RVE8sH2D8va/jVeRU+z+Uv
kprMmYZ5FS2ZUPNxQX/SHNgtBwHif3NIrxGHeze0xB/hwj0m0t4pTNIe3WVPBXpaIOtadkCOw8L1
Lv1xk9YgkBHKUFUeSpNm17mUDBwE6v9Q5SBFZi6KMEjYj3jpAqSa+TJ0Ar4N/NkYecIM7+6XBuDf
vLTUaqgrSxHBxhRT+F2eWMzt9wefgrwqHV4ZR6O4fLllRV3ClPDJBkT2XZX6yrar6n98PebuhwCG
dS+/o4rI2hO2YsXRnK9f1qFbuWdBMcCtocH23GZ94w5sH65JFmnFsiTOKeg7sUjRjmqwAAuuD4D8
TjvLsCm10lKT0hA/Z1AC5dloSz2IOIbrFh877tLplSJUHfgsNOb4xWN+xUJyhPxsHH4GFmfSUPSx
m6dKtbZK7Fy225L3ysRx7x24tFBsyOLEo0BwWMRkmnN3F2B+7h3kzSSTCVNXUd087XWgezpDnqKr
OnhE4AUW9JPpfWWjIvFRu0S9LUYID8xpEr9kqrJNz6JzEHsn7MHuhilmwgkSPLREv233TfHj9VjV
Bs3wTOPbrWCMePsE1VychZzv8B3cZw0mD2EKUmkM7hVIWj3MyRg5BNjDniYrH1KP0DIxcTnp+K/p
vtNz9uMIK1R4RcdTH8gWorXd/zKOzHB6PdYmF2/9OLEWXZXkOSBvQiWou/pu3W8nEMN+CDDVPju0
qUYe/lIyp6VJMNH5Zj9MaQzZxrAvl9g1WBfzxmcTCUACkUyjfayZMooOXxQb/Z1rzO48uKJPshgH
I0pCwRYFToIVHi9SbZxKqodBN3QezFHDnYbSRfIe5zPn3VgzsmtVI/u1VPzeOD/oL2A6hMA79fri
pHnqmj1by5P0+VBfXZlK9/Mawo1IG3wmiheST2v3BPJB5rMT+MS4oMyewN0J+3OhOhBk9KuKDE3l
J/gffqBpBi+Oorh9bDThLFWKTv9JGNr49V/fCbiR5Pl4Ob4wHNARegxr/UmfNfdxa089kOCLU2un
Pxuwlacrr5dGfc/LXEh3MiebRpkRoOfHr7B25hIu3/g+yNPENzVh/ssmq5CNjPyLAd1M5542r4TQ
wRkSamES/s0M252qvwJaQz2dwB/7IwQxqaeQV8gyAvJRZ/P9HgHFzeXwGNcV/ib0nO9WcISVhiUD
9TPUDleKVS/3RTWM3eNpLZU7zA/oXuwEBR152hWAWs8ekMrNBM+qYrpm5YZFjbxhgS7gGWv4nrVl
H6YbSdftBGNgcktVNGwmJ86yQwFdh7iNneOhECh9nRVJEt8fu5pSNuJm1awvzk9iQeFu8jz6Cd9o
QIAfFnOMWHdfgQRv780E1p7KGeFmw8bT8yQ0o16MXpMvSmG5tgLHsH6X92mnnDrpXTqIxLs4I5Eb
V5eCsbxfFpA5oCcV7gSHFcEP/sBiJC0JGMG5OTEstb0g6pSWCys4xddpLuLd0MXq55Zf2whi3Ic2
mvM8iM+MG7LGiwp1R61yLRT9Y7JOBDvS/4zxOrMRMVvxezKrzlrjICDy18NgVuT2IsNfkanBZYOS
58dz2Nw4IRuAHNZvr6rfAXdDcneqU18bTPI6u/Zw2XM00Q5r+KcfF+q2wsSl3yGuGA3uvw2MBK0i
5oG9yfeuGwrQ+PYWf0LCLIx9IGI8G3LKOuTbvWjC3jjHCTCmIFt8l/UtWpKN8gKyuQVqLR3n6Fwz
Vp3UKrh9EJQi88RBHxh1MBfpFyuiCWP7OkMljva3b2jRKBnwxxf0G2nCcf7lDIR4b1uYpBsVSTcE
IU/fYbyPZBrmB152UFhBC0Ca7lY4jMCDoVv+BWcYB8rhIGWmXrg7PgnKVMA8W/ylu0s82EvGIZkX
cJPqlMjWIjmcFCQssOuYi2eRDkKYv0nHQV3yDxC73COFybs/S02uBB7b4jeBqOHvjICHssRmj6tw
QuFXAmQ7a1YlXkqUR9DBDHP582UW53TDCuXbfRdeuUQX0yYGNHTXu4tGXhd7VHkK1j36RzApZiYu
KqcM6ysY/vk3w0LL4nvdK2JkGIw8dPEMBvQUH0lqaW8M4FFuHmYw435zMPapd3arVoTx1Ye9UDmZ
lVmm3dYCGwAx5zt1L75DWx/JONUuTp5EGfYwyOjsKP6uDtXm6CggGmpLgQ2mgjZqsZSN5hbGFyG6
g9dH7wtWz3Qnq3n/vrZ8C+6sJn8gtcWXkXHC+NwD0G44GSrVfymWyaY4y1bfKVFKoEVVmy7kWTJ+
zvq+enbazzRZlrsSqQIYv55KJiliEd1wHu1pwQPOrxIE1zePx1PiQaEMm4kY/dVp4f66FfRWN36w
Rql8MGhajvMrN8JJW5AtojfMfB7cKwf4YA7CyfxMo8R003HTRS0/d0WXuQFExvKOinHDFyinHUHo
0O5Ou7Cgy/vlnI61NrQaxps+T0oshIbgZzPTNOy6UvYsHYwWvkYh74hGi6pd/TNYBda5MyrHk9Q2
DDvsFHqQgdviuSQzjhLZ+IqjtaHHnyZIT7qzt5Evj709ZWvEZ4lhrZARqFHCAQYkSHoVarmV9k3g
2mj9DKPBxnkJLOYgl+fF/xk1trZfGuPvlBDiBFFDka5s0hzsBLKXr82urVJ1wiew8y6gcpsT1H59
4E41wqpW0PZF1TDsDWOmP2fjH/x7Ead7CcmwZveh8UiDdainCix9kS6eiqE5YoqIU3PvZYSwILsM
dlch1iWDi09Nd/4hmjx293mYKYSv0BBSy9/TzGbDakUf0vE+HVz7U0giRMkxxIUQ01szD2ORCqEC
exEQHfZ7DbMgayPc4ScWLqB7WoyLOVG+UCLzXFf5mlQK1TenFUDwnDseF0Xdiqbf9Su9TQdaMw0d
mfDM/HVOYg9+FQSKCO9oMYw6UKBoDJFQXSd4nV8y9pcrbYGaCxRShgkbaOat21ylws8SKa9wdihV
JNdEt3jaKQWXr0AwNohqt7CdcLYjW5OnXYsUbh7ts+wO5AZL0LHFvqGHp6ocpVUcYq5R0mPvoE2o
FvXxKAyEbp3UKe7eQ1a7z+VchYIgwwG5sAF2NMWTcPxBwTqot0Jl+4SAb9bdVCpDHz2yKhm+BDKW
8iOYnAOEnGmfNqEEnLeeNRJedr/VoAMirEam2EjdfYk0+Or9JqL3yn3SRmSTW047cbYQOnP69Lg5
gWgiBpS1RUM8b0oC2lHQ/88ZIbbfGLrkkQRTgCRjZ3AdVvcaFYsDLbk2Bd7nMQTntOIjC+3GTLuQ
ngnT7iyB3o2LqL6w8uUEe6NWxuqasBZ4WJULcZKgfKWnMIAXukjKtIdNH24PsIOYpz2uo3/9ZaBU
qNI8P1aOS+bVn0vw7v8bYAeYMirA7IvBvNNEUbGJghxfwT/PWQAh2btNTaLO86XRxF3mMlYfAMMW
JDs1m6puqXynQP47fX97vfcTFUef/FHTdleLWXdn+5ZZIjf69UPGCafhgU1tICOeaDsTUWwbZ75E
xK+TLNyb3Z4/I/JIydYjX/6prXm+9fH2rNk8mr/2TSMVEOhsS4+/sBK1DPibLm5mdS9TqE8QnkHv
nS5mhugisw5qZYghERDmr6VYR8fHjpts8NQQbkbylnEoaxE0QwSTed4EB8sfU/8Ab8Dy0CVqSUkG
NBxTPTyw+ObCBZHmyBJ3R+fcyOQnSHWe54UVXitFG9y/EXihbCtZK4TGKKnc2ZtUNF5Cxx5EJZGI
8y8Mj+isOlfzMyyIDZ64zlGFzEpYRC4bre16YZZW0YE1zty4mbgrBiagyv99wXB9oZL19dz/T0BY
UlAX9POtANbsNS9p/SW5tW0XYRoko9MBGQyIECmo9dkROuCiayhpx0SONUH0rNsflfGDlt/8mIx5
oze6krV+NcABiM2l+QmPpEtNAruUufnmKpO1eRoZzUs/KFh9NRiAluSqpMbmgeC3s5Ur3rk9oZ5U
Z5uTXQlY0J6geeIil+ahyCEAnfw6mzuuMRWdFERJe6Aw/KDVnX93xX/hc01Z/g/vYCYZyOIkov9l
nzdii/W8qoQRp0Zftq+0UgsOxMhD/lCiYNHsXBgL5OB33BW1UPfIpG+AQ8uhjFKacHmvBs+v8pIE
t3l6gByUolwXkF+1hE+H6G8BW9z+1IbNWHHdkTrTRtijyV4auGWbXE4EYmTfUquK1e9gleZh+zX1
ZLF72cVGsPCR/vtqFUh/2FunrzRy8vNyM0IabO/OkZNifW6IgpbGZo+uhbaF8pOPIbvIyjbYi1jg
ys2YvbmdISKOCYu5fJJektFuU0M9JSxQo+qerzQg+MdQQeupq8s5L82qqdxcz5i53sMjisZos7ED
EJDV6fz1dRm7o0PmayyeIoX+4IyQnBcvD/bn7dlqbbu4rBMo5dWO8+woJR2nG3wx7np42BRP5Ctv
cVEbjHs/j4NKoshUZCLZYki8kpv8TCBckNIoTgut+DMu78tBBYBT5lWrhy1jVZrMTs36/d5lo8kd
OItiSFuS4IhuCsVVUNOAnjGBlYdUSerlb/rbOdBMYTxrwawJ2x2LvEfgcJgjEA8nPqSJNf2TEMJT
fqhY9nrckJENGW27vFUwXVhii9hZu+W80gL012ReE5xHLTU4Qv46X9NL8GIBhbW5+IDDLDf47A2q
d8B9eAZwCZatAChOGsgOOr28dY3j6SLhxCZuuZL+CxsVTQ+KJgilJiVvqGplqpwj22GhX6eJSOE/
UORkYWGPM1DUR0I9i9gzhHWO0KXwLn798jF9K00mrxOJk5CYIgTjtXwyO+I8nkN99PO7rV7al1CM
/kSn8/yYN65MO+SBNhPwd9cq3bny1/ampUTYAa94Rxbc+QavcO/gc6ccnt70H1AcrmAGkk5G5j7f
xgLGbYhDoD3+a8AkQWtmHQ8yL4BNn1b7TPgFBFuRRL6nWAOg9+S/Czq03YkECgWHaaLGfcTS2QBf
tvbsIHqkAf0MM1y7D0ZrfBudiUFvdHBOEMWw8bk5WiFyOnevXKp2c1CfUZD6RjCeLPc1Z1zVSX/I
Q8pxwvXSWmzfOVpTJGGL7AVyxB9+kPefTYwBonNrw8+3ZkStFtDCiAFGt46JUlgQp5kXJwSTFIRu
iIP+qHsKTTtWFai4LpGafglVYlL+zzuHW6es873Clq4ih5rqDo6yC1vWH/Y3MycjS+uvFTTT170m
3WjN7pf4AsOpFOo3pvepGumHIi1MK7Nt5t1g4AZ8KRyTXy+R1TQliHEUmDJlIdNOylWj1Ravuvbh
VaUNvk0QAQQpa6SMEaulAcfxhsbAwK3RBm8VIruNJOA6fc9zPN/Jn2ncjilL5ROwRZvDY2hmJHaH
ec3yL3LDhzjdD39ocUNV97ayd9wIjgQ5IDK3hiv3fMs0nBgzw+tGxR14xJaD3WoXtFuN7rXDLWQ/
oWaAZuyM2+UpJNYtPwdkQ0DwccfVXXGQBk7HxCxC7qhoKGfdEuLFtgiehvo0DVL7WgMyX9qmeX7w
N8/yb8o5HCk9NzoQenC5MUksKUlRgCFqA8tgNfrX6E5IozK5/3RQ4XzVabSbmF+KJ7+gmsZYY+81
OYtOtL0/OSFnMpwgIPBygJkJ6QBRXzCIJYYRrYJf2o3UtQcqcd3ik8uq9v1X95BEbLvy7EPGRyTz
is4Kmk7iWM7/lZz36lOx+0TN/Q0CgpbXgKRUgBsFgk7UHgyreUjqdnF0ddC8A2VEuB809X4WL4kM
hitPlLVLG16DKMA/Wf+enxxdXyC0Z2wbDQgQaKtwrpu/N8omBLnY5WlM8cSWu/5rxas+QqQEnmvw
Jp/eVVbexgQhftQyFAF4rLhRD7Pm+RqVuc5ly9tEcU+226/qF1XEOBjTA4kB+fqw+FTV8ftOujIc
G7pt/g5nKtNOvlsXO28qaQmJUA88dNE4uOkTT4bYT166qKXls/yIItUKDU0MjkKa5B73Gq2M4+p7
kGA6e5M2YI49eO+8FW+gaES8h9RK56rGmU0B4/7JttfuJJn9cDJ7YxIFZoew38aCyjF2+ULrJGDE
/0hulk93xZg5VAb+m7MtS6XGIzoIMWYVXb8SIIsyGDwaA+iklr6n7joiCSw3h2yPdxJNC4vmHJa4
wiGygdBemmOHZrFRt9gR1KXv4H/CMR8t97scMtsW4DyFpj2vpTR0nj689UF+16sW4SPOeUcN1iXI
8KHmeo/qLvv687Z2IXMfkeOWy3PUo8SMF1lnSZOfIIRLvEQpHXfz4wGqiVkge0pc1jNHVpgGk4ax
X+JR3mx5bpgTrV03BxP07Oo9Dpl9ALUYzRmXvhzjVnqNk0/ibvErNzz6Bw4N++o7NBFznSUxZb98
LKJ7rwieJ7qy3gCR5aWDkpWmRgXkQdoyELG2MEAkBBmzLApzZOqFb0uw4tSGwq+rtYR002ruMIEZ
TrstjA1gcANPn0o2EbJXiOz+upOicysUiyke9uZh4VhBNPh4jJ12EOQuMSbcm1gGJljcO8QaN8jx
cYylqh7N3IEMT6CLcSIyHm6jDBIk95ITQV8USVIDbw/HT2zw0oW0tuptuw0FhlziIbqXCV0l39sI
ejP4rwxoADjUc7dikIN6S0fU7H7ZyVGXTLQorGEj+jhFS64MrviPKc0duPyN2cynCQd3kY5TadHM
PuxVDPd2it4PKvA6AWYyElp4YsqlpG+zsD3aht2XK08Td8MKZNsQ551cXgPuoCFMB3qZvtEyonm6
ok/QHy8v6LMbR7rFstKq1Oze602oUZFuRwWauUL9lUUaVRtf71coh4vU4BZKr2gyQ/X4mhrVfBCR
vvL45fiGjkHDOYr1MA9G6QDKge/0r3A9wmjuMBB2J9eUaSsZXpw5FNCfkEmAlLdQN4wBgHPTUVO1
uBvtOzet+/jlue9cnAMMH/y0AEZpVr1HdGYlNWM3yt65SDvwnnjuOwaDE4OEfRuN8M82J8WqOyyT
kNH/FoHk9+ISOXq8euxRL7rlArj1z45zKczM28zHHzlwDJgj1RQrPeVnFMC07vv8JOlqQm2l/cir
ZmKoWRQYF6eS+TN5HWZSEty/beVIBrdGe3rcK1hdZE40mC/29Bqdsrk4GLSehyFxgIRpW8LHpDiy
2OgIWJ5HR5iGo8m0qeS9VMPa3/riFlvB4FeZAD7mk8HmaHieL6pefxCY+lgOXmKCMxE/XeXj1DgY
gTJ78N+jb3LFMgSGaBe8pf4wg7UMvvikz7h22bq6Lk49vilZOuZpUlQS2Kiw2tORUFRMh5btZ1Jc
yzmWbvjNuOKeN8gV89WH1coA9L/RD+h+woy0qtJK1Nr5pr7/b50cD77tF2HTpYttbMs70Lru2Dwh
0aUu+O0ImUhaUNdQD+kArQ4lvipnWD+sL/bzuoyJ+om2gLARTAK+LUS73YVg69NZ0/+G5tD+jsRx
jF6XKL9m/dDAIgPrEnsn4I3R3y7jNxfNI7doylw/ssWDisZA1jLE0N3/c+Yq9xNUXLtzqJCFN0b3
MMhFA38RC1ICdHfv/7tuevr91cRKVUoj397aQRE3M8WyRDlWkzjrMVYnyxBrCk3q1zE+W8WDU0YO
A7/LSjONyeNGfoHFGwQTifiUEDphY7xRpFlUV82CAhI7RbAWLDXrsHTCXWa4BjIuWJx+l+u4L3YF
jHWqJiU6UFmLSXChN/h02UWV6VHL92sgV6hVIIyBlQ+gkxetbSSNFIwPW1kqvFy+jfpR4DNghuhX
sdtCsq6l4IwWL1SQ26Y+JPlBl2L/UTS1ueddNQ+UxvXmfVD6Gzpzegbbz44GIG90B9/cxvsZz3A6
dUxkCdEsE8FMFLsdZU+FzynUDPt11Tbbhxt2aGzwYOpawRUFN+mKBxAetQoN35vexL2qG4CHsGfx
U34YvpPVjLXyJ1DrVQPjcvZezjrHa0nEssVBDiDXAhAO0hdW09vP760swM11o7wccq1Mey4JNFzl
lDcOz5OHhHz3149lkGUtdBSdKSCRHi3Mnhe7B4ilMhYXoJTqCs+b+Qq+qgfvQffx2l07yrBkY+Mq
9JmNNVW8L3vc4a26J6F/6Ro5yXbP1L8jCzdnSevS/fpyeXQMEVmlN33j10rZq8HFXUn0MGNO3Z/E
Gs+TjVFJ1J+vpMxS/zKj++MLEf61HWGofTQ7V6XVDhsvYIA0bWcq9i4kJJ14S+a0PdvBRBariJ5/
vqukS0QtxOLf+0GpQb9KJ6iSX/BBqCjuWi3GJguD17AsKByFOjQnZOv0EmHCCCK8TvrxWmZnah3i
XENbCjwGKaalW8LKX/609A6HQHDQa56+Qhwm7xcHMfEr4ILDj4TDD38h+fK8+goweF1sx/k71BWE
q6XMF+ze+WANJaSjcS9YhkCRUgXB8SRhhpAVJnbYMU177FwmHLMMWSJ2TFJx/ry4GBdq7Y/qSwfy
MM/uo+sWOMYKdTps0POqabmJTp/r+ZagdfvJUYtBX1NoLKOCp46XAVe5FpyRr/TDocfQUtTYNPZf
+bbc4S6OtSI7R3tiLK43bPattiZLc95J2tgxweUdFA4rUUpNOCWaQJzMwl8z+zsV0sBgSkzda1ue
bDtEsIV6Cg2QGYiwrM66+1nWu/I3TY9a57Ma0/+tgaGCAiWhoeAkz4b/U6QYkNRGqBgrXsamOTCR
tQMeNu4z4Tn6dxc0kZLuH4NYbZSvu9NBSSZYAiuW0ukzhG+1SARtQCpT8ybiAg7j55e9KJXLl1Vz
MxAtmKvXu5/Eu6DWPgtRpJvH8RHpb4rvqiysUn+hR0HGjK1Fa7x7KQECwI0hPpflayXdOh4xOLKE
/hm5GZULelSuYzI1PkHPhq0CDz0NIJRjGaxKZV0bC1Ei2z3+YuWUdbeRo2qixcQeHhlIBcEPD0zU
KMpfHrvTGe1GJMsibbKAsXXvEWrkouRQbj2/1DfATrZzT2tYSvIR3d1ck4XW26xPQfYv3dwxYzED
/IZk1seINumHOAY1N0TVtA4P62B3FnHvcDgBN5bx3ti8NuPfs1aOM8FyCZGUybSZGEs0LY7VWjSR
YJnTm2rYW6DnzaSQs0JRiCasJgB7Fxyu143A2Y2IeXxz633o8GRIrckJIOhu3zLU1z/Kot8yar4E
s40KDgjEvlGRvXwARV9kgMcqz/8deeaTpC8FuhKAGqZy2czUz6NFKtWpF9jfgBJvNx7Xhkg4KvmE
Frrx6+8mbrsJzIzIsi8V/Ybh15MVNCB/59Prv/Rx+xoG8iwD7xcEOmRuhQQzCOQyyQ+51+39uRGa
aUu/+fpgd5EnmPLOT6DwxCDFkWmoKAQ3w3Q2mH/CEWz3YvoKCSWlsaCSab53FD5oe8mU02gy4RT/
avoAqKmQqv+EiDc2D5fwZhkB7BJyLD5MVi9opj6EG3jh1C58+3vjiMUHPMEMKZALKsEc8SjITM5z
yb3fIM0DkvfjLUS/rYiUHveri2NGbDAgCA4MYvSuHZpiomQdyCIPAQwRb8VkANUJ3v3ZTFa8pPHp
X/gqvihPS9BfkTsGL5auJLhpoG01SSIOG+/a04vIPNnC0btDl32oOL13ZaQX1Nn5SmPaDOmpeZSB
mHLEMZpn4crZlxBGjtqr24VPYf76nwFS58j07PBCjGwb8phczPgZfVEFwlH2QD8hzF1i45D9uQNx
pKiIxatbp6yN21a+yuo/WPcwGgMl9Y7RVJFRhIBhsEAdEovbqiXQsyy8kRcGrnJ/TzXqoNdpyJF8
PNzkLbjL52BtQ11pWuLDHdiIIz+Cw0ADQA7FBh8BFbI9DzL6JGfMoTXnA87AqhuYLVQbfh+bYfIQ
CtKOglRWlVlnVp011WBCuJFJPT8z3yOkC3hLSBTKT8517uLlOHtcCCbOgKChxr9Jg3OXO2SIRrHY
FYP4nNs/hkYUO+jrWuHMfc764+tzDu3MgfM8bWtdqTFCtVqDkVq5Uuyy7E7ZTkGFKa7phoYc1/nG
GDheb2vAH/1Cl1nJvIkNsDclZYH25dUVpS3Dp4QsSAl/lQMAng8bcuKTHZzU7lY7H+0ETDSA7GNO
CNWvhJfD2OUAIAoAuSq+d9T8Y1UK0bROaM6onROFEncj2BltxDgWPg5toqoGTOGNUkthfKTeg4Qr
WglqcOjCzvskjpmVtJ9XYB+oTPpeEyehj4R5Bf1h2aE5CBIWxbtRoV4ljinVGA7oPw4aN0tM0B/8
+JKYU/6Vr8K1y4k2+sCJQecFNFoW7oEscO7i5v0JJrt9SAtpdG1RR3TuR77WeFHujYeGMnEXgWkt
FIdwLxV5p3iruhHnhFAn26Hgl38YOaDJuqqOcK7qroWGTLX2V7coSkmvd02k5c0YuNU46JxCc1P0
tvirchvgZDU5GCG0mBz7xaCAQTteOXEJyOdMszCI8u4iexCiWKeJ4OZQqbl8vSMrNfJkGqwF0f8g
QeDMHHGLQVGyzUqB3NOIVwKYXrrsd2xI1BlV2EnuitIKyHdKPH9d8wH++aRN2lIITeqp5cttVdza
NaxR71E/8hEtYTdAN12fDK7g6R5NP/iOx1TqYpmkcK2pAC9R1A2pB/mBuLUfzf3aaRhUdyrxksfG
J4rn7p7ZwwUhBNefqupihMXPTekeaobvzWyr6sdIcfrlm1hFwYRD3cktr1EEI8BmQlYpsCrvoZFU
+mtfQ23xjU0fBzLYHagfhF2Ob5BY9SgtJgA9PYvHNYZ+tkH2FG5kcF0Gats/5IYho5FtlzJ9Aelx
j+Sth5RV31MYCjSdH5knQQbyjK/ot7S27nW0VCKYjcl2bAbfx5BXGKzWKDptzTGv1tLkhyJQBqn3
/cmORVrsqdwdq28m5nMYUqNI7AkgOI+cAOE02c1qnoxHJYW21V6AhX07cscHVzhkpJmr/BwR8ck9
jzC6N9gP2nPxlnsveGTKFiW5SkeFaN6hOipVJOFcrb0UdBFkQpaBlXAGSifaqdsiNge22Mcodg9m
UUfpgeEfuiGyfFd9aCFxb0khIdQQljrrWp7gh9b/jZxqtgaEzx6W2o98W18r3k3lZ+3WFwqu+Ovc
07Mx3rRDjqAfwjCmFGW2WVGbEhy8mUaas3nPGKzlBS4AJ3UizFtn6kEZzkTYL2l3QJXhJz5AeRhH
OVeRedNnEzlgymagykzcmSukSnEQW0pgJPA7oEVPeXRtBznkMi/lSgGusB00c2fTyV+t2/ROtNJn
btuzTpM0RLVPlpKMbT9CplD6RZ4ROeyorbPwEfaTHnoCI31EV6zdKGRQgX1I/5UQjEDjB6lfoS1L
kEcT66YC5GnqVAiDkaC7sLp5dM7DUzuduohX2j31maGCsYH1dTRNz0UiEiDgRGLmfPDVnUFZeiCn
bZd3hDx84Wjfmlpq675Co/orFzE3ZQkHHBzwR5kU3aXTEor4Ivj823SyVNXZPeDexyNeUz466gB1
YReD+MNWsRiGoFUCulbyDSUsFDphn3lmByU+TpZP7cE5Doh7QxSYsavdMK0BwFVoOi26j/ESuOEw
uvNDmTHzVr4VFGqG/XygZbpD+x9mMjZC6X4AjJathafCYX8CrN08MEEQ5LjgqAtiox/uKAmy5ALk
MoDemu4KNmWFXS2fvAtkrCcpG9/FLOCdAQOiYtJsH9o9upa1dfCOWEgTyfbk9DAAJ5Hk7JFQZqZp
zENOOa0wUpo3MIypbmaCXQM1FpCnQxEvba/wdDU9SkIVbd1unFmDfFYorctOJw1h4Q1Jx/L9upeA
QJ9cE+oY76mMd2nifYIeno/zS84GKbZ9qmDkIw+tHrY22SKw6zsTHWwSykchdF0GoJrBKJ8hWM3+
fu9NQZ4msK47gEjoTgG6qfi4uwW7cYmAH6EoIFGMzQc5DyVM1DpIPLU+3YdE4cc40VcCWUYEhAPH
umSZXfy6B8WbO7sW5f3kXhiTuE/IygK4K/mnEkE0cx9vl16qRRioE1MAnEY8mU7jrxkdVoXrgaQ1
Oz7HrLYw6M54R6tgLUp+CFc6cO89hyDNypK41oP0QUH4xy05PhsCB578aoCuzGdVC87WBt5ZL9uh
GohoipzDhYLAb69cD2aFBNevoFMQQwy571Ia5bBZuc5+7dWIXvjqGeQfStg+736igVCyfMWB2AqW
RpaagM06aQCYfW4xbYvuRHppGAiHRYEVUiNKEeIiR8LVEEeAdsFp7f3tCSW7cwjTLmfQNQ1CEh1o
I/ego3R8djE+iXGoa4UVgWEifVx07+ZmWO3K8wSMtAvTBQyrrA2nR2cFqh89YHxQcY0hMczW0ePz
ryTU28YD845jLvku/PI+WDkPZ1d1mfba6bNWyQMVoqo2Jc9tuFsCJaRafrm9HcaEhLouxViBRKyb
FVcSXoukdjVqIY1oLPqtPnzT++MF8sHiyW+/qxKDmIie9zk8h9T6EqOthedd+sK4qqqAvnI0MwR2
jpsY96DtqmRUjkg6qsDL20VKPxwbcs1FUJRFa+8V85apVfUzhdIuGWA4qdR8yl2oo5UQWrHkfmYU
T4KMHjEQAbFtzo5UI7IixUfKSoeQ/w7KSGkVfgLeus/qR6zfSzI039Im8hEsIzSzxltcK81bzrg3
yYBbjJHye5/MZD0PewqBNTPDKL2z1zC1Q/hZUTZCHyYaMiKohQ2T0QdPZZA1QkZPgNhJBtBqgOPY
Ry2mDte8JBMSinxAmhcTja5xh9cPtmYoSMPNhLwqxq3CYCSZTZFZ2rFmRWmhv8dyikRy67mVzLAo
QkJiF6X7iUsZcQH/+eRQJS7rtdC0jfHdVdQ0Y5ZEUckeH/K15MeAh5GiwMmM2m8vQo9CGZWL1T4c
fp4rHfvKTr0zCAeIM7bseth2V34gP7deIfZvaYLxu2YWXBGtk6t8elRcDoikVB+i21vpYLfC4+VV
ALxrrIh/jPbHdLqRcV1vOHYZ56JeNDWuy6L+rz2gbQojtmHN0ebEQzj0btU10FbOU4KCJwGyZyvo
Uptc4Pu7pZZjVCWEKSvUTlL8UmqZZngw/kfBG3qSGV1TpZO4DBsAmx11PcXkCTFCNKGtdy6UJE/a
gpvmZ/KOFnKzbdgZoWqM+a+Nk0nOWMbJgNOxYW0lkx+VjVa8EkGixafon14Y5nuZaApUlNPLTQO/
YjdSK/KT3z0biSdGV3LLbuLtuAo+Q3Ab9yVrmvjLVDgshmAQl324vZbwoKUQFAeU7mCx5Ee8seHa
vESEmqrh5CPjTGu/5KcdXwKzVvLm0hij0/tVIVc0q0V1oWra2RsrH7f72uyZMahm5sDJO94eMoaR
hxywSa4IDt6FMclAq6p20CNGVZ6HrajrfuwYlR0OTTPLKIM38QTlvCTKLv5UY2EytUicj1kI2t8X
rn3tRl+OsuR6KUGM+f31GNFmcvLRjk4hNazVzXhqGFkYTrtYDS+X+EQa/fivHzX6Ppw02i+SJjpj
T5cIJoKReIxj6hcDkICk3FKza7ZsMX0C1TY3AnvExfkYh/RPtytxtDhZC6ZFE+FrCsbvp7upzU7z
46i4j7rOb9SE50D21CzIOC0cU7PYsL1z6BV+EC5elmGIe4B07W3TJwlfksnuaAglIBE/rHcLfGue
PZXWEDPeVM+3ECnmbNgyZRfIialY4/U3qxBgePUP/yizZNvkZ+jdjiCnMS/I3IPuewn//6jZaXEC
CIAp0BKwJNPWbi7wrV2fw10LQuRWFaXLwACnj/7ybJ6NmoE88mMLgBKe4S/aAOHjGzigflPgneH/
7S8ImV2CcQ4aAJyf9N7T8BOwdVvFYSfb54+jlfuEMXHt9w5SQcFchv2YMJUM71mGQO4FrqPRIvhX
gy7y0UrVb/zs1BeB8uX3OCETdaYjvGvoBEQjvGW3FwB3BmLQ/l5dr43BuCqcHiMf0Z+Z15UZfN8C
oYVHmdaa7j1j2klkcESUTM3hnxyi8o0Lf9xYlhOq5xu6+z+o92lI6+x4XGv/j+PlYE4awMpQv16F
K+Q/kCQPFSZvf0I0FWcGyQne4tOO6TaYT3KTehKgIFnvLThMaZksj3EY/bKbhPdQXdm7b+SGSLq4
D1zVrHO6WblKs53phtcrTMFgUELN6CvRtKOrzGCCO0BNhaZ83dSkDZgQp/iv8gty/gVQQpyuzIsQ
2f4Tl5BNWFGYJbqzIJC9CWfq4gi4df74ObFlQVxC+hBCE8CWwKLVS3G5FbKJlV/DjDqQMv2wcy6c
A8uHnb/P3dgQcJwAdcN67uuJp2ahF+3EdrgEAlP5RPFOHVp/tZKwPDY4H0mUawTWuFh9aDBaAfiH
UhOEU5KS21VsHsDBxBKe05EQ9JuvBpfGg6unZ7cU7hYKN/+VYGtkO8ZhUNH9evtN7iatBWLMvVYZ
ZGYEL34T8gpBNJeX3uwvPhgx/DHDTaUc6BMC7CjBp6W2j9RUfwueLTtT06f1J9zJ1C+XmQuZNCsD
mHm79MsrstRrMJ3tvsuRlrDBmvQtxC0dxojRp7zWIWOicF1eYC2Pje3q6+oDQiBcXdd4RBWnMQ6c
v0c8TUCJzabGTvXonBag6Fkc7smtsfWTH4ajAaFuFEa9cG5vNrPiZBMrvs58Eq3xlXyn86n+TwT1
l0R/jAXNaUpmtKBIF4ui0nRwIUJSsI78hMLH7D8fRzZSXQ5kQFxVjEwSj5WbCOMmMPFYdOfh+xOz
/ok2hsyffjpVy+DhV2cpy4vslA98RFYHayTtRbpyRi5AchNB/FC84sXmknzdq1irKpOKyiSg6gq9
MMB4O6PvvULwgzZ8z62VqMYCHLa1OpKDuBpW1kzkc9xsOiSftA6gaGCPO5G5Hd6SwIcUcbEf/3sZ
558NQIledcO9Jn00AFpFYZ0PCBVSHA6q+RcUyIJNgb9O50PixqlqngwLkHa7D9r7a8nURG0iP0VI
SmAHYP4tFWZFoFx0v7Li9jqQsmcKTEU8XsF7tDMlng6BPbk43SlCNikr0tnqsgBLiq6UKzQ8jXUI
9lmxaVPAp3DxW2iZK9xL8Id0iGA8SB59MIbT2XRHA6dY74zk2CwjHXgvVMOhs496g6xWDAPgAi1D
7zUE0Mapx25R+URl44z4xCDg0vHSxIlAyNmJxzhL0kbzuP//93i7VTOIhgrbHU2OtdFsh4b1Wa+n
q9k5Juk2WBQchirf4AO7CKRkD3tuzKmTrtA+41dQC44CWcxPoEka25fZ5I8kbHQOXq8aO890VAyV
BsJq9q3Lqpo+/xlQTOw21ONVK7To3UiGX19/aOn1u/pC+WtJFJ6sgPWRRdUZoNJXayPatBOPo09Q
mrOhNGHr6SEw8xREwCecBCtcSGc/Ze+w2Wz7eaYFLCDoWrRQujI6mDci0WTZWZoSjD7+CIm7S4vz
MIlXOy0LwJZqS6uPBLysHmKklCao7O07btAAlfdnDsMB6fPm4mOB4rXOL0FcvNcbwHcvKJomof2W
SjPPVzhRuJjQOIPW9dhLJRZIdyBgocw5lqqBXVqrXlzPVtvSoRgA6jTs1qGkZSAM4y5bpEwuUJ4Q
150MdIHuAoLPeY/B5sZvQAVvMY2NgJxfBtaC5OAs5HadtUE0ibQave9qMChzkq9kXUxfQLdSgS2g
I0dis7HpxHKZgFXBBBNnHnB4tRsO2c3mUov+4ZITv87+g2rVHp1haK6sBQkkdJaaEjrVK//Fn9Bg
jLKnI2DotJc2w8Pi4QTctNIq+JZyrBWFZrokJmL6wgrvV18/9VvR0VS/zJFgPO5+fyz9uVjLrWcC
REp/3qvow/8KeYaxhb6RIKwRD3/yUGiGZXL7d07mXNubKJ+WqwsXOMP1Iiu64ZVaTRhgke8eMH/2
zw178RXYi/5UrQsCT7Ihd6ZG6ySEvFrKKUgRdqabuExP+Sq88qP00fFuoeSx0ALA2KzjGsZoDI0f
11PwU1NC+dW4DzgIqTzCfqEs2vSvBJsZghuQ2LJaiy6Z5fzAq+madh7mbXW2JTFFzNbEhd5lSlV0
+jnyFA8D1y800Q5BGehDNqLjDaXKAs/lgaSrS7d7EhF0XgDGsNjunjbiuf9y3U48t7O1ZFlK6ciM
5n/6GjAuIzUlDfj2tqzM7KbY4Qy7Ul548U4YPozb/Eq+L9ut5DflMeArOZJJSmCg9BRvqWOY7HlN
SRBgUpN6pn1GHaaps48Xr0b5aZMdbeQZWWpuf1MmQfZsmt5S15lU+4GfuJN1akQUSjSi1e0vfFI/
+dnX8pQIvPQYDip+zbum+91yb5l8PAZA64Q85o16MEFqrGyrikKQW1mOjw+Uscj1l9ve7L7yzIn0
TtW38COM3YG+17+x8tgPZOe1ztooNYcGulmR8XmR/b8Iclb4//qEUTs8+7zsMmm/iCA15qsD4rty
eKfX8qls4Ln0EA/8In7A24pWCSfmZ6G1mrwEBU3rl7JkqKc5r2Ym+lf4MX4vbGpg9rW986YieZAy
gnuwn9VPcrvWVt4J8E8cmGbtGTlbg9r9QgcSk5/h+Inz3CRyII6a2cqkPU8D36U5lnPXnbdDnTl+
yontzIHNYEgn2gA5lrUbiRbkXN27XVV9XGzpYVn/SMp3MrooNVi06+YBDXQs7RxLVoy1r2zL+UbX
saQOQnOOANofnek2xtbOi1t2OgJzxiSAHTk4IXNBa3xMn4EY6GsGu4zrc2gQe547zTvIAPlybnyO
/12m9t0YUKwccMM2d7/N5Swn0n6xwC0LEExhcTcvEEwwsqf5ePocUYBxXLH5gD30NAtk9vuEREiL
4wCKRihO7HHgz4bC+iM0VgXmRTvd2FZGQuA2VeLqaOTuFrGdozT6jT1hmKDiW3lCi6awICxCKU9K
ZUy6hBt/F9h7oK3PPodAF4l1Azyg1owoHVZryzh3Zvpy3MAPD5rKg2k7xmMV0+m6WbQa0mJRXb+Q
GUUzGRSgnzhFVSBSsWNXDKbR4/6J0DODL7BOXKvl1iDHY0w5OP+3HdT2p1Ghu+wqsG+lcG7L6Ck3
aK3XapSMk6UOxuCHqmYc6FWw26RSbR15gxaDgrUpk+xDKg+pZ3HMRg2QZLR6CCHp+dcw5QLPWDXo
3TMHzx82KUhBkJC0L4HZ3GZcAHcILLLMzToloRGonz89VQn8I3AIs08M7NDg3cWWToU6vosVaU6N
wWnaZSiFWUPs/Di/6e7wbjVH6R5oiznGxoiROKhJZGPz1AodlJ9M2XnCdvjNPdxO6FCXtYfy0fsF
PcWDEPNmXVRaWDrrZRlJMCiHvQa3a8FE/Uj0mw0j0mvh0c6x4jqb33Sfj+TMaBgRcj44onEYCSNt
PJd4zgvMhFWPQhL1w/S7/3aSXxZnFxY6MeKNh6oarGclrpSiBbEr1loOJWhmY/YZ7d16MmO09a0y
NQUDgNZLDIBrL1mfgHI2Fc+CAvkxXXIfhW2KzBf7G8O4I5HfffETL/XwmJCQGskvXfx7n08jNfYh
dv5bkFUYL9ikr4BDRtORs5u3279nkgNvJkX7zaZwVo/yZBLsqfF5wXwy6d1FAAQjsrF7MWtX9s1Y
POV2Cc+yTWAro1wjcoaVMoGmjbRbtO7tm8NdfSrVmUEb8yOJW+UWjriQPYYEmlhjnVe/X9yReWY1
AYaMybpaUy1+BdhkM6BZicH1I6Zz6erCGOXb0FCmGTfzMeNH2F3ZXkys2KU1BwvVLR3wSo5fzBY1
sZBbtmGzXvigdsbc7Lqm2tjY7Acs9KW6d4unIHs6F1+phBKsRZrU/P9tTBlQ8L8owZb/azwN2/dE
JRFulfUkNVbQ/Ro0f6ZPMOsRIueN4c+CLPO7uyIRRhTbQVIeGLPyhFxDBt+vHJ4grz34OnztFWeN
5XNLND5CBmSAwjRtRjuL4z58o+qcMOPDRzUOM9eJA2CNABLa4kRVUjpJf7DI0ffw+Er7fxjxuA8N
LJZzs5Rgqv8yqvCgZpfatA9QaaRV50fwhXdMLRY9VRebrb7n0s46ZLq3SjBbWCBBEQFJBRI/Ubt2
l3nPIrOJoq0/RG4v4WqKJ5TgKHABNAB34cxSSQO/UDta5JqaFEr5xNy04g6oYsG1s7IDo7zBC43m
Ki4wlj/WK5tUiGwrBdyeIvIz7ulaAgGsFc2FnSqL3U1oPyFNrfEKd1RQIsP98dFZ7Ops6RFeqseG
9w5W+/HLYeoqIcRJWZePq7VJrCwjrfHgPJZPelcvgtPtkE2AbvsU8QzsfsTUlgVX2M0JToRl2Nt9
jz7jEj3YvFFtQa5CHC5BJp+lbioJgqG4L5HP1TeygLv1QiiGRzTWgkNtLe81HOigVfCC2IR/RTlz
rdgq6VnwGt0N4YBE8vIPgi63ThncILd7kjzUTvk1TT2H7275CwDp/0mqyjcn2NzbuHLUts29NpTH
kGO3Fra8kqeFEic1ToxZxaU7vauV2tKLOtEd5W2HXRtT3ScywRZMwgYKu1MG1tys3jtAX0tjRMA2
KHgo3GONIDyFcRqHdShQYsV5DgT9iWVW1ISgwsS5A/Gm8b8VL3QN3sun/94J18C2Yx2yEQzC8cFl
m5TAJq5Bov4PBM77wWDWdJTFhZahOub2t5iKh0VkLjm5mN1BIW6em3nzO7GMELt1hK/zsuMD5hNJ
AryZEROtlYlPEwlxmmxVkGDcXEy7WzVDvtgB2/EJmv9KsoPX1vP77+zKDs/+48mN/OUPSGWRaOP6
ufwGK1CUWkoGjAMO+qofe8JFzASp4Nt1PQXgeXmAF4U5iu/DUF1oSAYDS5fkb7Aub2/Xrd4TXCsq
DOtS53rtOOKn0X+pcQc/29F1oEqaAW/HZXmgjAiqU8C30c7DiIze59EzYlrg8tCDuCrckHlnVw/N
1/5fJCPnb7hqzF2mPcZDpVykJJ86upDKIe81j/LoMBaTtzGwucCiI7L5LqNGVI3Q0Cu37mm2Twte
vNDYiWh08x49aJCG8ylWSRpDyr/1RgJzIypHom2V0u0xNctlrZ/L2Ob7kZq2nFy60dKgodTOhpcm
C7b5VYxvCMIgMOwp1ElSCLzJQjnZFQb8gXUjTb+HcacxyMOKlJGu/CDlOIUfZzc106WI10If4MO8
jB5gelvoRJS0xN8ElzHxkiOshNmuUetUXS4b7LFrzQq1bUIwNEY6puO8c0ntiPrPzQMbWu9I5Hna
PCUFCUmtNEKUwJGrEOuHDy8ufTqpovD9oK04OIb5IpZPvSupQ35MqxaaRvlX6JLdbmzrbDjNqO8N
9TpuDOPdwcVsa44+WL80BNWUdVtMajmS27Id87opJfK4EXrdJ7sYtcK5vOSy/7Z0bOXQ5jUoO5VL
BWjgY3+J4HSRplIgOPhlrBtF5bmrJPS7eD8ddxBw2FSJZzOghTcBQfI4yAxKPrvNg3D3qBeioJ+Z
8k9DpWHEIfwsysA58hCujQP0DRxxh0cd1GguIF+PL3dd7NqBCFCUaYnAoOHKOl14nGaqDii4BiG5
4owBqjn4OicroNIOvZzG3rb/6R1W5hjLYDPYZV5gYASSM3pnQ87hZnjEkLX/TXqkz9UPIORHXxKL
aScax3vRO3gn+NsLXSsq+IB3D0Znq+k263iNDT7r5UYmnOVQqOm1tEBacR8Br8PqLKSoUPRi/g2p
ftN7wggKG5JbJS5TF86G0a0Z3WXytpz08JgT6Z0z3ke6T4fGPiabb1IsH2m0fOYKztPWv8SgqzmE
JuJaoTQWbMYYHE35ns/IQD10jrLuNgjg1xFGR2Ci4vY3NpycsfPZm5Vhi6yPJB+OvzYrC6sBL4F5
OdMz6f8HOJUp0ZbgPoXIF5re7ePVwU57G9AQ6Ri1J8j1KFNbl/Pk7pPyRHoZBvuw3StyeQCF50Yk
uDuVCHxqIP7cWijL2DHj33AP60UZuDZXMp0qIykqssZKBqaTzBMd7rPJpx95uneU6jZAiBUjlF7K
Bj/NuJeWcRR32dns56+eonp5BCy73i9YBr+tP7oqaj1+7HpdALX8gXE01YK8o6+oq8yYup3IWpjg
UcenDyvKqG5+0HvpHXV1elF4wRz6qfBFH0mAVkLLvwF+MwfObICl43Ldt1vZyHgSsl05LPfmYj5n
CGwpvDO7jbpHMQLwktE2v6u9doRTPIoiBd/U6YKY4U5oeElLyZePTBq3h9ceY/JDqi2y/txKEp/H
KPs8xxpb4imSz5jbvbh2sF/pDwwoMYt3VnaLbTSq05y3UMrfc7I0i/WpJgDJWN/3Qm5SRFxU7V8l
I+3WFcZl3Qn5qTvL1nbK4FKfssCdjFy25lufepBSo73Fbdf506vOxLi34rEL3eZT0KgmqKyPc5iV
yOPznkBJtEM/nwYEEnwu5tIL5bKivcTgDpozPN7qgQ8M3WWRZXopL18nIb8EHainGnY4Pk6itk9D
9OpA5deBHD+6sqqAehDtpXpn416vZnJorTemAcpqM+R5qz+4LqEQMLh6TLx6aM8qDrUd3MCP6q0Q
DPkWrggNhhslWmCJNeV2iaYvmktS0yXpsGBJ7mpmC93XLwPk++RKilmbV0d6+xgPQdNToVi18ETV
zE++Mk5dwkED4M3PSOQ+hs+v+zecm8Qt3x4QGxCdfwCsQtvygKuz/VX7Quj5F1/pmeUsRQSrlBeu
Dx/A7nNgUqyrbbnujPkLGHll+/ZOtuL1SIpW8CiTBJjhW8s6hpBdv+Uf2Cgng/JF129z2ueRSytS
cQ0bhvvLoGYFAcEfltFh+BuKx6yvutM/ZRwyYSRZR00vfkbmuFptPJ9knHWDaDn7w7/SfWuMNhR5
XsjrU0PhY4tgUmq3R92RjG69toxqhdCdLsP8rGm+jyBRUf6q1+7KnF9vI9SsZgbdyMjZR6dwScIb
Kb5NOgiDCyZ8najGEEnP7QjBbeBEDBgRAtJK/xizmk1JjP6fEs3R2Pgdozh83eBLiseM6BZGGggQ
4dWPEHV+4B6cVFqy6UNjZY6zPFDSMWxKTiNsMvh3G76LnMoKTep7CIXIy25tP+R7DlVj68T9M5iI
iHmGav1F9zcnT+jOV+D5iqL17yfTv1O4P+dmIvVmj09LEp2JO7dD7T4xctGdVkGGjnH7qGlqtWEV
OeyGNuQyFY+7CrfaLtuqPQD+yqUnB4JQyzAluphxTGaKUASdcp+s6cN0AMFfHUPvVY/PeE0UfQvj
TBfNb5nDGUDGDmnXdMcs2RLb7unkgbAWxr1nxtf3q+l1C4yoXlSTKxeslgEd9YdxX/EeYrSb1e/q
gAhXb5vF6CR7MYS7ybdvmUlYvQZZQuePswljfbc2DcTMCGRysoUUQiELvnUrfo2qw84hSi1FQHc/
HumcQyQQm7W+h2TGSuxDhSgzIJnSvIsZJXjYggmGUtSX7QDbOTzvj2aC+9ou4jBsEanyU+YK6PYI
C2ueISEjaxPyU+juhrRfeMT+Gr9TSpmgop7y9KD97s/6MNQ/74IGi59MhAEagoEPTYZY4iQtfyRB
5vE7e2GGgKrOOV5VXzX3Ui6+eP1Bf2zCpQExFMYBhX7PGItlTbTHMdz2jpyr4ENLAwd3us3+rcUh
YPqwujXVjNtPSFmlt+fRTYui1YNp4GJ7vTJUO5xbIk9/xzia5AUuid7pQExW9WGWfDZxhlUoC4zG
ve7tZkwPcdvOWb7J5howPYRnWob5SI4t7RiPrSEbs3ztw64ZPQ2ycJaJGBUGemVBmmp4+neQMIic
SFlZbxK2pn7VBbvJ/kt44Zp0Is/SlHkwGZ22E9XYOjXLzPj7dXIwfychxNaFUfcstysE2AgEpABo
CXoMZ0uGwaO0s4+SOVpJ7zEvzPemlSx7w9QeZJ5zRRrESIhMcAQcs3MbzTmH6XaIhSYt9LhiOupL
tosDy3jWjtMr1rKdX+GLsE42jSFW+7LSR3oHzew75PMPhun2N2YtA68lArIUsMsOzlVN7gp4X+d0
iwbZH77hjipPYQECb5dow8A/X25gwM0T1EXmEBSbEtSTCqurm1LTfZatTwuznMW3lHhlU9mkdJ9G
sQYN8+dykDodOUEMUmV86YektiB1QtPhCpk4xuDKqO7o7hjRssEnjt23/awdPrg+uVmVSCspWLmv
JKyLTxh8w2/cgy/Sm1LmzVoFB1ZJh7jZBSqH7gE03sB6CdpjB8NOIuqDNHfd9hSPKS0jhJGG+6Cm
yBUcShLh3P4GyHlsCkExWLajWkCWpmMHlMF8LlLb9ZNCCSf7lsAf6WJ8yiDFxBEfGUvLXjJ1iVJB
ZMku5f3kkyGMCXYfVSuEaWxPi/FhVDejOSasngtHkpDZkVEt6QZB5Gsw6awLkys+j21qz/H8v6+K
r8tPDkXsoJ5Zcydj+3PiUeHsqU+4L20ta4M+CeXefoVetbVeY3bJEl0wZ9GSxWfmTzAfPn5P/ECT
eEe3YnDv/d0oSUyTwF+5YjQFcAmIxlp8GgJdS4OrgcUXvM+TZQ27/6//3DM8JgQfJN2wY7rpQwL5
ty5qKIwj54iWgLxhHHFmgrQviGTeVaZ+6EtrkqsLu0NZ7fV66n8kXRns5D4FSEPe7RCJzzIJkH07
bamd2D8UG7ynXi6r03Dcf0EDHazMxf8EKcajlunP1shnLf5EC1h2Orh7B+c4HVkdum2o3tKOjhdt
/jaIa4Rzx9HARPZbKJ6bJrKFXnwHXDfnEtFAGrzeCSlpIzuPpknkiDTPb9S8e/eksWptR0p3h8XO
1HXtnR49Taf2D/Y0hKEV+ZwwulpQ+7CPfQUVHQn2UHWNOFYnU/thD34iEr8T74OGwlNl+vH0ns1L
DpEnjSW1YYStzKdmjL50YE419YV12H0bFQLG2w6jfcSa7Ly4mA90xMbji/ctzsx71o3hyDybB5Lj
8qRnuoX/+1jJYH+nmFNs+WUHYxJljXtPvS1cu9GER5qyD8oKTLQTlhmCeodhwJ8sX9frF9Te/hT8
oqojh9+BmjxiBYdnGHFNSh2bDmveQ1csYEdCP3fRqznKTJ3AchRr2xm3Zi/ifpSWA9zTqE7x6kQt
V/oO5Payxg74WHgqwg+YiDhLAgMT4x1ixDn3o+d4zMmZverBh2lhgGFcHPz6VIEp/e9/PPHNV3cU
t9tHV3uolh1Vma2hTztPnS45F1hLd2VC/uIdnFk1mvJSfc7eqKfLgXFIEqCc8U6XiENGPc0W4jrt
pWgnXKt+3wkGKkYZeccxfdzjKas/qakM2idw8eBxHZ7STxxazlbm/BLfKb9CHGEWdn3apZ9ekurZ
8UZFUlFVX9GTuSSb6mWZN+/xyaM3mQ+SRo8ljIJjcS+jvEmvQTpdcHPlxtqogYYMyQHtb6OvPnxQ
rFEZyyVtpu/owfMY3tHIGzGwiB+sDwMyyfsyu6EIBasKuLLUsOqR37vfTrt1oFTpGDm/kwYxsSb5
eQLDdocYj0T6sIjLiTzqP1kJrsSjweo3NbAQ3uVXwqxCHWQxEXAZmCNuXywnEhmC/H04v0eqBbBj
3c1kQFmOCWc213rjnYfYN1yRZMnJvtUV7b/ePDiZ4uTy7Rfjs91OvDSrT3leT6tr8zS8mWozU+up
nZbx3zldf2ZJzh+qKhjjt/7Rhkcop10J1HuUgN805D4xzmNVN91Mo6rbHCJkWpFTXex7p2G252AK
RsZk3C6wECXbhQi8cuRjLNet6Rg0j3YXYnKD6cSbxqN99aYfGDFElsjESUUVVFweaaJWEtKRhULi
fkWholKO9pmlI+PZ9K40zNjkKuoMOuHSSIau4mLEn+gyOCeV+uwsRlNIc3y5MvqZtHCBucndBHGc
SbysS4lcuQveUmnMK9ve0/dYZr4Kq14zi+eoLpMea6EhwzpvIbWd/A51kL2QigjnsJkOZXxJnRr/
Tk1UGqWkn+/DyM+JWld+cN9/TUEMRaZiX7khj2C6D8g24VbG8A8kuYZVyS9uRmF66Dcukra83ZWt
AcuePdp2oUDyQ37vFu2rSHx51DAq1gos4/HKjltleodpVRw4fjtxny/FFgFvpQ85/mP15EbXqkGo
f2fouQvyw6AaVLGNQTRVDiTv4WxQ06CmsUmBNIIXwy+GMcW/dyg33ZXGLrNGtfvWOCjRbg/i7Bn3
GHMvOD3yld32dTagBH5+1RZPZa0fJNuy/xsCJIhSaykC0aRwYC0ACUh+9DHSGZgmAMF0fcT/pajo
uqBabmaQ+rESrt+nJsr00Map8PMvXCUjSewFBtvBMO8LFXC/rs7B1vEBEYKHLqIMiCoEL1SnAszd
tZJdGl4JA2oCormcNkivQIcq9rLM08GNVzzS3Y6HPgnjAqEpNQPOaKlqAVDbyPlvS3YwqrUXisyQ
a7qv93ZACehi2dLpgI32qUXiebXq9Ybwrl2JVdmXsLonN0XAF94G8c2MD+dSWOO6WHNuBm8s4Beb
Ig0tm92l2wN6Zld0PQGjghcIeOG7nEyUNQJ6+1pIqBfXUkTW9UGgeFtFCjqfiOkt+G0ZdLzJG3N0
W4R3flxu/QY1CwLP74A7RxsqyeGlUE/4LECWjHXE58rIb+xxKAYXhqk/eBeeCRtq+oiUK+jkl7M4
McSxrZz4uPT+fKfm1vhp7YwNYQk94QaOOF8MQG31qjGVFjlhxq4DhzjJo+Dr/+JqA8F1qoO6J3gQ
gBcwoqsX4QaY9EI8WpmeBmKGaj+ZzG/k7HsFpQtBz0w0Wizkfq4KusL81B/x3MlNxhRjumC/qWsB
B2palUzNIblI1ktUTpVK63Mm7yOS7mLkb5W2PpWukT3LJ/7qAIxPWumrQVq53amLU+4nYBTzpoqq
5YNZXteyLFhiMIiUeJgyySnd3S3dcyJwDK7jBnM3GyoSpnp2xYtOcevr+IU6Q581Fu6NNgHW73At
zJ4t9k9uaI9XPQvJKx8n6adQ6PaHh9vBBZGxumtHSUYTB2mr7AAXOMEJLXgV3t7fZzL3dSEAOeKN
4U5IlwwBHz2rj30Op/8gFuIAPo30ZH1hTEskv4//UNkBMxNH1WY+OEfj81im5rz6+HXuSpgykrnW
Q2a0+8jSIYj8Z7BqY5OVLZ0IM0/gKMJyHTbaInmyugNCXbZvTa1cJrtCSepyjtEIVQ9MQZqkbSNr
2+cf8zB4zi/adi10IhwSj/nAdwelDbwlWRmxf4owqig6/wGVu7nOBU4qENQs0ghGL4Mw+Ca9plU3
rtu/SF23oYAdHmcLYBapjq9/Z37WZuJmFHatfeskyyw/qELqiSzkkn6LqFXxpWrLpKSnewlTyWiG
Grf83+lsUTt3hlL83TyyFyI9wes4KKNFXtieX4ruGUQ6Q6QG22gejN9kt3XTqP4naKKQM8smENMv
HtNfqCGNPoSjxObb1/eU60vFuI9d9TMLD9t4KfGxsD+LdAgSTx2KTNQnPUW3XVqVXrc/8YJlkn56
UqJuyQp6C5LzJyo9N15PeOX1oob5kz5rIRIqfZEMbwt+A1PZZS+CPI8j1pUkH2v2bvE/CZivMUG3
0FMv1oBY7ec01IlBOA7gXmVjyRyOGekdk6dj/e4mQ2K/1S5uzHuWg5i676zTC6MWQZ+DaAckOnNY
dsqWX0hAJq21mXo0vMkrRY4RYIQxjLVff+RAlxHPqdmezKxMKGAdr7Yp9YDA1VV6qtyZUuc7pJCa
/cNdD3J+fzZshlvLl/H65VaiL6FKiKpkYVbgYuiV1xqbLWWzZ2ky0oM1eByF5T+bxI/JMVyPH8jj
eZE3vgg9G/xW64BEMumCXZ4kthzFGDKsig/g/43OdFia1a/yxIw6qf+lEKrJyhfKBvR/0mpDF11X
VouAmEuecYhG4d3nam7Z/dSHnppu7rea6gpMCDoc60eNdTJ26R8PMFVjnJmB9puCaWxN9WWbNeke
1gLk91T6V11/78iv6FkDKZ42oEttZzpYcyFGRInBIE+/y2ReVU7VMsljbjOzEsu5YdZRxHR+fFEk
fV5ZAWBCaKkS9v0wIqKUyo8U8qDnBv1DETJzEUMzrsoMhYj1GUQ6KnIY0AZjRTKOy76civK1pdiJ
uoudn0ZcVkC/iET6QEibDlo6B0UaOKuOsrJth3rlOXCo5qtK/nJ/jqvgZPUuunlYppov3OC5WyFV
zvVnHpkSEEH/tpt0oH9GBCWwC8Z44pEDvpngfQjvLELTn2xstLhmK44mI4tL+x75mh3rlPFiSaoT
Zzqbw4cqdxOf4bLAQRF76MPUfRVQSYinYRCSTtGofMNgbSnp+QEF0FyhMeDbv7eLTyN9l0kSH9Ng
rnuM1r4a69wJok9Hy9Xa+1wGQAYqs0ctH5InP+9/X4Qr1ucl7C2YCdj1N2tnVoAEaghBQs7gycoK
+2+0PhNJ6xeZTc7GNLNPyhQnW6zn3Nh0eTyAKrRmb7W7HxQi6+kQ2jOuA4Dj1Xn+6mMSRhX/15mf
jDu5cqD6LomRytcX6sFMFHgzOv9iVT8Xeg231udBKxBETZzxeGqkv1CMRSFnNxFwTLcRck/fH0mY
D+jUo6gWdUY1tAemAUmQxUVyfgADriDW/ta8lo6rpRPlbkRKiqmUS2TxR6drt0aHDjK77NVJ2gXJ
bPDniHdVe80v4xHq8Mupa7Y+8UxoxbZiKnaXbYtpcozyEFFdY9pv6od3A+xh3cAgM2svjxGLo4VG
Xzzp1qpQ/Z6wOZ/+/1+mH5Qhq++6MYuSOrNJCg+R/6RUnT1sh6+mzU2VL6teAm+E+GinAu5Cgx8E
QW+p1eUqI0D5oVOWH8VSRx18kmv/EOOXW2hlGjptka9ikR7plMBxI4k5llJTm/v1yFjsSHq+OpXD
9zdxERByfSJg5lzN8k1mEkwf7vZ8U7UTurDCaK/FPoQVtHaMFtH0LJTkpGJgvU1pqTta9xvLszQX
EClZ5xyb44GHwqig1nBbdcKd6aqn4IsTyYVYxA36PNv+WHR+7GEsAz+3x97qCBnXCAlj1ve83tEk
tbfinH0YDpG5Ao11tgIcj8zC6Qv+Xq/Q2dIIRSYhlOJjVY78yg6HUClxJaJBoceXVTdCELOwUetr
LcTx0LSprTIPI6hXG4JZO8sgrHaxe9WDjQODkNELEsWTJ7fKXQPHLv2dkNdXGiTanEKWdVYBFGKo
YNRWYfV0pomWgYJDcikGIcstgZmeRr+sC+Xuvyx1eRoQLVWPT/U0LcTV0YmnJT/zCLzzL2rvNDkj
VjRj5F/Gm3HrxdIqgmRBYmDzozHotXzJ+jteklZvXfN8hAJsEF3Kda/vG4XqoRXs3hDpcV2DMBs1
3mCV+Oz+jes67U+uv/Ljc3WCimn0cEz/RZw1BNGLgLkhlBhA1PN1FROX4eH0jUM42LKWNcIRhUc0
9gAKruI23Ik7m39PSTQWiEpyc2FqOd4AAhda/CVo+XMlbEQFzf3TtI28u/5j5SELbct8fX9lGaiy
LS82i/DeNe7VujnACMwHevHvLWEZibbu6i761E8YcClsYe29r1tFT8ibqGCFnGAp1atah2XSihL/
doxAFOVYcNgOAwOD5bs8rqX6v/FDn5XEsmX9IWV63Cc1n5JiOs0eMKal6696a45xNXfwXHWN+Xws
8H7Dn+6QzGFYtZis8D24iia+70Wcl/mMTMOofhVAxSM34eA1fvLVzcULRAwsAL7fxVNqJRt2e1qC
5HbatD87iFpTG5G5KyiVhJ8REuO8+0GfU46+WSBFYB90ug57Z7fyca9NSb0QDk8kl+n9G+FhJzbA
yUgU5ppk+5uJVaStFftSEi4CdYna27R6QPbANGv6XioG/3eLsEaGUwSXejH+nKipNIIar4OcKj9j
3c2d/4XKFs7bcKp5Gd7e2rVatuu2P3xou+GotP2QxU10snTzTuKFiLHiAuJZz3RihLd6P9G3NGAN
7r3ADul9AC7SRGoN5u50zIc5KsGwbFvstlj8dgILvu6rR5reSdHv3UzVKYNuZn/tl3Am8BjNLo24
FsBpP9BEV5u3lLuAw54zNJSJR5kBHNORhUm82m+8vRMIokapGJbRi4e/sd9q3guJ1/+EODIg0WIz
Lk2/nvaAY5IjzY08WY6jCQx7z77DUOonsSxO3LIyZtd0METiPJCzyG5XOZ0/SWFleMdZAVjJDLYR
w7yW3NbTji6/hZrS/25++rrM+5Com9L6JYT94J48AvW4XvzgW2DCNxBARlOJUPaN1i6bLKVXa5tN
1pULyYX977mpMHWOz4voTIYosXbubunkSoPSrHv6XcIUkrWhBxKMd3X31ZixPSh6sTnx/mWjHYPS
zbsGBLN6wdzopXFDzfmT34NWTg1HeK/x/yMdwiiPZizbMdWF60RUj11oQmlbdHxcN84elOMtDVlk
lIjnmBMCQQE4ATJp5btOKef98nPRJXopnleyMq6+g9vm6Q8lomXjO6tUjFEJDUnYsvrBd5/hFATW
un+J0ztRatwp1vDSsHpE+5QOhYidX4EPLcd7iWZ+mZLPPX8CvAU10I/R1umO3jL5Tipac6JXXgpI
oiO8iL2AjCkhaknqZrhqMjPz3jvJteY/Q8/dzUnqiBE0oFzDdnRDxcjRrZPSQlFpsHXVEFYUk3ID
62JpEzl8XQKIsIQ/0ejID4RFyBC4mWzE9m2SabjcoBD7SbPZK/XRxAFfkivfq/JScbdcEvFYDl/y
utDQnZsrMZubvh0WoOociCjCclyM2Y1B0N3odQKB/rJ7FthQakjHnagdVjqdiXYPfwIe8aoqdmMF
cI60BfWxDszw/O92IQTlj0oboFt6Y61/KBTVAFf0nY9XnK1Rktn7crqT6bIqOVN09vhsFoD6To4q
gdvAtIL77Y84V5CN4F0z3PpQRtdy/Vl0zOXxBFV3RRpKRbJu/DAdqZOHQEMgf8lCXOzVNC5GDBdn
SCzWdlRF6620qcxqTKrYq4MPQsgIB/5DYZ2AJX7+YTBXoeZv9eiiUGeXDMZKu/+slhpiyQls8W/J
7umL+pK1pR3mi7nPRd774O1fdtk9okIZnBuuaSWgapo6rrHy6Xi0lqsCU1fAJE4qbKu45Wcu890Q
sr3dypZBoTqr0ctLxhUvDBjoSmqGX5VPNs6t1ia02aHef2IHlSHkSgID9OIBktowbVLNoXDjGP1p
1qIzJ8VuPciryhp2K/5XQ2IwMt0io3cswwddfyVfffDb+MmqH+OWgs/to1ecFQSVNFgfHqdzg5oN
qkxuXMWc2RtdN2CZIszKaaDxvit/lyDFzcsVosHwtoyJXFXwElLmU8B9QNDspPqKlGoAOaqXy32M
CzPzpI0p4H/byVQzelRA5jZD19v9UNo3HdkbaA1P/1wNk0W+D6hgivjK72U81P4gt9YZFeO8xHZI
nPTBY6sbpLP+ucM93T/jJrv84ileFF6RUxoRc4mWMucQUYfsLrxa97kfrWytK2e2P2AshfhpTYcS
0/0HsGPkjLZvdc8LM7DVDvhUFWLEd0i0rIk1hS0NJLwT3R+YhqgQeMJxSQIeIKxp0POWiqIqUKwa
kBw6ZAQLkJc4Fc1qwSjLxsmPe/igQ/La7+/OKwQgYkHD37Wwj5LZCBB1u7dHT5/DMrYgaA8vlDXC
bGCjYmxXwwZC2rL2JksPoqH6jiynvh/OMetu8VLXuQC50y6qvzW06pSkPKNcCESTr7vwzcjuWzeJ
iJ9J+g6uOJg53q7K3XJyD1aB6tT4RANUWE84o4VA8L+FCUFT7wuL8zKzgaoK2ziuFBxky4ZGmVA1
iTrnJcQUUqmk+gP8GsE2ryX8L8ko49m/bBazcmQmSWK39KRej83wx6IkQq7JeY0KASYhd2PYe0sL
q1k3AgEmX0xZMZwjTF7E0awL8u1EsK2EOSUNKWOX74VHh86KDEHweJj/QEyUifirvy8pUVChMAa9
cbBxFRa4aTtVNepypEghpj2ZmTPi7DzEy161Vg/MEJM7LScFdrJFfC6q9DP51Ta3udrszNlxqYoy
LBf2zb01SR+oh51VjZ3TOBzIsQUT/EbZcSpINS6JjsRLcRjRc3LKEe9BljJgvcHrm5MQi2VSf63G
IN4XlGpFQhijzyl428HFm21nR0KT3RIasc8qMFiEdbI3gSvty1Se9YIW5PrKgwEF9dbWvJVb9/YB
ru7M8yGjFUjRWKrGbCeaym/uJyxTiSN6frJaHl6Q3uKtSk9MevZiFj2oxGQxl7AoYoEIJ7MBDUGA
UCf6N6Evop0K9Ti50goL2xdduLhzYR00rsmtBEmfMWUGkQDbIboVOmqVnFKgdcGpvzn+S32P6GGs
zTV70FsKoMxYoAKK/gzP+hB/pnwv8Fw14/iqKrrBrX8dRe3xLY0lVjHqPaaUNJcI0vonDW5JOOio
4ezbuT8PlK3uFsr/OpHlanJn1F1evP3BnsXKhmrE8B8ktw0GTr9Gmg+zLrRbSxOZcThz1lFI94AQ
zMDd2Be8rrOQImZih2Skc09zlBTLUranAtPckzjZbyeyGjd4b+vpmVivOv81miHD2Q1YWaRGWJRK
EvedLyzC2SMQsEu2fo/hDzwF7GUS1kkXJx/CjzNgasJ2u7/zDo07J2dKFPfCdbmpP4ONtuA5MEnI
ukgbN3SnXE5gssuEXma+dOIsNA6DSQ+XFK9ATCoZKjiDmRMiiSueLYDD7De1QoJcLc0c9ClTZ7xP
2DIeF0wl+VeX1Z9rGDGDj01m3+fHabm8wRZG1sUgICcoCHzUidLIvMl92p5/EDVptJBKYxsOy3UQ
B/GEaVNDgKR2uDWxl8uQd04tuWEz6R2vktkj4QagbVaTgzD6coiUmTMkmaXi3supgh5chfLko6bL
u93z3xwQ3DqHCbgbEvZHXjaOgTDM1c3sPo39TMoHwqFEb/8Vh6VC3e7d47hRXqkslW1NLY7VhBOz
JJcfKuEPnnzC43ufLNmPuX1QjPi3Y7APAoKm25UuYVf8lSQMRMzPRJEli0UgZVlogz7+vXRMBvjy
RTjszaIHXEuoiqUlw7F6V4CxxAKjOphic3qWzvL11ky3PR52lpB5KlHcmc0ya1KALRVeTu4eBQav
RFl2MLW8IvzWHvR04ESl6e5td6KR54Vbqr1CSsjQdWtqbXBMh/IBEZIPauGKaYtfYo4QtEKBDs2h
5ibG3Gv/JUgzgf5k2dOuBfY/1KfJOkhI/zxI9LMUetV4JnnygAl6d6nGOtfKrVeiwI3R4wKaYCaT
Gh2IIq8SsJtGK31mvXrH7607/r6xkyWCzkZPtaINAyh1M9q1+m4yTRrRowyq0nZDK69H5HV3g6dx
pET2gjKs561K/nqPRlMfg8LNkqLxvD/EI/nGszqK+eK9XtJtzdQCey7Z5mfRrlc3nXCcnw20VbsZ
LrX6PBY+VyaTEcsUdL/FPKEoaeXpehVfBmSROk3b6XyLg/KH6/AHX+37uJveshlD/K1u38f6nrWU
yD2zB7KKdt8bR6NMv23Ck1bhhNs01+Ifn2EZC1H2j77ThEcNDnv3h5lq9Y6qCFjKyNTp3pykZcGq
xNtOrkOk0q+ZnusyA8Z4JqLXrBDTu4MSKmgi5nIIz2E5th/WqqATcKiN2v35EBlG4O0wCvGPPgT9
jyfWODJlVRll9yitRbluYlVrDKHoQD4slAnzoGENvTIoqd+RKyToniQXGOlL95TojWxawTTCIQQY
x55+spXnD4isEx6NlIAhlc8779zPsTd1Pc9L9W+IoiRboXoDM78LiiWmtY1UR3gZBXJTt2vj7SWW
gBjQ75ZPzEwHVtPaycNRdmTtn40HYWslQgarQ54nAIlXggwmT8RL/IKpDg7JORQ/iJTb+bjTpwuC
9tr2RJ/kON16z4lkl27TD9GjermcAnLZ9y03DDiR1OPlRhZBdMQsTlCGAGpsNv7rtVfYVQFZHEeX
2CL9AW+9hlBZcb80+Ig/52R2gl6u7D3VWtWS+11k1/NGUnIW6bMr6yoslUlZ0Z6dLIMvfghescXO
ctT6cbO6X2xssF5/nWwfkFrxZ3Qis2AuSnawTflDpZkPbM3etnfcUMP8JQKb/m53qk4Ae//NYinx
ZKInpDlGfHFVK/lEmqPRx5mnFLU1LShKSr9KizLy4v3t4N4oR1ZtG7aA/YvF+HSX2BFoyAWxGnmk
Q870/gkQevvcPq4zY/fZ2gcel1MorbDHzzbwCXAc2AAwE/xxgwQHLmwK6SnSk3/7Uvm5gtt23Gux
CJ+wKAv+8vposdR7yG/b+OHo1M/8dQfW0PC4pQ4EyigT80gKiJoRh2U0z8M9JfY7RC+vudj5LKXG
wL2nVtjmIZrdKkwHYRHgIrjksh/ORYRk31499XWa/dyEMKbElo8mXDBuc/w0JZ5T6EMlft5G+Bmz
LwfNAL7P103VlqZ7dc0sqAkWCsN1ZtJhyF6tVK1p/PKo2GMgQ2FlmH9CCxnmt942YxwgeFDY7gEm
s93+waBkUVUO7XMTnF9lNN80Yn8Bldvz6RDYxRuL0gy3NR7XdU+GPCsJzNbyFYP4usrntLugXHdI
gImB7U4b3ZVMKeHjSMQZ2hNrS2kzNsf46XGLB8EVmhFhrS0dFcCxI4BwEYSwppGIKIH0w9OseGox
wugMk3lnrRlV8QeqFBbT77mG7RQGvXfnjgLACkvrMM/jUx03CnbCykGKqAgkcswhF2d+cUuP+SWf
FcFPV2DN/IGjMmeynrkW6gjSxC3JU2zNp0gQa55FKYC2MyRDt8k5aZ2SRLt6r+LLoBj66yZNefnN
qH/A4JAU6ygffbrAhknRDpkQbKIfl2BBqRtPgqyMZXwzW+eeTgUXS1ayzAmydqMh2MxAEED4FrP7
gil18VK49bLcBXCaYWLSa1PlbRHBB3q/3bON54jWdsOSZBL2D2JuKwXOUtjQrTWFG/LH+jwGGFP7
bF8yDXkEdxp4ugGnwHFmqLoOYLsqIjq9BYYJDo6pL4I4kqq+PWR6EJ2UpEwM8dR1ZGHSm0m+wnEz
W/fqmWnbV9hp+yR3WDOchORdjWHIUcQv43g5MTZxMvJq7iUGliHg6XGm5Siq80ASH6cuypU6Rxm9
uW17hyRkf/aVwYJ/nQUg6dzQcHknYD1qYEwVEhhcVwoSOBQYFjZX7/XqTCjV1VQpMhG+V5rHgdB7
nxvmc8lAnry87gpSvhswNZL0f3m4KAiODD8BXGiU0LhH/DI7Tp49WvltslM9CAI2X3It4CvY5IDu
BwMmLpjReOG6USSU7raxh6I8yH8jdFoxvBcFNOf6q8UNhJPM9uRCWlYgWZwbzly29RqPSx69OD9V
tbpWDY3ZhYtjBVyAYpewt5vSFIfnOYz8J/VeNRKuqn1s/32KYe8yjC4G17q2KvI2xXmIylXt+IdR
Pe/dkQCS6KD9qyoxPiqxnb0/GOyrBIqWZVP8VjRFbiN0jsiSgX1ptkoVZM6lpKuDN9+kZx/+SKO9
3W+n/sucoqNF6DTYvfUieh9A/DQZD+m5CDi2mfoYBUMX/r6HrwKspHmUOQloqhrU9YpU1JS2e/r5
SwS4HlFB/GbsxzcgjD9Q30X7oy1leSPGki8/LjFR2u15lYg8BMMM6MpfhzgPLcn1jsIU359bpIgI
/uBsssv032EBfaBXpEKyZQBF2azW7q/7VNy+hy/pOXA6Wxwgs7kshyuGPbFn0nv3xI6uG4xvjdtL
dO22VTXNQKjFI0PPrQSDONhPtERoqO029m0DjoiOgt/wM9w+8GsTqnNotkQf+tVba7+SS5lw7SBw
wceWv+TBkm/7LGPRg1pH6OB12iNBbch6KaHHPGpDIC5LSPlr2Ps0SgMCGTKs2uxjM8/v7/1QHZUG
7tF0sjxhJjs8k3ndB7drrTmU/ABRFAt4bUtmFUBymdnYDDeFxnQIHn5ea9uDOp9ZVrn4ISmaW3pX
UN9dsIAJ15HQ2Fyr5K5AALBwJ6DTyBO2hlhGcgLkph2mGNUrMSeSYiCplvwDGUfkv/OsJLBsM4Hk
xKLrodS+MIzqj/nMmsctNePWYZoEBsI3iI0P9VXNIPtpYlAsrWdG5sc88Xn6GCFk9Ds0U9YawpNQ
jMOrKZLEI8wC8nF1TfpCBzcOf9VtCDmLVxmUpWFK4tuYPwM6RVAZ+wWU7NFq98+qPWK0YqRmjvQd
y1RWwjpmmqDS+ulKO5G6rqc47B/jwR/JJr7gGEfEOeUHxDc+Z5lTaHtclyaYp/6L1KBKjQYnV4H5
aEGPcGCBoZ2s3vNYE7iiYXInO4uwGxOIF0zDJHY6yWAt2qJD92mBtOHF0Giz7KrHkQ64q7FJFjG9
Ej5Vag1W/FWyadJMIhJF2eZz8qwXbVQ/bV9UoXjfIgtIsrxdwo4HbqXfab8wiC5ooEdnPQQlqpwm
Y8s8sjxRilQN8oRDVd+FHmo1VgGywygLdr6Wibn0+9UPgWeg20PC+xH+5kwNohPe8rU/bwqLeUX6
+pMW6C4PhQP7pAvp/zWXnzk8jq1Nvc/9hycATSt9PhYKAgnE91hdvagH5pCUrOphfO2wtPIGtw0K
8lPYMVTTb6BElRvofYXbqJ962cNf5Dto2clohFQqGnJVWxRji4zaWjmpjzf7iuPDK0kzMIMg/V/q
/s4FwxyqRXIvwGRkvQ4W8tYE4bakP/3ms2hxxVIYW9U8fiOwU4T3TK8Y55Lf38qhwrwMK5rmZxx9
z+/rzRfUH/f59O2s5sywtkeJs6wj959APe33bz96K2j8bOd/Rj3RfStPM32FMunCcUXTRfTaAaPn
/hlVcfbw70Dw6F9DEDWN+O0Jye75ikW1Sc1L37Uzxb1ur35ElMyqLiEeCXPoQl6Zwav9rOFHq2NL
7ik+z4fC760QYY8d5Ze4xNUtn5OfodOIS4weuTs92+xy1rYD0xct3bvS6dGNTm13tj7jM8Ooe+LB
FTuiMemU+6FDa+WFNhz8k54kdVo9avWOjjMMcgQl8/MX7/L6ABpg+Go2eX31FtF0FB+uuXMlI9eq
srtXp4r+yVdB3/f6nK/o6M0HbwjMcTwAleAzmoFU1M2x0TfFjm5RmuBrn/Nli1WW48sabu1mlqCv
8KsR25+UWfsBQACBDaKN0Mfy/tnSY4psBnhkrhRxQvTA3OQmAwa4E/+9ZlXEUhKNrQZV6KdN8JB/
PmaJ7lZ5w0ozj2A3kG19CQ9yvw4aKIy9idtvSeijITKIlL5s+UGN8F43gZ8dNmTvuio//oQ2YKXI
JtZVvaMu7TXexJaWw4tuD/bbFv2dWEIBzJhKt72aE44BbfAD4zfQ6h6vF6eEPLU/VYnMjNygMPDv
bN8rZqKU7y4Jjte+L+cjd2522iMk6plRPXF1mGK1EVDAh9qufZH/yD8cKDp3/XWxWMu5t/ma3sq+
6657zUqsNyoT5i/TClpCZCDWt31e+l0kJc1vBZxkbDIW9FuLInzQz/kKe7QoxXmSHeCulomo7cgt
GVNsbgDb4owBhRqHBAO3XuGwhqefKtqbRrivrlXzjzcFMcz3ZQT6MDJC1yRYD1/sR/5wLHgYk8yk
+IgTYdum3anbhf07C65VczlEw4M6UEhjjliqrl12+aFnfdZ4HBftWWR/pNMjDuRjgLxA0WQkjVZI
e6I9GGLpNthN7oanT3jSp6WD4gURymsKPEmA9FvaPaFHAn1U/ASVFyx2/yU8+0jcSWf7U0cNq9QT
l0tpvq/BSMLw3UlENe2eYonSzoM8av+BmW4tKHWyL5S/mfQTeMKwB2khjtQv8LLPIYsNooCEfaW/
3Yvja8axT+PGCsKHW8mntKEMDKuKX2G+zT2oS0yyNNIwgAd9C7CbFGKGSVNmLN9+mpwB0E7l5PRG
wVpMYA1ND2FvjEWRDCNXiQGS0+ZOT0t1z8QaKb/yJf0rs4rCAlrvHmDirJhO2L7deOk8rYO2HwI1
rgfqUQiPkFq1EQGTo87aUKkXwIiiEi8bXPY6eFzm+tEgj2TJpaSqbiyEVLjNaZjgVw1sHKPTmDMD
1eq5cJ6ueIXpOPSoyBRFdvgVgeL1wt8H2vjA3GdVnApxoml3qGBOOm5oAO+qE81npvFgnjxYtT4R
kgHI/7FSvy/17dFLMnZwr8/5VWKbPBN9ImdXGjYX3YG/YJ+hO2KQdHFZaq+sXgABLJwA2AO81rt3
99ynubxP/Q55TwRIzNu9aPfhknVDV9z/hj3nYjc+9OfZnlYPiXxQw9Vx0qxPeRzy29ZrkRO7oLT9
AJSEd0IDlI3MkvFlil9vtqwDfxVnZYsI2CevXjmxxTVtWrva/Qu6V5Nu8Fx2vrQhx2M9h2kS+nAC
/QHEf77k3ubcpTNAkV++iJOQAbv/DTVE+7L8TFN/LDxDRIVwbVAbkxYZJI8vmSokOpL+aABE5u5e
pzK3z+Lvu9kZ/dGLYtCl0XkrlB8+6y9umF+pf69szd1npbHJXcbarBDvFifnlqmjHzuTvExkD00e
U58xhHQX4S11SVrYTnOzWohApjxDLLv7RdT0dFaGHxYNBBV+6tStMyGNtZ6LfCbOG8G0c1/y6SxW
R96XZcJa5YISX0fh5m4k+/bxxQJZf3MxPjRDimDHbvIDMiLgfmMW/5g0dwWDHsyvisUGovZ0bZ2c
ibhi4I3VW4GyomW/01BELnfa/WjLH11GUnq2gV9wGLLaCLAXhlEkZfI6kocUUQIwmYhMdQo9mTu+
EyWH0tqcyHkWWRfZ75MMES+33ULxKLZqhyXHKd3zlAmTJuNyhaLrQF43rX1yRcDJro5ikbR+7TD5
7yErXcwYh3EwLM7J87wHgtM8HyY76Bw9+ct5ht/pQNlULfoZZaQgE0NYe5zqAcbjRYbgRXA/jY9h
bX9DZDZnLZDHuLhIORtrwKCfxoQaRM5pdQ+ln4yA/7oGVkqSSlQXXVsyM7Vy0P7aZne1ThAVwsK2
F4DTbb9as1JOPh5K89DYQ9idTagI2ySUAHhTfMjnS32akaBmvJmn2Kl6qG2gvK8iB3vYS+2FRxUb
v1R/BgAYcBllG9ituCmuxSKcSTpOPVNyiWT0KQ9N3viYntCAfkv7NyvalVUDpjKkSXkG9pyUTNkk
AKPjWidwmk/l1fDBzFrzZzjcFYn5KnyN+yc3IhifcATqiVuw2tnJN/DI0y0ZILr7lKAhJLM83a1C
JApVSnJ09Wfyl0DAcytlL5/MdnXG0hKEPWVXNCqYMls03nrImMvGYViX6B9qJIpNkfB/nCx8VeJe
LEgevuzIS+9YNrpQqGBtBn0Zcw7NpTGcW8QyN68qFUEMKa1s9sKhrnyLuUjSQ8kmHttcAVTS025p
A/sdBRqpaCkAHsWk25Q9DU5AiJfsMSwCCnOiT0eOxgvqu3KGFRshoXeaKa+CBGTnAV9A4VJlvphn
yNVZhrW1TZyRt4BVAUamEpdwFfKI0AgadrbnmtTqakc4VLHewGXohBfD/Mk37aC5OfXjT1fd7KzT
sKMqXMKPD8MIvnA+hqNEUZ+jkSnsqE7b4Ijx9+S5xRsCfAj5oIZ0qGwZCA4yPL/Yj0gfWoJXBG9R
bpTaH4MUbzLpBobh88S2PSln0WE5zOQB/Av/DT9cYrR2vWeTkCdP1rHepRSqp2AAmaCicgh35Pjl
TShcz6q7vz0nIqk6wONuLfGvEA3CESwkVbkZ0Git9fLRTpSU2ScyP+uXpBdz1Jtzora30CqjlsAa
2cZlAEjjXwPWJQ5Yw0qCW7P9lZY5TPymsz8tDeg5rZql2wdndnJ9y0BGOw2u56MoAqAzWM0aM0Sj
n6W0vSAnqLsZvhf5ohEqTrwCq1Z/XvYY02dznId0oughZFQaMaz+aP1CsMV+Nbe6ol+GW3c1s8YX
bOSS9yQXI3akT5i+0UR3tTdN7nJ/py3Hlat4/oCyEGc6y5rcWxvSzS1b9ct4MTcE0zQRFbXSWGHh
E0ZN6N4d0ac/95kCmS1I8V6ns2Sy6LStRImX8WJS0gj0h2dnKYXnw0YJPQgvkgiiGuodoypszU13
5NVbfMRqA5K4l1FL9WB3PG0mqmI074sjdqC3XzcWBBW8dg5+im8I7qSW27MBaAbFj+3mXdSd1E50
xEMLjsTP9/xxJ6FCuHHad39xRi2qRXsZSizaPguIMT9JUbnH9dDiqf5VZmd/SA0mTp8mhXzvBVBf
TTTWKb2GGBCxSdBx/xNQC/COsSS2azEnzhSBnIvHR90P+5EPY9KlssxaQY/kwJlQkglF2lheWuU/
QjH1lxiVTixoxB0qmIKKrFZwWFVYR8wlEMHg9PvHUA53elcfjcKxJk1S7PS0uPotnGa1P+nnkTKe
zRf66zR/vJUiIv1t69vtQwIOX5xX5ON5DNkqrWmFxOz20/D6cd/1c8Io717fCQf+bAYg03Sh3vxi
jXmSpM4E/MDwaNr9KdKTDVWmBwRUYPO21beH5lUCDtkoswIn/eHanXh7V1W9rWk1zvAUaOdsPQuw
AFt9CBVnSDwX9mq5QY2cA2Yov7WtyRKslGNBqBgUeWGTjoAxu+/qtEtsbPl24GGnoqkteGnHl7Rv
YFb/x480Bs6cmFQPRMi3cKnFBGPjvdiPtb6SOQ82+E5Hh8LLNivYoPypnYI50BDRvAwRWp+Peirw
vEQnZMDXJ4D75QnAr7trJMxzNvz9ExseZB1Ec8Ah5Rbio0znNjqJGPDjFkk2r2rJpWER4Fiiu1n9
Al/qZjG6XIITq9spaIQvVpTQGoykCnSra0f9JCUPyGR5NpAQfOZf+abg+VhxuovLp/oswjDaz8bc
F0dOTPPOaUtSyFXTav/K2ANy0WchL2yLxbwA8Wd0btS7xfH9B+EHsP5vViOE4Q925luBKWCFo5Ck
XXUdSoTs47t57u8QAx2ErcCKqqokDQEvwMOJPbQzKnNGNVhBwBdlm3xpN3qHdR+gkkpKRICZjFyF
o5IHvYOZ4aSxmXPLOZ7v02SPCtd6Vzkl0xTbmrOJzqlfvR4OyilbVDBQMcrH3Y9hp1LAokNGPBcI
R1uJLv5rPlM4//DXEbkjllznj2wK6UYvp8YKI5LJf2lmkJp4WMyGdmj2+CyCw/ON0pAP6yuE+E+m
3ndeB8Run+AlqXvrz3EM6/EotvPgcs9SRDGL1EwTB80LA4RwFqn+b1qgydzErH0BAPAOAkEeWPQc
IC9PISyANYNzWH0u84GLfAiENc1j2pfFdqHJy1L60HXWbp/StWlLwAJg4E8N/+CdUDJlJzNbeDiG
qyyS8DhkTqex1FeAMgz5amJ3VUBCZDmcX72HHSsQq9Swfw2NO7UUHtoDpG2uTQuglMeeG+DCT0UK
+4GUKCRW/VYtljy7i6KracPZpbY5myTYAGg6yL9LGPJHh/zv5hHv9ZtuwT1vxDzIoSn7jNW5TLrg
pdIn2wOW0/RDZ8AGWzbyvzkX294oEl5cg8WqPUhYUKbt37UtCSau1z1GQ3Jvq/wVH8Z3gRNbCYd4
kS1NkaQZWEjouHfuTnkJh1heNA/15jrBH5XQUqARKGEH9yqgMJO4zAfMIFTX2OEdjiDjujNByjFh
KR/0mnLOtnBOxlu27VYDhJIABT5DNSukhj0AQgJCknpPE1kdWyA658aJWRzd9C7FatXacTizY39p
TXCZPbQz+3Z0sF+79MQ1z1+aQQ/LQpXhPwd9HuCZK8JLmJZsj+a3J0iQ1ZPmIN7JxMl4F4s/f8QL
CoKcybTUu40SpE206pSYBUWqzt/7zp1zJZ+YlyVZS65THv5plECMQO6Rgagi5Wm/6okPCiyFJwN7
709Rh5yU6YLb7W/EI2PFUtDqljEuYcKC6OE2cP3EyhJF3TJII/XUeSGOqCyTucYAFgEZRg4pQymZ
0ZLY1v/OBWV37MlheIxLJ01ZoniS8m0sCiqMU3LZt9kG8kZAgUXTlufrlXGOFq9AHLS4Cx6i0VHP
tyEoE97fuI/zFnDUX9d1QyxI24U8By9EidJSuvtcFojaPlr/3NuKawQBjCm33k2HOI2xW1S2vodf
Nn+c3q84ZE/VxNiwt6mGi5VMPH10bmqb/XCEzU2OkN5aHiNDrCeVht5n3Ww5EUyFJWcrZsxeSy35
eRQbR8x0fX+g2ZtHrGqh0N6X72LebSt5PijxxzcBBWGNIelcQq/iXhQ8ouYxrh3XF6GWTbjLub/O
ipJQc/+MAsfNblUL2xKt0gc9LCzhje7b05l2WNeqQwheItAA+TBBCJO7ZxbLJ8tps/sCZoWugaxt
3Vt1sg5hAOXYNLYBur+aRvl2hS/7bERIhoS37bSb2fld5yybXG+PAWGipdQgVYTmViLabymWW4jH
eyzi1jSSJPmoHsiHcHzcQvmeNom4dyGcuvs58I1VgUrS865suyHukBnmHT1TGDlL+kwbJKN4taSq
UCCoZBsIjN+pJxk0dfMiY0WdO02fEZw5L7OUQzlh3NfLyXQ6MKsWEyqtM2wBW6SumLwWd6yGHLXv
RX3vTl3+fjDC7GbWIW1nGI6KI06rp9fK2Dava0mXQ/mDPPYgsBJZSJ1JS+3sTMLfylqjNyzqt1eP
aseVLeJ0E5lbqYMG6KJGdilKTOcoZzuxTceV39y83bzF1V85kaZ2aHJ0Gvj9vYJyC/7Na/D+f2Xx
sfoWOlBhIdOG6t86nq/mS4Wll7c+UEmLyFfuMPBbUdKrWKWyudeH4jzacXeEMBsk0tyivU/p/ktG
pXvWNLs88CJoFTzTB09vaO/3K+9TXNoxDL+EM4fuKSEiHmkuUgdY7n+iKfOmHFKxZVNWRiqSNctz
2gepvg6uD2ttDvH8JKOT/IyF1HPLnqhkV0sKlYGj1XsvEQRJbh3WgnH3coLSjMcRUfa7MWGWe6T1
wEcEE+074LK75EI1jZeK3Q5wmnqriD/YImPgi1HvQPQfkEyDXLw8oNX/WMq1AF5YRlZKCC46t5BV
f5rN7Wf+0T+KNnSPJZKhR8NgcvFrH4HWQPS34+/Ht5QViNZba12UOxYOlmz8J5y3BFxYAvK2jCFJ
AYoASeuhMw0xbjG/RRPPK69ZE9J16ARBW4cQduAeffwPhEmwp0rBvdl3qzG+ZuGiEGeyKz3VaRFY
1EOcIGLyloHfllU41asgzeNoZStwEL9x4Xr+xGIK5ifvtwLBMeTN0dKRBLaSC0dfjzt6ptsKkipy
zNodMQmJf2dG5WOJLzkRDBSrJjqhfTIHuFSiF7X5esPSTgJ8F6VgzeZquoKhHMVChd5dTtxTKg69
sHO0oxsQFxiiyjnfknjRx7J8ZneTeFQSMLfTuO0ZDZrXSN7Gt60o8zKJqrVjZyt38Qz0N+4fFVkG
92OZdTMYHruJRu7e1CVGz2F675ZGgeM16xZ/ZehN6trPqXaSm83Pnqk8AEXf8moPUvmC86Y2paEy
EIQOK9zjayPcGE9hvdL97CLVC2LzXikF01er3vmv3Bm3OTIWxsYX0NmNRbdIMr7egnMt8yz2yiI2
hBNMKvLU+ogR1/lOYQOWKrgm4TDXTulFEMqPlp0PJzNMLD1/YCpH0nKjSANSYmpl/9CGsvK/TK3S
HFPbeEiR64LL94WTyZVNmFPywS+pwgcpHZ5NkKxQnvmslNZA32dtVoEaMWMEpuw1Zs4HGonJHr+u
sH1v1byg/wdfBZyRv+1K7ODcUcobQixljZxW0IFwAe7S+n3WJKB/upcgUxgLv4VlJtloXsdEZVLC
TNSQC4qTh/sytmTjFa5i9dXn2eBUEQZxDfhYyRThpKoT0jLAVuCZkb4uEQk62rHZb3qrSq+feXN0
DIbvt84HFl2S6lyOen0tEGC1DYVCm2odJATtHcavECIzS48e3qV70V+Kpcb1DinWAoLuw2JXC7Tf
0m3JyELm3BXOPNc2/S8gK6w6OgS+jUuACH5+C33BZh0hUMFP6PohmtRvd7sdvNOL4Fgh6YfALxaa
STpKAl6AWZ1tZ47IekYVaBANO0QFZDUkF5BBdgjFbi2pQpkw9emt9I1T12qF6biJBinNZNQe1rdc
DjGubbT1ijj7dYNhIIsovLgiHub4kDGyKqutevQFvIIA9d7HckEbmuxBRJn0aCEVErd1mybLW7s1
CEi7V3Rktqnql+i+VMAc4wWPC1Sr74RB7rhZG3XWi8WCVuax9SCf10uuAoUGZiXw0wJOWtTz5RLT
+LnEnQ9QpyAdAmolpyfTIXa075a4iBkNbfXeXjw4FkyIerqzZcmSHkfH9Qrayj+HQmi1Zya1J6xJ
D4WLs1qU1MAqkzEEad5FvEMIVPu2ue9z7uiwqKi/BUeH+jyjpJMFGZXdxXdd4PNAjb6ZrssIMJka
vtl6h58tTduiQE7r3iv/k7OrEu2NCNtgJb1zU8PSbp/0qMRuU8v+sEdOKloQJWiSqWlEefdTKUi1
Xj+F5PD/F4N6AHwVdn1eCJ8euEwmX1RXNcNxpK1WiD1Psmi5dYhKnTWszq2saaukyzmpB8IPN2aT
Ej3zH4a6y4ZPs+LJaLRs+vXs47HtxZzyLJsBO5S4FErbCt2aS1G4iLTV7ykXhFDCs/0uq+i09RXM
RC7LjwIbaIrqYIIM4IEzV6q2/wLBMQi6+efu+BUl0RLmOyZGvEbCAxtkIe9seS5oOjpyZxccQriy
nloFGko2Xenk5giyOylnwRpCQllv6JI+wBDEYsEu7Kd/GqSe+0e5tMgwOBU8rvQPeg7p+ZT2Z77R
k/6rliWe3UT4pAdNxDa4ANLVfrglsJViOxUPNk8nwu0pH0FV8Vx5EXI0Sh1P1Bezdpvvu6lSDwkW
mRlOD3SzzNJBBJcb3Ry0+zO/lgzTV5N6Ut/RN6QyJ8pC3IHP1HFJJwITLuYvDQKQpPwrQo3lqKKN
ymR5xQF/8vgnmXDVbnfw+pOJDVxWztjArVQ9N5HtJB7hoNPvDWW7v8WpMIA9hMtUN+Fe5gYmCFTX
3axSx8i6dblkZQAC1VG8o24UGl0WT1wS47uU7ceuTV3rC87RCx4Ajv0sm1h2c7NGbg3Wl+3Tk9Ra
zSEI1fxAK/FL8F2OxDpPfE1Bbkgk0BYUzEAo9o5SbGIwg5Y0WM9CFOgdvfsBKt1Au2KxJLDSIYR5
G1ALA3wlepGiH/+r0l7o1hBDllSxdWEjHYYP4lgAWu0PNUdY77LKhK2mHYIywLu1iHtcuGAqBDqb
y8Tvg7fgUzHGGk02gdRJWBNQeXeK1q4N2L0q2sw++H2Ne9KQtClSfkAn3811fd/gFfMqfVkO4pGr
ItvuT3WeSkkelHp5dU23jL9gv1ni/MtaxHwuKdQFozeZwemAzzOp116QxqxLxFvp4xz20X2nTVcT
/dreNsfSodYOljNiajI9qqd3F0LpGx2woD+zL962Kwzrer5MKExKnYks4OXqq7AoeDKz9W3hprAy
p+vz16XtpoNVhL7HtXo0WJidGag7sYl2wDB+C5neLy299LlpsTGVxHr+ZAnPgGDaDWQm0E6uunQY
zM+G6hyzprZvYu0QBjyCalRvmce/OCxmA3nzPHkji5BELHOlQ9ch1H3bxoTgoaqdYzcMfv6fCb3X
F+PwTf2E4UO2iI9ngjRDF4GJf08ek+abySWKDOkSqIWSxYfoNLj0j8FILGZbGg/w92TqTS+uJ21+
fO+I2nB5lwKNxeDfUmuH+rlKdZpPuNECbv5OICf8Y3OleXw81XhjlPofXZvLTMfkE7u1Gu7FWTv2
Sk/nNAnlSgy8haAgSR5HHyMiuhcfck8mOoyLWdRJ1/R2KOsL4VnC1ycr04xquAS3eh6LCU43in6C
Qme1bICST7ymaNlpmFat7SCVnwnzKwSMAXL4+XzebgLaxbUJu2exVNytWHlZDmhPyijyR1X16nwv
bel5ChZ1f1apMMZDV5P6vKzawIyKa/0rcFiDOxQluAreMK5Lx20IzBFbsRJU+AY8jr3shuoMu3hp
++GyYe87nmfzami3p8vXZdWIjHnPMgytjvfdM6yeiNppJNgT+gbzA7cw9VMLAnKPVdc+cpJ70TH5
kWJAVNtcx9OInVCoCrHeEBrPXAQJE38E4OSM9+m9UvkD6oJuB+4o03jm2l+Tg07Yna+QsFP5zg94
PEB6ZFX53piaeEclqoM+6Kmu8GGDe/UNf7scb+18XjSRedM5ovhVKwrcFTsbeIwQwIfValP+b70M
sTIhFMgcwQlb/oOjgO9qFT2UjYuxykp0oiZlmmKyC1khpBb6vPlp36piBVaTlxJK7EDQDYRloRwz
lDOs0XSH7NtZCg//T4fvHX3UkP2YXO4hP1eh8uSCMEGQjTqF6TRIQ2J0iJLw1+rpc8+0vv2TsF7N
B/twSw/jG1mbG2PWam9aJVPSuYTa2bNERWl78OqHQSuZm7YK43yp/ONwosoGA1kpPwvDvij2O6BG
HOUIZZCIzsArtnmdx084XWYjaqBuf9BrLZGB/7UItALeNSC33Yrh3iYvJo0Hmi4Gbqj0tBvpf5x4
HXCLw+3edny1OkX/MRJNHrsWxohndsDR8/6CDJdjUhwWhLiNBv3adOXxmhHM7v/Kk0d76zHOda/i
wyXLg+o8OIkuTFbbymbMIUzrY67H4y1r1kqLU8mCoCBzjMFVX3fpMRiBk436pIWd5rM3Vt+6FUux
IJJeJOp5oPxdF1nc5aaSb4juA5rl+ycLIPJRcabnY/C43Epv4vU6xfJt8qUuBwtMv7fcBGBz0BVo
BUmvZ4b0Phd5kSYCdhAETa2WcGuR1gn1uhnbCuiBOnVPRGzxLiVXSccFbSZrmZkGA4+yDNGbmpLn
5Ut3WkJUk85mXJnWXVov7RGuZVRCBkCOJ3TKDC8kCnufRv5lyEjZOwo53cJbU3adhbcBvT9+1tHv
uQ1nj5w/+SqTCDZWVmP7HU9YjdyZAOANy9hX6FF2ELTriGf06J4FK9NAYjWjpgubxgvnG/1SDuHC
/S2a09mbxeyfMF72Q2P3Lr3avk2IFncT/Jovd06aNOyGAgpgQS3pFL/8a/xj78g10Ppy/gZpkv0U
M+7jrzcKly838QF1mgKKD06ntTpRH+qU4g8w3zIKj8M5w/plxsUvkPVXEdJSYctPDKj2qq+s9M1z
pEYKAR0mhCmV5O9mqlNr/5Jr5rk8Q08z8a2Xin+R1ewrYiI+V7asCnXNsFN4v/ydqMftgrmhcMMh
YfXBl0pyy7Cpm4GR6TA8lF5sr4LYgt9h7ZeGc9ssX9v/8oEi4xU+WCAhPyK2wTdsHURSNjTVYx30
oXGWjT6pvAT3rsM47SNG8L6eUtM8MjU+4y/nprUMau9p9QztTnl6mnFo8gKMDnuVjbJfehGHjWjc
5f083YNgqeSseLRUPCyYEjML7/4uMlBUqqz/wR9zcnuaQKAsMeY3pRQ5EevPjuPWqOokETdytQ2A
Az9sIc3iKiNGdm2hlzhxAMFU3Xd5WPtUfG3xe/4zt6YQ0NeNYXzFhwvno85Zdq7w85z6jmNcGzAN
y/dbhr9iEA2C9zSEX4+OZEqdNbypbVQnghROIII/ckOmmvdW1+PTHGU+zrkHS/RUUgUe3JnasXxw
kjDAX41sQvgQYftelyhIlk/jqZJ70fD6Di7nlsh4aWDX9HKZ8A65I+bdhFNn8IcbCfSrP+SmldCt
8Z6NVWOWWXdZvwmYS+0gLzwLUiKMTbwrve/FgHGaCfMRupTD5PC7Ilv8Hr5kMqYxHsfBTc32MR5p
xL4IRj7Ri5l71IEbY274d34EacPTuymYEy4l4LyS6evBRCgdHuCc+0wMJN1i1v7pF8Eedopgg/wc
gcGxo55yb1aGTyApHUMCdNn/8fCqcFjy74rfrnKNiR46g8LK4oOne2YCyq6Qfs3z1fn0dbw2EUFs
nU4Ag60OVo5wP/IOGfVBmMb1AVbVjcLIaRqTFKKPAlYE2LslQzDvExNRgl8/TFMDd82ERb4l+mH2
NVPK1vRAArJNi1UC9JGvL/UKeXogFsUcak8/SWuSxybbkKZQCKkNYFT5pdqV71RiVP9I9VnWfWnm
Nm0+vX01OC4OajSb5Khq6MLF7e6Y9VEUnGR8bKB++EhRRyrm/lYR3bzz0+YphiVpfOgjjCnALH8U
n04gWYgJQGA86A9IacW895XVbKfvzHEnrtYOol07AsyIJThhKGUG0lW0RnWKBde1+eJI4oZypoO3
+S5gZtXEGk5BDas20iPiM2E23OU5hNkpDDS/XsDwId5QNjb/xccZbHxgxrPAcw7oRXBsDfRNC1Io
Jxq3gAnbU8bY87RTwvxLmp5oq57A3GoCf2Lb+NBPZKbLKQv+ekim5vaOc20pQYvgLHEP3k4ZfwM7
Q9IT9XJVwgxwKkP+WQXt0aj3zEdcmiQuqk/1vTlluuazr4Nlt2Dx3KkNbUD8H0Q4v/knCyIBPUJC
SDxJfqeVkauESzhO7lGY4+d9rfCgzaWlsimOPb0t/749kFsfDg9sehHp3pNkHpILersru9wxYkIj
tY1B2daHHSBDGSUKG4ZmUNxSHxpf6RLuCq2u/kTNwnQIJP9gr0xVCLVXfuXOWXji0tgNNI8CaRI5
zsE5JtpWacAtUugqMYKFaobOEYCXkbXgqA4UmLT9L0PbPo+pjTK71Rs5WVTkBNiWPhTXEMbwEGT7
XO7tCiLN7YGvNPfF7eIyyCFy5DVM8ebGU0Ba73zzwVK9eqgRHTEM71/O4U+O6SPsYSkVHhHIzGzT
7WCQmzCbkMWz8/VQc5+BC1+qtu0GYefr0P+2OcMFsEIwA30RoFHIxfLai497vUfbktDkcmiB+jo2
bP6pRj2u6jTP+xqivyq4BhRoO9yQSHQwB37q6Jo83DwH/PDTNNtGgW226iFNzHSmJIKSkLvgUk3O
d42UdzGeSq5QbMHuDdWSa2uIBENjp0v24hAV8cIMNgYODDQdSJZ4sO+8xrHtWzz3wcdij9UuqlQw
rARB51hCyR4P0OJIi2NxAfrHCP2Ohgqta4v7A8cvPXslOsanDT7kUXfsoxelMETqyHS8v9OUSj6U
XIg/HybFkPsF57j58P+QhzxDo07FcW1h5b6jofr3OTScRwoIfrSy/Srwqyk0CxhWOtQBWYQzxo/X
DXNCnKqFANLfdzb83mNGeQEmeGmTjHLHhDB0o1n8Oh8A4+MFBZSFalHGPW5rDbDhwYrIYPPG99Ug
JkUSUtBNAzgKBAz+aOp9KCxALuWTnpQRehcddptnF0Yjy4z/h/fW6uuaG1cr9ASLOlQfwnRMSacf
wfa6CbzCK801VHr0lsvNywiLCY57QGO/4IQ5Uqg1NPDMZ6IXkYETimef9sJnvDxUFKRHqRoBsc0l
v6UsInQL90gBo6j3PA0P615ofwq+9a5Lhfp+YCJWpaPo66QcQxDt42UPJzmuKTHEr7D5EknJyvL/
WcHEGdeyYJW//kJsUoAxg1g+Jxfum26b6SWszw4cOHxj7wcs/YVlgE19scC6wiPhv6fhD4WXTMcv
J7OSH3Wb/9KR+hDXIpReOwubD5cShMnkDgX73R0U8rVtuAiFdonWCuIRzE/IbN5VtoZafZyvJMdi
v2cD5j043cvt4eiBnxwNtR2RhV5cGnmmfKqmTHkoekPv4oagCcb3r6pN1SafpDq4bfNps/VH1RSd
gDwjSxFHJxMzpW1Aa5wXXyBvHDFcDU5iZ+j2rdYGJ/eqazBmKI7tF0HecmL/ppTzhpw55XiG6kgL
swD/9tF2thZfRiSwizqtIDR9zy4GNmvpEgieJdo3ZpmunU7iH/AUAPpNdvIB0VHEBnnGJQ+IAqgn
JKM09qhed0OtuHyPPMaN4NuiYSQLY6uFoZ1+leJHCNHr1svOaC0x2BpfFS78tGkJJmggG4xEiUCm
0gwBEEgooKSeFtchm8EYoqxZD7nMqFM7nM5NAYgfRGDLhcbZQeTQ7fixqY4cusjVuXTJlvH2KkO0
ait9TyuSgK/xgpsymr828mQ+gH3oNtBpY+5wV573uY/xpm+91XaLmvqTAV6baRj8ZwZD4JMMPtH2
p/nbthCupb8A20Fe0PusaPhJ4bWo6Ka3Juu3FzGP7h0VJIg95Cke4xBtdkZEWvlylqnOr8PhI1bq
HM24LhEYoULsZAyJw3qHoja69b0/Vv9YkCuJnx+HEUnfhA1CvgQUhPwZ80wO7gcCGj4Caow7uKfZ
9HH+OpwJONs1qri7RJxKsNzLGT8+YB0AE+ur0gWsUmwBojZr4n+6WMCIIto3UeDKjg9QBzt4sxoX
6UTE1PvABKung3ZdNQCGNbwxVoIRKG8h9Dwz+cg66BwbEnM+mWGloEOdCAx9yS3awhlZGsjle3Uk
0qNkmNLBu9KJl6WSnZORRhBugfvd8CuIlywzzvAdM4QY/9X3MN3Tv+rTFtQM/up1cZs8CbQ2hXWA
cGgV4M/wdaujg7P0Ee9+Q7Aws1cTx39XsmqviHQxXkjnDtiM1Ps7RqKIIgNWRZsRqh0dRJgQr0Nc
Jh0hsNZYNfdTolJN9WIYkj3IXR6m5g62rJ0sLwDrJ/kAALv9Q1moMsnWXfSnBmt2SjCNLB4qlA6j
dAJmxX01dHRgWlr1FrIgSCGZZUH6YLoXBMRzUEw8p5ZMhOxQiJQSb31vCP0wlR1B6/bo35tnWqtB
zyTefZt6275TOq9VqfIZOg7gTnXZV77OMwjA02YcY6ZEBCXdz4tcCq7MiZ4Yjzj3IMQc/6KnbsWn
iIvFRMmGJB896V1mBXcPALRRmOfS9It9Vkb1TgOIYgtumUt/owEf2RL88yw3r70BAjS1yIoPFv/o
8wFoIj7IE1jGCvk4fozwprbNIyC6G0vGQ3+pXComNTe+C418E7uq/InL54ALZAvtROUMFOBbwaRS
Q5Ecej3Y4uc4b8JFWfefUhMP4/KcJ2ac48LmedgO09JVUKsSnNfq5guWOfUYNXxxW5Qm4IjP96AY
mDiRcdbkFLrgK04QVjs3uFLEmcGprS8BYwxiUpZQ4yI88dBe41i/OiwqgnZoqWvunbMOcplaX+jX
OP2zX7mXoHAGgoluYWixjG8oaYMX6WLqT8W7VWlIF2akkhcgkTdWUbOeir3MRn2/GGpxe2JutlHX
JjnvkkoCqgP+E2PrEZdht8eWRlYgEVZ5eXsGebbf/rKGG3uMGiocB0K3uIN9oQXfzwfjZm05Y8eW
OIoMlYEdtAM11kBpRfwEnYbN1D3Ov9+1e5sWui+GQv23qL4r4/qPd9hSxSggKAsjvahFnPw0i+7e
3KrdFQ1Ji7ojjz8BaUTOyCfORYJkviZmxi+JspN6/m15KXyPRs5fBTYh/N3hyMU9v8JK/w/wQErS
apqHLw4DaP4TVsQhAgTL1C6l0VR5ENXrQDSkHY47hqjKJAGkQqog/UXwd4UObqiK80BerhnR5xta
oH80lsJe6gGnLTtcUHUh6MqnBGqGsjHhb0meHItBLwDa3GAAQNtfpz3LT7FOT9XnMz34g05mD266
N/iQIVYUzVyBNdiCz3zvJtc+7nJ4SI5YmclL9nIekNFHGEPqi8j3d+tr4ZBuE8CzzazHpSghBm9f
/Z6tXLFqrJ0gQHoIkLmLAhT+oKo+Tdcg26zQVyjn07PYqhPRPSZhD05EU2ogknHwtjiHEySYwAN6
hv8gTb4SyXoRZ08D3m8MPt58kbE/rcAhP+A8j+DSmG8xAVo1eSOZz8NR0HC+f6MjzIt498Hqnzjr
/tcUULE9LN7wtFSV7xiAb2fqGDFQdV0W/4TCnE1gtGewTZDYPqkyrJfDdb4CwUGmTK4KKRKYvNlh
HQOyJsNEzVsEHT2qs4ZP0FVF3dWLBZWXMIsSLKWLuESXnaq8iQKko2+732P+PYk8SXFy04qfPSOS
xM5/cv/rBcl8K3YjVjSsfl/TNsyHBeTDNq4l9DQm7KsJsLfw3Z429vyj6NKfnXe91IGZ/+E42ySQ
4QOaVq5E4KFemBNqCUGl0ybxjaGxaNBSJHbPm2hArdSZsAFYg6auRbmKWvWqvshUfDsLU6TjXXJ6
3j4g7lW8YFSnQjlNpMZFPoTWi5Yo1+s9eCqKayBpsoKYh9BkfkJQh7695SY6CcOFY7cOHhxQ8D8A
OjOzYRdw6sBh1FtizCHQF9XjyndC9PK/A9aoQUMOqI1DfIdE5Fb2tMLOTKQ+YFVJ/V171WvjbPSo
LkhUJN93lCChypIu4nk9U9oWYF3Br4+q7aHivC8LR27RPhMfi+FK0HPnHf0WiapHM4shw5m4GQNJ
YsAGTWlCAjb/Lpd76SDNJj8/jq2DnHQK2i+BiKAhQ3ByGQt9bkyXapzij7JWYSR6StSb3VWdjV5/
5Uud7zOpO+nIU5i+S77zA50rnJbughVEgyrVveAZdIkjdnf3SsJ3Yz2UmWwxnk2NzLktTfgQYBiI
7q6o00amvBvAVt7Hu37RfEQinFIvzNr7uJtb6uO0AvX5JgN5vCdvXEAqGZBX2djfXkTAVwXxC1Lo
Ehxm2Gd9aRMrD450aHqZ601TsoWziPGYM/VxGaCDXbP4//L8ls3x1fGTJ5Fg4yZ4R4OqPuKjtZYB
NBJNB1/sea/4koZE0dbc0/dx3Q7Rlw/yberk4PjQJKXTmKU8qJSxT9r5uckJMH742AZI9kvNVKtR
8Y/oMAr4TqUSMT52Sa+IZARMp63sF6Or998y3Iu7HaMJuDptcLYG88c5bM2vVakw/rE4YkaySx2p
8kSKuQaseITPWisYFik464IqXqfFlevu37J7QaT7C8D8EEPGm86OY3gh79ViOXOel3tA+FtTBTSR
mORJnioaNqrAlmTnTHC1EBrh3rsbkW0vRLq5IVzU6bDz1GvHWKmZkVU+RNtKmdYtLrTFrB9Vm2J+
xwZXxtCNBdqqXcx6nAFlxgnuZhRjdm2qItlyH524tVqR4xnZXt0dleK+f/UoKhU8Kjsq5i5WjqsU
vmEgtiDUdmuTXMeUsoQ3dcf7CpzddR3WYGF7DmBznQq39VubQRhOGFL92QXaD59gIgG3wygEyE/P
JywFhYsgkNeWsTp68EPWhg6hLGp1F7mFscsMMAXWQzMTD+km8FqWehlWurU9jGSGFQNWzN3Ctb3s
FxgxyAXB4MaQxAnIi8+sW4DmeP/OvJKiRupt05d/hauiKwsT2mh5zuMb6ckrQ0N0/OzBiZ9bxJPM
SVFVhzCLuW4zrzzooi9ez6vyMAa+fvC6FiOvCVmB/0oN7glqg/6P+Prke93s68HZ3GT4OPBRiKbQ
+72Y8aPy1Wr8xArG/4eJUmHmToCrqqqM2ir4OcbYquXGLKE+k0ECgyoXlHmJRU1ocs9cNKwfbrPu
aLH97IYUS0k5TVJt/eRpMdb8kYMmUVm7N/yCQFA5IR9Q/Wbs5riOIs6sUDI/ZZl2fD1ixIByC3uP
ICBu0JdHz4HFQ3p9ID9i4x/7Gj4sWZH8D0NK6d3/QEH3L4HPC8R5JGE6M+l5UuVUVaOoIaudW860
SPOMNIJpvNt+ej//nt4rX+2xYOnNcFFa8udW2pacQAGpkZOLCgUUfWPLkwNJVIZb9jEEED60fnII
2oJ3U2dKOiyU/gI5SVMALwMRJUc9nfQYpRFk9aXrcnv4PIjFGUtQVUGoUObkQboNZiLFql3N2MFu
6Ci2ShwOedoBPjkhTaqZZsPFRUYRA/oxabeVHdpHLBKMANAdQDFyR2uaF2bfj/PM6oYtOacljdQd
n5akOKG69yvvMAO1k+l4bcZnXiCt4G6SvoMss1GbD+Txy1enOWdMgaFkwssUqTdB3zStS+76PaNT
t/K6wKAK5gZTyAalYW5wSorNjifC5xdwQqm5NOHEX42WjUO9KTLvUAFzbdwZbrw2tzC1aqQsekcj
yiU82zE0+7qYBFOR9GS4YoPMZ0rcWHM+ZzDEkX1D8bHqxzuTJjB3/ws4MTX602wmZkG5Eo/Ze0NB
Le5JCN+zW5MK7UJ/u8XMl9mn3CrHIPFZq2Hi+nWlE3Cx3RlPJsyQ9jj/tCCgioqrfF187c0/+3L+
rf6Y/5rzGp38CuBoXFYOT34NRscpAelb8mFl0+B5DdzU6Nq2LVStdvartGiFTab/mH8nDuXQIbSA
WfO/m5i6kcgffuVUHqXu1RGMQ7cSZ5C4g4b/wPT7hvqevQDuNP6OKEwH+mNwFmt5Nd9ljrf4ShAx
3FUR+3f+g4o15BaNBdexi1p/jb+L5hIkp3UQFe7DFzbdr1Z+ALDOefzZEWwV5gM84xQ1WcSD9j8I
eEXWgYGywmgmtPWrQ9gHVUr3TFuY2NhcxeTIXfiamqdRXP/l106Ei+4FWpg6CyydwLvn67a+usPz
mdpsjzUXmhLWX+I/HfJfc/vToOOZFcs5w/1SitTmIBwzGYKsZN6jH3gE+89/hkRK0PzO3p6TekUd
L7noIpVzsDr4xVI0fGqxbcgc6R4WbzbB8LRMz1451fpqDOIsBJiQId0Rjxqt4+7aHeTohDm3H/4i
KSku0aEep+imgYgc4VIgwIq0Tz2lwAMvtTBeHXH4vEqDjljW2xRKlUZIRd3F6WINvfgNPlyRvwoG
pKPIKZR/C/uydoGKMUyTBX1EB4G1KWgxugXuXcCNrU0AQcPyFOrj8JIfhOTTa+BcARMrFEQr6jX2
2APju5NHGVlVdTfSNQwOK1e/rSPk8U6KhHdpnedPE/L9rnjpWL1heeYpH5Ii0wyLO9P6cjcEvSRW
VsAg7MC5UxWXkahU6Qgdk0PjrchtK61y2TCRa8+uGSKVm/qZjpv0fMjrlsFwdVmBH8tTkqhhYlpj
Ny0sO3Axz02hZQS7ofrt1nGzGQByqZFOPeIwYgk58SGiCbzRPuxktmTRdd/WeB1kGviEpvsrDeaB
BLEAOXO/z1LW+4S0+QWMcKVATmnWLMdhPzLX4d218EsFXC6dftS2TCmXY4De31kJX4RlYIF8mJHQ
wZnBY2YN/Kte97PNRzgHhBQE+h6P+tvaH+oElO73z6sg/FW22RnTFgimUEVIzy49kB8RL08y5jVp
3u3oU3dHx0SE8Kn2n2oR0uF8DObNz3oarjYtP5gRbViGKD0jseMujZump5RkjRnkuWuBMKMC4z7U
+++NZqSIbhmYy5ULTaZ4GofR31KrWdQDgcCDvKcYE5kY2RvIPhale86AB8VA+r7MraWBZ85aYh1H
v/+Y4H5/EYJI8/7NWw5dq2TZzTc/55Jz95P0pw8QF6evZZFEdPeEklsjszkyhd9CZ/WUnHblA/KX
yY1r2Q7b2Xn3tI0Wh9l2wlIzI9UP9zsd8HLTunIJ7Zk/6olHeETlxQYmykYhTetlpvGV3+GTsbzO
ySxdEIpfSwjCzTAphtgDjW+vCnMmGzOXvsn8JeJMNQgK8olRaDSpuffUk6e2rxlqOu0T1a+pBx/z
YqQ9wQCqAXpaSNrw8xOMvQedDo5UMYuJEzLqAGWQ/fQd8hV5IBoOfgK+f1d+77lGjkSWf6tJe/7+
wJwQMxmm1eyEvl2cZTHMHLfTwEmf2s4CVY8h9ApGKYsnaPQNo7w7ueGz8viIi68taf5df77WAwbH
xA5eqpocojt4l95H/JrLMPS9pFe8LySlcNyUJJu/fyiCZtJq3GhdRa8tJem6GjZ+v01O8LQ42IPm
byXZRgZ7WXqN+YCRAp208RrC2/MBsBh2n7Qx0jIQ+wqk/omqFmeJj1EV84n4ehMRMn3OmUDZcyse
G5YAAp3H2m17jhfEaP2JBk6a7PX77iphNT1+etnXch46Ec5a6snBKntqPCeWTL8qcKEp5T0e+Yfp
PfzW8LVY3zT5dCuFunETWTzudeIBu49XOxZu5ZJMNGbME3LwbVx6+BtRVHVlNUQi3buI0pg5+j36
y6RiF3qTGawyHJQOoJk7vU9j/TbWpHGYNty2fhCDO+xKqw9IvBi7ZRN9xNI4SwVu1OV3u8qvTEP9
AyXy3t5Wx75Qm802VAjtDgpY5krr7ifXBdHldRrl2kHKPxjdqsJqkSLRnX56OY4bJOsJyI6TC4G3
tfyP5TklHqKGWmSN5qshpUbz0knq1l15v24zKh1c/8yOvrTdcgVtAGkQTQ5OtXYkDJZknFbFOCPj
mRDq6fJNodX80NnMoYpzNaz9vgBnBH0MiuzXtnrgSLiznjNGPC8D2yEVvDLVBnqMLKKrYsHLDMXn
ElP2tzjmmd0slkX3BDbfffC8trFGkxPmjK+fTXJRQrUd1hZGb+U0hS/1HnCLCXSNDVkQTTAaUOim
3LuIFJC1B781T/5tI0qGrfzuzxAQZlz3WeNO4F54kwbFIcIuTfnKgoyRRIi3lkHiYT0JE8yjxW5I
L0sChA3BVxBh/8QeP2+qGdSGsW1SArCdZRh4H+BEBADlDt67oKXVAkNSpqH6JNltHztR6dQxDY3m
SRjYVk9jzWAdhEcSPijpUlc3VuCqdI/O5re4f9G8++ZW0xxSRJmsXiBP9H18H4jyGg7ypm2xlT91
VLxhjxOyNkZ7a8OuE82xwJlZf2EudvDHZEzp2lTbVsEVbhksRdqTJCchSrFA/TD8wT5EkL4vQ7/d
shmtMtEdNz9Lxvza5mUXW3AL0q1etx0bbIYjLHAk9lgek2Ic5O6DwolG5/ZQ6B5UY83b4swJKfZz
Ak2Q+avcEgk0vXDGlKb00V3dN5CiCnEgL/TWYRulWP1X/4VYDuR1LnFI/a5rywjUJj+JJOPalFfQ
W8UQZqFnrrgyids1PRGVSFZOmwUC2KRXE8RFyJqfGuNJGuxL922K78xqdH/TQ8CXytfPgsuzdPFX
9GAarTFKS0oe7WMEo2o+RdoFABnqg7cxHV9wJKmyhr/xf1WEa0nFGYbpvI58c2vtBc9gY3vtyDx5
q4bGstlLO12wcf9xoX+4XJWmclqGk94IQgOI2EEXH+jfTO0brMvPvdtxs+eUbO2Pc3TK7UunJStA
xeMd8yj5/sZOweChGiYYVoPsYEVEYGFeL/dszCzT3CERSDifEJra+R9gZqb1EfJDsdeXybu2s8AX
0OeTXT76bMkNBLNL7KR/Yu4K8aS4+MKzVk79M1QrFa7Wop6sXIRpEgtEqJKLZCdiWntcH1T3iRVD
G4jN5KFXXYOViJMbFBwKu+4J7i1sKnXT7A9sECDFBGqc+/o5ftZRefKzXvCW7J+d+6VM1CEfPyTR
BHkr05o2qi0dYPCm/TZ2A4rOak92QAVUilXzO/x2bOEij7DabC4FX/GK3V4vw0UGuaMm//N09PGd
mCZkf2mJ0u/Ai43ZNgbSSkHrS1vJfJQ5zg0M56gyiZVT/pCo/ZyMX36qJjuISWlRD1oIyJtO1Nj0
XnGByAqg4BLNxWJA2dPDR66lKaGgDksFvwHTijhDGFDlES0SbFLnTblHzOpXB0wgPhreSEX075/1
Sj5fHbXrsODkcy4h9mwqM/sMGZD2T6+VDdT4tpPxgx1dO1kCtzVDRki0/qZ3Zah3ZsRuRRFuor4h
kgC6jCwaexcAxNM9AYHbeohmNtCq9qvg+iH/DBbHW6V5RCLXynThnlB13RuR/B5Tru1LwI3775gB
lrVX4Mvg30aXFfBGd+YnYdnYH+WaIaT3Dl9WZoXwAYof0q885nqU5v9bxqmjDFqI41zk50jyvHEN
zMGJcqzrZu6TuIQSIIxgGQ375KQ7eG7ULBMeV6pHFFpIKR3AO6W8MHHxjbpKRdDngrhwKIPdbA0m
yxYy/CkvLVsZYsB6Wwt+dnMWqZQmlqXko3VryWyG2Th148TfXlTmdfsfl1i2Cpvd+GhY20x1LwwQ
pUJB+IwMjFGZiZvT9MxKE6tzW2GCUtKYGOFEIersIAdtHYsVUbvJNAwMz8Dmv+vF8ttZdoxfvnwh
I1K+HR/c/ShYLcpuxKdX7pHgPWYm0yUl16Rw4SD29YCPP5wPB0ptb033Dy/Vir8IM6Dquy+G5yWD
66JiCiB4PsFZL4L6BIFdV7nfZ/JBbA8NaEzRrGAH2Mc/3agexlSO+l98I2h0IFr3zQpHbf9AmV2G
sphUQWS/kD5P1J7eEalgBPkOSFqAO8RU1QjiUNEEBTFLnxV05OlXxRVl/ienUO/WWhAJHkh4g8yM
SwCEKgQNJKT8vfadMguRdRu0LL5cCvsOIGh1nk5xKe/yVV9MO5NYSWte5WRE8ZSoCpreoBei4Nr7
T1BUKzhnRhzY9wNLbljGdIc4JmgcD3VzcoCP4a8uQ3Q2jyUT1rNWvX7rxKlC5kF59gs06g958KNN
8MuYhEnWFj1FgwMOqMnaxwh8RaZ1INKCoJ6wRDbPF0MjxRx40YkMbkYbaGXy9POBnRwG9sJKd7hB
hfgOSk/jFvqCr7zwxLD51cN0AXWT+xgcOAPHDPjE+Rh2q536HckIKzO3GGhuois4j1zprIaA/lDR
TsEHKKaQsfUO2la6AWIGoizV9tPNCUEXCxt8PUIKXyJ1vAj15capKdAEPG0ReU96RdRydpu1X5HN
24Emvyds19VMNiN34J7diXGJlcArD/e7jq+oScXxIcXkhDuVY3GRL44n6z8rURkdVU6U+3J4V5XN
b+IfvOyHuVmyO1pmfaxczYrskvTgZ2qr85UxysCZcMIojN2OzErVJ7UCjO7PD+kWWHaIyGmlcuH/
UmW+ZtOR91rTkJBtztovWu8f5X2xmlfuxcOja9chW60SctdwUkFbNcQl0c8S24l/7DpkntZaa6Sr
cg3dFuQQhRW8Gq2DdP3M3dKRhrHBgid602AqBrKKFmKaZ3mETsLt9eCGPoWq8qN0QH2acOdo4JWs
jPeUhOzL6YNNy/PErPKtbNaCSjz/Tx16zyJirlVhAzKEjUTsbSNM6vWNG0yTcfl3jvPOCx0UochL
kVdWzZXligXmITpvcAxTo6n/UucOAbT1X9dzp6yeaz3fmNP3ojX/9tG1eeYL6y7JDAxXfyOnmmWp
hwM8P9rlAcS5X9sWao6bPCVgjbAiWmzQKgvGc/RZroL7xIs+wUwxpVoiczAMrqUP2lrszwSrbBmZ
H4zYIiDqG3Zqj9XX9BMpv4i6UsGYDgveL8lLE5EtoldhPPBxjt7Hsrpcb3cez7w6a+QBs57i2R7a
WpXNJ+fZjreUlvW1FSY5jfAMGeaQ+rdJU1w+mgpZhsMBddc1XkCER2NW+r1MEPSI0xbxerQLIOx/
3GCObDXSnN0DTgCYPe04X0CAWbl8fUuw6CqdaW6I44JnNof2rtPWO/rIECpso5czN8za41t0nygN
3llxzoBA8lNHPKXSJxJ0+QeHxfGqWbP4GuR9dRuqMIo3rX07lgphhbxGASR36e0Fz7D63MNq4U6K
H1gLtvDfmUlLhDZyXiJPVJHh9+1bZuC0AA85jLvNGWz5weeZiAIkE/QlLZ5xL6aTkVMkTF/sv2KO
xI5EMk1x4IolMu0TfcnQB8jnWEJ3AgW5PAtOokZE+O4XDLtaBqf+ia+KVSEMkWu80omsCF31OvbJ
5uzA0TuTHGZ0A7g3rzCNSityaolzhp9w2HOBNMvnzXqezlaOPiGhU/fjuMXKwslzoy8t1KkXiRE6
vrPMec1AKaWMW8EEFlk8oJnhg13xs2fjys2qi0Db92c73L4dvFT4BK66mrFCFCCAHJukzrUtcFGf
qD5847YwMOoeypllmJQ5gRt7wzn3xWhcyiE9cn1ik8ma1T3B4Gv28VUfdWRIx5hFRKwUhzlAovpG
HGAzKZroaf50mORX5oS6LwI1kvPPZ3i/Mrbp7q15Nw6X9bdrZZkzzDq6yJi03GjmrglPPNGvTe27
d1U92tg/9O2tkmIhBV4y0Yag4ikGJQySiLIXYLi3K9BXIjYJUtGWfYiV2JDrwi/3sembPCoGbXTL
6gpmfdCSbhV9DCKeUMhOPnQVJpvXi3H9U9mw4GVsbTZkA8s0G9T8CFYQ8mi9prHWDDULr+kGl7ms
liHLFz4cC6czXND2vw1bSbhqn5HMHECgrtcl0FcQOtqu3Gn6UsPnZjj6L5EVMiIs/n7nzVhShRqv
Fk1FwttwcoVhXwulS2VLcUtDqNaU3S5wgi68W9fh+oXTLL9v+v3SmUdQ/RS87gvDbcrkfFxe4178
UIXxuaahTo13bvtydycWG4YjqnRcJCaHdWEiqpvCnLYzrhWPMu1bdPPa+mhJssPtJxFTYz0wVBEm
rQPybkRoNAvoW/UyjpVmwVgNbXfkl8LJJDrMf0wyIxyxQ05GO/rb6ajeYjmWmzVeizQ0xgOX6xAz
RITrZggvI3Q/Ht7NXQZjdlVvIUrORQBByM+DFwiYmI+ioFq97ypMp0WM+S1/lPJBsMM14oPRhila
G9HdrDXZgNaOB1nChc5BnRtA+cWCmD8zSffzC73Zd8TqoxNgVg/ZXLeadVxtWhMb5oQSB7/IVov7
Is+xFo23+S/dgNRzQpcezL7VeCLtdK/e69l3bKIPkJb2jbnZmGQtthtiYZzxNvi0kMvI3LmqMZN1
gZq2jeYjgapSAMovv38n2JVYREOHoK4DdoUuQdZBHRsuicl1rGrN5ldfLD4SAl/5M/ORRYqjGJbM
v4EfObqNWVowot50492qLnG+JO9PM6fqv8p5LP/d/bPeuWBfoBrNScpOJcul4fxx4VixOsXB7r4b
6CsLuzdfNJZJmWLuB9JjBPz+Dmf6iEJl+soc68wJvNraKEDzZtwoxBqMjmusJykNDe799Ht4n2QK
90vVdcEMESybvavMombx4ZHbKuqXMLkX0GXtdH5/fDvnn6XJgseTtIxZicp9rQFIpF5hATpoFBbY
BCCTHOL+5gge8mt2YbpzK2ePUGvZ0Uei2vuhgGCvJ8u2yuPlZn2xFhMcc+6D5PPjFkJRTWoruCoL
tRFrFmlsS7xeAuGlHxbghrJEclXIFXAQnLTj0zbZNxkSi1eWU4BFVfv9tVd7x+5cnvV9SR2Dx2Wy
dsW+v8bOpNX1EPoP32ZfT9twBfmujT2jZvj3cHkEKLnjojCWy1VTeeGJAJRe4d0b+nmeTsckTayR
EOfgVKKdliWfDHdXhI/IFP3OkdklPYH0ZvzBuEvHU2hVcUyiMTVxjiffZFclrJfdS2wmx7HCQuFg
NRy6/opUWp5WPRHh947NCM43Ln6S5cZtlszLVBc5Y2n1NAfMhG3bnpq6zPs0ieNX8OMuPNtUzTZE
hkqAQNGVtmptDw53HPJs8iGt528EdyC9U2FFlIrwfItq1ERPxExBdqxYD4uQa/ublZVoDMEEseOX
Qzw3Y2FTb3KI/JegzzbJxDGT9KrTZuPfurhAosIN8QVkzBHYe60Vm6c9cLwR5BCUXCx/JbtT5JPd
DpSZUUzHDVDie5572rP+COlPqjExDJqxPxHteEtEGq/fYFRh666BX6UfJE1LUljr6juVHUW+Gf5Q
bEGr98Jft67oswmrMH088fsLLjLab2YlYLSC5ob9ZvHP1buEliVDKskN1SmZ8CB+RFHWjAX7p7Tg
PXsmT2p+WXG3/RBN8mB+/8a59Xf+7/kjo9fDiVkGgLXBM8szow0TyTmXZxa3ch9T7FV6S3aTS0D3
1AMeQpBkDY12BWubbEdrO5F0gxImn7CIGaGGzph+f+favMaxY1Jm4eApf2rqxkiI4cVvu8JnxywW
9PlFk+kBgTUjaIkVqTOGxjf3h/HY3loxk1Qc86UwnAZfJr5QG9oVsG2ZKo8GUI+kHlVC7gFGKDP5
tS1a0b+W7Jukgn4awWAZUvplg5X+Aw1eScS7nIjwarNedcUQmkIyzvupUEI+V+4LgjQ7S2/78ciT
FdMG5S5OGOTwGfRnbcTGk2F61NNeIC+hFdQwY4QqS447G83cQU14byNTn0aqX8/pCTLndIbU0iYm
ZgGC/q7MhHuwlpBPecqOron2GtJwmEEhY4cW/tPjhwlDrspI767JN5LGvXp/MMLt/yLnl23htSVW
Q0Lds96BswY2pvQbq5qbygRZ5ukP9VnFRud6zLSDkVwbXTmTxz6l2BF57PIdZFsiExTOYdPYEstD
wSCPdfDVnDHYdc/apy4N0/KQjOnhsYHdJeY4/dJ0Gm5ZbNxO3M01VLva67RPBMLRli6XhsAIlgtd
Hd+lNivfVjqONAooy9DQTTHCrVlzPBAv6/2gy/EgXPaim4R3bVt+9LRxN5+dvBAaDFRfbE5PPvYK
9evOCPG7dnEGRDDc4epKDfaCvklulDadOYDbw99oVMbC9KpVGTb8SMiQirQIhq9off7W9er6XUpq
DU/fVlqqnXvu6HF0C18zCoUn3x9zLJQ2Uz8Y2EwNLpZRXJQtXhcs8u0MOahbFVsrzPHcbcazFCME
2Ew/71Ns1E6tH5h/ezqk1sW3xU4xVJ5PgQ+KYxx6swOaJPMqOG7Ro0ZMIBKSNtjDtyyS4bY3PS6j
IbOeRaiDdSPoTUQbZGy+cSZKeUYziQVajzpqR0xREj8NYIcyvuyUVvuKbPs9zs0DQ7RS3Ppxxej3
PwrysycdN636brEUFlexBJskvkc1dl/TxKmCDHYIj03JqynQEwXz4iajUU+77GEQtYt8h4gaUl+d
6wKC9R50d0ywYNeRG7Mrw0K1Ycw46bC2fx0FlO7wuL04ox0yk/d9RIz9f0uWLwb48Xs3d67eqr7r
Do6lg4nU0vI3sqQXyg98HiX3jzeF7Xx6/EhCy5JAc+XGUyczKlelQu44Tvxk9YxwgfV0CsP6JsvF
uLEugDl5W4PtQ5gGTgw5xFsieePwVBTutmPpP7XiSRaueGVlz87/VuvWD+DrKY2Ed7auK9Cvbf6P
cayPUWd4CoVHt10VR3/3UQUXAwIviI043ZJcEj7MScHSmXyoKwrPrkZ5Gk6Z5wweAeT8pf9JYiGI
6Hng38f/TFJvXoCdHEeEJPkjXFn/urqRu49XYqP+B0XSrrlgxypN22pShD9qk03xRCppyWuvPlMN
TI2I5zqt39XyRG4Yiz6BzNLa7tUWW0TFhxYWl+jOHRQptRvML4WVOAAVZP9A64vopCQE6IU33EX4
ELYqLl5Rj17LANQXrmjvLFmJiq9TcnabO8KdFtzPZlCiFvItPRUspBvzrKVFHZysXy5yseVKZ1hl
EDKC2p4YQgMu5vnub9DrpyjcVwrnKNB3JXdL72zycMKxAMzB+d3s1b7/GemdV3lAVrZa+abNJj94
E5YxojMcmrwXZOYDJRyaUcjDnrb65brw3m4cYTn9TgRC5FuBnNXHVbRoLMZHX07AAzQh//qQIr2o
ym4+ceZLAaMHbry6o9A5568Kn6up0snlKK/8o40KKQmdIDvmOzf/zq4Ip8cRYz3uiT6PW/Uvz4CU
lBBwXDVrcU/RoCGpCfePfkbbkcf/h/zIxHGTWQu5Wj6Iyshee9I8UCNzFwu/oJjpuGRD4r4iqTwW
/bA6euVWovH9WcfpNiKjTN6NUa0kMgvMGzkOta0fFteZLXrrr5oy9Cnu6XTlp8UBlQ0F3rTBmKjw
JJ/kKJsEbAYffn7mVtcSM/+Vzmho8Or89KMf0AHdxLb//xE//gaPSAL6JkPIQzk9FPL34+txexGj
vAFM/3N4XMs/eWxkjTQKux3IW+E7vZSdqd97FW4EUBhZe4KU4TsImAj31VyWLhLQO9eZ+QOZZ9s3
oNyiz5cNwmDSTf+NMcjyJl68IieOhWjBboVLwG5fhYekfTWlkR5T90FlYQl8+xOKtPWIrcxZ/J2s
/hkCOLSl/VSCio10AFHsXyPUXvQrDOZhn3Vk9tiwXKSxZbKGd02/3VWZD9gpa6FNrqQr4DwCNQk1
Ur6STIMF4U2yoLqB5qnEQSKnIfjowUKQXz1+PDk3xJ+3KS6Yl6r6AiKXss1tairBwepOkQ48gDeD
DcP01EAk1xlHXJsdzHlB7RZoQOf3ryzOh4mWTjOmnGEbZp/rijJkl5x1YanGNIYxMNPVqNtudlT/
WWgqbT7tdS6r4XMHvqu3muhtWpPsBX/CBwK/39Kw9MFrH4m4+P1eOpqzDpGjxCpZJ4Llb2m/C0WJ
yYP/nHKMAxxqHr/yvG2Z8NuKTySwWCi0r6DJ3ZAiq6SFTsfQwKw8Em57l3qb+Qw0EM/P8AGBauNX
E9sLTg4WTQtbTJsmAeRqn+lDVemLje8zWzlPD8rKrft46+SWLA6rbdfGGgxgFyCdCTS2MqEW10bX
+hqLXeqcegaj4dJfg13cqoygmWzb8xDjSLRgd6xnmOvqTuiIjPl7EEyhXEWC5U8OZvanf7r6MrnU
xAQLqeQQ48MPwMb1CYHfmIGbD3qn7Q78N5XmWZmL3EaWAOsaXvldLrkBCcSmZh2rrhz1tuxOCS9b
OrPp+b83OiaCzLI0xzVEt5AmL8D2EjmvgmCaCnQJ8mrZfVAs6foPCWsORyc9kTkG0UaXbn6SNE9R
m9VRXbfe43ln/DvLUCgdCEN/7G99VCFpVtrIpdShkY9USmUnLWn8FRYnqT/ODCGIIyAzAF9wV35+
UX1v9PlPYSOWfJt33LbJOQv7hO8agmkIw8JxS7zG6rkx1m3zYJVk7MtLL9cUucXhv/9WMHNAB+KT
gUIQrnMtEpzAhNDOw1cyLXXo59yOTM1hIt9FwuOCZy5zb0TDkeB+0HGeUsq5Fk11NtqJwJFzEaK9
l6TKJ8gGdn8HKYQhSGryeihqnsRvKtAufaZmcOw/ZdPV0G0tETggDd4odySwimwcgdUQ17RAr7Yx
LJqe7hgr2Q2v8j6LljVMp2bdOOakazse1gO42tsQk1lQovHfRENKTCmkIJlwauqLEYeg1hhSZ1HZ
JmMl4rYGIVMvuiSlTikE//nBEJqipVsJoZ4Mu0I2iVpHCp6DMDrDV9pSeX+xsFSM0gN6mFXKa0Cq
thgMheyKNZA6TrPkD0K6B+/8p9nXhFwgacwJn5jI9q5yshvGTtAOawAPtQslqdtxsqlPFMgT0agn
NCAuHNwSNn+fUZvVcSTTJvZY9WmgF1n5bfRI64hEuRt+vsUDUQIUmDwsXQe71S/37md+RQXKpQSK
uW58Iijm27dofFYVTxUQwmhopOQvxkJHunjSe+edz/KAlVDi7cmrTlTp2U+lR6uytPVXovZuI8Lh
6YiIWwQhDQk++b4LpSpgoInZvgLG7zZ8cF3qCdmFe8d41NSuAu97i5gz+0N+TDVumTCENF9ide4d
S3R8OkG4p5Bq2zVvpOtfPDgFLc5jSESgYEy2qFjSVbwznKPXy45rV0NIq+sHfnDuq/joXeAUPp1e
rGOuPtb0PT36fTdbHzvMYhYK+NGO1Rgyk2r7wE8NKviiS31CL+Z1tiTkQdMR3k0J+7f3ieSYeW9A
cGTL87rGmVrYepN/3uOI4vRhR9biEaT67VadPDb3RngOfz0tHA3vL/1pqJJ/jIpzNAd3gbukNoD9
VUtsx0tf7s1Zj6OKakY9Vf3QKJ0E23gc/Oq/uGRBPDfJzhpl33Rev76Fg/gsPg/2ebtGVXEi5fkO
dWNceRguSBhcIElVcsthYsDoNHXVx86oWgSDfQIokLCpOKaWtb3xmrN765kcKC0D6aSqk35zniIo
sEM/iRv93OQyeaz6zu1mhAx6/x+tcMuMt1Wwui2ialI8whVj+bjyYtKSQ6p3J42hqEWNawe5mAib
dRlNqLH8/tpOg7qhuhQxAA61ZBhOKlvRWNU3H76WMNWEsSEuBguJ06kLrO+dkSU0nog/HP8YDm/W
odQ/zoLPuTJXcgPDQ9adfo2K6kS7wkcS8r43BNzkonBwbDbOmZDHF4VBV44XzcGtex0z2xsY/ZZ5
D+92Z+3qwGRRrNwqjQIr+oXjzfVozwlT3E9sWlPeRzZV1WhlyhvqLVnqZVOYG8jSXvMh2ZB8p81G
pgrZcELh/uN9H3FLlbDiv9JJDktg3nybnLSTQVmUpK4VB6Nxz1ksnxZC3UhJWLyEnTY0NLQ0Z2cg
tOUAte4u9q/9vctFJddftsnrl4fu24KxGFlua6AmUAV/TRLv8hiunSzMLMUjZ3snpVFyxLBPi0gm
KxZA6tj4Rj5NlI9PZNo5OqZVsHVgGyBNhQVFz16AlIBn+atf02ygEnbFzSMETyDzTkokktAQ754a
BGAbFgqQEmDE16fdQVABIqHuv6fViXEDfu7lWLK2FvPxMnnXGEOWpdS+PibAToZCT5i0Ob0sgggv
4jYiYqbvhJYasrHvjOUPlBA1xOH/xk9MvmRc8ZXa1syNetjRjGSvBzGpYw99cYEndxqaWR6PNvtf
tsp2QOQ/SJTzd6lKMIUipJXN/BsYf1/vv53KkEP5OKlojA1/47O1lev3wV8NEIvuIB6e77dAVPsE
UeMJ8NBiCE/nzTXl0BPBqK/1U6nvF/cbgT38xfSv6SXn8JcbrF1s9MGHSphR4v1vr1Odhu7sBYlX
ktIrmUig7R+tnSKkgnwui9FclBqhdJvjvrgKOvCHIOQN6myKJpglLi6MiGfPmQ1SZbUDJ49Il57Y
BT7p0N6sdBHtSiy9M3Zvi5drNvJkWU7VrXw3+ZWJD9MoB+tDY9CwlfowoCcZWY4+j3J8jxmdiOrd
kSCFTaaiiSr+GdOnh10eVFryKscUY2yaDqVBrMDlqQXCx9RWzFQnsmJOURfD64R26akF8kexw8At
4yU0dVkIgEFq906u6KHvV2xdtO608ResA5P0LkojIHog8ZZYxCOeMCsO5FH2ZFEeEsqtyXgGVxrK
I80DtW2erzrksQc2yHhCiDuO5CRQ4WwZomOGEiDNn1V6gDuWr9gu5YnQabY3Vwi/6EaOJz6X3boJ
MXNeyJKLfflzHjzUN9bVvPBa7ljQ9Azq6Jvq3iTZbeqkhOk1AbR2hgWuMyz3aAm8IDThUKCJg3+2
J4rCzKWJIL3hpnNe/ufk8QJxke1VfSo9sxUtJ+m/6FcsoPtwsweRmJryTf8BHTje0P9GvvcUGCrk
SWut4ymubWWRj99WCZXTmRRYcNHbdZ2MoRjxemLwRvZKqYupSA0PiKkbGKoPXOidXNfTPEkEbMNx
uBGzKz3XQozKQZw9hord3IDnXj18YTxdQARLZEFVbIK5mtNPKSwrOlIXKr7XIvwEs6/sirbMKkV/
13+EArXGDgRQmUmJs+l++3uZavv3XZo3pQ0CTV3C7F6r883+fIvUTAGbSQBcgzR5HFdTejzDDO0x
6Oj3rx6fUO7Vp7+u+i0RXUnGLJVNe0gigfg4t2JaUJ6Rd3QDQ/JyFJ5bHPEYefOU1qslrfVYknN6
l6felVmmwkbJCBmN6LcLNsCT9F3vfauOdJHBQaJp/iyqFn9dn/YYU6DDZ53Suv8SV61a1gk2Wh75
MqGoKApTKXEiDPfnmkDcAmbGtuf00T2YiBwTfBhQPPcN++Ld70wEVygNN+fX76Z1M1dpdwNb/+lj
T8ik2T/Ki01mJXd0qssB3od/Yk/NdjYdYIPMszqSuvGP/hBJGAlBvH1AERZaYN9ANr6bpqGxTslQ
BLyw8dtUZEa3Hnkl705Sn2hbe1HF5DCOdz7I26wholFOIJJ24zdmbR/8Tfj4HaDf6gocQh2Tn7vV
m8bN4aycnmggalHYx0UHTxA74b3HmPDDWxUE8IaJQAy71XOeCKelqT0NdD4IRJldAzkLGbQ7PW8h
LKhLY/uDUJmtF+Sg8O7AgHXqfDqplQzzfHfyaIdNR8wGlgerV/yO2smGZhFNhXJ76qSN0/6+XydD
4YRu0VBvaV0FQHC0AmMtcwsU7cHOl5966sp7KhfidQ6Gfmog93W/T85HNQN9RJmuHMrAJhDguWuT
iq74gukWTY9cMgcl9+6jXZ8MmwK56IoJRNP+0y8aSAWZmqKemyCu0Nepmp7VLJPEAZyFykbw1M1e
vd3ZerftwpuvM1sfx1tbYVjj2gDDNKhyipY89O8sR9c3dfYgZ8MtbLmJD6SBjZIuxtmlonZDtE5u
31x9wury4TrmZ1t2W1n8P0BALMPhLgPbJGyA6ir10CM6DTONJ8vSyJEmEK8kPP8qZ1o7iR2PYvdP
ZIVphYbV3sLkZVgwhTSUXw7ImMAaDGMyB40H+WXxVm/Gt4+5HFkGzdm8Lt7fGHCkTzFYB4JOByOj
fYWUkQWzJJAKxKwEUXFWE1XM/7y31l1pdi1zOMCNgpCbxlUZ8YhA9BybnVZB/eQ36q7AMUWH4VrE
YgwYloQ6pUbkBV/L111dRjB7eChcw/Zx+wf1qY3f+8LzrcLvTqF8usKGh3Y14UAHPElM076vOLPd
Z9HO0jeGEaGTv05taWP9dsU+X7JxSTp0sxuWcxP2VQzihciWtQWuo7xy3FDk/TiACv+G7Qnymr4k
4uPhRu4bq18XEVXjDc9u4YC2UwUXmi2eDjnbDFiUvkyK/Ya8pc2+5CfUHITSCfOvv3/7bqdh1XDG
LkIphIQHqEQlkyqTo6QU90EAH1FL0ObIIUCIZAc2lyjom0HzWkM8cPHlzTfKdxBxM6XdrzBkRL4q
k7Om8LyP2/zs+AGhYO6NYF79tXbW9+7BAhgNABBk8PGcdaxdx6+fzenSmUUcPcAZahB7oj8oFia5
+40oFimT+YH2f1Qr3Flj5FR0rEsymS0RR5O6pizFPlg/sq05Ty2oNseaHMUUkyEQuJaYYcWpP/9d
yJlnz+UggtLaum6poAwcz9nmy9Fw+Ao+8Pc/WtxHDKyAALSHgXemMx7MmdENlwNwtNrWuMs8jMSy
duI2UkFxLv/955l2Zq/zyw0xLvqVDycUG3aAArdNr5bnMoV0wXESArEugyUZem33YQGIQpMdL7wv
5x5gnQQIk4SoG99EnHhc2kPudnYAdyJECjsa+HbkQ8mjBkmLK9dIV3pCgeix2hp3w+sJdB1qlapR
gqR6UQIXySbodMfq+ln3V7ysWjCoFmQgQ1I11ZgA8sjnCJjV3XNfMUWQsw9FnShMkMkDD/BK69/a
QRokc7Itw7coo7LyfHbJ6SsXciJw1VqpUngk7PQGpGssow572jniaqBPVcpLscslwUAorXsKskgd
ElVz0xmLVu6rmjEX6/KJ349o4pXmsf3AxFoIZVnJDmpH+ycuPSHc7middPz5QC989mJnEWR0Ecny
wNAlZ96h39+U4Sgmn4BozYOJtasIO5ond27TZnqNFvKjsTS6D6aAsVjKd4ZzXYzwttEPfEfLNGP3
gQSMTDh7oILo5Wx9kv/QJUInoXtGOhky5vYFkOJV1H02+/bkhfYlaOjHG2R6TLA1w6lILH+rrB9M
Tz+wKiZJhyfysoUQMY5NTp0iyC/PPLlm0TiC30uSKW48in+xibN5pFXc4Z6xAzLIW2OW8KlBHaX/
75EoH480udgI/IXorZsDaPUpkomcRtDyVkGRdtTWT0e7o0cIqj28eKEcrIT1fJOaODsgjDpbbDaZ
UY88iNwSJX8ongUg0Jk75AGjJ13oh+Dvnf2CIjK8iwNL6w+8ds56iaQYfHYm5F4R4/uYrMJ5OFza
pzFVfnKONQMMc9OzSzPk7lddh5xukKsA614Xg1/PBIoAx8mp9fxf2ZKrKvSPni6am121yJFKhEj7
8LJhN8KLs+X5GOJfdkEq0o9Mh7C+7uEfvRSjiveTLW8fK7LlOhf9xXccRko6sJC9rRSizEf/KclX
xM5JU40qcJhyjD0P2MDpxNaslN7ktW+RSJzjs524MKAws2b9hhSKbQcfOX7vCkiyr86XTgXI1sOs
VcRvaTiKn7eWUMSYRZpYRgzUzEdiDdeqRSCEuQfQbrEoKVc3CzKq9NY2QMoRQb8OgywCFA/N6ReI
urucFL+DPnP7a27sBmeRxC3WUUMZx3D2TTLV1QAxJsnw8q/p8WeNllwhsHU9z0uyzWxcl9EfmJdo
qicxxyPVffVNuRGynIylv6HXvgvrfAK/3giKrudIzm2PsiiMZC4gvCKb8zhQA9HyZ7xjsXxgNE8l
tbINCjHoWBJM55AW8oYmkQpjlvJ4qNmS9IKLD2wqsMj4B6yyXhOPaCdiw3y9sFvqviEVRGhtSawa
Ivvy9nzIW83rJ93A04yvaRC1o29Hy3vvUdDMmBsZDGjrxjcKJDEXyZ7L1Djgc5qA6qsqotrQjtw7
Brv4WhCM6+kt5yG1zHUviZTwyOdD78RtXtHU39Mhx7XTS+p8EsgK0l+pdwsv2ELhv0USUnnPFkqe
4kVx0HeQHq7Ip4S483odK2MZQX5yrxwNvXg0WiU2FLuAWHfYiUWDhBJMxi4FBnFLq7j1ZKBdTif/
cakjy710RwlUwoIYgc7g2FUxA9HFiH0Q6wBxwO/HMzKbg53Zau+U/0FUuU9tFCwWeYK1jMYz7uHP
up2JKt30+pwu7oDESmeYP3t+aF2xM5VVxbZvecGTiBUtxLwDhH3v3sREGxo+NqFghCw5SdSk5Ls+
Vh3laiIk/zP25XSRP3ERMNLdc0H/HO4CDAFdmtkjc5qCvKcZXLHWu96aTEx76oy1s640Xo8sXkLJ
GP25e4njaF5J0+sczdePl7lvrYybdPVat57igEDH4jg+gLlg7BuFWp0isNydcBmPZjRk5BUdk9tw
Ww/biu+YyIl6iraA0woAxH8EKlPL8iNKBeR8ZR/QPayYBZGvNTSRGPN2UiT35ILPUWT/hl66Zj1w
sQCEv3tiqZAau2D+wn3eo+k1GZfaj2BNhXX65qjgt0Ywu0lJzd3k6yl0yn8QgxCvcoUXs5ePRNIg
PgadejYJwwfMUrL7YNeY0p+mjOj7y3b8w2/V9VOVJQ5cNfPlSTK4tSordDzlbTSLLXxi+eBdiVS7
JKL6E4g2dqaZJiPwLz07NwJvrCe/fnmkR1Wl6fIvXP2zUJ9fkoBB7MvyyE0lVNyR9qfpAxZEYSh/
Wa2OYbx/UhdBsF5VWulJHugJL7XDe+hYuDVUe74qPLYXRdge48ld9qxGfE9GKMLN2LIBHjXu3YRH
NbQ5rJDFWV1xQoQHDqObsCUVEqML/d7akFGsRIyt9TrBKGEa3yMg1WT8H7B7EuOaidsJ1SvxFC/v
uk82lcXS9gaQuUfRg4oearxdCK0EEWmWSgq2kRodr4ZcSr4GGsU9Gg4+FAr6OZB0Qpv5E/H9C6Lm
2ISwiev50V5lDYaYgm8OMZaJ4Osy1VwP1MVdufWZvKivXz3I8iy6losXDY4K4vd3U0fbPaNLrbft
rg8/N82jjbp15NbEeAF2A8xCTL127Y4uzoW2tHFPIwn1PW9i3D8A5vM/W02vSTletnA5zT3L0DL4
g/QoOL6B+dRT7mxlEwTbJDmN86J/GzKMCcApeykwRA35/DTEi9fAPDnII7smOHNETaAZd0o7IDzv
Hk5DpsoKJ2Ylm0iSKO/Sc+9lwj71MkNMEZOcyfYC8Olv4lH5n7rD0yIKs+ipgCJkEGnLE8b019VJ
1bj2pKijOJkbZ0URFXjGVA37xJZuUiZ1Va0AbKec9FzWmkoSbzmHmt9ehYA3iYs2CS90ZFNq07N6
vox6ykWMSss9IOohcY20OrTs6OmdfLTGZjshIS4JTAWJcBqJReaf0pIpwAyQdQP/ufUczTudQnOO
yaNhQ5ktXmzKgGBcal6BKb8wVV6dOqcQr/BVzEnCeZ7Y08OmiZRSnQFeQ6X0klHQ/X0zvXoGTqo8
uPLdSxD2zTYrNvcy/G0QLjUXTZRIELVdAD7J9DikNIEVz9SsUs4RbAoYneXYkecYItJGjRwfIhgI
B6RoNYmHATlzHnUtKSIYDQ4lVMsGNl1nMIiXvF/wibn2wpWKWr5dHZJkHBSEKcXAMpU9v2MIbSyW
9pCFK1AxZMtpVGQvB7sStCKX7qn5aLCWpNjayL4B0tRRaEQLM/4+6dGv8YCfs/BWHKmBvPMiPBjf
PuWz9kEdI6cNf8BTu2a4uf/RYj9m7Fao4I/vlT1wrN49Pf0Wtbs9Ym++CZyweqmyrtXKOYax+mGI
v9Mf8ANx3/2h+FY5o9HbK0YvLJKyB2Kj2ATv7gp+Fyj59Vp357QhRVXxpWtD6OxvYw848NdECJFl
nE/5qH3vgJ64khgVibYSu1lD4ELHMltioZgMms4+hCwjh/lvv3kpQ/UknsGQ7pIljjwDZZBCqFLu
/FBn/dYI1pplSmPe5KSsc1K5c28k9/vFHEGUk/G0ZfaZrIKxN+RW4NhEYDpCOauaWx/zvRmAkiW/
R1gfZbSxDGAjT/a5QmstkYWdCqsV8H6ure5fQIKQrP6DnG/mmwzEX2RAUmarMR/rr+vnTjHCfjoO
QEr1U+Z1J7O5cKUSw64YIeuw+MwbH6P8V8YslJCinqbLnL7Lv75VMEN+8ydNGZNtRUk05oN1G3y0
dUg/dOgXvZu5b6qNc8dqZjM5h4ohIwUSZxfjpkVAscIHsrA/E+K8SHGoTBCPY8go3GfaKZwfEnGz
JTZDKPrqTeq3wwEpNweBHJV/0APNh7wg29lAkL5yva+WKuko4ogzk/JFTmocuGte/jfyuHPQg0np
i29xpXXsX3Ipjun9fw+FIBAuPC8FNwbCj/dfYpgl5EPGudmiQbEXLQz0WdodA8niK8gnW1E/hE9+
ZY75RDKDis4hwX/bPwIZSqdkdpJym9w/3NqYwxXPETJjsPG+q9mH052bLlF8By+wO6bZa6Z19Bfa
s1lDcy0QO7yzlizcdej+v7GgEk7T0wDRojsue/kJXtHXtA5H6ByGo5h7vg2y6rTZMkl2B1kTw/Au
B/6bGV3la0KVvWvDbcK9Kluwo3J5bBzJa+Hb2nkXtP44sMDJToGPuRPfDJfACBYeaVQ7lYeda6Km
A2M0vSwcOTQlBd3vNX9yLwfMweXOaj/5kqOIYCWN5s1vXKq0IOcBt5HWrYezUkalpLYAqoUm9Clh
dck4eDq0ZRlrhgWj+wNEN7e00ENq/aIZYqF+3xq+rAcO2BHv7B6htGOfuPpokO/tR6tyQc1B4l/m
wCDfx1OUoF5EwxaLEXkooa9aDwqL+VhImBDixc6BfbylVzoUZLtQn3eQN3Ni+gw5qaMC1yLmfJKO
3lFpjeBH7vkXamZx4vXToVjVo8JhxWI/IqlzLIecAnE00CxEpwxE7TRT8wm7h7u5YWKciTD6lU9I
NVkTpMwduBIa9PtH3kFMGcbQWsP4oTAD+zOE7zZv1ORpfMs2SXwj89O2C95btqFHzYKmhWbwguy7
giCmvTKYkoOAG5wGjbIWkqhUObd962xAyRNpAiWC3TnprbNeML4b5IDV+70UTM9Ka+feyBo5VWFP
vQcHjgqiCLIj7NppgojB1eJZuLrikGLow1eCqPPplNtqi3bEN1qehtxsKlpH4M/6MBHYbPa60+Vb
69yBbfAnybaolmbZ66cpKTScY9MOq1EC9h82zdX1p7u/KvRnQPkaafYSIvMD983BG7rNN9N/omFT
WxkSD76ejJAapQIt0AvxsXpAMhQxeT6ACUmxnymnssmJn0wjkr6V/pKlQ2TW7IdhizuPP2yMEVIc
XoLVrD/kIBNTQCBbmNGULeLeK+ulzG08vEFv0tKNv1pA8hu+Q8RLfYzWIgiOXrPepRuRtZrGmrsU
2xVw3dkjefDZmhBtuwuWAysuaqkEr9WxkCAX/mzO1NMNAubEfeCC0piCqAiJMIMqSQr4CKR0IfEy
f0wUhnXWoJH57i0kyrjspGfb9l+lGQ/Q113tS5JEQDOsWg7i2HL017rQTRXIqacSSHm0O13HKZ4F
8X4TggnNaTjGNseDtHst0NEwVEj+6D0j+ptZhqxScpg7fk+boQ+hKjY5dDErHw2tr696ht/b1X8i
PlI4aMzh9dzT/aqjZkYLhYoPjf2d/ButTMWghiU1X7dfjx05PUa7B/ZKvN4K4B5/2AeSiH/SnxYM
QQHvukfCcYkAD5ct+YjdysC9r8HJfD1vn3BDnWbivIbpkjBR9Djc3/ogdK/jQp9RdmIYrLnVqWUD
q1BJtOcTV0C7sSGL3Un3Ir7kHNi+MPHWXOFofsMw4fIbSEqB2syk+D54IHQUR12bE1wJAY+WaLQY
vZITffCLgnMjXbbXvemijNkxV3WkfVD67mIr3C+eSNgEhKExCSFNuIi8Coh5KFck/VK8/AzGJ5CC
iRsh+k+q+BFNYITzdC31XLXIZnMnTjH8so2m0Q8kBtryzBP9yRrcKCEVJ4PGYnWv3AQQyQfzMliz
dXIh8xI4k+bD4aBMq231NrDurSJk9vVy9++Okg0zYnKyiAt0/kibr9IzMXkhJd5S2aWFr0MKVxva
H6fMsj3LtuDMNR6nC6zh/EbN9nMnEwQX8aZvvpV1TPPjvhflXhyLzr3U8cjlJzTCLy8kut9DkYlc
/18MhzbkBCDF+wGFkyhSH3rAqDpodTgKlZRoUZXnYiNsl323AfHhjGLeCc6vuGsQ+EoOAkVZsOUT
Iyrm4aWzlwqFg8Fs91JYdJ6CcVabzh0Fa5dLtrIda+RXTc8JjkN974LNFHivqkWCdGFiRAmsLA16
Xl1wZYZzc+U8I1xTTMYUOHIYvqeU+n/jf0sx8gPZDAdm9O+u5K2oLPWUo75EOEIMMCtAXkVB2Rjx
I9WTlUbTLbwZbEYjoRj+Q0TD8HVUUBBHi0PE459keBfHldhJrJ47WADmU2toNEQFrUIh2T/fPvBV
uVdMI1PEE2fCUHIL6LuDaj43eelTAIaCJGOrIQ3zchCUEphBG4Pxw50YhIaQlVOw2f2jSEO4eX9C
JeC+uf6FWKNZfGViDh2MlyW9/GdvfzJouJWyKg/apToqmthrBNHbCEV1P3TQUZEfzb6KcDcOCROR
Vg6hxAF8pmhcBSm7zGTD9IuVh8MA0uhypflUrr0x1hLf8KNFbqz6vSGLNt5hD9OSVtFQyycUYlic
1ZGP1sgK3iSdndVub4xeUe7jarOcr6f7uf7fq22ztXcRU/k4xHsF5FpnQMo98hUOaOhtVDf1mq06
47QP67FJ2a/ViWIE875ursxXCHCEn6uzNkIzSfGoxocxUdRwKdYEtA4Wd887Xpz6zTRx6O09qAwC
bj22pODAAuQ+kPbNZEA+Q9RaJSLDIyTu48YvGRdAGdwCBDxsJCqjVjx8bYuGOkF55dZL6fni5Gg5
48FqaRW9bwhHlKfvpoPWX0TrsNEnTk+bgqTjV6189mykTD7UOg6Ws086tUBaJ/Vi6Lb4mdEADU31
SFQUbfaT2+23OGuv4Qs4h96/rc28G13WvLcUwjvyeWUS4wbbWHwSl1dkVLLrdnPScF4f9oIKW9zA
FacDI1x/p/VOjNBfKEJ/IDCX1BxQMe+lsWP4a75ks6nsjP7E0d5wnvzu4lCpNXxQn3S18ww1AeHN
J4RyyECFTmNvhCXVgZgM3ZGYhUu7tzxT9VmgJDtn8vmp6Dk0W6tdaUDP024XlN0Fk8bq5pAKRosE
6IyCXJp2Sv+qA7iz9oQdByuCR9Bl88IjnwUasQ7QOJusDbray9nVU/lDIeLba/HC9YFdx1dhphCD
FJHDucnvZIrjeqneSnyvDkE78oLsisN/bP4VUKj1C1auaFH2m9QcZL+/LBr6Dp8ndYY+fG+fUbME
qlvl9bMvBcQas8B18LWHauo7zcWQ/uXONPc+5Ae2llwgR3gu1xjQvmMyfDGqyZkxN46kCVLCxlkf
NPuAmOj8fs9C5dIKVtkuPHa2NMTPtsU76yoOpSFmcv7GeO1DKlOs4kHfq+avZf5sCXzZXTYiz0fz
E5UUKGFp+QLTRx7//h91i750YO7u+fN5GmQoEXBJpsW2MGoNipUzBK8KjLWSSW88reLvo2f/Q5tM
o9P0s4eTVqxuzVXQlrPUosPI24/eJ5WiRhXCkN5HBj3nhRgoIyDQp/2AEDnzWAJkKm8Fzs+32s5t
XouL0P91TqWbzw5tLwMF43Va/qlWMM4caevAOQZ34uQEhYZidq1JIQ1+Ooc9Uaysa+QOxPO0t/DX
h8GCfjaxwwNq9G85BClLDGSSV7F+Tz7omtIFqh4uxKVHK7oM1sLNbi6YpyRP6FYZvmcLMheHS4qz
3rElOKpjXNT3aQmrbcZtw4hjN+VkyWKmgmWEWrmUdZAlXnCkaNvLUaQ66JyY6nxSpmItgfNouPTn
quMBedfEFyH9Xr7cZklqQ3E/XejAVUcgyw2A+X7jOc2EBpnhDlreY70zRE0UhmGwIjtnSdRMM9mZ
OrNDyJVa+wpdQn6ozSzs3+nc481BGjuAUZ0TOZqR4YhdYEa31/K7GW3RGwfrvhdrAX+9W/r//8mQ
WyrD6FMJUiZ0I0K7UYViJRhVsGKlSt2ikHlnt+2daDhbdxVGLFf3oJTqQuKA8A5TOBDJSeB5g8Uu
zMKcSjp4H9LhVIzkNcDWgzqhNRsYKM4i5wKJI4YPVNFA7F9jX+XjxCT3j/JJBt4vWRqJJ8KvMejB
3ITE9FS65XMxtpkTS2HDGBcsHyzqxWXaviE5QTIParmHeyCCShs6T7bWheqKOOlxhWWtH+Xt25DN
iiJ5L5X6c9NuHYJ9jgR3ia/qJ4b8RXfgdW/ZRpP9zdTw5Mgy49q+bmGSNziGCSHBFesmi414ppRh
+8nrrTti/CGBAfPX4byGy0n5qtwdB8MFHfcb6/gEJ/g+tSg8HD0U88yb6qH/r8M/1cRse7i1I0oM
ag7kRfOpIecVkbkCJRwMB8bxl5+Blu9ic8RGRkJzFpJ9L9OWH7zc2DWa7aw1DbNf0oGCJ6DSzYQY
cqGIsavSH3EK8Hd7CPSFd81cky4sURs1s13OZvE/vI39ymTAmvwOzveMZ5L7qUYrwSAYU8U8nveB
zttbgnHAkvAsLh01e8Walf+O8tZKtW908Altj+txaRLI+sxP2+MY3d5EM5xu3A6f0qYL5gpYwPlB
bMu+89RKFFegR9FUSKPcq7qmmu1xkZgAN8/WNoheu6H1J6XZsxu1TXEJrjqwI2iteNE6CT4urb5U
x4csr20fF2d6x49SJEGJ/NOala2ngE6pfoHnfDrLf1HR/ZuOSv9Pe+5ScR8L8PYH5SruNkgbj7X3
VveI/406heRQNywj6rvbFD+lwbuMtQlqwOGf3uOzJ++BRVCrP7Ii+1Bj1sapaDcxGVPSKeFq67/d
NGYFxpFVTxbYt6fDqpZxOTYLSa7lTNCMHA3/E9chfNnQN4+ucG77FGqfIbPHz4QA1EN3jY9iU+QS
cjT6rvoDw1oRCX1jNbV4fiX8CLoatRebTYEpCoLr6utlhk0qHelAyVsbOIjtqE39ZTYGAqGpokv7
fkNJYA8c1jVK8SW+EQke5uIcMRge1VdSt8+o6D29fZCGekPT43rEnDMrwO8ljNbWHmk9/WWkKRk2
foaJrrjidhQ1MeJZ++JTftng5PUjDLq04IKrAMLXV1YVaM7DwKGcRyTtqs9yb463dem6vI9gC7x0
1az51LQbBe5fQnI26igh8sg2rBXL/nANZXlxFbP4lNf6dMYzmFjPlUnHNB8Ij0pyH2XdYdevfz/T
OVSwPY2NWH76XE1ygxFVEw9IUiFOH2LatkcoyoYd+VqKuqnDUb3qd4icq88gCwIR1Fz7DWQyDz7n
bextC7pQJjl3+67ZnZTiKrd6fmFkEekf8JK7sLJHYcqX1UueVyIdWJWre2OVet9de0HPml0dxUzY
Yj/s1k0sTCU5CwzQ6qDsK6WbhdHaSdDUBKoxHepDOhqP3eoC0UuXZM8ZMZuscYFQYQV+5ls7qwRL
V/lL4ZdwyUd//m3E7mbqMD16eRfEBwXOEwVMLCdhZ9ZT7N1SiMQmpKfMUNZHE7AtQ+GDo8Rlb9aX
jSP5rkYyX/nz61TboscbXSX2ueu8orpoHXMrqs2fwFdC/vSKFbtbMM/DnlRKo/OhZNjS62o4yABL
UjBTEKF7OwycrCkhVrE130UTiFF54dv6oe8Jv3E9n7kpxPNx4dlsz1xGKoaLXXnF2tLVQXvwnaKV
7RDica4WIoLHkQlvzqWXO+WUvjPUpnIHB6xkY7H4WnVrc/yyjRgRtvPpkVXfKKk8IqH+DbEC6DqZ
sOK7KIbJfHMm12hgxo8oibCUKjtXFukqJkh6xj+aCpwK6I3DaLmEd6+8WHYtobIQJrwhljpJhpS1
ybeDXMek2guj1vLmiDio2ouDHMrw9zE6qlLqxw1KnQz+SOsobnj+cl06TcuoUB8PdMnZSN1DPp6m
sjYS9TiM0DM1o1HQFNZmKZ1ogbjgx/AlA/kelD6uRSbGTeqaSUII/EJ3bAtSpslRXr+e0QJsveTZ
YrJpd40K/IQtAk2a9gRmjI6JLoW4YfLoDWeumCWn3gDKYG1XBmpDEeMCPPOdTC3KrrK0ObXZIqJQ
nAVnbqk+O+egYSGHcxR1Cc2jM57ea8MOZVnYuLEC/2TEIv4MwE0lAWDcfu8dwqaz7cjNsUoR3zbD
QZ4JByzmCNVMGGFF4P16YMYsgeEaFpK2YjYotjVF7dwE6qQf/PDPABChwV/8OhhOLP/94K+h7GP9
d3wJkxieV8pleCyhqDCLQGT6Q/OXTD+3BUKPOlfNDTvvKmSXqJcVpDidlyVjHDn/MAdyieFn9cAZ
RHUmu0EYqYwhsdaxKdHlu4e00MipSy9KYHoIE65OnbHKNVYWPjr+0brKazFA5SIrJ6H8RXSXG4v8
ScIF0Pz+DlUL8pjLcJ7x4gK9vXhh+INlEHsY8k9m8ueLO8U0FHZpFSjMGCTQ1TM6tmTu8Sgw1oMz
A//NlkOzV9nWOo1edXJXbqyGImhUeb/7pTZrdtmczQRWHqF5/xZD++flF5Sk4qjtdkpa9yTKReBx
qdTwCJcBe4L3KkY7eEMWFYwgtoRs7UJG6oMuVedBNu9vYTbxL+b8zKp/e+LiNkM9yA3b0+C1dxn+
qfVLHK5+E6qN1cbTDIt7QcAx7+vc0WFHKLfCkCFDeXsUGABfpW25g2PKAswWMjjcoURrTF/5SCbU
MdRs62d2dwPsftZgGvrLO5I0G2cmRn3jSq16So5UzKOWcbTvmPi8w8AC4t8bzv1CgIhO7kJ0dcRt
Kv82rhEVIBZH1CCsf92jXio8phQJXf1qAfVKqxFlcf6XdWOAz9MR8Iq4s1fVVP7U2POyeuO1woS/
Yj4aEaVfkWfB9I94mFh+D++l05KFiVGpWDewmxdsuLVAqtzOofXSanhsNzpkgnTcuzQ8EdIwiEum
wH8KVDt5PKp0wsrDddZ2hvH986wT35XXe8nxn+ZDGWFrP1VFdXVqPXRCv0ihIsvtS5AeF3fG0WpQ
a34zx3gSR2Fc8bQWJ+20hsz0GsUDwW0Y3C1Vi943z2c8gPDGtUkoBmtdsmQlGNUuJiIOG71Po1kK
eM1sn0h58YJjEjs61fEdwugdlB36q3WbekMVffLn0uvbMtVPcnNpBPnPNYz7QL1E9tTBiuRdeJiU
k0GBEPv4zMT8pQUS/cYQyGAELxWA3Hs6saddG+g6GebvTNGZXLyc4sA3B9nP4+dt5AGGaYXP8UW6
zyE6HBtNFNDhElv3ykhZrqbQ8BQUkkDlRbwic/2eXBH8iFjaTTGr5T+s7s+FvvUqKOv1gSW7fuj1
Z0ML7TGzhaU3IohJ3wUb3BoAiGxU9CBSsFlW78dXvvt1LfVQTZ+8rcEcchIhBW7pvsV+f3CYX426
Seak65m2KmkL5Efm4pAmyj8pEPbbl/6nhZQ9T/HlZmy3KVhKlBUSr4wEhTLcfRLii9QA66Zg6BY6
UR4wtdKlOzIYQi3hXYR81CFaMBc8xVMwAve8wl+fmEhv/gApglv2sGkL0lyx7TROtRGHEJ++LV6n
O3KFCW6Q95JN4Ujgit0IJIxzUavpkUlvTcI17R2kNzLWRt0uaDxcFmS9xSYO4DHnhVAfv1VlUPck
JoUrtMloOYW6e0uykXlAz4L71AjtZGu6p18/7GJRIiAUUi84knkBTgKn3zU/msoc19JjazNcPxMV
K3efsLH0/QNReG1u73BqEYMsNErZvCfjI+CzIe9p+m5NH9Q5wDMDrdjdfq6qCTenu2+gYNC5erCj
yOSp0uswYXDE7ZVLuq5et6ckRrZLVuJ0mrXyrgG+Jtr8WAmziP3mgXNHd01w4PXK8lG/GeLndkO3
1A4U/UdM6L8YqNqWLRZjbCTT/B9igE5df3ZZWQ8BnDy23ChPS3xApgqBZ/zgQKPfYc4erLkRnr6F
xLAOkmp1knc2oc09ab550uPQxG+JJJJ/SJQBSs+cdUpPwv4dm5bDKlzJruH1eX1ZDr+mLmaEMHZ5
sFVxa2MEZqeXrhINDRwO6k5Lnl7YnBUaefVWPP33JllJ03AQxMXlH/egjryXDu7KYxxaq4beFct3
2qCwGml23JzAjxb7ZcLYgS/5bAX7uChrIbeFisRCdmNCtx7bhtrNWXHhdFT7vg4tEzD7Ng6Qxv+A
BXonrU8TLfGFu21A+0J/ruD12CthdrE+PcefbWWS5tBuVd0zsgmZzipIghcGjSL++p5UmkLEyHnk
4SZi5apDIjqdtytwv+mBth9DMHoqtqrVIaqPGjskTTTrw6rkbWVpfiHcOft3+Nz/+yHcbZXxpILe
5emm2b0OKDtitnWhTvfdF/zAv24gAWneAlBty93mEAjBSIkSuPalR5+L5ia73g8tiqe1Rqx9ViSS
2MYA4dAnFKtZMe5HwZv3VojgoIUhaoDVQ9+bMBoOJAWPIcOyzkb1FH+cfK9FJW9cKoCBqWmOg/zw
+VjiirsiDdX1FYMW/nX60i9DOkRnPfZ+VWcpuy0DGrb7DRZ8eXWB91WxpQqio4R4oLoasqE8Cq1L
oDI1h/URcErWaHTGqXaSjBGzSneXmwdmftNIK8fJ+5rBpTa4g91Czjugd87Tff8Cc9MvtrZYMTwH
LslJ11xJ9l4GfQYXiH6cwOmC7flpFyNkRxIxkn8p/XwNH1ZElxCy+8xoA1jcYA4cmDgo1DGfGRIJ
LV1Ldb5NRUkZhUTadYapUankhKJD93AWZiaqeoSXpKuUxpAAVAFbxt0TSZXJCtGq5vND+8Frh8PZ
j94t4X81/IlYKOW1YldIwVgc5Tbb2BcAsJIg1sYo5jx6kUmPMIK9xS5/icS5sFsFBwLxfwDZig/d
FN8Az3MK873ZQzNw3FDTcMWfuQPk0aePnqx8FPwrkwGKlqM9g/RSbHlNSFxfjHdSmHBZ+rrQIul6
eFGom32csrFSJpmmBRUT/mquujCKKI3LNUS9lEdx7lwLX1GRrsG6F/VMXEVCn0k23uCj+L6Yas8c
W1SN6vA7KoHnrRL/hrDO86FasuCywh1rk2k4mxiHT+9fMtFN7v81yV9MDRYOHrMc/iZ88f2MTR2+
Q1w88uirJ/Al70af8TmbuV8jDIlqwEOTlMc3oFhIfr+CqC0M5c5PxD/R0xVsObRCAaE/te3d693d
DGhhCBbXQrhgSRrIZeXwkV8I1i1XW0A6k4q86ZYp3yAEAqzucWPigcqTsgLMUeZ8MPOZBUNrera1
7uEPPDBYBP892XvQlDRJVuUPAmbLEfrVnwAbW4dBa713HRvK3FvKVBeNXPxsxkQ6YUlIq6pNm0ss
FpUPXEZBqzOpIqAfJnBAOSjgORi0powKNLElW8Rng8V/2PwgjWCRJKWRjXVs3vgEH2QYXInkk69m
wkia/y2ZbdzsfH+bSI+w9PHq/bg6fAgHbV9tl5pf6bnVRbYhohug7BwOWvsqb/aGy3UdDDVIuPAN
eHhd4EyYd+22/xRiz1UOPPa+fYbQDgSESqNGLuN3w/ELyAEZMF+bcYVFR1jhOrYYbFFPlBJ8CP3+
IJYHm0aYByYFo0ngFYXePOqv78DI31uqT7/sv2cCrN28wexFy4b6B6l5GtOf3alyFBxwy9uRM8WU
2o/yz3ChSyrJiGjB4qv9t8fol6KwuH/VQdwIWQlSL56exsnw62AhcdGeIuGK7926s1TZ63euENa9
ku9dpLeIQ3Np2N+YlcIMx/xTmWJXycpLKMWTUC7Ys529QpAlUd/4BV9jdjP/GK+XW6V2Ed3/CCsn
if8m/hid9GcheXAdOQn6wLsMB1b/zF3ShjlN9jaMrpVGTE4mFETB0B4mbo15oyZBA0Vq9X8gxlgc
V1Pv+FKh1Hz8QjmdRM35psrMh+b+ISaiTHm2iLIIdfaWgcl3m5FFs2DDQ2O0+DH5uECWoYgMsg93
X4ab7MeDsNHCPe8rpiiQmqlCsWjDhOrBHKmjCCA9fcMUF2aecIaRfsP1Km/eRDPHYKbj9gWE1aUp
Dui+fmNO9frXmCWF4updPdNGK+U7yHozM1TLk0Bk6UaWArEtgGpuoSY5BSCGmM6lDZZrv3FlqVAP
tPOr2J+noXOR8Vdb8oFDVmBAMPxdiQbETT2zzuDLqUYGIFmw34CeCjg+lmh/EzOLeHc6jt2Swzqo
9y242Yoqhddq/AY6J9EMz1bh3JNkP0MlTkZvZGVyvCsvImzCBPp4A8E3OW3mi2EZgFZ1Rn9GkHKa
UeerX/5JvJ4M0vFfIibHxDMz3c9YXZz9jbnRiyl1shE014kVv1Oa2lBgW/UsaD6EFz14Ak3tTMDC
qdSgqihqLt2HVhNNN4uMe+9TF0UpEYrYymMS2/WZoltY+d+BIhXvhRDDU991dkGv5/Owl0TXGk2N
acAaaD6YYgwIEB8FqbStbWMB15OaS+hg0k+2KGjQ6OElsqba2SCKtwkkdYJNu+qTRvSrwK9Cu4+e
JOVvZ70Ve0JUH22L7srOCBsNWpzYV+/H/6ocHdhM1jsBKZrMZGXl6CSsmgacUUsKezQ797e8zl4o
t51+BWvJIKRiem2t4rhutY7208wrWuUWB3kW8dNydQ0+dfHsrY5yHzyxvH2wkuzoMqKF2rvnT01N
OX1nue7qTzmgVnhx8mevBV3hHP8Fuob13ekQx4xvHC1+XZ4neWvED80qrLQ50XlTQ5lPv+qRo91m
q/lk5D4yDgNe20Oo710tFX25BcGa4pVtlfvbkPmAMnQJMf4Ai45K/D0Jmew73ZC53zjVbOzFC0YX
HapXOwjODzpNcabf5KaQu7dU7qZuPAD5xukzdSz9meSt9kvs6iMmOjtF4wldV/SWv6SmUV/eVfZx
58Q5YeLQOUgl7tMw+kus2YyWXC6mrGrzBENp3M/SpcYxvXDve4iBim9+FLjGh4XtfWGKu4dMgmOV
QBCUrZ73od9SncEdGZnHnTDmKUXj0eFCnz0bhNYQTjdfYd2ssW/s1PSKKxokvrHqEDG1zBnXMrsT
AKDb3pGGcJvBgYUeSkFHSBCyQIYUOP5IyX9miyYuda5HroPeuVozyaJYS9MvLjxINtkmXBQqUy32
UC6Ie2zyGWzItHs8hDSXcwmLWvRs7vPlm7eZpex4KlELbQt/lpYBN1hYY4Oyr8pxOTFFJrQ2gMAz
ECNmP81f8MIhtoB00CxbPLNU+0uEMOI3M4gSEWFzqx414QQ3qZOK1NmLYFyMuzaiOFi/GldNWWo1
xl+5CfAqsvX5biYc36wolHQaNXCcGxZ6CwwecVvvy1v7QRvnrAtER89bKUZjbzYeIPMJJY31FbwD
AxHrlE/o4UzuVk8uoB6s0aJ6ZjZa41X+wln+Uo4+2gJh5KWd5dm1aQlD4N7A93eFGLnzAJCbMINM
tMu6SQzRANn7eNSYoYm4dbkQtQ8uUDzqSZNqi+IEJ1AdfToOAfZkRMcGI2dw5N7pmbdYvC03IAs7
q1LYCQYmP76A0MXQBbzWg/ZiaPGtjmfWbnOpUS86ohRNRItvdiaxFNaKCdlJeAGvX/ORM3nYfRe7
/HjkyiOJmvkP4+tThesdea+MEpqFkFlRCsTUk+kicuKe/2PklJD0Tx6BC0gQVfD1NpuaIwzej5az
qkPvinP0uRsQAUO5CXSLBaSUL7lTKMFCSKeRGD6oywPkqYEw1vkbBvXJSDf4D56ZWCtXTUOj4wj+
p2OLMR9XWkVE6WEd1ErVEDQuAWIItOYwqQNsxfeBDRM/BaCgdYSuI+VhS6l/S9/n37ldYYFQWqSF
8ixs/CbKdLrjWRgdk45dGS/xnJEIT923BNRR8clnInVbv3a30DldXkv0ziodOS/6/nqTnuRVj8x7
PECQvClmucqs4PROxDue4uPzhLMTuT/kt8o1BeaR1XeNcQKRZhcY39YIAqso4+CTh49vqZZJWa1A
ZNo4cU/k7Ezu1mtINjXBuVc+5E184g1RUTKWwMe/liDjtooxkfDYohwxklzTk0Ou/N2Of5Z/BpJN
fTAGMJHkL7ze3D6A+9PafcFyYwy8v8QpPJtg2rl2BG7qSRYKQRKZp8rZxHYzHiS9vhgR9k1z/QQv
6Wq+IexJbjGu94g9M/rFvOQMmGyx2Q3V+D7teOJExSsuVnD0FAyyIGOjgh36OxBdVfwAqFQNBVUM
/tDCYc+oKJW0NbnwxpLfot6iqKKtmWgwGkrZ/jUZID/ZTXADv/ZyOOtY97nwxQBjwhwI9wODFFgB
VV0UW9d/g5fDzyONFfYrisNAZfbLRaol6E15nV4CZzFihn4qnIvn1NQYC8xbXlO1H6tu9B186H8M
CNgWZoVJ7YqH57SpwkbG2mc8A3iG2Zbe8X3pw11n9iRXeKr0dnPriaia2ie5jtUhMMMAK8WImNxb
HXVi42CtoOJVHWW4iKyphnu4qJ6wKzTUZAq7jfFXZ6vtrFRymXE9UYFIdKtNb6Q6rJCbEBjS2ENs
JCoTzLgBdug/Aa7wRh+d9Ug3bXu3pTi7mPdAwTFbGTc22vG5Q344KrS5d1Fqs8f45/CErX/xXI+I
2n9fAgDj3b7bRb48Vt3w0zCe1P4/xtxmnW8CfCUDGtHmLVHr09phYkGEA3++Rs4KHO7UjTDC4JNg
71sGDmzlCZYbsCW3SaJIWzirN4S23D1XeXr/Im2B6eq5zgCrhFkZBXG1rFYVvqfa/KFM3SHldewP
1IynRgrZY+YMyk981bRSlt4UetCjRY+VM0W0i3/EXOMrLjQi4UO+0CCUUdp9dURTWm1vDpzcA+AM
kVtiF7J5jINGZpdSsFFCMqsBI2ARoyOnNWbm968yzALCWZROphWsSYJIpzlShNlNh19QFHs9l0TJ
5Zz3RCQ4ztxsbam6RkXiBzGwQE4bGxick3RtzQs7pazcubvLtGZrVPF241jLLiSONdOWE/KnKR0D
ufqXd7BR4kNWPppF/QcX4n2fosh+VtackWIGoA+5MyLsw6q5DJVZndqP+4233arw3UpoI+bYu4C7
79CIQCiZHTKan7U60mKZavrQFWh1twAVDLuIm2g2xe7rVHH4tSJdKX8BR195u68QxbPT11H357z4
q07yg19hoaBI+Rt1vx7gx6Z2brgx7AJphd3F3+NJCSlxxBlGEsKIm5vdbthPLhhtZS76jxU1Qs7K
aX9IViP2ZDcvmtxTaBXbDT+Tq8LKTFwk4sQCIVa1bbYCkdrVaUjvOpH5FlBuP+4LXBb/FJBrD5H9
sp2WQnOQAJB0DYUzmp9WR6PndIgeeSLIxkWs44rtwcrFeENWIx4ayfE9ADfMa3hbmJSE8CVv1Ct2
RsdwTXJidKtcfSDvZZVvzovzJlN8k/p1NzpGAlrYD6T9our4/wqSh3Qw72Vrm3f9SZ08lWvSZMBN
L0S2jw52FqfRpG+zVSz7BHEPey6oG4xcTh3qDbBYIygLAG7248qZ7YPFvy+ArPG3FGErEwK09ct/
kCAXbbURvJRQf+JMtC8OIFX1gXaacGAvxPvTIsNNx9LUA9dfZiCmqiwm4eMB9esy0K7zEsDo29s5
WmfxtujgpOimZNMUn4OMMDIYMvgkw4eI7rNyz7b7lEnw6tkiY0BPiv6sjWr55yySFEUBPgbi83fV
R6mcVHTI+6Y1a7Az2fH8iTQUk+I/Cg5h/8RJ1Kc6QpbBLw3hzFSyJJOsDNUVGo3DQyBIhqBa45Zl
vl9CCSJBT/D7QJBEdciq7JpRFWP38DPxb2feSEHpTLrtBTslv7nJn/O3J2Du4p4koozk1AvwNS4c
LTM+AHz4hmU02VcpBLxaQuCKzU4OC+RfYwrvBMS6G9WvyRScSXaf/dDBeDOllNKHNiC4q/X3UFjV
IZL7TWS7IB7lZLT3Ll0qIqxQf1LZj0a/RVffcOJ7CaGJ6jT+5ywRS+Bb4dVtpDNVf0HmUlSjOe+e
wJyMB0K+KXmFlfyIt0CK5LPOW0zMyExHOF0umk/DHjxazuSrIp8i2EQ0yKF7X9d9uYrLKkLgJbDc
F8VS+QVEbFYiZDl0kmLdakD/JqxYeMmLaJ47xnqpCEYKI6vn5j4FDRNIgaPS08pnlsrwgXZGWJVY
hZFS0qe9/3wVt5QUk9HC5EUuNqxQJj1P7JRFrsm4qE92CZINTaKjBwzHADTJ//TwzZfeHRHJa1a6
rL6yrYC1xwavdd7Ylwk1KttibGV2RY2n3oCJmfjUFz2teJ3VEca0uPZNEvc1W6jDP24xguewtgh7
KlhjVv7yQN/Bz8Iw0/MrAwLVJFnSXMNaEthK/jRxGfXatCP/fad5t9MBcj4bzkRzbyp2/+QyXKxj
iaGiYNZQDac9l0w7RQo/rpV8V24wKhMFpuWagfSuOktz6dJC/9ViX2eFoMXS6WiKv9yEQmXq8Iph
vOE69VrKPvFPhgn7afyfeem4dNa6tPnOHay0p32g9M2rMJBkuwQT1FTXV5s0Tm2tVKdLGH3m8B7q
qF6+e7wq8TESdoRRe9dAn0jYIi83TKCKQ8ev4qoiWdjCSKgXbk2WvnxLMFh24KAER3wzCRJGUjc+
3F/1+PpcOJBK1cc5K5zQGJcT0nj95LzabtRjcHp6M04G4cKtZLq8dHEo/t5+QRQcm4Qy0PYfgP4f
cgbF6yMH65DfdFBwUY0zMpgxeVRmQeJa7v+gg4p3UF0So4W0hl8m/0jRUXs4J14eH0evHRClby9f
NUq0ppn2F3YsPj+oXOuvuUSPnHCTnFG9gFyCBtn6TjPYllBkumwqADLHW3G03WtoNmD8LxQuLcaS
NuBXOGzmAVEBFDv5yYd/W5MpgyTbgMJyje9VDX5kPesroR3jkuu+WYhcm7f/GHUtwpBuihQ+z9be
04ybuy1cx8lFuHIrSUTWh5ma0HRNCU9b8stDSYSCtJgGIIDR2nspmGIkUbeTvmtZSLLf8vp2+Fzp
vy8E7weOKe/KdQRJQWcDzyCEWy32w+ggREFqrDyCqOSXIby0UyiC6rNFaWBMHRsqft0YHtQwda5f
22+Wb50ubdR0ws8cwaQb8VDYkZrNvyAdu3nRl+2oirWKADI3rhmHLtKYEnD3UVvVR3pJjql0Spls
LRY7MKNVnFgVmVJabaal/yNJXoN20JXdjEnXoQ9NSSNs3FTpcdgKvv0xUBb64qDlk9zxOAB0M6yF
Vv8Kk9+cFnoHglgIJZ0V+FcRoNhbkiTjajAc7SJfMH8LMERNP7/NEkWYRrVcLZ6k/Xbw+AcSYsIE
cIRHwOiOPVP3YaCTrsJnnwQJo7+wFwIbv2vTn5Fy5beUbBaiucLp7bXTHdwY2x3CyhIwZ9cDtGRB
L41rAPaMIpUje+E/zFdt2BHa8X+ZCNJKt0JZQqtUF2yJz1c3iXYVWYN0Y/vRknHaff/OvDs1ehGB
9zz3hrukHvecpfO8qPlytdrF9kI/sKBqREkYtDe4dhA1Ht+yQuTGqGC/h0JKds8sS821rtRzyE0e
QrGOkH4sA0K4l+HPSIdsnkDQqOIPe6DNyiRIyJzZ3Qn07MS7Hu2imzCmMSgLFrzoDYYMRanpKV7+
eI9cRHA1M1fv1J4HyyeGgPYHFsBa9OrKKdnhPE12IV62D1ijQwsJFoi58wHnxgsF+v1c5zzcZ8lP
X5Q01JntUCl89Ig70ZLpgr4gZk7kOqBG8WNbXlAPKvKRBZT8GlQOPMKMo5eMj/ma+kEyJX7cf3S0
mU+Da5LcXmisAEuoy9f/XdhGO61SzT3fL/weW4+BcpdNfqLHJsZdfTsK8yJDCN2riqsrdMw6N6rt
DcATok3KHDEN2RtQ3/TUeUwwAJ+7F4h4hT82Jlz3WQa3HIb+WD51VkCy21bIg74Gye73RMQSZmVE
VhLDFaLxI1HG/R9hMpOeDiiB3YQ9anWz5/JxXIWXCTpbnPsyFJB46+UC61Iur+Tg2rqHJ+VFT4MD
DdKpOAfh0AcMIyfB7GWcvGJut+SS8AYgCrWuNemG6VhI60q+3/tEz6AxWa//4QgvN26+whkb1QNd
sCCvtK5GURJ5hsEkC9qcvYncnZvOJPCVwRhBis9jxykwoWMgnq0TuGDemi1aPuFWALTaT535Fv+R
XZ5HuzhTS/22+nB57/svg63/VrJrmO/FPRjtx8DVIjGZewwvTHggohdRqL2u+pHiif6pYuPqMUkN
OAKMQZnDkCnBWcYe92WNdWby49bIFGM/kOwpa/fPH8QmFLXC7oNqtHIKaZtxBQSWRv4RnlnrvKqV
gmK5VuoEMFBYubyziJMxvaKYV6Wj3kS2N1dGUvluzfSduHpsOBVEsQWCsByea0h8ZPSiTW2BVwAE
auaGzSe5NQa0i6BBHkRMYlKi6Id/C3pwmYbfw4QRPV2NP1bvwJTtCRusxoKyskrbGcwdpPVvsh9w
HhAuQ8IIqdN6510zHPfjA6Im2q2WXrsfPI0v2kWU2VfbZdmch3Zejo5DJYQdf9X2S4LNMvPcZ+Mj
Y5Q1j7NI6oLqLfX81oU8ozJJ6ScdPr5FGttehl9akUUSO5/f9D71eEoJ9UCeJ2yjBLsUcZEKTK/0
+FiO6zm53WPhTt+Ss6QW/G7xpS/Hg5Kn7upcUjh5EqPeTYrUiU6RYBIvEE6YONqZOALe3tQgPVYe
KqQFtKj4EHS9SxvGHhvhYJ2Hik8cAzUTC3kh5zTmSe/94Dw85mzUzhZrHGalAvfO2QT+cmaf7Lkv
0L3xqPz4k59xkZiyfS5sHjLBK+bZ5Xjcj2ksV2Yv3Wr6QDTfOfb7Uv6Crw8+lCVL3h4twnRu/TzI
MNxGvZQlnpDDr3lzG71SkE9embyMhAnTeQGl4ykXtOzFbbW76el34W2gFybg1ymxQz7wrX+NS1If
w6mgr/4GfhRDNA9Hcw3QD0vmrFAp2EPuTltAs2SjRLmGpzuMdu8vuJt/MnPsrPq6athZRnx2zKJC
heL+wEkDBGjuVn+RwQWdAUQ8rlFS9JcyalXUgIgOj/RRhBjsP/4qpxBOe6ofDjWId+KLd/EUzEkm
Cf17XIX/vZ0oElKWqVMOqy5zpasOQ9g6op6MMrTm0w/Ef9yrXpeWbj5IP/jWwaIBGKQQVE+2mK32
2MCXdNwiL3j3BIROpIXib/8LM+AAflRiq8OSWkvMqzYTVBgfns8YBfyXfdoYXQs8TuedkPOIuTfb
3zjMgVGnp7xR4W7S+4STQ0e2eAqMgPyAoITCQ4VM5CODBvfmK5rd2zxRDHFlba5Qz915RNiu/jBb
DWfGcs+OVNbta+7a2HAKPNo8zBtswVflG2fXc9dBdYKkdE0HSudVMU8DckTHXfJWRz1TRPBq0pJ8
TVpdEWBMYR2pdl8X0RLERxLUhunFDM1zH6xjVNOUT0jE7Tk+q4F9TBtb4ifnzrYCtkCPadLb5xNT
jidb1KToJWy/aZlxEj5OcmVgiLyvU896F7Tm0nr8sCsihER9Q1EMp2VT0fh9eX4w5gyFZyMnUt5i
vpKJSMXEZfqAK8YQgXbMBowyuoirYZg2L0o4oDjnXEdGw5DpHzgc0PNQLMDaXg1Tx3yf08rHJFXT
JfovmKiWrNKZYgPMuOCQoanC5+wEZHwNQ8z9ITUTDXYy6+mCuw1SE6++bgjEGlBe0mbgtarIJ2Rc
QPJdMcNIHNvwcZIoj1XvFkiIozAT5zXAUbFBiNj1u9tcVFtIdcY3cBd1nOfWhb4EPOY5R+oczXdv
v+tnXwhsUGpNS/R6rfrqn+I16D5ktoIV5kwR3a9kGV43Wb0DheMbvGQ98huZUFslSawPHf6T2t1J
b25+DAqFpaisTIMm5Q4HaaVc6nC/ffyl09OrcHyHvuUhUcUaXej+ugXI4zvWeMc9nAsO8wfVviSE
EBo+jYr9FJ6YBZJu4ER8bQJo6lIGH/oQPkf8wcyxksFJez7h4ZlSmDdmiaocvkYG22v8D+P7a/oV
fzHPiDzQLuv/p2f/6XbxUWT9Za8PdLUG8CfpWT6tPlZsGsvpc2g11RANpGaNDu6e3Ge8k1813Xe9
bHsRwpEcMT+8VhToBKvTNMNICEoPN/MOsfvMSiAdCszz834bus8S2iWTEJ23Jk+P5GXyFiKlQ1r8
oKdVV5qUypqDwePdcyI6DTY8DQV+uS+nRkY50bGxNWFwO0cLI+csnGJ7QCbBXAK27wsMUbJQH73y
f7I4i9xsBibywXRQSfvuC42dFD31tmnjQbvykiQKeQSd9mnL2fgiFmnp3VRzTlHmgYPe2uyLB2hf
lz1aRNnef5T3TngPnVpnqZjQlMxCW5SWF6yqkDSR4g3kMxZeLEkqnxBKOZ4ZvZuVpQDYLJXZCQ7n
HDn3sLUFQPgQ9iCE8mn+LAIGaoaQgfvFyVpDqz5lCgSXBYrX1pjo79hqQmY1Yx8EUxNXG43pRrwt
JGfU5lisQ+6LjWIKRW8cR3Pu+p5rLtD8NC137tUEI8M4BcRMznnBUyWJ+0iNIeQ4VOoO49ZjxFk7
IFYqmE8Wza+aDg3feZZPHWZ0hWXA6O8nUeuvxQ68EzZyFyyPBJtxcy6SBjy0dXa72ZtRtOyBeU/R
EnY0swf5s21lOypaGa6C6VWrs6W/3D7J3dcQHo5x+zgfCEQDF+KxR6lR5am9UfWy/sx4AFqnTFRt
bXYi/SUQ+UqFVA0I1RnO3XZci9O5aIhj5ipPQrz7sLXla/l39O0ia3DTi6QM3HVMW6BJKDfMR/Qu
enfFFDIxbalU1dgm9I1VsA934MnSzN4bKcdVKT+UvSA2AXov5x7pXwAbC1GJgjF9pKBiCjScAh1Y
Ms5mlCguVBdkFoaG1iJyJ2t8O/mftM+aqiRyj6tk9LlMWxoCpYkpL84RfaClac9mN6NEk8F4IMhi
idnw4BeABcLtyaS0ayq9N8iiJBbqU1UgARMNgv4H0KStlB3AyHm0vdDnGDevFcPj+9XgJDHP6eLi
DBUHKAZ4Gd5oQRaNaCUDbb840Ik72SkpJmacDHKOacGJYzxSpV7HmrwKAi3SQ6/blOhkesgKEWlv
CvpV6Avtbv2MerSxKWhmY0sF1xkRWaoijLmJ7+IJ5iGL8k6bQ7hgd0uFyT8dUIGZsJzFwd2aDhFG
dUSzVoLg77oCzfNTR/aXy3FdwYzA5cDheFnDlC9wIxdWuYgsw1iTsnLR7rKKWXi2vesIHXJwuCxJ
B7HpbmuXBmmvH3tdwRnIFEOqgAqjMaYfPLzVTueezv6K2iCgMPeJcfmnwcUOQdJVx5C44Amf1ea0
82WGp+mmlDByoXTxcJm2hS+98U3QvyM35akkLtPIswebWtaiuAlla7BVCdd/kkZaUPCJ/s+Z4VHe
e+sgk3sMOgfve7NadHzPr1gR1l+P762pyw8dRpluzsLY4omrPLX6RlWKUEyyohGsw32wEzDVgfc5
bOl+oQ9eCJM4yjs8ndxgF2ccEJuVO++rCun149W0x+gDTz7X9h4+wd9UfQtc37VspoM9giTwGEDi
0bzLflXna921WOxBoISct1jOwTRRcvk5iE9Ri3QQl6dm+g1R11/RkjwrpIrmGgTiDJ6RhtI3Zxnp
Etuz5lvPvEF6g0tJZHlX9KA6SdzdYpxNwpx5+sCH2in60gkVhnIZZZijlXsgH8jtY7iPxd2EcI66
iS+if5LYxM5C2QUdsJIzV0jUFRG007YV3ugGPHLHX2Xi32Lqc/4hdc7eB/czJcp4VMY/nNccfmw1
/R8U1ky4MPUgsWqd0W+6+VJGmKPjNF12hCWCkKe6ci3Uv6xSUH9CtFHCAZ5DQ6pSWouMf0m3uZ29
4dX69Kp47ciU7vi/Q0MjW8PztFtNkLk7iTCdVIfLt0VEUMtZHxBPLNgP5TDdeydqwgJJnfmoH9FJ
2LtRpeh4TWpqCif1UOIeJNYJB6bpKhyMshWZQEZyFrWvpOYokKSTjyNQ7Zaub5uhOV6D0Ge9u+9A
UglOrfDOMvFSSr1X+C6wKZpHph8S/bYMybJmeSBKDk5K/FxaWFFn/KVkZqEUbi05v/Is/chzSvar
MUCqy07ygnYXtgtprPkm6vfzzZwAyUAt/2iYnO572F0N7cii3gDGQfrU17k4DieJg2D5ytiKRG4o
TYdNebkCf1q6YZIbyWr/D3DvvgloGkQ7iS1ajwQsvsc4PGec99XVyb08+NKPhl0W48ALPEijz1Jr
XafMweJJjBMFPUZVAeYqJBtw39wT/Y9wa9z1D9q6gqKm4ldFoVoMqr5g0inJTl58Rh6phH2mISb6
doLGs87FoZrrApeevCfBl1VUjTwaSAd3y/M2a80JQ2MIO0dAbZ7a4GjbeaFp4MYVxj4wOI9dn6nN
OAZqwsZSLcDvUAS+LBgyc4t3X4mavaEIBeDI+lXLi3DRS6eDPCCQAQoQE7GGGO7vODox7ozTk663
uKGJtpppxplO3FebRUvz2vQcTa8JTMlznlWZVRNTLOb9JywqEzkWZ/j0SLRwbaqAWCq4gdcSaO3M
ujrYX25DZwBtjYU77RrpAugGPOYuKVBqZjXy9Vcv9qhCwKRdz8MZA2jmCgo3qWZxo3NlYL0ccROh
2f+6ODnpboPynanc17Uv9naixpR5hVfLcNmEg11DwuIE/ObnK0OFtVv0q9womWwapCeWBzkH7u80
kRioyotSoZSfvKg1r+Y828iNXV758cMyZ9ksylw04+pq+Mcjm8K91mavOSfcOY1rh/a0Y4S5E6fz
eZ82nQ8/g24v+VjMu7so4sJQf/6YPrDc6wMK8AVNVd7abE5rsjzr/5HqbQpLxAWrqOnVBcn1LAW/
GE5r4WqMwqTC3C65/RH5nu+wgDI7BKvC5y7efyRKg1L184ehUu420E6KzHWVNdsDy8Zs7vv4oULp
WoAYBGCgXOzduIvWHxxyFSAl4k0yfdiOwkHMXq6/scPc4ay7vgBMJNdBhJ5w+NjXfrCV46knZ15p
p2eKayD/EmA7Q02iqxoZthP0oXLTQFOfT9OZ03qmDuCeNWPPrWWB35et1atnHUOrp3A1ZhvTKIJz
pbNIDnRdhz+FJONzmyiJ9cRNUiQzmZQED4c3PM3EY1q6gFXNTq7/B5TjqkU1lTH3cAFG9vt0NpYn
aroqBxYmaji2DLwkcafzHlRtBwcETJBgD2oY57FlOjnrzrUS/Ry7xa7Weis0jhKbkrG6vkHQIxAV
AJdFs1ZYzB7WvZ1xbER0xgkO0tIxd0b9dsd2kQc9f+q2WsoXVZ65YJ3yK1+eBA/SUoB0/ge7Ne5Z
Jxbn+gJ0PfuPRsBQceLndnPjvn8AClqZ2c7T08dXnX4dkg0f+/1KSCabu92PCJJy2w8pd//ffpH0
4IU85Xvt6Hl2rqJLK/rFD39izBQWa6qNFx7PXFfAqLBF4O0pB0R5bu5wXFnrTWSQySuF89Ov1FSe
Pz0TFDw9umdpiBwC2ViAEdBF/B3aqIbqYhMMDMNLkUxpwTlCYTxiiCPQUVxtYUHyhZIwjG/29ITm
SWj5g5CMdp2fDfo1YnzD+oXhVHaVSNFDdIgp0utN8OLLWf6/Hse73t/lQrhCIIy5fELcuU2lUDi3
DLhH+qVFzajItxJmJT8hIhAbZf2Txw/xQ9vCnRQB1aLG87oiaXmwU7BMKFoivjakwV68OI0AOF2t
FjoO534sjZvl2SlA0aAfBuh12O+5SiE6jr2qfd2ApfWoZBSfrHDtfDS/tF7LhLOpfkNXDQK4g5y6
p6lbM495iFHH3tF1qBzcxh6FZr5LiNQRP0/mzeqZ8H3u3SF59amWZwf0Tnc7B3Mi+G65K6n5GhjY
kOLQYTFYi/tabVKzNM9WMK6D9jdzPBzjLWNaEAivpbsXCxOWzhom1e7WUL3RMrgDNQ9+8MO4OXTF
NE76IhyREXKVMZ+od/EyS2x+w9Q3DBBQvC0KH7pBmD4OADG1wMocAq5n0U1/XQwdkvr44fFRTUvv
A5tODxs57A6qq3HYTuwfl/lDG7eDSoDsWL0XoFX7WDpXqQUcsdciURL/SpJ+7KHRd0BGzWSMrB7d
c8p2UpJAeuM3WqfBxOZ4ajZyOySVqZXO/r7r+mnTGsEqqswvuOEzprz/SHzY76LgB+LWdwu0jy3P
C0bT4AsHVXo1NiDCzy6w97bJu8UzUaYvmeJlKKp+s+EzKEg90dTCblfkwrh3sR8p08qETybuSomI
t/mR6pLFkVknLs38JZOI+K4tiUhsH0Fj2msrZ53Izsn2kycrQUqsxtUqjOECfMOayMpK0V4Sckbr
FujLiD3sEEwNbnyfy7VPphCmysistKjhYiIdJgG4eTzqo3MTrjR8Z+2di9OafY7u6F52E6+dgFnY
fS/PdGn21LvxIryzj0gSCQ/WeYhE8iZax2me7E6mYeF9f1nN7isvCRN/AEhcABw55wSPNJls6YQS
EWp5gN1ISMTL4kmwOI9c2ZVoKEbuyl5trO5DPcWKKYoHW+6d+0+B3GdyKA1JLDhVBhnZJ6EH68Zo
Y/g9eRnYx0+nrtadi1WkFY3qDka5Ou5CSYYSAIZlLE8BzXqhLV8XCXLaqm3FRtuNjTt/ISy6aqTR
IPuoxZh9z1DeByZ+52GqZR4+KUWisG9w0qOohSEs/7PNHGOzgqpXqjwMW28b3n2/gOzKNZLMiZz+
2flDPPZTqCj6jzNN9eZeyYGntukuJvzRquaiaXXg2yjFhE0k0piJ2wORVAsRJtjDET52mXSWXqy0
XGleNv5LXb/HU4kgs85J2kE1Jt3M4kc9h/WetnpprKshibFFQOJJirAghnnUFnpk0ZiSoCjlCNWC
f8jkIl3jgmgfe+RucoeAzcAJMxy8v0IpQdSusui/Ugn91/qLkMW/SprM1RQxSiU8gMEk8veb64W0
4XXyoLQz3M6FTLnHioxVn47+Rs+zYh6sb2iSG/bZPoNZN9ZNw2n70EhgLAnSI71wgicFu+2TbRof
/QhiX40zqCuuRzN/uQDy1J1axm43LXgxinItWlEGO93ad2It1HPtTmJWtwOvxWnfIyS1NcOddlju
8XZsWR/BEq//V1cN4mj3vOwHwtBmTYj4ZshS0l5U/2ZB/vb4RVmyvkh4GSpGbG32XWKU//0AGV2Q
wp+Mck0lAv/VX2q0p7OWlEMbPbIHtoyPMuD1DZ4OVxnuc85aJDg0j4qL7fXAGBHeJWyW0JqauDJW
JWvARsY+WyMiF/1mJaKcaFQl8YT89iDuq1rglGCl59AD5H/rERFnmrfvLA53s0mzkiZV9loVj31Y
riQG1ddxay6QXabumfNLerl2fUpX9vWIhh+9HixxORhf7x/+1ZM9vTNRMW18I2J5zczrUsRl8PYx
6XYn6s1sl0pUgKFi2B7I2RHeCfaVEAHnrJvotpxrCec0tPiIhGYXEmC/ft85EbsTauVjqyQ6chWl
37ILWz9HyDrvwasmBvh5WmeANLQ6zZ2iNEmVRGqlFEwdd7eHVolnHRMJPpYl0ZLpceO7NOspDp56
PD53hAAD+goJFv+xgb5MnIViklE1UHktYTJQ+B+1xOVHjQoEVShC/9zl04PgY7RxmLixYf50TlMr
bwG1xMCo0AnIs2Wa7Vhl9+anAOJqgLc82Xd0ud9p4a14jj3O56/DPRz4h4HALA0f7SAfGYGx8k5S
d1RyTvH8g2Ak/LCYaGGKHwCqJS5ZUoxRzuMB3dN2G1azf9EPOwnb9dzGBj5SlSvFDddrj679Taw7
PYnI98TC/Meiulr8DeXLGxZnRFOJmJnMZp2qNRXKwEogNYhfyYQ8M5JLpRBI0LdVOdnCEf0PjBU7
WChYzBSgzqAOdnYEp3GSyxUB2WfB7zJQVb7xWKiBe4vpHJgs8dEOxPknsTE0nWdLkL9jPvS/jhgt
VvTd+X/o+BKrRA+FTLFngG6++2MTnu8A42P8xiW/6oqJHzvYmY6oKRlY2UHtAezMCRNGWBU9xaPF
yySMNS+zL9wa17G+2FwAmzpR4zbvJYjOHu4oLIGN7Po4nD2OPjurZL1cNbJJBElBEZvoz1t4IoDH
Xr98Suw2r9oIfTU/kJhoMeer4kqUzB4dpVJZYz4gE6pPf4orCy67hKPgfjXe4UtSKYdMRKCw2nXb
mdD3WhIbtWvLTBj68YK0YYN/pgmMFErTSeJd0TSqbppquZA8uWhxiL9R/0os240M5Mpvqj3W0H79
ml1AYEIvnik6bchofPohZnsVXtjXfFSvGuWqiCMSNTjRsG8R14KAU0hFzbIpOC6GsDqlS659B3oU
NPUa3DQx5ITe51gV5p2xg1SZUPZ/Wpra1jMSp/eOoH1xSFM1I9ZCho0W/tcqQ9BxRCtSBqXL1psb
DnwI2ESNNDUe/YnIgIL/sCHxMYxiYpb40+QSERReKLBJQYlNh0jJfgJUtXtVYpG33pXUbRrja+Aw
skMawVLtVVjooWctUiAtrN7JO6GPf5ABPlnkVouKtq1E9PjHP+6moHbtc65IQuAR69H48snhsiy1
2HMB4rcGUE19BZvG9j6l/N/aiAXFKV1fXMQ3NgVbfJsnhyneIe8ZyM5ou0GPrKGRLYp6ZdulKUfH
XCdgi4Jbvvyns5S69e5jrif4bvIVG5Ucn4mtEchRyWS4XZROEibTYWfK0gmHtaOhu2CMrgHpd5Nq
xrjo1TwFdr/eoFcETFLAwEmTJRt13IQ59rxy3vBiLo1gc6I/w1BQcntBbsh628Wu7ZzjVGI2hjZk
IqESNaqWeHw/AyhN/v7AicYIF5ugfCrELpKtEZOb3xhVehcej/FHyHObuGQ23Rq6/hPAL+CJbaeW
Q+ak5EzIGwUJreN9LNNVYGRsHu3JIqpXcwNiZIDMm2kz6FhV6EH3PM9ko7MFSHdAuy7EWdPk4DIz
B1+5wHYbyLb1eS7ogPh/LxzfgHi2PnCuJ97Vd8n6s4SdDAflT+YAE8el2Bk5cFvec/vTqXS4s5aY
8984qbyz4Q0TZUA4+tugWWIZAmQw92ldloj9d5SICSBblr2kHvEL0rSomjifdjdltUBMsELrPFOD
1yKDg1ScKexGDsGU3xEXoGyHy30IbU/DwPiUU7+hBlLOTxeCuMZlksMDSbF74rp0gPwVtvVq34sw
FQy/LJgaA2pHXPkH78Y7lXvNhBHXr5TSbcfYIcAj4cpxZMu06Ta4hPEuQOwfTHxnQMxX0gAJIb0A
UmQoGpOU/5nxaqgeN7mFbUMEgwcD8jdhT9445MfOtG020/DAn9Ad1i8DaYSC/k+6r4FhR5/2bcNe
pBpNxjd+3ZvSg4nB9H9MDPVjAgxLZgTFvNiOUo7PkNog7dKL5hUhhy8KQ4BDDMBUI9s6yBxPB0ec
NCCERa08XgsRO5LZVQfdByEQ9F/RVUcP5iKamjSqb9ztds3/zIzvESwaJdT7BgTI9Fr8SQQWpedY
hP3ttBLvSKXR5nyoyfuRH7LPNHkO1r1xbvrcm0pBzY+WmYsCLdxhlLwtZtwyJ7S+z4qiZueTgsan
27a3cjmx9DNyc1VZF0RgMbKffohiMDRW8MbukkPE0UpCXbTw6KrUDZQpOlI68dUEmsjSXrLQMvgn
/neIEpAkNX2yBETiCdcH+nKr5P2S/g4rc/YXSdE9b4UWPAh8+JHa58rJcLjfNLky82QDUQblTWk/
XXetmyKSgwk/VqvWY6I0DftPgUY9p+r9F0puJ6PVauC7FdRn46oG9Eqe25F2+Yws3jCHsffKryED
jqqrFg5k5+M4iTA4kFnG4Q+XMHi72iK3R5cr3gcHjWwkiIukLHnrqtbcw+t52r15WwDww/CodIOF
i3UCMpWq/vFud7My/LrGUe3A3+GTwjMaVdY5JkYv+KKWbHM1l4diUTbGhtdPKmaDTiUCBPCUq1Tz
ZaO6IGvDv46tPAvi50RBd/A3aePp8DUb45k6Qk9fWt4DTEfaqMhfv/g9GwhQ9rlR9mCws28CrBoB
MEmaT70Nzs98jo4+Go8D4kBKZm1e7Nj1MPnL5417BwIDK579lQkFtuK3pX9MLjYIDq/DFjPvJ08/
AOxwCIHxxiOE/tKh9kfxfx0H7c+6cLnlSsh6Q2FDtKVN3nhvNHj+0u97xT8y4e7erHhzcWtThyQY
vzXy6cmOK9+6lS9hG4z/GRP8bnYezePjtzQnlht39kuAPqZQEOkATsBYZsNOcPYkU3AjSxzSgmen
xt+so2lbMx+ExBklUapsYWnJMu/QPUFTaAyveEB4hyBTXTms3NGjkvSejxRI71LVBysDdsAV0jFb
LVqxZ/ecD5ogcGfVunWr9O5BzeTzBgh3LpQHZaKrOAODC9VZvDgoe1a5C1py+UYYBhsJJduAP7bf
dhZAxhUrP+UPx6J9xOrhH6a+t1l3WdkbrbiLgBjMa9JNe/waLVkMfxyEXxkf3o5qRRhKe26oq4Vx
fCmZT3I1y6JpQ+E3JR+dhcw4M+ZAXfZHKInuum6SlsXV9mCTcl2VOI7QY30QAV33NkR6QIcj6W05
7j35vlneQX63sgvSS5wkokT9TNF4E743zGAJ+2pBv9vhEFw787U0+P5qMlVNYtV0Zmp9tcZgohdG
eug+zdXKdQ4/bSbho+PFeroHXHHtMKIfhglfCLBY1mKjREKlQwj3FQDBNpWG8ipcnt1PQCL0qRP9
LRYjeYE3kwn6EPpbwUe6SZuWudgjsZ8lTcd9Hed3RoJOwLnxXYPEEDlnm6QaLsFW/AT7S4bjlgS7
4Uw/IgvWayiohRFEXpgDijzwQYWYOdQnXhIDSHB9k6kqQsJqHkJSiERwzin0RP4rtqN8mQyEcTgy
NuH/B2Bab0ZAB1seSh0kYK/fOiu2jioumTaa8xoc6wzrDzTZcAhPPVIiHceBvvi/cD4PylQ/8nv5
ADMd4wbISuanWvmsrPh3QAODPKYkLum+RcvjMoJx7eIyUk+Vb8fQurr0ZBZrwwUED+6zX+yw9nY6
Uqby9fFg+UmOdY7eaHA4+8CykbZRuXrC5iB9E+P6Az5iTJfAeo5bOygWEnbl7HiKsXXzEDrK4hri
6lhw0v4gtH/nqpB6+su3vJWBOim/ESGENJkxpLiR5jvMqbS0lQeDDiVnpzaDpTJH3vR3ZBaSOlsl
TWQ/W3KuNnb/7FE3+oFpXI/2UBsMmlYo8a7JG9wCezN0MAjApphEMbHxzg0PiMiGupTR1U6ocitb
KpZPst4hvqx6/dZcD6EfS7OgiO+mmRckPLebef7IH4TaZ9CzfyCEVjeEd65lrWxp6NSs90sCjzhU
LZQMdWE2RJiYu/rffwZkfUuG+gDhYqkMD53xpzUQc2+F56JIjgfd1/8lQaGMNG/8mD1wT+CyjRmO
KJOjhBiaFPbmFxPp1YkE1+uI90yulfCrICR4wEeV8GShDSE9h0drIp8OLjMESYjO0sUaH4CRbvoH
CrPT29drfHvOnYIAPeg9fpUDjgMth+HpVG5pk5t/P9dES6A5ER2wuDK9Q0sXNF2/jz+Ihoh6zUbu
jNgdY77uHrBRsCPyYEc2HtbK1Cv7fiRkGNP+nTtWSBhjNAWeZvppwDOjClNgkauehNXHI2XEQQKM
jBggJ5Xr6jtfock+XUNEkirT8ZOHP8U1F5vIf6Pzl/f6krvm/y8+MK7eWHeJrN4U3Q2YYIcTPV9J
cdoAoN3eVIwXa02B3NMbkHN2863CeWhUA9VBib6YEf69VTfCbfMn1zcdd2dxQiAkXQ4E/f/MknPt
Sh8tZob0qiLvpVHLGJqk/MHfeVkvQN3A6T4GbLCujmgXSRS+jaHRpwwCbrk4pg2ObmT7p1MJVmBY
r2bGiLIiWHIJiJkVw7PhiaIzCQbTU2FTyhi1M/+3HS5Y08CePxkETF/SM1EEXIik5qXmyY5lfKs4
bA6xa6USxy4Sn4Yj7vDQhUih4CGgtEoD+lHL2cWd20eOjKPx1E5J9JOfSAw9mFWIdM2YZVWhBbjl
Nk0vQQbYfOBXzN8mjy1KPGedL7wLV4KmtkWDHg6ed9U8Ds6bUAaK5PBwRNIn4eB0pOK43YZCLtRh
z09Qtb47ERIAETxcbaAFH6VzaEVAHuV1QqWWWNFGd7N9hnMZUJFlfWsfEDKAEGhi6ByKes733NTj
1JmzntQgcxhDPqHy19hhKavq9PrVhvScQejvqpW2RL/pXWvevQ/jV1bWdA2140P6N46nCBlnuduo
8C8oxYAiyry6aWxtmVjluj2lag3Q9rFFbOQG1OH5hfpUa+dAfcBbj0RJ83OTELbOfgwXlRTmQLXl
ZekOM3mL1KZ2Aj/5kld9CBLpcaDI1Dzwrelw8LkqYCWIggYi2p8F3qmHviXCKpW3t990KWAj+j33
UfuViAGCcUXcEE0on4EGsmOGfw74mbQW2YnTbifFKx2zlwxJiqD9BFsxlLYmMK9YEOq6PhNMlNvJ
nShmmrF1FpNumC2dx2xF+IBIHxPqDYwqZuB7Mk4NPNV9zBS61ruaSNqzrOPdcy2EzumSIrmvVuP7
v/HmAxozsoXH+Iosvi7ae9+l/9z/OWx0xS0/282EsaRBA0rPq8sbwKNshoCFL2pwrEeV4yV2NGJR
lSn/m2gpdzAsJr5Z5K73kYDLbGzttQHGlMWatR1V/zxHrRZU1AHO7r5GqHzs6jO7ArlBCWW+ar/x
JWrbZoTB510ZyZc6a1zZKT68IpW9CEtjB7R5d61vJeVP9SsSZptRfxxR5hzA/6yTIGjeYPVRgWjg
/C7ChWGcaGtY07dtmN5DRvgaFEoC1ToaIssLegLfGGVlvqhWkVQRGoPAinAAjwIQZJDbLDgegf7+
fP2y3WGlE90/E3S9CU68VpPWrEY/9O82xAJzdxYqqdlb62Bd95Oq/2+Xuh3C3je5BR/qxJs7KYTs
1f34Ld05SIWh5E14CRo3k9WVKO/OYtILNTuV29TliIM4IR7iUQbeDg0CFJzIY8hA7doNDg9m7seR
LkGcIH9vuHBMVwEdaOSlTIuTIvJ5qjCDlSWmvVpF7ldtoLu4+BsBBd3vPzoEgK6yj8yfMuyC+pTW
Vf0QCi9/Nvia9RNfOxgORWENAXHZGUhtoUMLhT97p7WNjKUF6WOCeMPRz4+zQNbNg2kks3yAdPVG
ofUmLhmf9UyewVV7F28E67FSI6xKWh2f1w2sAclJR5t3+LbaCrTXpE9cuYqkS9AaaCwqlo+wAtGt
bL52ZaW2xFo0Lha27CNhGWXdtMJHao6ebmeovPhO4RE4gA5+HP5n+hofPh90VFEgfFAue/Y30TjD
7z0wWK3rmC0XY1FfXtAbhuTilPoZd/umE3LpevivlJAUE3qSoaob1do8pllMyZ1x/tIQ+8mZWjfq
K2jleh24rGyBJQ6ZH1jePk405v/Y1sly68oA8LBO5kAhK8RpK9g2jjsYYQJJOCAYvf0X39GYX1Z1
lfrXXkKk7raAUqdqH0nsQ0u+ieRo4DC7a5rzhFnGai2K1frlY0/HxgrdWMKeef6B7Ic8Vrh7m4ow
9PY5NCPrj0m7Ysx1/3t0l3c5koVQd80+QtgKbKFRmsrg0nMKmqAOsIvMC+2X8BoyixYD034/pU4A
5qX0XL4n6P18+HIgxrUy87fqD8Z2vNCaJnySMFtnktZQ195GO2qV6Sa/LJA+0dK2X+VdVcJpuAmH
Dmi7ThCv8dk7LcMP1TiNMxH+TuN+tW7KuvC2tHo9dy12Fp9ByIKtGWFs3GhQSIjKsmT9HS9VVKC9
yc8Ho2rfwOLjcjA+Dksv1P/3qp7hFA4uw9cQu9/zJu81VOjMQPYQuKyquc1ndGWzs+3HuFBcYsZc
VvbC0wmQ+1vnWZpsja1Vvxv4Dc90AoVKfVDrz/eUb5aFX+CdHSp02QOLN3xsjmOKsCEwTLkQsp6G
gunGme4nL0/jci9WRcXdZ2GPMzEOTK9kUVEIuY0vud5rNvOsIf64WAYato3k6+Bpa+narydHm2oY
GyK9eX3mAYnkJOo46n3wJB4LwJlvqsPgFRgnAqhsDCR71E26wQkpXpdzi65kc4RdSRRGVrsX5skp
5UXWC0E1BenX0NmWtVMr+B+oo1W3zGQKyQ1zqwaZ5NtTQvPsp5ByIOKm8XduIpeW2VhsP/EWvc6a
YeOY7Siw+7YSWhnuC2fWZzISdaOd2SLeLvXvRzEqRG+xj9PqKrUaZTvFWbkv8F1n/o/G1USMndYV
eC9ahS+Jo3C+KMlTSvBxQxuvPRL9k5TNOwfNDb/UdAgrBzJWZcfm/SnuKMnzbum7jNRHsQdGatAC
OGYKlTBc498vg12uPftR4vO+OTkMNieLKq2LHqzYsyg5MTH+8MeX+FMnYXQvoLn6tsyFtSVxdM2m
f/Hmv+678gR24zVFn6YLqA53hZK4/BDw5IBCDEZOup9sj8E5t9GLzsd85uSz4ye1278YLIMWtB+o
WHh2jMyPjPOQrD5T6ecPp8mq/6wnqrb0jfxcPi7dda2SnaUUfmqR3hToc0CQ11C0LDvNgChUS+Ae
yysWQ/jAC5A0NGFal2f6xGkrHNLZpdz+3ExY4uyu59h+4mNCtxZqKYHOgyjSsuUtpy6AFqT8Zw4L
yT9DY756hJybxP/SjgTY9ZhovOyk5RzThoT8XGR9ctgZhiH4ZjOYUFCDOhYVQ9sgSqlxxseXGF+v
AqY5jElrN/PkKD/4irS7ypQUrw8+cA7qgb7c+8TarNntouwPJFDj2j+22O9L50tgpDE/EETpzEwz
XZiW5smAeMZZQFNfXJdzkqYblNNmpOwYUerNr1f52YbtovTA87YkAo5T7TY8X5YFliLJXpoQ9qmH
gB4h9olTsZOM8c7N2QnXNtAcAmjGdB+P+N+xMWeovRKODlOZILTlFlorMVlSXly8JzlDOj8ps22k
x5bIbvkWWrYaKlNyn8vqeIxiwfQ4Akk/02yqn/bu27Gi4gEXk5k9j5yl9LHYi3vWpPEy+xTt8Pd4
7n2eXb4RE0N9/wv7xtnJ9goPHdFlImFELmn6j5PiMlrwPVeZS1sdLmslNJghzSG4TUb0Juw6nXdE
pzwdVWLoj5J2ws7PsK7w+SEDB7x8oXicWGKj9+VZ04Bt3OegPgg9mbrmZ+JXp0R9O5X5K5xdoPFj
CmDK0BvAPU6jxrUPe1C+xf0Z73Dtum9nyGJvOwbbjVymkjQVfyynzziGhs5aBD/EVo9wKT9OAdXl
RyK+ydjiG3al66kuZ2DYfIat0UKWflwREN7FtiMz/7TBTGEfQjaUHA6l0BcCKusApZBrrQK3z2Hu
0x1Qp/jfcbEu/XzZbUaiICmSpjQx2+lkykwtFq+uxN6LOB9+xCBfXiDikk20ssyPiYlyy1B5U4HZ
tQX40rhmEhr4fonn9xcA1W7WtKk1WKTyaTA1tDeMySQEtVteGOzvVrq8i4UQxmubKv0RU5PmHVGB
d6ctAzMKiXUg8nZMbJxKFs54yqYsMqCPFPkWwDtYEpz8317rmB7SYymuwdK73Vw1Sc1HM7O67Sdh
BejPzdFc3riKRq85lTuzdiFz9REhTpQlFMv+3CfVew2bNS6XK4RSuIaLepkXUK3T2Qee0MfycDIO
zMuByR9dGFEUq55uZjTwBGSpijWwfvP9n3gMQDNKaYMlfLoPAM1Wst+48ajbLAe+Ih8RswLvKpjU
rtORLbN9e+GFTSHLuETre+zVSnXN2s23sCtn5n0am5q3DMzSQpFXtwRCvVz/lVRY8avXm6KrJLIw
A6e/wvGN45eL0JHp8jVX1CQSL2hkNYEF80/VOAFO2tCS0Akal7swfaek6fBIscOCXbOCMK42Pn+s
YfuzwacBGiyBztFd/bOwqre6VYSGnhjrIswP6Vr/zHZlnMXejPs5CTSSF1P7gFiiqUdFrFoYnzXA
KRJysmvLylLTxL/jdFsThWqcB+TwvFgbHKczBg5QkkiDF1XBa0Vkv+dJuCU9AdSLrCpJ7IWRE/rO
dFottiaWn/ARGEyugVovTPqeYsR+pyqTgJ9TZ0E4p14rZ82ywqRoPNdOujektTiL+EW3o2O/E1c1
me1ZDu7zzpCYkT2ZQ9qydY43cE4/6PytIO6zyuB8Yba3B/yqR7t9KhRX9QkHTeCUuTNZ7jQEahG8
eVoROExLhR1IAQo74wi4ijWRhTyzXImINCAVyJnbaHXZd2EXtzKBY7uWZ3+CcsbFPKoOMZYADN4u
v2d/7r+e7QZPEcJcYBHTASetK75hVN7/fCadjJ55h9j91RnMjw06MsHTwEOE3tHKS3Wt7E9xo6Wr
YOn7keVrqeGAYT+G84IZDAD3peiXUM1cKfTukDht+Y8t+ZV+78y2Wl4E6DUrIzg4HSlOKyO/1seO
qPngJuYzZhtsVlYJiWbzWOrNdmvTL7eXl4Eqo/nV7B+37YFg0lOdgodRgAmg8xGybHDRz/BD7Zf8
alkrYxNvOdFEkqVLXutqLC4Zxr9paDzqumvzMB1opIDx5PfKrn4otfxNB5FIKx/HQ+PoQ/QZzURo
fE4GuS5Om+1H0mjkPrh0AY6ONqqYjYIWn68pZs8MfyHYRIB4c5EfV0GMkQPStbKflcNLooYEJEO5
NBnd3ITnTNF0SP0owAq8SvAhU7Gh2yV1RoV3g9x3QK083RNxzP3yilmwjj6k+ggHLHANf7T3JPp5
R82PFBiDeIgI4P9ai86uGRb9ZnHrPXACrIbGd/V2tdHFbXO+gJOiQIqOvTMiiPEEJg0iXlEAzIqr
xwTaE6AjJMpOIlfRChKRDaponALAx1m/xN+0CDlwSLbIVq1jBeSp66qWfYC6qXezVuyBqav2XHAF
uhwssFG8USMSWIPnbi4lATIgYlXiVHg4c8t4IkGyVuqdrBJLdg+hRaKcSdGXyZ/6SEhBqR3N8215
UnyrCyBx1mdX7tbHDcYEj+cUjrPqTQF2wrcfJYygN9kNM41hqxbIDp184WiCud6ywF2AY6DmEciH
Eg57287mcv96At93pqFDR3iQAC9JHAzF3rK6wlIJuQxf0wreXcNNat3EVrWiqNwptt2NncYqkaH+
ScpGkMtA5zVUU3kSwUp8zGlxr9dfCwxID537b9ZmRnSG3NnS3DtSS5k6H1rv9NT23kWUZwCoeGcn
QJMCLO06cENh+j/Iqt0QkZ2CWui8K9t/HtXd68kCbs6zTT6TRHeJFHVas+av/LNj77f19HiXba7f
tUbCasXrguMjE2w364NeL2WJNPAdCO7qflEjoVAcUkJ/Lh6+pgD7cfFDaDI8UjtT+LHhCyDHI3ZZ
nV+DV+t6RSRbh/mFWS97xSDv/w8YiZpziFz3GMrjaAbDLV9C9x7S3vvMXSzTqQ42WlC1lGnQJxFu
tDXH4jJg65c+bQRTWx4emDGiOZSkFCFO9ugAwQe8inkW9sRsG9aHvyYJUqpgrUsy+8AOY2cWFLPG
KXPs6NNGGAujgoxYZnW+wIphOgLUp4yi1+Q+xQPpy820Uvrd4q5BcpI67noBYgUC9ZDIR2FclWkV
wXdhKDENDgJDbM8X6bECvi5O6lJ0g2cXcUdJsLJvHkMTux9NoxeXO71Acxpp+tYFE957UG/DA9WE
NmKXoX02efSCbiSF4HCK1N9cw4XSU9osHevsL780/H7WlJf9PFygT7lPPrqrcFA0lfxJI6e0gzyu
Q3/mypOHF/n9tSJV+JqqkMPthg7IJgJd3ZfHthUcYaeRZY6vecrP2nXtlA9wjnRGGQsnqqojFY4Q
FVTIkYHFI0ajvBA4gK6prww2TrYknYy1iydBHNjJNUe4b2wWBUWorzlCrl7RSIKLCZO0LTrNY06o
kqocYB2CS4oBXwtnEg4+2aSrQoZ9Vg+RilH6MPsGGz3/1oTTWeWOFo2JuDP2ScYkCtIghejCI2pq
PALaapn0HDQAijXGWmM0RYBL/guXXj38Zte2Eh+BbiZ+AZno/Ue1s/yTzVXHhMkVNEDpZxC9wVef
M+mN/SKJ2H10p3iGtBQCkitfrXQh5qWMZThhuAXgz/DXR94ev5ngf2NxscPUhF5Pe7DIYgLzFGbC
n58+gYtq5R6UiYZYwgrxS7aTQn0x9uosRDjfurGlHxLTZEv0XI/+2W9FAzBMiR7CVbNuCSP38lOO
wojGIO4e1WfzT7gR73Kv7Tngv/zI4QNDjiyQn5g6hzYnrnMSa5sngyu4oTleqv7jeB9njvjaNFuT
ghKVMnzyiHTDLLWAa/aKB/DYpaNc9xsDr5k9M41S+N/0DFGaSz7B4YsmUonHk9XkF+vr7BefrPMo
CviBSb3tAfYu3ZH28PX8vQEJ0nLLCePdGA0E9dqtn1AhYY8vwMxWk2luCbjau7EYQ+HB5DOSDDex
r0NruNOago+gIW4j9FTmMznDClkcmtMVnW3MHA5sormPLPnCowXjpnKnUckzCjLF14XkX5n/3qdu
CAZEyxUoxUofKOq+/S/gtEwgBFCSJVqhRYOyVyS9kDXfqMTLLyIuXbqI8IWtw09CkVwAs9DB37wd
nnrNxul8YtpL+ps2xkKIF58ow+TwAXEEP1GyvpcAHCJLIuw6jH21f/QVmLbKtUtzWuJUBsdSSaJO
ur9hHaDQKrJ6MMS0YaDNPb0YfdDPQQ9OKgmc49bpzIPYXFRyfyV+ahus6SN26e1cW7b29jljrOzk
+ues2mQS5akSty2BZDQvIIs9OYLmie3M642K1ouUXQKq1VmXdGKvsPabTrwBVGrQHYGWuRx0kwzH
uxA5JTxtQJGehkb1aVejYzBBKeJe74GXUkcUmKr0nKw/j3nXUr7ovUfFvnfRwWCVTBsx45g6FXdH
dYSrV5mk7n3yQ124EQjAw9X+KHETj3FdSkUruqABnAedErxpgz/jY98vPIB/q7z3XqvdOXzhXumU
RY9RCMiGcOFdMg7LujYDZ2o8wedme2X3muLmL+LniwN/zGE6naMEYB8g/sPJK68CZCl2bBh1FR+N
S81JrYIXIoHbevgv1xH5c5ybknWBzfnFSm61hjQPGyjEC4iOnZeddoDSC3uFz3bOJYnyz8xcWUZm
FkFILyPRu80ipzUYcUXD4IypvjDPhK/VQ2yVSIIQgZRMd1rIU+ho0d7+3fhoAdTUet1ElzAq0rcu
zrgCUjoApOr/D9qrtsS6k0u8yisbyWPebxsuCMijsYuZ4O4zfkQ5/CQzqsXxjEf8uUMkRtols1IY
/GwE8QHh9sjvRWPFSVSkpzXuJaJY8ENKxe4n7P/3W8XDL0YSKyrKhQu+uab5akLAbdqXEOnA95w0
98d3YyJ3MaJ6mqIkGjOA+s+FT3bRIomrhuXEc4QpZ3SWF43ddbMug2quF+XqLuvv6tJz10OCtPj9
WNI8/BHusgOmGeRYeruaYAMRfbP6OkBIAIRmfKGnjryyI0ZFPOzDfJQV4KQAnGUuVWHCGBmQhlIv
q9OTBkwbR0jwj5tcFBcOveXkT4ZcferkbxaYOC7ugya3jAYpPcCK2Fw/gL7vrgiKLh1ecSF8Zvur
KP+Pf+WIzvk/rzFJDZBw5hlCAJnJDBxa7VIV75GuCtUmMKqNnbzmz8yCjXgpVgxSQ5hTtEkGHDp8
xniKQWSmpFmAV+YWUJkOZOzNX6sihBFQNty753TdaWJMyEeY8gAqr1QDR5SF8X/TqGjL5CNzTFin
c7Ks4XgNWK2DHLk849zErICHIdjPbygj2KqYEKAxmtGxQDo54R+0qII7VVt6XPcjtmkrxSrgMupv
Ufx/wPok6T+wKaC14qDYbBUns0qk3cYWFdevhMevl94Ik5NxHZehBoQPD53k5eClNBzpEs9gsSgL
pCK+CLKcXF3YVNn99TQ3hT0Cv5JJ1od3kOEv2QNo4atz+nPcHHCJ3mejtqbT5v7MRYX7JLAFTl8z
69f93KBIgdBKqPqYsdzPUH/hZeBV39vqkgFxpRBcsd/4Lcpnlze8JHrNrjL735a0vj03Ayun5pfr
hY1Zmo+eZus8dFaPGoFUbPR1tgVAdfHw1j7wvz7Ewb8urlGd5aFum//gmerY/SS+/AGtHeW3fwCk
sKKWk0eIKqq8Agejw/bGSYvp4M40y9Nz/aiGC3Jsa9g/odmH9Qsn/dM2HwL37BH/r2UYBfw6JUCX
i0gu5rWPzq4tWmdHJ2vRUQrVa08TU39NeDvmSQeUHxFidf/dN+JZ3Ya1yTj3SyVWg3SgwwXPOfOE
pro7sHQ2+bb09nkP06ZwxBen4fRrLjkMOo5hcqMD/kdc9FJkf1MpQ/vAjQtPLa708Fg51yFxLnKH
gwc45rihJ5FW7W75TAuc0zXADxN8taF1X2PZGgmr2FBzT5+QWs82yaMqA2eOtFiJpaffFtoSGNeJ
3Rb+YcUhRFBMvOpejM0RJGP4WQxWXaf0Y5GkFcRu7NgGURQ+7gfy+O2cO1gRFU7Nl6Xq2SXkqwLe
n0MJlygxu+9zF7gg0WBMcQ/qqy/qIZ82eLAX6mEGJ4XONYG7mPqz7w3n7rl/NhechqprFVCE6+O+
uLYcL8cfswX2CDY3WGZMeBQjg8dLkwEMW53eelbnzRZk52Zg4ruWafighSNj63gMFeGJCGnNpWOI
dhzneA2/7bZnlw+LzPoiN9rQDFVY8kmfJy+HmIfS8p2qYuAQ6i5guIel/lc/SombVy1Z1yj/299G
6HOIpLOpLL4RPaUD/LeUTyttB828EeK3HgnCNuHWpji8qjp3SjLqI8R4//nk9r7Jln3hnesg6BTi
8HVCXu4qyqvPBB1Z7eAOxFvJGaW37ioz71ABhORwsMDIbSfKPd/63CUx3LK/bGu934ufWdTUxAw6
RlQRNWagobTVLR3aSnzwDRw659E6rTQhREjQI36dFLf/NyvT+d7dl55TlsXgnvNyWnqbECv1o3fu
MRZ+rjC+bo3zEvV+yLx73fiJwVXIcUug5S9/ND7P4kL8dE3FmtndPYMF5ATekvgPRABfjUgByrkn
wYx3TCDLUOEHypYxWz4CWyB13n8vlajHw19EBKoUHM3D9A0U9A3u2/+aNLPtGev0qsI1uR1bACOy
p/U1wbQAgRDHmTvAn5lyPlGCFI2Zv1V/p6Ew5ilJ9vncVTLWoKbPEpZB71K3UMoSkmqJlNbOFu89
aiCBBk/kf/pnTpJMi5RBVgUE+BT5xtwj7CZhXbwGIlVnvlQJ9ALzs8oQZukfhxq1COmK6gD71pk0
/SpO/oWMx7h43VYcKHMqCwMDqbmi1xUzCqHLPHKVUuBE4Jp+vHn9fKT96SQRNWAB/ViY3Y3GI9Y+
TChQWhzAsvlcYJYFEiHnUZHbJbi+h+TvH18AF017uEo9NCic4hUx4SIDhBQZJG5va4mi17pvETJt
YE4bLlE1w/mWHWnzJ4KR1IPl1qaSzwVWI7pL+EmfRorG1fnWiyexHQ56G9d3GcKC58la9Wh0h9wU
WzLcK6akdeheTKOS9USJxpG3sPaTty2uPfaAIaMtHlKGIvkD6EwpAjvkp7Zr5ni+bu+kilJ/B590
nghLDsmX5he/lTzfW5KZleUieLjoy7LwyEIR0uA/H2FaErBr+LUt0lweoxgzXKhBRwxYSIVFZ+6X
xeriYTv5uxFYc+7N2DL5Gze8bThQfLJjwks5Je9qScgYw2SOkgoKBwn716vxlAAVEWXclouTG2bK
va1IDb1ZIkzXmAfZZlpHArEONgTumHmIV2hr1IdJq9GGrCZbM6pNjt0mklz3ayG4eAikVn88LV+H
hmQZBBvLN4i77gyNYj/54UbCEaFZmuTrhhsa2/9DEbNu92a8nR6CsWovW3qZLrwecxHFqWTT5pPX
9RZP093J8bjqDkTb/LZFX86SSnPC6s2bRlNDot7Gz3CanZpey54tNJ7VGaDL4FYgp7RCqJQj761h
UWJG+yQJYGFgc7neVCM9rJ3le+2DPXSFY8IB8dOfcQFNJGuSeiDrAU4YxWVdKwuzESB0QaqVtG7D
q/upMrCefbHxX4fEWdrfNvwD3RP1gQBpULFKVOCbZcmvX7j7MIowMEUzYxnAsvUgR2Y3ZhIXKRta
oZEAg1kLZWYJGION8JKWkV4rd/AxxIP5/GwbL+OhcQlYqm66SGvciPGtb1vokVndf1769Rk8bqxH
IbFks2s0qxH3WjTijXLTymZYUZVDYZNZdDn96pujCc4wK197aZitCfgBzjhrmPwXUvBr+kp+NAVL
m6lvvOuz/VzWSClABIBuPsDCf2B3HUNfaf0NxBBLZqDnElhPwKJ6x1zWjYvHFAVg0HfJFFMcp15Y
/Lufze4TZ7QEhxQ53OuFyO+9AG6fqP3p2bfkZKUVXImJW6VwyYYMpY924XpQa3kyIvP05hI6W8tQ
NYAMl2WGi80yononFYpJr3ENHTuc4idklnrbO4ErAeyZp3zqmVZQSvC9zhkFix/SSiqZwy4BTZix
sj6xVr1lYi39ajruKp2a8nx7+ZcokFtNwRkV+JbyhPTt7R/v94SnehJN9LAdtH/lRHhfuAvcAjKJ
iilSitPkO9U1VRzzeS5UTAohvkSG2QOoohomtaSX5tnCp4dMKshk12dbbhjJE/BCzBSruJ6VFUtK
qH6lxk5PDn8G5kn/nS3nXLNq95HlVQBuTUOYNRvZSaPWEwC9tUbCCBD/Ylw2xBiYzdlVAT5OA94Z
NJ7BBr7DXmHZtqVehbchaZnLs2LQFVJxsgJoqoGo4u1qSP3AESQYCaForUWKJzYivv3w5+Uni7gc
q9DbSUFkM/gFpkaFrK6npzdN7PkhrAH/JaJRAW6nknv6lp6C9CSRJvWHBHEhwjY+LAiQK0AObeCJ
GjNggmhe5c+kwYPUWIu4iGqTjl+u7/yv0lrloUFd685VE/QrHWYorL1rklCdR9fojpHy+gQIu8Yx
YgfcotoYzWSWUU3rbqmJTV+xcjmgeSSYkFW7bANhqM9lvhvIQRjtcKykFU94EZSp5O00sPWb4gwY
2lWBHAA5BFyAiUPw5ps9/wiNXp+Oo17/3lEztGB8V1Q77dUh8eViCPNlxN1FFJuyJAIxhzAOeh95
NFcH6fpZmTLc3w/8JieAc0ihJBWv5UjOJYiUvdanFqcgzDtUUzKmoK7hLklznaPEbJ1LDpzDe3Az
c5XqkSr49WTEEAZlh+IWvP4ORKguNpGNCghP4w1rUNKRKU6uoCK6XS4b2BFlTVA++oscNshjByFa
65kRUBQK/vB3pcixrbsW+GqX6hJlG2x6153bLiH+8OeeRfaCT+g/uyLT2iefzEjs5WM0D+2uhk/3
F6XyzCgq3sNx3ruhHuLnd/LLwKOWFgvI2xV/6yfUTHrsQUMQLiqZYF1UL1xcyUmXESCGpGjbpe6a
Wiktp+jQ97H4S2KqiY0QMS+sM7rM13cD4hCkWMjZyGi+0luS75I8WxyUhyKnR+7quNRiVrHQKqCA
cO+48hKByr1CaPWG1NKj9l6ANRJSPLmSZmrSGczk/vqhIiCUOnEkKF254BUlzJDTbroNlCcDoLVe
C97VxELFEu5/1ebLrtkw3N4xtwvmPvRadWtfwg+Lj61xG6i7wfbqm24iqv6mJ/wKJaCIupwDIj6Q
CwqBfXIhGFMgPNgM3pfAFkKuzl/QCt8UBLEbPUuuHWwQvmIr+1Ul45LovFQoe0doAMi2FIs8ZtsD
mf691kDH4adYuKiqkQYfkyS0p3B4C4fmY+UHT96DlzwjbPlvap+oWt3juZiZEMD6+Fuy9KLiHvda
Szrqm15PlKxlvCZlxCouKLU2TJKLt88fWuqrLKNrU9M1WFvIxUnGlw8K5ppaGFj23OAwy0LX2JFa
hYdxnF29JWRP7dxswHxt+INEHDjA89+Pmeq/j7o6lGF3lMJdgCqwSaaLXOF5A4L31eqMUZKgPIaR
gtg3GUyrG7x9qpk5cNMcLRKk+yG+GcUh6oTpLq2wea1KUYn9ye1fe3NmxvR4n5PiBLbktrBfwbXQ
CxyYRqAj7l64miyz6OIOfWQ4/3/5X6wGNK0m+l2KnkJ5m55UJ81Gu6lJ8YURqjLZUms86Q41javk
rKWpt3Edb19mQkCrbsFNr/VYyF3mGFCiTEOx1GNj22uEmD71UhYPPYHsRBHOyVx6hS0JGvtIE8ud
qFaEa4Hg20SiRO8yt1C8Z4wDKr3easSwb69Ix/lFx24KBpLSLE7b8Q588i3K3uni1Tcj99UvNjQo
94C1OxB4AhB8/ORWTeKZZpYaCTkzhSMpmaR3VD4zQ3Ds74zhvZ5dfq6Rfhc9d8giELaxKWZWYqw+
wSiFOshiYdGwjfwnjw78c2E8ArwM+NaoZq21HcwpKaojT3RrgQvNIImSuRDdMduTLqAbA28nY1WP
M/raPKCRzNq2jWDPfQGS31VG0V4Yaxko+x2ENBcaXcnvknP9rDMz9optJp1yk7ZMwNeVXBeqvCfa
021naxUmtx43UjyUWo6BKrBMpNz7026CK/wVEAAxGIHW6imWmhGM0QM6ATwztS+2lp8aqlWK0srQ
ANdLedYhmSFQmoS8YPLftC3oiNbeXMbv5FjgE4vy1OoXy7apsITb6LAidhoVKFLb2azmpMV8XnC8
mvzKxf+OPEqzwzXGk9dAa529f5M9Htl7hXxD+waAj5PHbxgcpzfm7oaLzR1gQAs4hd/UlgNZb8cg
zLT9bbjUvtrfALfQ3/+3D2hIHqQ4uAhC0frQMzBcsYAVtFu0u8RYdU0V1WZD2wU6kBtOZ5dVCgrc
8LRtUPz4ygU9lfQGKwz35jk3WIAYlyLhBYr+AUQ203kUnr9AsIFUN/ZzTzw3p4BDQPWDiwVhbHyC
vfPl67QZFIxjqPFfW6SO8rjc1CcNmnSb/uCw6RIQcn+sdcxrJXvBalx5gPrlEbqaJQdWkwhXMNeu
pWzA05Nyg4HzT1Xh2HFLlK5ONXNRvOCheE8ofbtMvrSQgQmMJq9PQFIAXLiidZF7nNR6qXXfySRh
tEWpS3W2CzZKQkUd4IFWYE0F7s1s/fUHwrD3+xiYaEN6XmVKhcdgQ1qHAUdjDMC7OSAHhQAhEUxv
YD9VEb/8Bq46d9IXoaowvp6fj/VaQuWg8MoexrPLzLow2ZRrwFavxaP024KMRxU2qrYRGcZBwvbG
DFfrd0JQnNbbiXQCKCufq29Atf7Bak3guDkicVkr47xQb27+igi28CyxMJlfqXmUXPeCcGMZbCnM
IJVdPYh8gjJ/7ua0eNDgK3TfMjiufRzyMllyZmJB1I/Ulg06wgZ3AUsIhxs6evQslhizaOzR+ZU1
OpIXzOsQi75a8sR4sAYXyVtO0OW2WsG3zy9wR4UF9DlbSsWw6aPKP5ESFvxG+a0nvRE+9uAfc+d0
5GWvpewIatMk4EuigZrQZ3DT22StQHzlUBVVVBE2Zzc20pGsbFWn6j/x6mPF3xQYPz65bKgvDiNO
TZjEok+MDvBWGVRwKp8bvMKish/H8iAsIwDwdit0BlMPFNnnDKE386MBoedpNNTwdUlOonBbI0hN
nRMjhCoxDoixJx6Gz2RJwcc3pFcPimKXYpojioepHpn0rBZ4gfioNRukl44CbgR+JDgS+JDbcD81
1de4jORcMSI7y8sMWI7RcVtWl90OrLOfMfj1A3eToryTq29WTJhjL9aYe78puv5+yQ1/qZxBAJoJ
9VAHLYpM8JZDXQ5PdG2y3LnqqyHLY90ZtjJrCg9N4QHkWDyyAgoCoMsyyOncaIl/C9a6hQXhs03V
lC0/AKoQqEe1UryC3aam/Kuhp0mg9700A/FskReo+RJDLK3iqN47MdzmsiTrt/3xNpOoa0dgIDO0
TNyGuAaipQ5aa2CxqYix0XZK5c56pmQF5r5LopDUh0aMrYA2jgV+b9IreeCwACjpbDPeCsCgfDLh
hZBGqT4nPaYJj74iNfmLHEpcjkBfFLNPAAx5VArfZmTJnixMCzepWDcOYC/nm4RhgjxVBjrRo7rh
2OefWk5aPb3gbq39NV96uoRosVl4rOqLMoYFMcqv9cXRJb7vX0zcdDVz/eOpwHp8mPLA3srUB1f8
2oaaZH97xWjOh5BnIO7Sb2YpkD4rsA+UsRP1bIaIz/wNiN+4Qjvq8WfxPlGQ9CqTuOlA3uTmBNIF
u+Su9b97Ux/g+ZWLluSai7eBAcOewwWkXNlmqzsrYmw+aSXAsfY2PgR4xXwZ7NRIY/76CWG4JxbD
HbP9EVGaKzcRvf7ly1CL+qs0emZBTc98TcbGVY8EPrzTka8mX618wrL6sXcTp+13ma15S4wenF52
MXEZSU/CPgAttaiLRfBE7mp0AAVJXc3i70o7pmMTV2rMfD/9ljE2tkxWqysfe++oomAqUBYYYin8
FNeBUkX3Vct2/JyQjbvUnZCXxIh/3On87MuUgZt1JGu1VXyViResjUZJMUSgZ1UNh6Gh8tVVG2So
R/H/SC0JhEAWe347mCDbVdeq+G/HYuojIXXxaIAUU9b5L1joPd0bz2ar93GhEdBXXCy/sSC66EWq
Z+dHzXex7mx/rWgJ+nrfDGJqUeUYSXGEuFpixLiK4Ux4omuhgvhzYF/MGqXw9g7as/1nAw7esrhz
TQBA/TALVy1YF4N/7VeN7Z67/SHRsE88y9GS77814VWlYz+eS9+yVQ06SbegZigNb5vw2CWtVySC
BSDP/xCD4G34gmeN+Td1Ct4VjfYP6JQSufL5GwdQvcv5JlhiTvqyJHOW5nsnSnDon8KbQGphesuo
A/D1796XA27EdCt+XWIRBVNUm94pDoTnCR+XUDJ9q3wsyfUVMhghUEYVmm8CeHUANGMrSP4ESQNd
6qeNNi1UArgQ93aO286QJSARucLIME2dGyMEfBNOovD95+UbtBjriAZQFjbZzfkkPC+sgJfdOKce
+1+XaE2yfiYO+jDnqlzqMKPkl6J3YFNrSLviZntw/aQFxjeccRjRzGO/mwIBluw9zOGorb+W4jQF
Qag/3NiDPM1+CarnFMZk+eMDj4h/064y4pLrtDxA1c6w46BH+/83bC2wQsR8cv/21ddzAXV83ixE
YdOJ5M56jpH0uCS7MchZgv/QYYgm4XvdvcN2+1+4n/AzM3iiOCoR+3h+X9laUFe4YgZ6eXY63qv1
fBGYKY3aMXheBt18WQId0NQJWylVRD1gfRWDpUGfA8cenI96qEf+tNhwXOoC58qdphIBUh0KXfut
2mmEdb/Cp5kKdKkxWdIq96CU3VDm+vmSRHWRt+MNq1Flb71cz0PjVEZud00l9mm9IwxVeQPwG88r
rzMT+LzDaL4LloAeUDm/2MLxbv9tEFm0hOIoDivMyDAFB8cEaXYlj9dZaoC5et/rbSwxfy/Y6iph
ckJx51oQRGgb5jTEA62JelWIeYzK20+965CHycXZKmwuIjT+EQFAyr2Y/ALDbIcROhfVh4iYzIxi
1v7htbf1Dx23yYRR15s3nlrEBpVmAR/BfyiDcQ/S7YFEkekE20gUnSVko9dgBllZqA7l8ybhVwfj
YJHM4fYQUb5rrbHLkmZPuZb6DFR9U//xkrvIecL4ifni9h1B2mrSNiAKXFkJCQF1pz8dHLDH/XV2
0PGuFN5R3pvlyOxuYF6oSJ/aKkNictfh7/J5EG/y+0e1QdN7GLLXJqxaGZsi4JeLG8iKnjdl/bzA
BRvUeBfI7SAnsStXafdmp95Ca1D4ceFbchtY5amdFmo8AVAnEg1fSfNdMjbBJ7Rmh8p16u2T3WNi
5kIRFceA7ul2thV9t4UUbLVXX2uLVcXUaOaZn9bUSAfb78UlzcPTow/wgtB7lsoQa+/YLAqUzFht
AVE6jPfhtJ1POq5OIn3xBDYaqYf1WcNBiR98c2Osrx0HwYsLxpzRXlgYmG0+qozdAVue8Zv//3UF
QjUNj8eWOxhVze/8DQ4WNnpYV+liufjqaG10BpI25CyWB3Jfr98meh7AT4gTSjXoFegLCTy77q7F
DfMMG/9Gx4KJAfNHAHNI8WFmO4Y6r8kPRcD3NCQMuSDgY4Q1c59Ykgf7X58OLaeLK7jcWZqTHVXZ
Z+YmhGQaS5AQ7qJrB5qKtNwSZ5c2UX2rXT6ogJrR3R4fyLNk3BxuUEpr3Sfzt86WwoXnMy2+TK9R
Tm43uRTiLTRoQxTYt+CEDhhw3SO0+K50vNOYE7LgfGdmgfHTumIjuC6ILu1naaRac89/W0ySMrbO
4T2oTIm6WluvQ/iqxFqXV7pKN3lBH8p7Vh04MPO8S3KQ9xhSWBoxtPwQWlc9aVSQc1FThZhwT7VF
qsSRg7efoVdtzrB2YrQi1dX0OUsrnkyRx7TE5i3cT9/ng5W3CV2Aso0tkh5KfrwGDTiudC1cCNbg
OdkTEXq6+of5NCgQZHHI//0iyeRvaiJZUwjk7tO/tC1yVbcLfdEMH0JpoLCK9eNkuG7t3SNBEgnt
oH56X/NhhcZwoSasUaFFCcPAFTjUGMQBf5SnvTwXlnd1543w5MvdaK36YVdC4HaQAlZBRQuoSFsZ
05d61bEqahVIUCjI3hpeS72bCMFcInEjl5t0AgvD1rwFRP2ZdO0DZ2CaYLDxUyTR++N58t9ikjfh
HS+GVan2bfmFdWrzh9wG3NU20STO7+3y9QTHerL6oxlfd3hSztce0nr0+DQzAdpBr95Dazv84neO
wz8upWUE2D8gaZP/iw3ZDjwFMwgHz/20iHEHBGUvcm3bpilwo+a4+vQgiVICAxwC2U+jVDOTE42V
zJjvpxInGZ+W9mWLEdBswkRldGy2CPy8M3IQDBLU9pCZoNsRbdPCtY8lxt/3fUKSSY4gUYWYnDCD
Z2bmhTPJyyRwbyO2ewx48GzYHAq7YhIlpXZjjde+CjV/uteavf7YeYJ5lKbLeoziVALfo2cJrLBQ
Y8LzLP3oXgAaCBrRky4MI6qpVPjlgSRWYh7aZPdbPq/sGXlSW3oxA10YzCFqkiRVz45Q0LezwHaZ
oCEZgi7INuyZIy1ujijcYA+VMvN0YEEoCz/dZAGvbEjJOaH3pozqlbLyl+dCsNcXw6P2+/ANQ/4T
LSrE21OKvvhfnvvyyIiLKrt0zbxlR3eB4PUAiQyObl0//N9ybs1s+Oe8uNtF3HSOghF88Z/lMWwT
0vzNEQR9j6CBDHN9Yv1nu0XVO7UqmW9lUkBoDO9mBi7VTvmqz+Ju5ATyw0H1gsCdGiIyhLF1Wa/M
P4t8SbzsnOqOyliS8IpMG2vVt11JwN4O8ud/0NKBDMrkeQ7leUn9zHZ+wzAZebPCI+OvL11fZ/sb
7QtUXxqwlJYb8zGsfdl2vKy+xMYqAz9Bj/4x9wTe9MTCvKv+14s+tJztzU55kTm3TZ5vH7I3/zpX
k5el8l5GII0HRpD5dC1otItgWt34RywQd93/JiBIoib/M0TOvPNjfY/h8mX+cQ1AWScRRKJSycOB
NrOXAaOlwVABEY1ariNJkX53F5EB+Hcbfi6xbv98rvAxsZeXkflaaclaBL5vjRNfm/ISKdZgea/r
t031SF0r22YXwIvFI2ca1xdH2tdx4i28oeZMH3T7RvuPC5yEEpI1SOcflH76YC2/HhxMaiMWd1B7
weqLZcBtdWMXsAy2tr68NYMWNbxS1QYCDpT7yTjV+6Zh0LdLbPh65V3w+9GoMIUFYs/go88Vexxf
aIKzj2WUTKboAdtuO6QjwLJfNHqCtchDY8YTVoKVnOVcOiadXHWX8Bc2PzLVPXZGo0wlPoC+LABW
or26An1ytODK0xECcNYvG7ZgooJwKI0KHnJOlKbicyr/WwzQaG5fM1WLncMsSNN8T4bDWXa3M20K
Tp0v8R5lF4+jPdsU3C1MseEmc1CJgqOrAqrGT5iK993zf9t40jmUIw46bBnSfo2VhlmO66bovt7D
tQUcImn2gOt3pH/FhstBCsHBPr3e+hFpHazFU0Ft8wT1rMxP41VuJXFxLhaoQyU130g7XmLd0I0e
9XXTwWHguRRcADYGOa39K7Bgu8Yp1W15zzx9VA8O1Dx+aJlDzHGrDzmzSve1CBLYcntmHWOfZx4s
in6yXhy+2nzsoSgb3v8/BkCFx0GC8/ABDUxEK+qgpqnj0021XL6JJlM9sBab6DocITusWvruDOAj
q8JHQDTPbRMKn4HLYSMwLHEr8FbWfLWmDUtz+baa2jiyWdeswsMxeRuLXqNV37OpPvGUEriewZ4l
couhxoWwbEmV2dD+LHDyslEi1LZfgf6sfqeb6/PZq5raMmEQEQpNJ36LR6YaDOqLbcG63Ce/SiO+
8BMzLVZc26wPWETCIqjCExIVjcKYnSDiiDa3eMob8Rv11enRJvQDcsUYKYxqLgS23aYxXTEMZu7R
/50Y61UMvBIFpa6fDRpDGJeT/he4lFUjgQ0S5ktEk3vk1kZYHbaQkPfkoWrDeE7MGdUI2m6oQtqp
rpEG0vahky9nlZT7O5dfDzzAkB6GY1zbphIAmaMUhMHPpbrRcuhM7ixX7HUQRY1FvdywbcOX4fNN
oK9L+cEq8D2wgRDg8vEHdoMfaui0ezRAhhIJyysjXZIIH8UfW/+kvWOQ9lYtSKqaHSMHweGp8At6
sq65oCg2Gt1dHpX7/YCGgMsvRVJxI0htQYfLDXZibeNitaS+y4tjeEhBBBBfOrdjm4pQA94DwykO
FO3R6nwQ3pFpunqrUG9KEcka/jnsSeSHDprIcD1SFAT6zP2kes+qE5wGL0uzsepLAf7MiMbicMgJ
x+bzLH/E2sljnjceTP8YgIo0Hp6ducOErvZvMMUhZRmdvP1581Zz/A/PtXxKKnb0uyQ60W2t4IgJ
Vf2VwWjTy9RBROPuWYbSZwPk2ivuhnZrlzm1fALrcBAnpDifnHDqDO1pk39V+LOea91/3AbHEDpF
iDG+ffdgcOSc1LxyWx/7nEz61ajLnZS2XtfWMMI9mp29u0Jy8E/r5I+n3XPGJIMpTK8MgLJ8pjli
j6trOQD3A2SibzR3uBJegNVLw9zAxBYujj/ieAvLa9+7dzRGiMDMPC6GJGHAF6nwsNbxwzBsVJJi
m4iYYF9kwy6zsFHLhVb3bjPKruIQv9PbDsDjQKgCVKlm1wBVam3geXw2Z1pUx+Y0eK+h7257Ty14
inm628o3EOYLnI0Rnu3s7TfHRUJlkn3XH2mTSVeYeYSfo+hh2Yn0/6+qzFs3UIps8gWdo6rX7Xwl
udDfCb4vIeWhW25spowWTq1ml21a5bFxXQdTWsS3qL0O8KKCpJNt2lQwm2RHIEYDwFLuqQ7T301n
b6HfYVCo7I8JNYrl+wPL55Xe/j+Cqmn7yPRDAqvdluT6lH8KhBbcV2IaSbkLoD0b+9pvuTJpnhIT
tZS5MbwnbmS4z5rJGxnYpxk4XtRcYQce0wlRKTNa5GYneMtPDjlYXRhn6r0IXZ80RekI449P8BKH
1z35JH6jZQUsgW3lRyArkVvfKETAzG44CdZAZZR0M4k/WQriP3MahZh02IRpmtqiWonPxJKkDdXl
HsSeYlDTmLvgZu1VBw1CrzZTisYobo8dvgMI6/X7zZb/3YUL+dn/tp0S8VlovR2SKOETGhsSWltn
+8UP4DrubJ4dhfn/O5Kmz9YrK6+zYGwn2gxUGIxul0Jbi3itFfwYyh9giwD+xy6XKYc2BB+CaRoB
LuPh94LvCrytD8G5MLMwVwIjFj1mRLIzlbUVSgIdGO6oV1vj1IpuIC3ZQ+enQS+BWK4hcavqGIp5
VPSBT4Wxra+FFYY+8ZmoQ+wW9LtP0Wd/71j4C2kUR9IKhra+vkiQDUiZVjLxIVCZM+EcAZ4jCHqf
9Bfc2n77jbejKl470PQ5pBR0gdObnVrIOOfMQU+NrsvdQivYr+PIIIpg10+atTmui44QMtNkNqo7
gLxG59ud6s7j6CVOFB0U49PljKOeHYyqxbT4zez0esvLOl/xuiMdvtdeD3/zie2abrp0gIBaIXSf
xpXsa06DIMiQk84t9FCevUKrXqOBQ0Ef+YptuVa+0O920zzH+B1n+iDG3f82NgqY34a0aapW3KQ8
mtaMbVdb73EgMM6bcbnXI3tLBhUF28LJttOgP7yf/qxiJG0YRuzaBltZZaLYvbT4BPq4sKStBYEy
8UD9fy0zZlzFrT/2CLkDtKU/gRxUX8+gcFuRxwHp5enlDLxdka44zLmWkaFqK2TT3xLF4PLfpndO
dFM9tHzUDtgxx4Xubls8wGrLxNHQG+ZNIQ+xMCZeLkok7e3ebU7mG+kATi5dK5voq8dHYEflkRqL
YuQzmjtnBvLI6x/MqcvgsfWu/NPrKtiPyM2qbaNu+yEerJK6G4rf0Tvg4c6BR+zJrU9saYmCA2Qx
Kgoqvt/x46d+DFNYDcmS9SxH7q95lE5sx1xsQWEUvBklUfmbo2CGrdPEz+d72mSSGqmsoy4ekPlG
N+CO58yXCLDna6OVPri63et8uVieGjtiQG66PH9mdYA4W05aM5hM4hXQb1YMzbuOS4gL8IsMNeQG
RM65VSSOiXb4aSBQC7LfpiClBQczl/ro/M83PfqC3vrEUs6Qoc0EB4ac94YlvqdyqHHfJlpPWzCB
smV2yMTABMJpqOTX3tV0d7v4syay4cnIiK+Tz0Z92oo00dGeWCsFshnZDGzTI+zO86wJszk8a0h8
K5yxseaNEN0+ZdflvS3yJ2FJ9RJHfr2YQacPYFp1XH4pY/hqO5ish/dpItA7uNybr0mAFrwYO/Dt
9p70l0k5gMT3kMbZ/k26GBuIB7Xbz0SLg6liY3bFTzP22PGpbV3rMr1R5h8lhuzJ2+DsKg1V/rQ7
i2MoxkviZQSJ8Q4GY4nE9c3RdD7/aQ0yku0imKmkDciCi24EJu6sQHC2RdZZtkioJhvpLzsENtxU
zq+ZsUhYyf2iY4bY9U4fotedVuEckLH58xn+V66nqD2/Yns3vB/2KOYTE0fJzrCPtHlaoJBKoKjB
LtLDefKieY21OzPoKA1eYL1oDxJ8PMWRAv5ttiQZ5V/SEKA0ftfJeIEvjR5f/Jd/lzs6JoFAKbJM
VVYUAwGiyg3LvR7ZtgcKICzMCB4edC0wGAeiCuHxgvI8KIQMGYr78zNsQEqTH/X9klEpB8tsZwj2
2H4vMYG96z4MRnDbRUmZvHjdfOOVOMIv32VDkZZ0tXRxJYdLeQPJ6PO4/Rdv6Si2TiHjhtF6L1BI
Jkxm4KGivflTgH1xpSP5+rVoKMYA1A7FwpeGcKpQpsfwSBQTVRxqNMF07PgmsI4adu9AkWotBhPu
UbR74CDSLUft16V6hpnxEYipD2bW0IJJa1YgJBs5h9vmZecpOCrDnH0yxIBhaY3vWUnLoD+Oewmn
s3A58RIVIaujUHYTd98spVPJgwOvT3qw7TpThxhu7JINrQn9YSQw1s8C6XczZ6sRHiWIOo8kfzzs
fpbNucnTJdbVroWid8bUrs3+O+rbDYDRPytur8sqQLn1VW1BKf3g8uU8QJI1T/SRuV1EluS+pQN+
rwbAhbrjwNzfhyw7JYWhC3mkjO4BoWvNWIBZFlLFl6kSUErPuRuodcXGPT6KXLG7nI7ZOwo1yTPK
iQLpNWIY0RTwAKqKq1K6GH8Nn0Zpb10GD+MldAmmI/OwgrmylL7C/SuE1KMCCMs6cn/UWUnxOWZ4
Q7zTuvRozap0WbZF2GovNf8+0lZKoGjiXJ/E5bL02x9vg+gCEsV8DxybAUYBJweiNSXJQyOKgGVU
80LTtAkd2szbUPu6j1KEZr4ki11KaM+ryHmtcT3EiMaMaSre3v0tTozMAc3q29X3kYh4BBnL8ft7
v9Y4fX35w4k8IRft9C8l3eqP6dgn34OAyqvBWnEdD1HMdSpP2aMvad0KNw4ct+pmzOZTKiIvNPKb
4oguv2Tamc7kb9X5K96wUAIO2c7R6PTlFYAjh+4RZaGTs543JoRE+Wa7BboX6O8oFRzccebRT8ff
KldHDI+f43pu9TaPJp2V/XvnA5dTrgLUg4gmnUjeZGXmWFxfmwsKediWE1+6mROjGICoreg4F65Q
2pzLYWLWjBK3eOQQhaCYl3Q4/ETqngVIAamSy0bJVyQp7ykg1S1JQP7R4XU3ns58nC0Hb45+9wge
k9guOanjCqsZipmQQFKXDaCgH6v2JkKHTooGtYXGu1ZZhE1Mw9L25ShvIpW7Cw7occo8vTmp4NCO
S/j7w4s0ikrayd3Hq3earsZkPkRScbzT8lzWGUdrwCaDboE6k8F/mBIy+T2GSVbXv6P6QUg3PBxK
Z7skFdkNdx6cgBpu4WZMKbX6hBV+ZwW20fwXVYM8l9054cmCKxKcGz/ivq1iF+DS967hh3/tQpcK
hNlURhJVViYECZS1jg4F5DH5ACCnFQ9DS2k7OWc7fdnp5Gyu2nfajIt0JNXpG/AOFC3hVAVsuozu
YPCzxiOBqJEIq9fEAKcSpEvGk93mQKvqcGzFKPmFx5HaXsk5ykRRr72dfwExcBI+JGYFKGvypsxF
PIDbf0z87PQVAIMw2n6cwVx/J8dWmkeL140mxkT/MpK2x5rrWcKGwjPCVGtEXbw/TfpxXkcAm2NP
wiuUv8xVVi6mGBFapwN8F4kaOXG2Ex7fe2oPNDMB/24Z+UqfRLxLhZiNGo7RJhtcnjzT4kYgZD+d
UBlVg4aFTJdyQN8N4WUfnGwWhB8c9DcIBXmPA7XbujVczkPhl0ZU1RToNrwfmJJggCqgjcFi9bd2
ELNOE06tiG8EkmSBYEX9qo+8X6xI1CrNTn57KeSxRyq7zlNM3dNq4ccFGvxPgH1ypXqJmlh689Jh
2vcXNOR+oxkZQACXEAwPEHZvCvIBUtdmonXN6dm6bmv12W3jwWgnUwoFBt3+yjA3qVojd1QNxsF8
LirVV9+Ak+lADM7ydTys3jAMK31VRYl1iqzAVm5XpdroS2m/7F+oEfHOxJIsWY6fDvIzMV4uSRZb
BnmKwqBvZTKm0x5j/MTsQf7JlYekOTqe9fdGODl3R/HQzJlwXNlxnKCd9P/0DvuUkf4VjASbXTLM
gO21R5LLKr9bc+RIlSywiTyFf07GQyi/L8kwrSnne6UHiSsFWFZxIWQybTBoHTsnoRYBKetlnKEm
YiDjCg7HgK+sWcwGCd6Ulx+rk/XIPaBzCdeHmfvvuTbR97cb3VuquR3O5axVNhPWinMxgltZjziM
Ubc1faWrYDz+ZN93stU/xNbQHLDYOvTVwXHymao/W5Dabz6BoUuCh2RH5cKKUq2CkFEOLlIsqgHF
hCl6hWD9EK/P9oiCbQPwZja2YsIQx794qvyBYmKQo2Meg4pKIKk4CczdFqPdZAkM4aukrSY0+KcM
a2Lz5EAmOlySNXggTVgE7U4cCM4BM5QlzaGbq1PxjSWCdhr33tmjAqj4HNDKM/PUuVecBDwXGQus
8UkROFoKaJei39gXR7CI/USvIwTK2qhYWCYPiL9Hp2Xo7nBdeLqdI0uWF/psUqqg+nqDjqwNZFsL
tXJGDCN9qbUyMeYvXikaB2ByvYxmTVYp6vB1UuDJpVJbJERnnyirpbg9cMPE7FovW8Yq+yotX/Wy
fbLhJBgmYF2C6fn/o+W6/G1dkOTt9LDTWlCrBUaUn+XIS93ENUhsqSIDalySeICO7fhFTlkeNjCl
PuSj9btRznQ82jrqajBMlHGF3vpsLOsXUkvBLL0CNgqpKP/DBb+T8KW2gM5QHBesR0rP9fnzNPSM
ionc+qB3peE1XBQNGrJqe387OdddhAFRCbCmk3VNGxVVgIXQQRBSwtoUL80wHQm80b+NgfavTnUQ
TxwI6Xet7W/hMBMn0Bhcx9RJWBzcYSNs09sJnuAhiu4XgS5v/wdKb8SngV89qiAO8KqSpuSecW1n
EFHK4EQerFfyAP2GUREQ5zkV2uiY2IGNmgzkw0+/t7IPvqrySp1Xggjlv8FidbPBjWS0CImHTEW/
UZ0N8ViXL9/G76SeP/3+GywVyVWCgmewAWW8XJ9xByqk09NHUfOb39sfEMAZN0T1KTV1QzIpInwM
moFQuvjL72NkkRYGSqKYsq11DZXl3S8iUjLIbvX4Z66Iux4XJVizb+CAqGQMn9t6JRIGMpJ2OUcr
CM0MmzFRLv2uA6twVNcq7shXvU120tHfPoMJxfi2peHjWaGznmdDRohgBA0Y+cp4rSYtmMBk0+hW
WDgMRRv/AQOTkrJiqhLdsCBxLU/E8oGx0DpWod7Djer5icymg+Xa6YLBm3rg2xWdQM2pYxMPVwgz
oLgA1yGnOE6oCcukRYELsGqOLTpsPL0i15Vy3N19SNqwD26YOOt3QoVL+GDqA1ZRO4fA0pM7U2kl
FPpDZ55efso1OR2U33HN0KEaz0H+Ss+WsvVF5G6g4hn0QBiA9le06JEmo2fqkA8MP1rt8ir4WCuQ
bOfFU8+Q29/Lk8c/466FyE0DQvIfvNu8kLfhhI1aEoj8NHZF9WlHHj4QAXxY9DSHDfDS51YgwfTz
UvEjJZY/z5rwCmt7pA0dpRW0rg9RV1zHAjVneNm2VTeqWEWe9Ys1xfzr9Wj5KD/sVa8BBQdFQ4Op
vdhmWefOCvEc+q8pM8H0MSVJbfr6uWAGg603ed1Ll3jkHI1nY8j8x07rHjBeoC7RKE2EzFlu2Qlj
EUy76rBs6DToIiem6rtQmyCSUeOr0ydVqV8RlsajegVRCmM9brw0mAoFw8uPn+lTcCpOT1hs0Nhg
jCD72BfW0feaXEcNECXpLkudmG/Lce8uDfLMebJ6FVoYbOt8Varo2fQhDKijNHC8euz2B9L+PWb/
DG5/KI4IaShXRwYV2ULOvGaJxZGvLmTKyJoapwvjI1TE9iixBdEJ7hJ4OmGCz1qz2aagjcgsALcn
8o7h9y7FH4tk9tjOt5BdwcrnRSmYEVj4pibYny3D5CQTyHFU4OnRO5EK9jgmtbZbNAOH6wEOBZtf
1GLoa+XWQ6e4Ti5yDcmgqnLOJRZigzvQtqvA4KVHZqskD1UWwt8nqq0A0CQED+XiOddijHdRkxYk
o09uSQPsXRW2e+fPO4KmDeRTQBmJ2M4mhsly5IMvqWSszAYMYQzLeO3yG7qufsdrtk8NUc/ugzgE
0LUa9aoiicRI6QrOY/2ycXloe7MNNN/Tzd0Zqsv9uSFvCTAOriiOZx2OYqZ2iK5qZxW3jpeUjS6j
ILEcld4DZqyPOm1I9aV09OQj7zC1bsQf3F9w6BUCUgeAMPf9geZIV4BPrth8hdVAVgfZ2P+94HGn
CRfnhEJX5/bBrm4KbdhNJ++DC83dDetxrT6dRIgk2AlV7kfptYyE7dLGu0XAAVQEaoca4lavkJ/3
RBkRT9fCmwKDzyLp7diCr9iLpk56urP9gNThLi0oNZZ/8tR08T5KU4oiaLztRT3IIXODLlyKK9qy
HXzERxgwH3Q7Uxe7yU1frGKKT419pT7nGWDqgGmNyVwpUtOGmCXqivVEevPmuqyF2u2RxGGgD6gu
yuWf8EVuJiKgPuiJ3/cauvWg4wX1eBZGDTlwK/Zwhy9cZwHcdmsvUUX4vPqH2CrZTyy/Vtm2VRe7
5nZONCmkgm5gDhk1ppSDEJNBdRW/+ixv/jv0EweLb7imapFm3mcKyOGS0/c99nU2GSxEwM4wQAs8
tzFFGEcvIbu1uge0U85GGZQY7Jg1SmyJLFa0FD+hKhvOvVK+qlVJGTVhURmY3pO8QiGJRG7Z73m1
JBKiD1V1j+TrSfP/hFc4tdFk9n6Oy3J0d14znxFywZPg+KImylGuSLAPwzmS4drAnMkUoRzAYq4s
0jvKZP5rrSQBIv46m1hS0jbA4cbZoSQjogrow5MCpHXSDVpkVu8ZnprI2c6C3aoGeCOr422DQGTq
Bq1Ij7XCUPPgYr49zlDQ9rKD514r/RY8xcCqnNkUIYpfMuLAMeFJ7WyTfRQ/qT4mqn6ZjUCpC3Ke
yTZKOIYVJGbnHCQ6UnKF3E2gGv4zz5PTow7j3POx9JvMlcnl0JolZ67LRFUAUJy6EnXxgsDuWe1x
YGuKpw+mj1GMFZ+y4wDwTvIJtLy3Pi+iWzavnIQbYMNjDpnjU5JGLNaL+alAG5Lsvs3q44br1b/a
WDCfWcl+QH5Hyo0qtAqdLq5G7y5ngmvQwn1H/2u32nnAnopQNfvj9Tj7cfzXSFx/qrEEqB9nhOB3
5MaMz2s4TYskdQjQzDlOufJo+sUiUbBGswiO3TSP+EbVFy6S+6FVUNnCvqSsq3HvOyfubO5uck05
hIp07JMRJoEXsBBJ/x5zFmquBAIRduQ/AHQxweRvBWIBQzlveQCZbE9hboJna+SOsnofWNFH3ZNd
QTrBcYFwSWTg+gWrF7FSeMznX4CRg+3K3RHWATStfBxeCVtQnf/ih2dNsyAXA9HHN1xItbKlkr/s
hGXdDVbuihImM97tpMVGzstOZLzcjOt5Tib2e2zqG9DLUfmZ2vXxb9uw07ncVgIfdjFy3UWRt8I/
YxnHuEgua2fwmiJsdaNoMZ8AQ+n0VRVQTbOUBoXJ1SxSGw0En14lT3z9GhYoe/N/XJQCsygvKH9A
7cPovEjc53gwNegOiMgoStNUpIlIfGrhHziNvLNAPNOWkeRJVg1SbgLBLvc3dNGYC9I2otkM62fl
JKl7o65NEsLrkWuRLUOSiuojHMPWh7sjezWSulfnPCHYhAmbFQinaym3gzAnpSzAO27wrUeMFV9U
F9/lG+iMsCjz+mr9gw3atv3xWpYSpO7TS1wXWEw/QSl88g2gVXgo0InIgUrGlI7IAi3nQ4ajyMjj
T+nuuf0n3oFkkDf5IxPD/x6i0FewVMqZ0V8h2tZ53Jzo9ZaMNx8lfrljpq9MoM7Nf3L+vH48JHFo
OapOXT7aaZQd1YQqJZ5m32aVF9T+kbamRAaO2uICmbdUVAHniHmu6oNnZRTZdjf7aEJLVlm2kCAr
MGYcgUeyWZOdbv4TU5bjLS6JU6P3FGinsLxVAbe6zxonXZDew1yily8/b7ev1CzEwbFNz+JxbOd9
NK81gY2QJlC4+zvn6MQCVdBXxkDVzA+2OTHDRb6PBKrJhM9eomGakam9hHxQ2MbRfVKiicHP1F3K
X/B+aF+TnCt6UVznvUkmF0RPIh790iByr4yG5IyQRYNv23CvbjmdOl2XgLzQahm1fiZG5nbqTamD
Root1WWWKxfDb4BxYeSe89UMyRjYZAgjNG5AM9Be829Bae+HPxzFue8sxCtdyqamDrkmLfjacpSA
F7y8x7quUgyGljiXU5Kk8SFr8BQvFbe6d0mjKkKEasJtyciQncfBqR1DPI7VCbpNneSdUaJk/EAi
dsu9gyrJ0h/C/U76podqRo3CWnvvDafgPeH1VAChhL0JGzCab8xu5EYELr6nm88Dw05gdqjMLBx1
hiZ6vCxceWO51Wr+KVvzOT+5a3a6G23qt2+GGmaTu9T2EnC5zOvzs1jO76hstsZmwGYuQ9u/7Fmd
/zG7yzRLMXdgwdOIVt0hG2Y1TnWdlYF2nolVNRHDesQYihNCk2Ovf42j/32BLy9EwJAwALAzl1ol
yPGTXZ9X9p4MksbcKo2OM4NW5wYiX9qluuq8f7m1w0edoeBxj61ixvVH21o7W0QBQZgKSf0rPNNR
AAc3A1jF08BLsd39j9D3o529f9rayzynfyxQsPNjw0DDCQfcq7PDWbz2Sgo71e8XMWEnxDMFLU+j
XDg+w/zukZkDYaMpJRuFh61nmZLuo4B87OS0CA2+xPuFwplt64DttN19nuJj5vMraLK3VLOft3Rj
6BEpY5NK0B7NH1NsMkpJpWQQOJQk2D0v/MC0komVKUDne9xdKBumep8cdf4/3CENLWtNfu6yToob
R6AN8QsvsHWo4nwW4zlnZ1DB6JYx9clxYqWwAj1mP3WiopGM/59E849sSzSNcpSnY4Re3fnShwyH
AFfqzSoAhMuNGTfafjP25GMRDiooN2LAWmOP43+1GsY8fOiQx/218Iv0bw9hPpfbfrYdHJyIn5QY
PIomfPw5gd6Aeuk36Y41iwOwZoZUAkt8ShqLA3gH4cT4/PVzjPMa0gGO2/BcwJysvzdggVXMevv+
OZJchcOVitQVUrtqiSSOmz/eVZYzT3dRVAzoT1LSawePNdrdB8FuGmN7MZ5P7qZ2QhefnnxJovVi
rwzbOTL6ss8C1Fi21Z6rOYW+IeaB174u9EJytBZdWtjw87McWUXBAZAV/+EkxE6N49sSbJLMKE38
N6G2KYuaHemZO1yfIscAOMYC22Am7RbDmzm3SERyxLtKT3RNwdLwO5m4NkQjXIPLm3oSGmTwSwCx
IOs+nRmIq5JnTTnWRRBuZyhywzJXff+RVo+Ch1akRiiLiQWZd4AIc9REIqjinwW2y+1rcgj9RqnU
ySIrigqlqG/nHbu+K7wvWSPw8lSRurhnbnwilPEJQQvU/OLugH/rvs854FnqAteakj96r1lOmSUY
OyCIN5pG6pNi9y2eqHflb/79TJNR8ZjNyrUvVP//QpNQVEXC5lBy23H5kYNP57huzNQ7Zcc8oQVq
cXBlWGGDHZp1BxmCnFwSx13Czi3hDgzxXr62/ZaFzaVkxgusoWqUnzqxAe4XfiZQ3Va1pekR0khG
FVrh2NRmZhGHyjNHd1Qu1f7Psw0P7HRrDUkL4bRU8TEtQXwrakbmQyyQOUoOumDCqUvU1Vq2SX5I
ZCx9LtMkHzARc2g56FS/uv/e6uIwAEgtW/jcUYNXdtQ1r5ThNnTRwx7paM1LFGHslMy5uDNBtsxz
ffq2C51tl6nW8/206qzBKFaNy9HvbflM3t1St+J5FgL8YVhd4WNjfpJPfJIW6VSQ6V5AKUMwQtMx
R6WBD+UkVZHvnkEe+DdW+aDafB5JUwYgjXUpogLsfBz+hkKPBkLJu6sW/owpSmzQdfqX+3wQqXWi
XE8p/y3qf54Ekz/7fXznGI6qN+T8Ospi635bpkY9lst0oyvp9KmdQSvyYZIsRq5Fq35aSJgB6GnP
IHeaqvejW1c96aRk2zN86Gcb0CDN5jS4ckqwr1GKCzxRnpyitIKfTHYc5G4yqgZFv/7+J86I3j9Q
c6Q3Bnfg9PRyJl2R/rGbI/HPE43LQMvHqoWw364Sgkob0QoM803T9JiCuA3JjkXdVGTju9cUXaNv
QPMa+JOsGtEOLwhG7ka84jzbvio4GwzkOEC56YPNfYjCdlzadkEkItfGZEWPwSHYl1C1azqMOmEB
7V+ysw/30mLNQvgJhYJGBLMNuxRGE3pe/9EuE3mZKRIheqN2lsjvnGYefGx/cQiA6ZNO+9WyOiC2
5L1xCWMUhF8ubF/WeXvrlW1J3AcAvYLSpQZsw6qKsUt59LhFe/lSF/dMRaE1K8C4P3SBCvX4gK2B
0Q0qfmOH3HWLhc5v9O4cbaiionmzezURiuXe4PlDzuGtH4bsAu2unxSnU8Gk2ROcWiYfQNIO+TD+
4Ie7B4j/zTyeqzxQBLKa8ugbozZVldK/H29VH/2wamCJg8VgIWt3iYeFrFe8KmGqiZF+hNma4yjY
sipI+8Y5pzEx8YUp4OtmBaFpeQq34+4++5Qd2ZK38dDgLKjXS1cffmdJIFC0T3GZiDyB9apzheGv
qEigE3bAWviO/hksC3RzTLe5ywXsYFExPBdYwhKY7QjpkbfxJzpAB3B30FZd3yxqewZNqB8piWz5
9BNM92rGK8r02sRqnY0D1E4bGjD8GOrW5tPNt73HroyAeBlEcE4wR9W43md8bwONUo92X+nzVlFI
fOi6kYm2lOjHtED7fIooAEzWEb2Vi3yPkLpvPwKpJsP15xtyn+VUZL/2vVS1rxgCcQ0eTUMw9dsl
OZt7/Zk/JeST+UKnIkbH1bvbhWO+uH3SbB5FzzPzfLuP61eXocqbCWAgO1xyjIE0LZYqpZwJle5P
raobpqEpuUGzMVwK6PVGDo+zs6j2o3YO9MOromd9ulRCUS0kFNV4VS7vwPvXgavvdkRYRF27Be9u
b7rTwsxj+JIWObSD+zPBrPTAjEZc9+e7r60ZeLQ/Zi5ATzevZtGm9PS2ItpBZ7mDInXJjtvj2BPT
oY8149q+oCXhECj3o47VFifvYwS89nTAmM5/Tac5yCQpjq3bJphF2LC73hmposgvVg1Dx2tSkBpJ
7m0UsAzZhEzJ8csnFyu8VKaYKJmgsuKXDUFIjc5kthh7V2LTg6RLe13n+OqPMVyOFOWqKoacGYap
lvyaTZOZpoRWIAHT7fpa/tn1g0eGLYGdeG4ilKMMyigtL7qKSSOgrOpesEDFhA+ZyZMpuLtqHF1Q
rnJAu/nVDKk+DMSyHFKblmQ2XkR0PmL1GVmJEg73xdu7oHvGJX36B1L7I+K3lWEhpY7Y3hNIo2j7
JUVizPo0Xp0FePlYbOhzrB2cSBNu5fNeZz+CmyxbsfqNpELd0C4v9Gj2l8QwQzXW+nO20xb6E0qY
GjrXYDy6VC8j/RuZdHAEyD3Ez8L3F6jeBcisj2YZ1K1AmMU42BJqenMV7QhxefKo/RcnHVYVj8Td
T2I+nFEEOOduGJ9CtbLLg0v/8bF4zd8xJMZOvVZuy9Q/wzGDUCnd8VXDnDjxWGs4BcYZlqQARJ49
hIxYzDB9+WpgUefYRj6cIyKzTFNjCfsJxSj7MImxYCyipP0vFi4lxwmLtiReotHLDzSc+P7trXW9
0hQIZIwQvoMjAXHs7ZdqvVStwPiyCNioTF5OUZ5remojaFcUI3vXZT/jA1PTr3WOcjCgKg5M58VJ
LofgH/2IUbliPDitd13tFuDO85fQVWV/yyxr0oGJw/WRNAUqaTA4L6C5Dtdt7aboqCc3Tg41wpbC
WScBmqhleC9JfOLeTFxy37IpuD75xd76OkTPswKJMU0gkDu4N2mB/W36WP3KKTU8Ij9sgPh4n3Hr
L64fB5QmOH1jee1dbyI+DE7uF1pdxZfLXRzrsBbPe1eexTVmZZHOOk2oI0RPP0A3E/JOQqxyJX+a
0p/no/GTqNtMzTNtBmpQVbiX5+do6GNcoDvlW3EYxNBWK7KLdlIXd2uf41eRH5nWGVNuYZn/6kyZ
6IKOrA7JLbIsB6Ze8azfnuwu7Kv0Vag9TP2/SYF26GW/tdwwcyXkkggkd7bzEbxpSQitQ7eh52wC
odV20jh2C0TOT+W5AKHKxe1S03taKeDIulLJKeIqfO8HUEKadW3vXShNyF2oNIt6cgPeGUMoCpqg
L7+GJygGnni3plxBDnt8RM9UMcBuBeN2eUg35x23u7gmHiteZjGoW2g4NHKiRj6RroWtjAijcH3t
/vAlnTb8poihU/8+hvknLj3NTMv4Mz04hqkyf95GOXsqHIw90V6336oWlv9EjOtzPWXIRkmYXG4C
FX3EpzeXDr82XuaHy0UTDO2I1FCT5T3VQ4bGIrEfKJMWPJ/PLMQHMJKIyYN5lygZ179QmQfp5KAI
4xYD0jRG+I0i9kAm/WDwWlJ8QUEr5gg9irInZeDWASGeyPHR3VzpNZSl7MtHRnt2aKMtsqRy1c4S
hKM/6ZivvghYLP3pjBiL7g/jOMyJfOh+iSY+JUS10eVXBYTitHSwk1/5plL1IGwaGuSn1WG6qRUT
tPj/r8pdyiSa8V8YKKliRROW49BqvGQxINRZ5x5afbxyQWk+QJoSz+3fEtalKS0eHPF8EgRqyonR
pgwptC5cZK4s4VP49O+CIwM2BJ95UyCTf+qaJ1Senh28yVrRNgOS/BMsYV0jXRCQoE1vK9o4tDDD
li67LDBb+3gH84eJr4RCzy9i2KzOOYs4bKChLOqv5a6sD77cTZfK15VjGngEJvCfD5v4ccTAOKyw
FPX4GHBlZt2Gc7xhYnAmp8Nmalo3lH0wWuKoluuxta786vNUfXXvz4+O+qUE3qedT57qjM8QW6hB
aPWax7tPaTT41N6rkaT/EnL6UjtSBaN/uQaWMC+2X+LaA5bYrWngA5dxSBBGFeF4QTZ7yllKRXR5
bG3dg+Lr7yTN8axU+48LD5NCd5lF3Bu7cXTwLUoAjyChtDSyYjaKjNAcI6w84UxNWL+SaqGcnoaZ
ZHbEGwRI1IOWxs4uNPeotJfCBfsiNNKXG9z7fx2QUOdXHNQjn43+dqrh6ON6w+YEV9CRrl6A5CMh
IdfJ/rHJpCDvSI7b5R/D302Qp3pDCC0HN4iRpuwcYCJv0XRgSzK8VMMXYU8RGazzHoyDglkewRJH
Fwbbi2y9W6fszlqO/fekzX4l+/Ovqi+sT03jlQxEec2OBGrrZDvLOutDSfIrrdP+h8pNNNX6W3Ti
zbFYGqtFVOEZRrPLP2jWRm5fAdTdkN3ciazZtFSm+qSECkzVUoIp2l30XmJe2+HCrzdq/E0+WWxt
Qw5WCpd+qgcm0QJts3MloqpnLnHCF4+d08oI6e4YEJ6xTHuVll1GUYPKS/62Ik5SZORVIHxyS+e8
cZGSzAs3xTgYyE1hrADUkz7zOpgAEfOLSJ7IQP9JhQMol8EoRXWGq7UnZ/NjjcHB0yQnvToVGtHv
7joqlFAxZyO73LYHII1itNrapR6uIMsxnk3/yP2RU5oSrXddmNUYgRvsKSuPsUIg8X+Ku8S6ASNp
bMrbIaXUOJN/OE4W4oLx22FEEBKRM7GEEkmeEzqqCKLsqp8ci3E96o05usGIgLMUITVW/dFshshj
PgsmqMSVaeLMWdY9qLC1NBNSLqpamc/guClQZOCH5ZR0ZGDOr4KXrFSfDA+2qDT/yDFMLlZtVudn
EkkhLJbO5COjN12O7WZUJMkeqQdmVVdI4SjdvLczhke360S19gDdMLZnQkH4BaUs7dPcMy2RUB5D
yj7775itOl0Z59qR5SqdwB6l5CmHl7fea38i9M+RLBBTungmhF6YD7ioqnZAX+z9w63hY/6v8VdX
7ZbwYwzoszahc4Kl+DUeMCOseeDFZk4+xfsTUDhLiArkcZiqScQOtmbhg5HFbFE01fcmFsBzuiEr
KFw34/5Vm2YH43BVymY9fyMETNWJym0gelZpMuc3JPl4qdlGL/RaRk7OfbCbjfgQ+5AJ/VS5ck9N
mCcestRJRdL9wVlomNTZNGtMxMZmbyfG/1GY1VWah+VM4fJLTQ+jzea8XJ9c0krFAu5zPvTWfdib
0ayX4JhwIdKjD5/cJiztlbvv6pkYYNQeMEMxtSJIC5gulxn2bkZ1liRo2G6muojVx/vvAlcHgimN
fbVudtmE3/xxlfEDO4pAQT3mD8/Xr/aHlmKWvdyzBuLt2qeHVF6eGo4/y7kEewFb/cL2mv4xXfNH
xjAeoHxtcXfy828P5JRHBaJPLp1k04hdKRb63OhjW7QlkS5/ZcROjsNnDx+RHEu5/GgoQz8lIFHl
MQZOYDxjKcrQmacGGzdbD7Li4A2NiWuO+qaMNnNFTT/qv/t64sEq7/f6dLT9+b7LlwGvWVB5PfOH
wbQgwHjEtkOfjkJrls4LCZohepTWgL43PktpikOAJRG9HM18seuOreIjyKpm9HkkE7OJ/JamJsOk
VklFtCUGX0lLA8M0vZvGtB2Y+YrZXvrdDTaBPsUldynsL6osC1Af31D9jxDcKviFbZuj1dBAVvl3
Ge5KT/G8hxjanhc9js0No0VRX/INwWa8c//VHsZiVq1yWe4KT27BAcaPu9I/trbk+3ZRvB9h5S+2
G0UBHxpKlyCJ97aDpPo5INZnUv5FBLknW3IWEgyRjVgBr0mF4TY/GTPjPOxZ4gn/+mAzYuvLQaAy
kDrz5DlqI8/D+DMLDIBEkI3avtjtMuRsPxfayGL00jBd4+REo7nurgO7Prbb4VOEfPix72aRcR5I
ptqAtjWY+LyfRahjDQy1Jh4hTfji/uwwiNqsdAPhYAYagpy03C7NdIrSVPU+886+rUik+k+L9RpU
pqpteg8l1QbaErBsUmOti+f6n6ijRB6WW2hfKZhtsQb2rhmCoanWnN6AoosdwGgNbTLJEdhIaEKi
dQANjX+VaA4165fLW519V34wwjeARTATLC/tr/NxrqE699VyAoCNlS+0e17R8HxpHhWN9eAPJNao
sfY64GrZkKpvGmIX99/Rx1aK+kfvK5FENUZ7gMdFw3ni440SMsLjhVx3evdgCMpo2XsKjquNUofi
LUdM0HOV7ZaFKL+mNBCSZ7K/vvMHtHSA8IDzRzOOcfxBaWy7gnv7u5N22OU/NqZH+wyGA68EZChV
bfyXxIcZT+VLC1FdToLK7tCOPg+Xcqd42o901WOmV2WCzFuO+O/R/rKLU5wmx0HQpSC0Uw47MIJO
EANFGA7pOk4tRLkJ5B40PhZn14UKeL4gGGYh9/EJ1+GBbOmq+Kc9Z3DxA0nF1o30jG/vma8WuvJ7
TPFNd7UgKuIUsaHki/5EjRcyIazkMxx4hVaN+1F7aYI0fysnXbfANxoqpkh/EipwDb5Gw/Vdsrjs
9NMalaahaYeyoPnumnc5eGK/wSrXabR5qrcL3wG/T3vVWHQ4bguQXt3hpZP1gBp7Ut+RVqPlejsL
InXyGQSPETY44Lgbtq8qbQ12fgf9N4Xt2jRCNNH3wDTH4kJ/weY1bU/Nfi7Uh7nQ5Na3aK9bjY8D
Z01IQYi82gNQUXMrjEYptDzP0C7z1O/HIenrAtyNGyYQVGCNBLtxRfqBitv/xY+mNPTxgdLJtcZC
utUymjIDsrqwvPL9ChQnr+9U35RSbnLoGrI/W+Se8YWhuzqqs9I/Daj5aeKCgqNdP11FOaV+HCye
ABKt8JPZ0XA2OTG7dFpDTVJ8iOO/LibG0AW0BW+LsMJq2rvKSCLGbrV0UgBsQSDQDOoViT45L1CS
rAP7LJlOY7iIzr0HQKYMY8QtmPY9/QlPcKyyLIdVTTz26JXjCCQuds2L5O6EUCOSUMbSua1DTAfg
BYE85Pm4GMozbeqpp3lCSXNAoL/ANTeGBHlCH7N5aFoeX3Faz5N/ITOXhnqQGyb1CNL9aQiHQOfh
Q2Iu47OkF9LNp7JJbxIBNehBwZAgD57bRilJ7wyacJrZYuDNxozokcaOdFn9tlRY4VkcCj9oq9+D
/nhU4VOLifkKXawmIs7RtCmJ/myVZb1ODHWZ/b4V0TdpKmD+wvkKoDWn7+Nbd0utS+bImWtqX/6E
7z03GQytX4yMX5HnONVnxfEwCjbafC5lGzi/D8pD0oLNqQq+svq7Rf2pChGnhB2UjCzMOZycMpVS
y5CP0LUK0SHnyCNmoAygLTGSq4fn+QH+w18ZmZv11+k6hcZY6RVy9WY8NDaDSXPjsxkITv2uKGTK
dbYaV2X68mtTVSvbM9eXgmZej2VaQ9ULWPmgIToz4yFrNWlcBrAwrPZDfju3PlI7tRsSXc7APAzS
WzMHLIJtIMZ6MQCndDa6ClN13pj3FEdvB9COxMwRDFqs3sgaIj3XgR7K8nNsd3o8U06zfvUIGLEV
fGaBhK7y/QqBKjs2V7yMyHZ9GZLXwYilE8caobXqC6TxiIN5RtUPmhlN99MrnhZdhRHyJtnuaOCD
RjX/enJAlv2gUgk7fHo21mLw8xQCcPE5I+4RanMBZigM+h2hrLWK2jYgsXv2a8oWlaZUtLoRfCdt
Q0Nacf9LXw4yXZp9EvMH5EJkeieUHlg+U5QUMdDSzBHW1MxHUXJ9GaprgYi0Xldbbc/ApELvqFVo
2cek/5KBCftfvKhXW28DAFBUogFetHv1RPc3XTMo6rWHm+jpNfdHy1UgCaqX66SR/q2+26/hcCu7
swB7uBXi9beBqueNLLLtsWXLGAg8i0UvZ1itCcJRgLtZMbnxPICk9o95SM2dq+xPGkTKF0KnKYww
hvdY4PZPYqjYpP/t1qrfqffOGOayd9ipmAOFx4oNpO0S9vHJbiG+Hdx/HDC22LvsevEM8dsRLVNp
9c9mYcn8LvhXW8nO0pJPA/c0SxyKKZQhy7cKm8Ab1dhM7pDg+UHIEV+Sev6IYKrzvzn5x6fHYUtb
wncleCFQVa+f04wsuwvkaM0/fXM/q+OyurAGUh/H/IVRRdfkEYoRQIr9ij9hPeJrR6tVK/oU7w+F
7rRcgVHHrLJsRL3cTeGl0MIU/wcHkcMJxC+MCWLXqaNTZQXB5bCaiKj4Q4NYcSRkI28XaG1Wo2R+
41YL8dzgTvfcTJ9a8PMUILSLPmIEgjX7TeLDnInZ07WA3zw495lraVJmaOx7n1P2p4Z8S6y8Kc2M
ZQrfwDrHLiI4jiecKjknA3u1GsWQBEtCaWEgfMnzl9v0byiJ+lrY0w4OwY4LhxPmOKNqrFsk4Z9d
1W/utOxc/Q4oTci5TPrUbFb9eQcboaXfU0a1doDk+/J8GN9qbwx43hJ5IQnp9csJfZxMwz5RN5RM
VrqaKgw3pqbcVGTnSsoc/KzkH252YoltEZQu72R/ofSF0Jm6iVpwtA06GFNuGTS9CPb9nGVYXn6k
PIq0++djVNukpe6Xf+6yTSSrSu0Kby89jsLuFsvAbNBqHakg+TC5MZlUsR+HLm7A9gFKdNSHEC/X
VxUXcmgAHaOCZs5m4k3OGsqVjd5VWYNRJlXaAhcWExgP8pektgwuB5xuq2+HRyOXJdhprNpzvJRF
37njRqfb0HfQ7vaY378NIUpNM327cb3hzhr52i+o35fqQuvXw9iHfWn5Ytt+eCAVhPrc3qnQD7yY
5+TPYbsMfLplC6uctN+O1o6bzKNcUSw/QDBk6aY85fwG/VPL7hT6bMbdVRLAYDmF1pybeYRgnrrX
KwQlf+pbKsPhGdClpEqXKEWgZ6uLBE4yqHtM0nyajVNshHLXgGgV4W5D8a9mjaw9VXaWVoWhBfvM
a2eRrRZHrdpkQs3kq6+Ezh6DHRq8rTZO+6iDnfsk1Zxv/VLClDbVI8ZdWxWrBwha0oRBWAVZud4R
n5m/FVYZ0Szq4T1y/6KJckVlg/ClA/7uJ5XCq4SzAfXDt0O1/yGLXZDwD4axmRACgTQYSOSUCxhb
xjy9fo/eYM8Ptl9p+yGdITLZ0m43//K9EelbFNMTl0FDXU8ZQ/zgLf5Wunt2V1mWTPJjI/u6zu7K
ws+kCcNzXotYVf/Zs7jEuQi1B/nwa7x7DuyQnPcpyX9ruGNN15RP6OZz1uTcmap5n+PtmdbPgGnB
MFgr09BBxWbZTwYIdPm5PIyLk6CdacxlyY7jgUsbk6CYb5YHh5u3BApuKjwvjKmWlPULNYvKU+Tn
3sYoLjNtj9xAhO9OJeaPUIvB2J/ASGOif+Tg7sJFynY9X2FFbyAzc3azXGXb7pr3ryDCWDbOM5ZL
nqvzpptP2QEwz+tgPk6TU5Nc7q6rjxgmCGr2BuKKpEPYor65VLehQBjFYHYLUmO2EAwQh29wfMJ8
PfLeJSiVgfnHZ35XKAvpmjW3JlxXkHayxvGKNAW16Iv1TzHbD34sFZqVP0aXpWVa37jRFGwH4ctu
ndIybdlm1bwhOPD2JgIq83LVAmG5wNK56uoFMGIBpPZ273F3xf5GxB8zfQGSCaoUzi5RHLqjcm8L
HC1vtkOY49up9LXN+Dl+xHUSEaLXTibrViVJ39GFPyP+d/5VwVX6EfsILsoMHvQwxNpHSSusLilA
XZgwB1QaKzT8AIBpEsZpqtS+29j7nMr/Oz81kOHwxduRW1KYqN8smPalz1yU3CbtwSL96LOi+8gW
sFTjaFfs0dZr+OVyU+TsRc2/3ul6q+Aj64Ew6qRw0MjuRS8qkWXr+t50SMeIxEGDCeToc2nvbWqB
06rmJfRHQuNrUN3A77dAsxjDIn2Rz7vTSEFvAA2L1zcLIhWlHcPIoDyXu34fYm+RiPxa2Cm8D1o/
h9RASW7Po5P94IDTh1r1ZB8AdPUj3jckntbxsdxl9enpp/L5KPsBNi3p1Y1W9gXeqN0E+eGzg/tO
b8lVfSenjgZ2I2uMTsxSaVCA0TKk40c0DoVAt2TP3FChsPQKvsmvPSx2DT51h1Cz+jk69zw7FiL+
UWrzl70AeaL9sSrSnMkU4Gev27ScT96RTxsfRAlOCbiDBZQtStzjMQaBXJjZbmGVqC8eZGQhh6Bq
pbTyQjk1dou+8HBjOyDfe+mcb34O1iN3qStlYjhwTi7Y73cKmJlWwssRbjGLXAxm5pu/2Gonydtj
XhvzAOvCREUSXfXRtcgwJZ/b44ZJlTle7JI1h2fFqQKuEYO96YiH+j94HMdOkYoJx5g9shG+UmPJ
T0cNgE3FHnKm+8YGNzyo/MQ5gadotZqxdMjkSzLQ2Ais13KMCsRsPmG6uFTw7SQ6mnmC1x9PYv9C
c9MrOahqu/1AIebQBtSuNWTrxmFlqYcHad/V4KsEqoJ1JyWFrw7dkckQcX2AM6lBEXQDBBIhStVp
W5Ki8i2Atz8d7K8Jy5Dea1WfsYJtV891MT8d4R0g64BYHDDChxPRvpvSgB3uzsAUn2dhGilBgVRW
nGBxQ3OHDMbXDMxOW40wTlwiaCbURlzWhmZFE907oOdawboTarcCTwyH3y2rGcG4bsxe2/2Vl746
2ATl6gM+mWqvX71wjDPMX6AsGtfz3tFeHMeuWx7YUYNrhmjj86TJcrLbfblYdfmxSY6ePTiKFOQP
Iao9syjO2M/NpofQsTWjBN1rLgtonaVtHJDzal8ydsJNO7mMt1rM/+8GtF5Bg9YIOdv4zblQX//3
p8cNzuXLQZm5t2TsimNMp2Mie74rqwCQ8dAZlFviIeFEYgggulRUO77pNWH6TP0zcApeVtMlrljI
+Nycsdb7/E1/ahkoUH12ftKt0zyTbHzpZx10Bmu4Re366CLO5FInRO/hV/G1sGeLjC/U+ISJajKn
3WBWwkqcIaL3VG7MV9NPnEz/TP02oMtYvbj9jZeyIHweglRRJ+4p8g4GclFEGMrP67jYuCf8hc4L
Q5PA99XXqc1LCkFc/MHG+vkJZonDBgKcPL6hjuab6y09INF7ExRUr22m2rT93B475en/VPK0fLW3
H7pK6Smd4fTjyssWfTkfBZfkV3KTtivxwDw6g5xGoKx7+uKAFUo0oHi/L7Ks+JjZTmuqCv1V1ToD
jseZYRZxpjAXX4ndf3dOaPHFzOVw2kQwhNp5awEUOHghPPYxit4PJ6KwIm8ZlNessHUByiP7y0wy
69XE3AzI0fGapAsqtWn88+RlRbLivLV/trG+jVGtF+h6+XeO/asSNFzFZ++1bMMRhZf3Mi4ClG8p
Lqn1yuja+EBPbY7m4KhG70r3+xON4nJwehpHOvKRzRuucBjxExwQwzAh5xowzo/42/lEWNDH09Nm
nCUlTQ59CB1NC3CcsXWpgGXTq//B5ktNyJICVF58czBxw6yQaaUw5hWWeI4vmuivHyqjudm9jinN
3PLOqxQrLm142E9l76E8ZqK75TM9jRokdaXcUGx3v1NdWeoYD6k+a541m80qk9tjr1LzQugaXspB
bYRpvCqshDDMhJ7UENGcegU6Z/bHaYeBIn/jRD6pwglWqBCY8SxEtSFEq+VX+MPoqMTq1nViKHVC
P9yTywzfd+MryU8Y/RS87xkw45nNQzh01w1pGHS52Fwy3W0at85WkILrOpMuTgpuvS8SXDldaU2a
q7bHLA+kgp8C9R6JihMtLAbUJ9iZw9MVJuw1XwHl65Iv0ZmJU3+b7XFr67fWjsB8a22asU5MbqIe
Fer7EQXtYNPUJ9oJSqU2jCAdneu5q2SCoQKgNZvJcES4+U82lpIHMpjihV57zVx4P4cxfMxpm5W4
quKe5oAfVFgcmjtyTejacSEJh3mNQaG9FnuQwaUkfXIQFx14+P23jA262u2p9r6WTo8JaimlJHQo
8vj/nbwDn2tHljZYuLKLeT6AZx7w3EDP2yOoHD1tGtSdgvJsE3YhBiWjgSA2IyRmVYKXZKzojpDF
l3mdi/iVZCTG8wijF+xvgD+5p6yASnCWeWfql7hKdBD26CkcSqGlWUw65EtQRqAaDQnBhEMkjfsN
KascOiEPR/VQnb4niZDP2kqPlHzCVgVbc+aynio0EWhyPFLXZHgL2qKwAMJ25NdnD2RhMXKm8Myk
6nFR7sz2fNRhqYxDfV5E3OmZqBBO2lgUJwsUTimm45h+khKX+WEcYm6kBb+GmftGnz2XWSEwNOt5
dN8OgVnDnRyJH+JLLB+M7qWtbmFlCOEIwdhPOPFX2Pf6W0DOsoKYLD6jx0Qm4GnXRCIg/rIprfr7
e79Rz4Eie793YhDNuBLPRBv87OA8/XBHShl3h6HNbiCegG/djgw7S2chk4hr/otgOXiE5/rJlJdF
X7/7XLFBhhhS7FW55Irw8AkpOXozzBkGQGPAJSme8wKWl6aBVznwvpi7TTtYf8n23eLjnM8/6IZ1
/F38UZWVJpyMm71WXIjb+3HOnt/GKE7s188nav+/pCC67796h2Zh5QgTzvGnwGaWF12jmnMZrWOR
AcgKvUIk4KK9QJGEMTxXIt+4sS7aaW7LBCvZecmOIU7qs5Q/Uizra2dojyIJ6WOv4Km+/webvSYx
W0BA6OCqypSW9vHzoQuR/Urf0wen8a5vveyiPfj1Y5qirXB0PhL6rziuPR9BMhL5MGAvdPmsVDGR
0iCA5Q4HtXT5CZHP29e/Iyof7bnotf9+soHq+fDXxy7m1HC1GNRmfrxKAFZQnSsWLwf00Ez0y1HC
JL6PDWDOr+onDHLDwy7hsZBn/IxLULA6hKLSCKp+MWc7/g/gBt60vBEOnboIyE7E3e8uB70AZpZd
ByRZ8FBf2sbgM2K2qsb2baijFXll+0F8zPU3BNhQ0jQIuE+3cSmMUB0OR8eNb8v0wa69PS+n/tWS
HdYe+GDi36m0qJsjwRqDW5b0N+8no8kIZumKsI58R0qW8SXrzdJiNBiuRUu/+enQKCL0vuNEk8MN
cemYtm1rd3LdAl7qhlCNHiYs7qCc/d88O91uWXJZMzsDWFzBD0RBOp9LH3e2rPnp+ox5a5dsljGr
ujVwHqAXhq8AttSXQSsk8msIDnvuFYoZpGgw1jSIqt0kchr3rh8lO8XVvfxTqNEWYNs7Dp7qSx9N
K33+H0PhEckWP+VPKDF2qaAPoPzgQMVGJhX8j6ZjLOLuNDi8R0RziEG5a4fzm76s3QAe59dKOdTj
GhPaibEQFiE3Jpj6HHiynjii+gs9TFAhTnmLTmulbtF1TFUY/nQFw1Ev2xLEcPctuOR6TEBwT6GS
//Ig9Wbmd0BgCC2nYmLbO7VmR6vc/YYdUihg4l8vszPHySDSaTSk6lAqwTNvoZoD/f7z7YFjU0Lf
yxX4Nb4Cz2rHxO0Oce3mTfWC1NFvJHYj3SDI/F8XenMJhd6aP61w/ckbl4Tl03BMePPnNnEiCynh
Ur3Ijs5hqwiCmRVMl7mogWZljZNZCpCyHeJYnkMabNbImHYh3tfuA3J+ZZ5de1kRn/oG0ufp9qXC
boTTvEKjcEjdx9lAdCmvN9uXaIv2lFu5uwhcJk2ZVsAIpZsp7pZJcIJZzi0XGu6duQEsNO42WVMU
PriwCRslWwu76AwzIMyHnD5Vx2SFHo71LvNDiTbOyfsTHJkZWJ9xfZezWaaDJ9mHSIZq+T4jBlJW
PzvmiWNOn4hiz+KqRTo+Hio5+y0MpJny/J6q0nPXk4jH5ZRf5IK4h77eGMRUibTSmN3t/MAsQNOp
xF5oGmvsnBHJhhvCFRo07DNEvo1K8apviOMlPExg4+Q4kHKvI87NFIxbMXq4Np87+Tu6+n4nraOf
B3bd/PQD+r26b+39x+Qs3lPByWVOLfyfs650V8IMDbU3hMxGXDeeGrqjb5WiOeoAbTWVTQhJhAjX
niTHGA789a4vBLyeemjGErANcgfY69VEUWP043+/5Q00HQ7JtQOJCWq/XyQ3scV1OvNOQkGz6JIY
eSynNJLQ/5oSFkdc9T5ssfL8B2tzPQNpfGeCc6BVupq/9tqJiHcLxNxu8JQRKnIcoegNpLE+LDdJ
JVzyiwtD4qYcbY0EL6OroI0T7tNGKt003UxM8RIxYh0W2Qlq39g2jRuBAmGmQ/FPovGQ364A08q9
JEiUGEaiyWhG1mHl1BdiP7clRzUG87U6VY/QRzJqToVIS1ugHKEPZ8YPRB0F4rlU4+fXtIfyYON1
6Lk4kwgBCXPRGYJsBlY41m/bWzQrUAtP1CquGKQb6ZA4NpLtcRYDMsGfCJizLNyJqJ5N89s2aJhL
rFyF/LR6JDZXaPxjUJeBZWD2YYeiBeHWi1hRoGL4wTonR80ScnnjEwhuBSA3qOdXNMHLcIrOS8AI
BPgZPFzGhlpAEEoYSwR7msIZHgJHbSIQoOPEFQqeGFRFYWvz836ICuWpJFL50Rn9m/zadCbi6Qjo
qiBQZjcQD5shOdSO7QpTBS8ZERFyRwtAO0iCo3/17ynIiVy3oMsg8IFcQ90YWWVv8I7oa+P8BPdl
wlnNSODfGLbTewpGCQ1AnFXuDcFNEcWZ5ofjcZt4DhPtUNdrpNdiWPl9LtkrcsIJs3Mn9Zq8/WCn
+SYQtp6Cv5haIhVliWi/wUf+GNTWhQJiyOl54beOGVybipVDGJgrhROp4FAQRS3bc8lhXIS6WQPq
e2r4yLy3ZX8c/lkTI4uwxrNrBIlZCybhWXyNH33k368rhYKEIysyODEisrzpw3krTo8PsLvuY2vQ
fuzvkMqBOF/t9Jc1bYXtvO/ptK0Myhoq0/vL+Zvu3BBXSIGfvXrI7HmnPXbDszalz49RXS6bL45c
POqcTQosjqrbcv8GcPT/y8OA5E5wCOlWsrvbRWMh9hKXNNmK/WImRfKGigP7xiXLjdqIQQZlgar8
UgigbF+ckNcEEc4LrYF/gr7Bu2Wi6KtQEIhLUyLM+nKEEZHtcf/dPZ8WYXVHUDW4IbZHcyrCQbY2
P9s29Lrkdi2E+/34le0g1P54Geqi4tYKZ8IzekZQTyEojL58bf4h6xMOtUx73VyRoktf0Ozaz1lO
P+tCCeao3XSJ6rLonkm5SXQRnQTzKtu0F8JigGPXqsZvfnzHjpnJqhXb3TOaTG48njGsPv/23U7w
IgjMT+82xPufXWSXbSt3iChu3sRB1Lk9g3LJByUGn/Vsdpi7zWdPB6QpOC06S/Po0N7EZx7y6lKh
QnyivY3BTzdT+WDjo8hYPrq9LWAY4JCnd0sA+Bv0OXkXtrBRXxowX5PWLyDj4CQRp/MStKK2OSWK
4dqJkxKX+ssmCwBMd/ZXMw1IVzbwqdu0jhQo+6jR2tyzWMtX4NgK8CrTqx7Jj8NKCZl7Ryyqcwfq
HeVQ+zuqSgks7HGgc66UYgq9OOHyqvgwQl48HGuOQ9Eom9JKmoi/V3JAmWNrUuO9+u4KaKt4lu5G
YsOdTX/1BAFSrNPCBcBt97i2UQJrZUvqABUHBlgosmKIBb8PxLaO3UJpluGnHEfTP8fM+mOwHy1Z
uAvlcXVrbvfzl05RUIoac/8faK8OJd/1l3oPauAn3JBGOXh/t6wd8llnMfTsnUSHnAjcoxEpAdoM
vOrNGrOx/HxKAy6KvRkgMHZ6ZcrZ2xPgwE0mg+Ec4IBKzz62uOrr96fGXHPIqfM4e8PK1MPTfuPg
AB/cicXTtHJeKFOU0BtGVvgOKhpuXHNNjv2A6I4jc9B4oD1JXcSUuGNDF2sWQNyt4dIA7Wgq312v
R4NH7NMgUBjey9fpbNxKFBvQ1Dvj08TFjZh+Iuq3Snc7nCKoB+4Y4so2j+OJcW9g/VVsio8nP7yx
PZoEv3UFuysyo8dmlHgtlFUSkwpGwa7e2ed0XFqh8iGz/4OG1T1D5V+lqdzd0alEfagLJLCEnOBF
gkYIlc/bUJ+S7lOhJCf3u7RRNj7oJ6BzJuub5LhdiYLnqC1aGz1XWchDLfuP/4Z3W64+UQnOEdiX
0vxg38N0vXYAakuzQoazbYweMho3fFSuaOAWOQ2QRLutj9UUsnPtIBdnF8A0QTWey4UVLfflzs2Q
p4Yl9GSDoKVwHfeaL0/IGkdUaTVD4xoCwUE4s7StOfsUmkn+XGngXRRBEonwTbxna6Ul6brycbzF
/YQacbeuTiJ7fCsgs4joY/Wp+tjcZ347XQjnmUJSL45lHiNERvpYN2Up0PJkiISWAXP4csljtaPS
H3wDAStSp7FL73lidunvWzo6GCBvW3O67ItnhOXWcBbsFQ6WsSDC1MRvJ1wC3uJAHFgSGavVKXf+
FemOwufwDcJsgEX5X7DJ0rq8NysqoetcYqskdmSnFOKC8rUcg5/LG15GOg3gWLef6+0J5GYVH8U8
8nPLUetY6vmqTDY4K07GTKP3M2D/VdiCgfTlS+xpRmFz7cxpVB3Hv5WuIuFvlW5Ov0C9WHnQifCW
/FicaFrcQmJkKrbKASOhvUI/Ilk4FXufjZeEEU1JOaJ8DC9uqohsaiynM+GRiT85FET7SoZcXloR
xVEwHFB2YvFbGMoaqm8QvHTxuY5MfsJhrAi8gUlpZ5imilz1dRLFApL01B6qUzH3dztys+VK7mN1
swOrNEuIAcoTftlB7JLknSuAxc0r0TDQVrDcWoAGCG979X9+V6Zxkp9PNTSni4cgOCXqZgg+Dqyf
6xJvGvrS+GPePSTmbHcdfKtB5PjkxSxhlJ7RxO8H4Oc+HYmbsDzBBrP/5Nf9/oH+p3HaMdonOKC0
HJVv4FUQ/DYZRM2SievrurM/VmqQPIQGmVrNlWNQa8+Sh+JpwCIPCNFZe6W+Oi6Asvl55XGjvIYQ
vo8M5G2rivMlqVHfR4BQC22VLAasE24ThjeM3DYlpKMZODt6HmcCcomFaeHhUB5A87VoC0frCXR1
1SC7W4SEi6y6DGs+cHBvjPxcVlcpm8tSqPUDYEB7uWqEUj4DpaGoy0bd5c3NhVgjIUyl6y+v15k0
D+ruiXdG+Ti2ZE0wH5FwZH/mOI5DxVcDqkUWAQFepSTEnA3slnH7ZOk3jfugNPMv6G7b7QrfHzyt
6bjgLm5qz7YHxIzh49vUROiiBoyYZsvor7vrvW+YdHBrGCW5GHuzkYjzBcLAMvKh247TIBYjspCM
v2+IT/nWdC0Ar4EuVZQX/UFZNOF6POyFfE8XdNAeiUjAFWty6SbX3AjgsmF+gwNcFW84DOok53QF
AOhL9OOLzYfd/tCtGkwbbXH2tB0HfmIyDjCcPCKTbcZhxMZVxvi3OtvWLQvbUmtc7wsLGFRKcMaY
E6ciu/ulNSLD3X2Vd7jbrifGrx4OhHC85CkYMxx+NWvKfG/fAE6IarWZUTOTMwUEie7vK5Cb3KBb
P0rQtTshIGqJyT2bikMVpvNMc4EH4KXtilWH7HJJnMOenoFAViER7wJSZstOP5JhP2KAID5bn4i/
IxS3Qmn6NcwG0ZYnenx6Ix/u5TzvSM/gy94Is6Oc0VcAXi6+DFb26P6/KcwW79xFMnvsU0CFK+yT
J+lp6GTgWdbCiYz7aPByP4yFKP73xouUp6VX1JA6GRHCCfYHAGIJl2gsS9m0YeZ+U+fOM2zWlLjO
bVTVEnXRSTJ5TpUj41u9BVfx6Go9x/yR6V7XzyYeEOvvPWCT317WuwG1LHDM+K1IoO2WD5KJgrfE
3+qcTmn3QP5ivbUNXufmipyA6Ujtr8r8tE5xFSjbgeG6WFhosH92uZ0CFmRuH3jpaCk/IKI3Bsl0
75woAR3LieWFU3ml4IxJOeUoLsvszjZi+xVsQ1ISjkX321pMM1YsuxRCfm2Y1clzfw8Ob6u6MrHY
4Psgxj/fSQljDEtz80W6V9nkMVdJ5cyE/DgjM0eUhKpbdbhad5FJRSoeKU+PlWkr4awXcvqVXlkF
Lb8bmnk+TVJ1MOeD2E9XaTTqx5Lxiv9h/AvlsGHvQ/2YcEypWJw3GvkPpFyoYbFivMYmaH31d4bt
n0muobgEC5Sg3SI42h0qV+FdHooBgsZjEDqNv47r/XQVzqiE982uAtrmtOMVH+kbyNqloVXHZ+F4
/gCnEAvy/FVSbqyD8tWpwib8Q5EpTIuwc5hRjTGp+QR0DUzyZBHuXHe8Ynf+SasFN3XXIp427+qg
u5EXw64NYbbTsJfFEJEZ/lv09vfTiBaMuOxobGUjRpYS/s4m+dchuCHD78cWuYpIDr1oTsKcw6Xm
qJ6Tg0hN8NqtP9qtOwTF6GR9il5OBtzX+CWqO2U1xzFUrrDtIN5yslNFexJ/I7GXVrKV8+APRgz1
SKPLOK0Qs1yMyn2K2qZRjxhmwedJAAdzQcyFcGLq5SqLt5UBJNyQsF0cgf7Tjgc5pZbJTLXS7xDQ
Q2yemzkqGj73PtUa3ZHsDaXM0SE4wkC/dgAMr/GFDjTi3jUq6Qgsw5au9idrcjTrwW2xtFwk42UE
qr9w9gkMX5/9EvB3lIj/lRh0PWScO6izR1gin4eDAR2vt+Hj1TBJKPPIjXkAC71V0uBfCi02fQ/t
TY+XW7r1PttN8R/pVpiKxXLIyF/AHLskla+YRIdI9N0+2CPzOcvdmOhcYO0GSfpbi3XucXuqbvcT
joD6DcpPnEselgdIrjte0KhAwvA7ruMTbReIRV1aJ2xjXLNPLJhjKOHej1j1uwzXCTY8aRzbSEWM
1SoR4jFkxJwCPrKkTkHz3xZ71oxQST9Hdmq+yo2Vy9w4WqTF/FwjfmL7LCL2jtg/6BXFTs2Qblvr
bm1Em7Eb5z5kTBT8Hc1+BwxevPp798YCfBl1QuTJGhwIIxZi0JuQkruunu5ZaNru/Y/mBHGNZybF
CgdjmSegbeYwTiob53GHv52o6Sh1McKNEHY6X0YFPOMyfXpVYX3ZsDnkK1oiVCPC9D2bVGPO8w1I
X80k+YUhEWOzqg9+xfL/Xpnbp92xVyGOUTebfVol5JwS/6bfpXLiCMCL2k/RE+JRMw9xgA/PlsKe
fyj8Cfv8TUQP/ZlgTbBFAC/FXJbXK3OTL+jXNAuX6T2C9iyfB8x/73MeAkWocNWWm0kp6hqBAHhD
0KW/PHjStYFbeb6xAGZrsh1GvpyR79QztmKKqj8Y5LQfGXBHzMK771wfrwELqZow4yAqKgTcF8cU
29/ddvZ8Eta3DRXQVur9Pvv2pFhKNjk7E6rRMUAHoMbFNBRrwquX/IpLbaQFymXiwj4m1xiZxrDc
7eIZpodbN3U6J4ZdM+43V8ZdJejNHK2V1e2G0XiydK6h98iti0jWBBONtdQ4pzjSGb3h/lkHGTSc
UDB0frMXuQTBSMf2kC++1h50Kg6jRaAst30vuAnVFraKVD4rGTG1PhLRj6su7a4SIRzxwgzGyDL6
oywTJYeRPV65okgZXj9SNd5sxlw8BkK82QPkWRrDxUL35VFL7RNhXN9FcLZd21YWmIh4GLrVX6xy
veLoqS7BqyoT3E7/bGj6LhE4OD3f+jt3zm6uyUh0UuM5hQp5d4TsPQtYrpthlzMfatUwYY++h3Ox
rZ9G4Ugor/sEC38qdjOSx+Ersz3c7HD++iWES7LWgLGzocjbQIXPyK/EXoWeI63uFj4eRIWwj8rJ
WDPlVRRkDf4ObrZQlA8yfstAALr19QYGxQ5frybuyrB3tbHT+rWmQoyf4WfAYrsMoAcOBIPJPolj
8ff6TlNi4mk9kFj2wgez+Ap8VexrUUJgIQMwxRLvlsALCZko3fTwh9GsS9xDU6HjeXAeYG3xiha8
sIrmTiQkLMb77C/sPmpUu0pThjOUpaGAITUpI6FRc3W+4H9bACGMWAfiiBi/JPvqI2B/evMvdD21
ydTgACxkdrnOzay5zS9W/bzogjhFheFqQ282HMdQZwtOl5wNlDLroUHMOPskaJm9QJtj9gunkwFo
2jT/S7KfX1KQxGjarlgAksYW46I7vLdDxjH8HUNp5E7mG5edNJl2WtjAE87y7UdWtpkW3CkGIt5K
Z3effwUvh9c38yXGjShwszjFD0YnS7MwGDD6jWe3d/HJRoRSC5KEf+WNWmTuhYacyO+1ch1e0P4P
PH1N3SEqu1szxB2W3WkRdyuJphLaHs/gG9wKvHtftyfn8rwKz7Mc7422WAzg5UwRAK32iKJxQ25J
L58PCSrnV95aZI+pAx9xiU01sE8nio3OR5IEw3rPa5IvOqn9XvL4em6MgMonqFxHc1ZEixDZJpt6
AdQOCxSTZFTMJ6BWwXIhek0wgY8qTsCXlnUi6dI8jxj5CvoyDV1MdSlvNpZfI0H2lOw56MCtGRxZ
pP3BUzdAgbqq8T+OYV7XLgkA0kNGvY9/sanmKfHait3wJ6yiU4fQse4o1bempZrne8j/bIoSCofL
Y+y9jsF5N2spJclQhaLdmXOK6M0RWZtwX9lGgCg7yxpxcR4E0VLZbX4n+qJwqifvMCFDepz/ppwD
/8y/oo+d6NbA30lwFsxviglkG5WQw9KwRHA+bWDk8PhkeOpCiCCGI8dO79tqjkuXXl2HKqyOFyXm
KKjCzbBsMFhaLS55qMrpxt+clb3TRDhcPvY1RNnnmRw/8rGeig776OrQzPleo9tqYz8L9R56LCis
FvEeXNdDqjF7vnfJ9w2+fLARA5DN/PSJBiEvoFzg/jA+e57l/Lt4ZV2AX5PsC1lTL0Ij1aieGlRY
lIjqde/M7r/VKosZ/Ntq5WHW8s3F6pkuhUOJlfSvdhYNaIIacziI97Nt+B3Jb/Vh9WKCVEcQVRNs
ITL0CS8TbPN/m+XaHdGxiu0JYxE7LZfFP9HIodEsNEvfs29vjlC564H+0hIF0t9wsu8PfaQrbyDV
eS2giinQ/ySj8dFMKH6wDOSIa2Es7z47m8z+70EILQSMFxuH5KGXrH7/S5uFMes/S/yhMptDEcjp
ETZR4m2T+jM9ICbh72yREixvDGzuWuPYbtl3AuPhooR3ZQ5x3L5LkmtK6H8Smk/jXMYY+O/C+l49
U8e0P/YZWit9l4W2DMe8UtKDBdGkE89hQXAx8QNU4znBSUakCelVhc5fBFdoJSp4hpt9whbMB2Uq
TCYUF5rTRYz3ks66fTTDcssy2DTCmVAoq2fIWI0dvg+o8HhixcBjELO8qXrejsrF0aisjGY9wP8B
gkiTQK14Y3MsfaRBFtwKowMoaEk80ZHSm+4m58yVJ53btJbDCQbG3AuFy+TFKS1D/7sdEqmWbaBb
XlfVpxJHtre7/URo5CgOORBeD8VkOQpdJd9/DNCM9b/VHb2EHkd2f/SISCpI2kXPQPeyIGWnEZR4
0YJoOGF5jt+dXIDbmBXX6qKIge9+f6cVKMfo+z4kKgrMsmfCaAjdIkVFR+NXa4m12djY7jwRa37F
tXBxnetnHzK5x/p/tVvnIvbDx1Bi8Ae+9UpBlvkbX9wHcAMIatp93Jb8oJeubpVs4/BjSP1wngGo
sMVgMBh6Orsk+e82xbt3T5sddOrw5xOprpqY4qARhdvPtnFM5jlBSb87SrkLhaCWQU2nyFtDJWQA
AIEzQj/CNUHCRMNRsao6zXpVD3OMShxCwaIdPjfC7LQ6HT91QGdy6jq3UX9fbQJ9wWyBPtNn0E/B
x1oNObqPWu6NYCc2wY5jHyAysT5YsVkFA+cPiauMbYVuQ42opq2lpJVAAVfP5JRKbwipF+/8rGcX
gZSyE/pVDMlZa4MyLt0cvZ2Hm6ysEduX11NTUUdy97/LrnGp8zVS05qhLxmCUFvWUXF+jXDv1qXa
VAC9TyIFul/KavNB0wWtoqBoOrUF9QGnhNUBwT+sgRlkd32YlWF63KMB2MntxLRQXEfl4JwADKeg
cXwgH87zD1XjAksRk6X9HsLEDtcWH2dbZoiC6qX23GbShbtzMtIU9UrQfYp+Q5VTmk6bQIj05b3i
AiFbGuvmlWmqcrd9w+qHWAr4Qk4aP+/k0T2E5HNBWoCYgyCtGZClfXST9/Zr8ozenKwdpaDrTMJa
t0XYgRORBhApwsaquJBfobbx+t3qVkX4QPGSY8OtK9HYCoGMil51ggv9RzJ5GCAw4HThzAFRJj3N
1p9cxAEeXktfdJ8DJw5VXCGvZeccOZsNT2ttqSEaRlmu4lu4CoXQWkHmYkGKJ/vbQgU/zZi5zGNR
IqjFZzQ0nD2BuMktEQJkwXy8VhIQabjeGBah/RoVvrG2XKXwNNKA+PX1+jR6OdF0MjKxdFJxH4my
uZw1K6Z6JGnqB9R93v0yZC5xbB2YoUcxgd40/93frZCTnD7giNLy3WlSO6Lmm9TaiKTglJUb16YT
dhvVDGTYbrh0GaxyfOsHhDuDyub0TxkNyde6OW6kdroDpgmMle5VKhKQfZY67ea7m7EY20BFe54K
amBHyM+8VR1mgkKAlNq5PjAE6kmo5yKKLCLpC89RJCh103XrF9Gnpj9Lyc9wUkBiUtcLqQED5dIF
34zfMqCW4ZdU9EduxWcHrrTOsmyzAyp66cozDDKzJIQv9oDvCLVwFc0euSVn9RqoYX2qGxuEGj/9
3uzNzTHifQYbiZqsLt2ybdsoJJ+HKtNdxKETP6jO+Tb//8PRkvtNn5VnacNpcO5RAX76MZjCMHPD
wK586Y9SqAP1Wr9wSia4bDZry+7nIYUgKwq+Nn3v9KJK2gmGx6YFxIe07/svGcf/KY/ALx14Pe0F
wXvGOixah7umi8jkD/neP0dsAHwCf3F9dFniLUgBO5SmomkrDKaBH4Bl4yCTkvuqi95ZMbLPFDBf
KrC6Vi34B2nQqQwqSDB26onhXnqZOVNUfODtutXgJXy0mPJqU3JmESJhyELBXhi3+IJ3qbg5k2ft
oebQrytM2t5TwQ4OIDM81QCXUYBo6OluYO7OGkdpRvZnnXwWItIdBOkZdHG4QL7/LeBmzF/5wjIL
+xTdMYnOX4/8bv29t+nW5IdHNlOu63DNr7SH8VqPnB6X9DnBMLYOTgDDMtXVgYnB3tuWpMEqL4Q2
BTgFx6BqP3jE0pY+V1J/K4QgcWHNcKikH5RYAt5LUdJCWlSFJg5Ae0gjdWTjDaG/vXi8W5sOWDfE
wyhoqQPRB1UgOT4UnGz6qco9D06mgYlUtDewclNjF9zMEGVp4uA2hxZUTYG5QtoHD/+30JY7qsn3
WcsNiSbqFGsOPez4RFfVfxrNu3ZyTnuVep/ptPz0zUhTlNlv6/BCnX35YNMaWEmkxOaZ/0g4U8aD
7KlvGbQOHexgNidLOWxevBPad4V9ziKEjRypntAnkrGpt/O0yL6mQjdkAhJNeYPVr+0+idHDzLO3
6qiHErMJlDLIqaMRXUGvMDIp1jwbEjwzc1W/djKqDflp2V9MMcw8/jjyLA1V1c5yWmB/IMFN/aMp
fjhvgr3BclQKA+aLKSHmdca0qyoIJY7+JG2xTCaE10M510INbrdoTnlPcZMIyvaz5w8mdOD1Sm3g
XeZbMg2febYtXEWzS1ZMEwxN5vPQDK6zk9a2dEXbvrMjA+cMjGZ/YpUW5sxs4TFX/V5QKWyaQ0Ro
pZmq7runj/Fx4NtDQLj3qnkuUu9eXWut2JQ26+6sx8HC9drF1kPGyOTveUq9mJEEXuDVAJkZBenD
T132cRIB+blNQYHpb2j4P5MbxsDcH+spQ/SUXeShVaZZbXjf5aP4NYoHgy5ns89j44NFDrps32Lu
Um02aDOYTbCN/hh66m9jSs9y3U8K4cWOAlezhc9QMVnD5TeMfsJdcgwyHX6jpTzYNnO2b3B9JqB7
1l0mMRmd+dsx/2cf2o4KZkZqRkjOA7uJXtxSr6+okCcsQRR2XLJHNiBYtdY/IJAHbZVdkcv9oyiG
DpTUu6UQf/Mpx8lptyFayJCTwroyjqlDG3DsEmrzUcAOuIgOULsbmLCSCkObFxGKPZmS3GUONM46
UwxCcuwRLf9g1WbUo8mN4msMDhPV8akgQySl9yZtj1W58JTkBx3Pm+ebMvJ8FkAXgZQuxWw0XH9T
F4VfOiJsddLqxOWZFcFsqKMXxnWWyNfChMWEj7JU6VSWKobUjKkW2JWr2UK9fANIcXh40r7UavqO
V2ryGgEldPGIYEseLVLxuNC/759o9lJymNeLRSGzJ94nj1tdWLhv1oWGGkKRthyH/a+bZBKfMEaC
6D5tCvh1+y9cYZWRT7v/qvwZuOP2QXZ+oV7zKBSir1fY5XefOMubHFBXYwYZaHenUWqIcAU/EgW7
j5qnXU+/IJ8uM7X62WVWw9rmjNtxVckYqKR44VSGFNWY+MorjJFUtesS36A9il8j+L/jYNn2teie
1Not6o/qfq/JKhhPSsT05wlAa3Fjph7fIq0nsz3bYv/Qmf384mXJ9ik8wPK0x/csmZIYRwCMAsDT
wZZ68tBKk9oytZXY3dUnQuC7NKrOYBFCQ8bjSJzY6mpQ+UoiORJnxq2gI/RQbpcXIN3XS8U6TTEC
0ToR+YCeb/+tNxxSSDVAjJ64rnxiBUmc9uG1h+6ZJWOeZ2NeuRM3ux+O6ehqmuZix4u/+mST65e+
rhTCHcPmKacA1vfkX7EuSTyB6jIX2OpgqDKPoZlbWTWeaWernfEY52FTUlx6NsTqW84cbKHH7RV/
mJt7tv0mIqBPYJRFE51ONTlzmwlmqFUGqf3fRmkiVkkr0RK2kJQlex85hX1omTmeH9mn7rq1U1/H
aJiW1na2XVsk96Rl8H842AGeGgazYLCbT34/tjWSXT5wungYQqhyLGxIRrfQMgV0my+sulhdiymq
cQFLBLo24JuE7CbQlVyi4LjDWlRnkjwXZpsHhBbXU6QJur0OhGWlO+uUjSW1twLc5MRYYT/papf6
S4Tmu24poL/VgyGWxDOCaEy2arE6pcZhBfWsfo0fLOS9FwxLeyRnjsYKjxMgvCMqCgIlo0l0M0X4
XX7RcetqG68hRN9hJubTmkFmt+yFzNCGHU9QInREmZ+h4ISR3k5575v3kabX2WJ/KgDkdO93I7T7
UZ7HEazSgs4ye+X5ny6h2VzTXT0NPmNnHf8i11tyRsnDQyIB/4B4D84j1N0jvLcGu1gsZEA11oGp
g65vi5NNld3WlWgk/N8a1YTAleH6zFGw8IO+Lk4NLy4hTT1BC0QAaDtYBGU2k3pRRMOgmVkttbrO
tqzNg5KvPMi0tBdtDjyCdCrrYuHN53v9NDO/LqI9WhDFwoC+EFGRfJmIF/FDXO8lJCVxqawY3MpU
UwKpFYqHe5eR4hbW+3ypSbwDE9LpxrVuV7eWhGYuQIm9IOVQsCsWe99AaqO2fl+f49NYjAHsPDCw
5FJXdPax0nF8c5kA0IaB9HsiVjT79CkhriiruETsr7zLq1b/R3agAqQntotiqucztCoDx+abM5n+
sU8YvT1eTFwmXwIRGT94PNgTrNIbMBw5CLTemOyRPk35rQKdXLwt3o4NT1Kn9HlBlSydIIvUvRqQ
13R/Fk4p8VGBZng08jpUqLEpjorsHOVeubCs6apnO2JtPq47ooiHR0rmb0aAe9cIFd78ySIiOOe9
wMvj5QvLR4KxeDLMLpob8cj3lCWBqvtEgd1hP4Kdrwaerq1LgTD4RvEQ1Na2tUi42jo4s4k0VCzj
06pV1ncYzGNDzbn+W6nnYnP8Sh8IN4fS3A+PbrrjcFY88FddkGDxuI5LlX3Fs+9QlprVhNSonOjc
Vng+DLkhQgnMnxIMIN40UWstleErlVUDndjufWxZzuXwg1sxWbTcywLIWcA3faoArCPGd4X5iRcX
iOXcHnCPH53d3orHMfkijKRSuSm+UdFxhD/W/KxW7itqmY+iD/QgV1lIeaZSM+Rh79UYSdSuBJfI
H+Z13y0jt1ai/H2hcPPY+d80jusbbLX0lTDUZqwOsT/KJcKzNDj+G380MI98K8zjYatclgyD0CmL
Q4+dBo5cFTNSgUcVbVaG1zQmE/B6p4xfbPQafxZEa9UHbyziesIje3/jW/IUtzB9tgbFDgP/T/LR
ZGp3WCx55GKRVHX3IWNq7HpKGRSl+F7awt738IXz2UJJPrYy5kk6AygskHYk6QYVEW72N7fXMKGQ
YPHAJftYEYuQ2PUJCm7p58ANbnjTvTQVrYd1BNs4u7Xr3DsmmU+vUey7EVSVbs8vNuKlnM3k0UN9
635jxhiRzwhRqGnZQwddqGSyB0RM+kVhu6cCbL8J8dB3yIgLm9nEfZsjLkfZvfbDuSeupO8E5hzj
wYhGRBV9771PiVdJUAJFCg4XinC8Vv/PidwaVaNAMJjLlQgz+9xR8fx67vshw33etoc929dHCsuj
hULIC5wTJW4oAhS3QSahytFD7OctCYEbt6KQKHFsP5Hw1mJE0DADCWjKQ05o6o3BFtfX6M0rIf1s
FWjhyzYGJk0BB/qFOuHR17Yt7M1Lh/TsWC/SsG+fpOt0XWaPnKyxNaeth5n0IltKQbagUm+Z9UQ7
R1r3Q++ei/SgrothtG6AyrRIQqY+EOSkEFirDlP1lrshExlwY6bk9UCSq3VLcJW8Ix4oSq0VExTl
QusTZdvhBGvn0QRW18m4UNuDlNLiTuZPwLqrLAkwi6tZgluxBFGsy4h5k1acEWqneQVgcZcj3Aev
ZD8cY7GCufZMsWtjMzSffh1iPx0lHl9PWIgmi1W+JHcL3sha3U7QSJw6qh67Z/AdUYX6ST4MNdAj
+86MGFtoD8YhpvQ2RzB3NeS1WAXf0q2Duy4VgDUerOxhyk1hdssL+VVXVn4ksEPWa8z/OknUUHBQ
rTgSq99k9P7JoLujP6aiyQGIdBr4eSPP/tSlfJaeDM0jJAPHj2FJgCc0V88PTe1FuuvWmV1wQSYV
YhXqLl0gRHfQjQhUIzOw7bfxJ2vz3hWreYmnC59eJXuwvdPZ6XEDmvssK1hqwvJcFvnc5EpQCA3U
I+UBQgdwYPmOIHjhzrf4dg6BFVzTvQB5SlsKILtbCnpB+IVbFXDzNh1M5iVGSNOED8IBUDD6nnUL
3MNPTGkSRtryTD4azJj2BLbc3NfsddYlXhBLwWl8KWYB4B25y8eX9j6LS1JmAQg9hHxQuNEGHt0a
jL8lkl4GSSwtOCxNiyTxVs224AOEPlEUc4AWj0p8shLzJagWyx1RidXaw5rSoOkip5YYqDahWKaU
pwJSfj4PgJdthngjXPYYanqFPDtGxCFMrJg2RdVQX7hLjPQlPSTJZHPtW0Tlqag/P5+t7FQjN0c2
KBmzG55RUWGibTN18zOO5fYF+RSGKK624R2dAd0Hk7pFjSD2MPU3M+ztHdKqyFzHIPNbAXAZxxez
4a5tLMVauW6urn6GbYfocYJ1tStvstQPdB0qgYYI4AoqPiROyGgKVzVmtdpKBi5/DcaBzfK5uTYf
ER6PUAqif/dL4P5Vqee/1h65RyBe2WeL7Z27PORhAUBsQlO86pHR9mUjXhqyDnqa9RnVKCbYGkBp
vHVIL+ehLpzPJGNBrflhiq3mQygO3YOjbU7cqVc70U0U7LXNpg0ZULDPXGahgw4mqvl62IZvpPTa
ze61eWVhZwo8amxImYZ8xv8qytbQ9vqh3K6GABkHo6iDD5a0esNIy1vQ+1xYMUDhonw+nH/CJTkB
P+eojN/3Vru4S1DW8YurJbKwnIqL16Ywk0JNI/GPUZy8mMDJL8sPAbb0o2CAcit57eez9VYSF4o5
9QwBYB4xFIni9eWGUYf2MIjXaksgHfSuHiG0SX7bLA9qHzM3yWnK0MJ/9lnY4OL/NH5fy/nWJT+Y
D8mwgK7xZjGpTRXPMUXaMXXGLzx98OhZbc8WPjxTTkN+yErt2j/sjfYdrc/WFS+fFyGbX/bujSmP
zk/eGRnVGE4JG2h2QOYJ9CmC9wJ0dj3SoawVre2NKwcQu3SZU9Al+D7Vz52cJXN+SYmes8vu4GP4
S9Lz33F4OoYJuV3w/jtjDx5vQi3vW3PUTZDIQbGSeeS2mXStSXLvbI8W63CFllk45ehz4GkjQrAq
lB+2tHQptiLBJwYD3Ke3c1q0bRuW8SQoRrOMx2+9sN29TzevcTQHNhdl4dSZ1phf31N4BzlFp4Dj
shiRJAR54GzJ27s8vJqywZOhbFdoM2WirHMjanFNogOkgYQCPXVAjAvzjzB/nH22nWAOiN6k8uU3
XImRjKGmUG3BgFeI8KeFtbJjPNuIp08hYT4MEnwR9KpoYf2NoMjuUwjbA4XzkG7D5DB1BfwmkL+v
QP6JwZtNFJcH6TqWVlFFpEsPP/1Nl8fmZk6fO2nP3mACfbUsejoPDVxyDAQNHIr3MB1P6c+LJDAA
pgdwHSMpy13BBR43Oiqwy98mwb3vzA1okhCrrNYlVY1QZ1AeZ5nGBIVmZJYRFfaeNq+XlrCQ0NUB
Ut1QulHigpUIn5PlG2F/NMjGKZk5/efoZpKOt9iP0JrX7wdcQpTg2QdHCuZx5GadT3YbvPeq/Xvi
tehHmaR/E8SP6UogXGCYNgs8+AAPxcxJ+iWjWFcJtDmsfihhVTgBBezi93M8lXj4MvDppmypY2GE
BpjbY/ETB9e1dCGkQnw61RCWZaBI4BlC3HreTWcha1mOSVLLCiEGPLsBkePUCLwkGXeXQYeapr2+
ILoL7S041IlgRXVaCrDBEYzWyOZuQ/sO8CtdHOqnMRhQqU8quepXHKdZsLZ4K7InL6Sfmxfb9gHO
sPEaUt4fJ6C6W4/yGbn39npFueA4lNQbXfBff3g1TRps5yrPIrYFgyy6IFZftqQSJCOAz6utHa6i
O2/Si0eQFRltmSRYJPwnm0cEqbOW38vgOSEziNE4MwWEzcQgg++KyS7N5p2rGsAmPc79K9pjcSDs
kCoPvud0Yb0hTJGVNsnX7dBuUCvABMGqBaIXgtLsbBDlOZ4/yY9OWDr1/iSPpvfv6OdT3BU6R/ei
IpbUzw83HZ28Wh+iuHcBt4p0vo2rYn+IchdtUh+jjhQZMhNStsBrUTbPjCRv8FK0m3mRi8LmNsL9
Zfa7LS3XYA6HCI83do6AUoYyeCFryXprfmIMwWaPdzji5IF6e0NKb0vKtSzSwDSZKddQEnY0cXia
dnLIahQurFWIFhRs2lshNZlr/D3P2tGL13q2bTUnqBOuczqsXTklpAU5IyRzshZv7a2fwjI+PlGG
USpQJRqT1use0OpRs+vmqDeyMhsdDmYVo78RfORwM1lE73SjHB+i73bSOuZZPTmTm6W7e2l7kB0C
/dbyBXigQ8LBb+wds24igCxAhFcYpnclW2j73OgToXsQNr0+aNeYgCrBnC7YhPhfYpsKrFPAdItv
Hlgzih4QshAuKyRypK10WLIPcjzGTxRDgSJ+hZ7wlDKOLI8eO9zIcx0a1xoMxyWKFKZfHNnsWNMx
Kl05YR6jb4KRX5Z3uzmkyTpq4z6xCx4emiEKJR2MyK7Ha343iAH1oODj7l5Yaf5xjeUV5HFmg/5B
wk1VWiqNUPCmtmnc3Ckvq8WHg1NS7mNkNxKJKdlgqGtzmR6x5lX2Np+MadUtJLEF748b+02Ebfbq
kOlpuq5vYVvyH0qYKz38ef/ekomIyNV55rPKbWzcqxFVtBaGqggWZJNDHqqGf7Iac2WRNx0cf4M/
Hl0zGyx4r+3HWFqul8hBjeLzBpfGw9kMRCCR3Oow1QGKKuifnrv9NIHBj0HV9eLXwIa9jOJXO4RO
lWZbZHSKxIecxPMBkIJdB21yqllIcRVNjpnJt1vuLq1yv3GkbtXoMyaW9IaM1wuNJ22svqWUJZpq
YIDssHZsuE6lHH61f1v9kufi7qR50yBO5goFcV86mVSJEm02geOLlWs6HSTzkoR7C2/VUcii2A/l
NKJV4aEaJGLCh3KAsYo0tDxG9tyLHG9GAZmb5wh+QXk+FPV6usL9qUjM+Ybp1zGhzAsnJPPgioKI
K7ce+e1D0Z/8MiNT/ucNKzX6qJAdjJeC2g1YfvRA0dSZWHguFaCPYta/mK57a9gAmFVXU36cfqJo
4yiEd9wI4gtDMKOnJNvHUG0EoOy9vfgZDlrU22+sYFbwvIDysQ+kP5cK8lbU9Fmx654/Irqp0gdQ
qYpMxvj1mhcZoUQbTgblKpVCtQi1ihdcCSlSoUVAQN/EuhFg3wAI6A/eRrg6/PCpeE7tlrbKfueq
7bRiPNZA9xf/vRps7/DDtBRAqVzA2nULM4/D7eeNtzXKr3RStd9tmjabe8g2+/cCHxmtgrSYsJby
1tiy7eKYfkbFWwOMsdFvw/EL/SomLR7uRK5Z4UJ9xlMZYefNhgXUGmN9d3vRouUTrroqQRGRfBqK
fWxM0mBlTraAf0oiZ9YUQTEuCxn9l4S1wfE0q0vYHQMLBNwJNkkJKQsSnZZnRPx56eCpcvq319V+
NkLr+jtM/HnTLyaOQcUa5uLdJ+Jb5z10y3Sz3lC8Z1OKSd5GllthNb+2LCHq55xtqKHWoj82PKy1
ym7Oeq8OyVC7f0xYLAo23YSJRb3QOpiYw7ltz9W8CheG3jVJtEBQlDzWPNqGC1q42qJekLVjqyHD
3AEzZfKQhOz1iD09Bonh0Dnr29x/GiWEJvNnJp7DHHNp/E7kvnkcfxLutMOTrMdB68fJmt+xCKdT
PvlYP8nPzt0z+R1W3LK18oMvbWG7BNJgNOMpLmrsON0cHwEknzCUefRTlNlhyXzW/xcSfBURBLDZ
xy1ZvHIb9j3WDkNZwufdhL2/8NLyA27lVLsufJZ0aITTGGAOEF/DJWleO5/RGI267Rqrxads1vqI
lCD8ztH5nl4azx0SVt8/A5YgfM9a3Ug74vxlHUwW529rpgq6oltV6W3jA7SYJVVtmYsjnRhhXwtT
gkf4qh9usAT5rPShSx2SRhbYUwgseptjl7hID2gS3ClVyQYMaH2vYHvy/3LflCro9CBN26sbUWrY
sGVaH/f/8VfjHRBfOCbORKRMTKeY+DT7VEvkPFkyAkSXy1n/P+76DRRXj7H8eEbojUalMX8u4pbx
gvCyYYBdMpW6k5NPGkQ7WYM++3FxTcTbO6JynORjDeV8jSWbKCfXS/hSRlfZ3A/rf/OmJT/Qvuvh
TjaddlT2JSvKtFE3l9k4waXyfpn6ZCcQxa/mLWH9cHNex3eUnwdfKzAkSzriinlFCxOUjFliK/dO
jhdnXsIGnfHRbG0z+VD9C8cczDypWywRGnEYpm9QU0lpgE/EgnJrTiXXK+S3bsJ5hQjGlArAz/ez
rf3DVsbjiFDH6GJhwdEoyPS9sF6GxhaJwPgnIWM6WTfWPRsfECLOzksw8gXfvgdnX72S10OgLR0E
RcLnNmNFDVXeQo97FEULqF5z0txv7+4PuymG/1Nb8bPVUPU0Apt0tJEmPjemZvQBJt6h5CGiWHMH
EBG5EQEeD6A3xs5QW0W3fqlKaljcaJdlG7gzuekMVXu6ii/hWxlQ1zhbdEjGcC2DSs9Xa+7174AG
vKyLiYfwa1s3BtXnLMRMR3cdNlbhvfp4Sb3dkjopUFwl0siivSUt/jmLBkIF+RNFC6fO8VTk7u+i
tvcKTZ/OxQgoOdGt+SJA+vlkXBxD8ywMvtto16VlkoufJXu5OvnqgPRKyPEdj0pbdRBnj0zsdIv7
8Owa+9zm2ueQzADVfuNp4XD4+xTuMlIZ9r/rOOmLUVVpU3ye/15WbRsOdycq1CdwLfZZvCQtJTWz
xOtvKQ3HBwocx9TY3F9NXsD/IJW7mSWJ0Pq3rREZepeaSMjAc/IwGCjWbFxiJ1lJ7ONDrQKXzxcg
xdcPD/70pmCMRwrWvOyQCidvjpKgzeZSb3gmduAnjNNziOeOWPBg4tcYgSw73MqyIJlZEROyUXV9
cstHVOZEMOlJAvdlJ/RO0StljLU4d4abLe0bIx9a6B3/1s0EXT3AkWSF8CnxFi7dnSt1XpYuRoZi
BQ6x1F23RCYeZXOQe9o+D0jfc+RWbXlwEcX37baGJeq2qz+ZQNflFa9BmH20NvgInFK4zPLAZq6n
Esi9G5rp9CKn9b8thdKZ9H6n2cbPqqVmeFgRVIN3YUUe1RzODDi5uU4NO7d039zxldeJij7guG5H
s7/nN9g/gFfmbGHEYKzXNbTZ1xnRzoJd25R5LjqN/FknAzbk8Xd668eemRoxznxOaKVfKbtrQ+ON
pwaGiQgzwSaxTbva6VE/CIZwbtsaEC05o1kcp9HbwapVS7xyglPwe72tZaifKePofxRE+DfknYyG
HT/xMRdjzs0eOPAhzvkrxNquQLcOd8rudGqBq4i3sXEAKkhf3nLtW5O82Tkt18CM3YzbBpaAqUIk
bB5/ZzcbfxrfGzAmlCypqzfmu3JTARkGAxThbNPWMICXa4cb0ZKozXxefB/fHJ1KimWyl26uFquv
QU6AklrS5u0dOlQcZRIwZax/gp6XYViVhnMYfvq2RkJ3sy0VTIr0IZJlMczG9ZfUVsSoabwPFpZA
YmpSl/nKwpv3xd7g3xXsi4lUSAca377ux0g0LrB8uAX8hVTAFa1VnLCJf5eMZfB/X/H68Ns8AvDf
LtJP7bV5jH0+6RiydbuI88/Shcj3P26ufziYqzFfYidXUcIENY6defxuFArqvq5Na4WGo9YMV4kI
k3c28fEC2wGtIqQnmbWvoP3NS1q1nMMTIgGSRKfDXXlAUzOCfSEGC+uA4TBiWcgfJVW+yWdae6Bi
80cGMFSDxvb4ygdyxFeICX3WviyNkCauccKaSajBFyzW0n4ijwm+7xYD63zB3nlKjknm9SJ2ztzm
Ospg59ASL1utS3Ze6AQT6+95Zis/2/qaMnOZJeKrRktmH853bHg2PoQtzgEr2fW3upv04CDogkHh
jOB0FDLKXcvYuD16U2B8rG8gB9f0K6hZuQ3IdHiSOH2q/VBmJAu6RGjtQAAUXo8p4y9QHr54WcHe
zCI3NfO8wQtUOPXUrUgn70Ym+1pbGfeadrErmlFuXO/D2OCiql/uoBzwcu4EvOfAuszxhYCvDpvJ
HFuDIVp0wj6e1CsyjcVq6VKV0021wPPDeXle5HtInnon5WoB/1Yy0PDScw/SW5q3bQ1zXeoNXvuj
lKf0YyAMl6kZS/739gM2kslWdDEe3iD/yqKP8ywe4Z5RsSi4TYg4g8aeOS1dEWL9l4CWITELvJ/N
PqboZ8Oy8p6gIxOlVp1KBERCExx+ys8F5QVAFI6H/+N/brgj2QVNxNNbO5ukmK3+mPVGTvkWvihL
p0s4riql/xE3KxrvA8wZF5EjeAT2ganOBYM4nZ3jaBPOeYE1nsjNO0jsNalPHRxhNSk9R1upRZ2H
AJ5tGKg3SdI9hhxfHBPB+8kn3cPOI1cWlbsEp88MuxMUF3tgrqJm6VAyt0V8Bkm4YbNCPtIQ998X
hpYx9x3cEqWmYbBl/BRkvM0y7xJ8kz+0BWwr9kXpup+SUBzuyH5NIbpXmvXKlNxnhmPrzxxnRoVb
vZrLvzB0bndntS3B+55nddDeddpoDtdBAQy/zoh/dJyXfE0PJWqNq+ZrpP/41kILNz9TExJXgZH5
Eu5AH2UI8+XdhDFW9DsLQfhTna95kGQjlFOQCUklArlx3Od1RWE50KIaQOvC0QEsg8Z9PVuojCfg
lsBBNlGk6nYtJGTXny0oaAhADye0PdMQOsumH2HZ542Hwf1M8lETE1opG7ladMFswRhdvaSqXVrE
ikDazXSG1EFAQ51p7EIEMUJzeklpeY8RqpQa9Z7ymRLcv5UbsCmiP68bwRgaR0JAIrKjkRiwFN9+
xQ2O91tTBwm3S97m1TA7RVPiSenqauYrNpvU9rQ2niH8cXylFZX4pANma2olkbGznUXB2rsUQgE0
jp5/VU3y4fTykP1mgSVvrrwEvQ9M3daGCjoA3GbswzA8LBlkGf9WN4a+oXSlmVCa8Ow++5Kpzy8q
GAE6JqkdlDn6bADSkJTZrGdtUjy8frr3eRSCyzng168AVmuWMkVBWvsY1b4uSUox6igGHKltlHiG
RoBNh5QnuQYMmyh84PWfkKKATP7+kR5Tv8+F9QHhZk8s+KufsaayVKv4HfvhoLCC0g6grrVVLZrv
UR94yd1ioVE0izwZI3IGlRRNFFbBNsw+XXr4gD5vGq2VClULpv91dpecAT9NrE0y6l99P9EobLs1
0bnt1FcUorRKf3maS0qB3brAW28pjAymchEjgiHJ6SRjVX20L4AWcl0RmFMU05OFkIVQzk/lNojp
uxoi9BkByxjhM5H9rqpEO+S+6n1SX7OsC2NgD57nDzMgCitu5hKThHfw2dPyQDPWFreKbsN0DB+a
zObJthkzxoU3DMBLIr/tyYtrDutKFi1H5UXNquitarl2vPXYgP80iQ1tPv12uvJeHah/DDbTLJY7
QuvuO0bybIBdqRsDjboF+eI9O7tWN37/3o22yJAJ8933M7BzV+pUrnwW4ot5LRnm96q/s3szvksV
3ueLRtJUmu8QOcFBN025aDzxKYZ0vxAh7Zy1ZTC5WRu8z6Whk/QBwXj4KxulCXoto7sQJd0NP6zz
uibjujQAFUlRoA+4gdKMmtEzGv3fib8ROZFp0CFI7w49LSJUmtp/SeVvFTzKbRQyssKfFtCWhBah
IWeqSDfA1KAGPtKkJ6NtgERSTiAAqO/7fN49gdDKGaP87byHr//SxLHXqLzQAYp2p4bfNpiOa/Zl
H1Ml8jtGd/cC/h+aRBtQL2P6PKDYQP5yZnvRL5g+4DbDUMpro/3NIMvyp6r712IeHoT2/QNybjA1
8Jlxo/L1pGq1g6JQfZteUC2y4ZwOg78En3LepuumQjpgbCQHQsoiJygKxIao9/xGuE2zRxuMy9oJ
Z6tuDU4QE2t1yftPvMcMW6YM3SB3vjyQ651hJ1LNRN3+JQO9ribBg2bQSdg0zZa+v0PKSoyw9K0b
o5YedzU8VHbniXEj481aBnavx/LY5cYbzv875+QxAzTQXh2lDQ7C5+T/LrBV6Byz7GlxU8N7t/j+
N0R6KpFm5xzRwz93ra74AA7hrE2N55J2I8EYy7jtv9oSBmesStuzao8Fk9QICuFvnH4RqlJsQoPb
56AmKcViko1tr0uDODsENuu8AllAgLz+Lh7tg/ltlXAix7RjYMKQveQhTgJshvUJxspBoxUEasw6
0YqM3Ql/D4T2mOKY5ZAvOHeGyMij1ETMR78Zp8+wd1gHHmn30cxS1/un9XJqpPS85ezrQNcRuD3W
W6hAWj8XyI5Bl1tzbkbb1oRDR/CMngJm+PZJpNwlvBbSju0F6vKBewLlPjot92fhFOlrFnHgaBv8
pUGaWWkzrj+d+sMB/zxNWKetwzIrd9MsGhyJM6BF8ulSml0eFT6v27plHstiaR4z7bNm6W2awx45
ZofeK16ifK/p0Y85be8vqjqPMweOrYeWpU1GaaJhqMJucWdshtI0YRA4wZAXFUGwWJKlxvF/tRi6
qjuDa/421/Q6ReqMQbY8LHvOuWZGZeVH6bqjY4B+pOcoVyLbFqT/rf7MHh6YfguDWFXAw5pC2lfZ
dnlBQ6uTmo11qeUw11o74uEc/XJyUheydlJaFwI5cEk40syXnamVg2ECJ/s1I/5gsih0ZNuzWzRo
lIyY09YMZK36Luq9hZKcoRkFZ+zdEhEwLtJeA7Bwy9bnoZOgh77KC8mVh1RJN5of7pY8eCKFKrx4
/YHIb1taPRYvZDbjlJzGZ0SNrMSwf+0ul1wNFz9obfq+i1Z6pyqdmKh1cAVlWk7mfPvbvZVvRNY0
+e/DwU+9g0QDf9nsXKylz7/QHRdCz2nggq9R1V3IDDgJs7Ce+p2i1kMmhx8KOACnWsHoV7Z3M3NW
MBAU2DF4xFtuUqd6mGIH4bg09L7RLOuaNu1EOez20CFDQe4M8jZU+CtdcEe5mugCBDzt2bske4kC
OMoYEeW2NremGHzmhaX2FTCTsTB/j36H7xxRQt3NnJFR2SMiKw8g0q7xG0DhrvlPbjjPI6WyvoT7
1grihwJl+f8+GgpZ1l1GPhSHKCUqCjlODddnjyY2lLcasULOvNdg8hzLaYl7adxeZ3U3tTYX0Erv
QsDDYaBEX5x/AyT3d2a0kJJUDsIaP9FNozuoBYWzPm+Ii81RgnEUXa7FFAnpDKjC0rGMfVhjL6Je
lacVRudwdPdZ9rwOO6LXrfjx27vTctQ+h9O0m+91rmCTg1rV5KnhN5bWvXU9k2K+LJoTwPJnVqrU
2O0xPVumS2T9jJyItFJTqvcVVH/TRqqLjexg/O/hfYaE308lLc1B6hBHAAEvk4ujNYs2HUk1UmWH
uhGh0bZBhMS6qSmlSlF3N6touKxxlgUwrR/6p6boZTqSMXzHJsxBOePc9ckYpoepbpU6Crn5HmHl
b+3DsmUBq3JVc1m6ECoIHs3iZKI4EwInJnEjDOLMYbdNDXH4SaLRq9FWGSjlwS4f7d47PuGqQfYu
lPT+JBNQQBarSb5YAFcPLP7Fl2zeZuOhFuuuOY2VC3znB60CpCHSfckGRkuUAk88i44fAnZcN12/
NDve7Uol6OQKB0oTrC4e1nBCDPJi7jadENg5/Mp8vRXsZYZNBle3j36HXB7PGUdkZ8q2zPrTSH50
TjnsX6C6hG9F3hVCrU4z0ik3s0HdagE0Q9K6sW8+pDkpE5lTqLWcmMQXMK///GHBNt5H4olRhKX+
PuznLcR/IZaqZZy7eMjxTmCF8KtVTinUbvp0L/YvPaTamA1KyYJYgJP/nAdMYVOTVRTZ2SkT0lOH
2cu33Va2uZEQnjfi65mSpVyJalrm0+X31u1l+GW6P2aMdWCi8oPMx/UwLLaSY+ldrfyok7n8FwHp
PRqgqPuK/DB/WWd09oDcb94LgccoJvNA2RIFdrP0PBpA6zmugGWgOsr62PYPd9Zz7uNJAIYBmpM5
BuRorxOLS/C1u+nKCjuAIxCkkkqrUYrk3Fi0XleNpUh+l4Gw1l4WMyRsJbitvU+bkiPa9cu3oy3c
gmHOxECfV+c1+p4WX5ojUOACzWh+JOEBzFCAmWJNvjM5IVY+tZhwQxE0WJXI8B04fYa87rCH7y7A
3JmEYYUhEWWrAQj3itok7cp0CESxyiXY24ciF1OdPctgIvvGE3DAwcnGz4bswRCgx8hKOKMmHESy
hMnlA2e63WoLWDi4mHW8l4ItegBLO5limK0BiT0RYt4s1Cu+uHbboUExbMcKHqOPJsNK0Gcksqaw
3SYHulCshvklt5M5qosmvUSJeVkRvFEbINn9CaI1lhPQQPafBUF4WLQRf48ke341VqCmRwwpoz8m
GgQfz7xMy8rRa4wwKCzc4jE15OpR32AktBoUtRY0ejXfxL52ATDijli2GzpmQE3pO+LiyMNw7Sdt
+mgwS6Vp2HtdYnKjdBYVXcF4qlOPp8AF/8hd0/cSmNnXYzQZidn9XbUbBIUF0hadV1SmPT3hdrwb
tT+47YS5+/QZFcJRL2DWa2z018dTf+m1ZkMcCvGBSxhq3yCOiNiPJxUa+tkwBCy/zA8zBGQw5GAv
GGxB1kXMlUXcL6iW5BkR2H5bu482lzxURiwY/TQj4Z77izdNRSuaw1utpmuD29EB6BqZvPZSvPD6
RGSTOCfu3EyCgD7mA6/Qd890ikwGqa2UGeOjyCIVK2yLf8jSD5hKLQADWVgLAtMK2pxz6gRHNFuG
wKToH1nTlj6h9csvK9pQWuQPaUD2y7Zwh507PgPIxy7+q/l0aH4LNBpQsVRaFwloY/5aKQJMXnEL
TG5ukTSC82KOLHcc5Sq6yKrvgxOINhe8N2DTjKzLpWLkGz8vIJ3Kl0zcnZvvVidnJf5FquvBaftp
U5mgdxMpWBH608oC5eeD+B/ufBUkqfW0kG6fA3hAvi8vAer4ItVuu0sBbrCCUvghqkA9G+5HTQ6D
/mT8FHQP41UCNPasA9jaGadLeGQL1OqIRTBirWmL5RQS5s3AcwKdyaoKVGFnuNdBz+pE3iFUzfCO
TnoNX3iNqrbS+36jrKbdXFyDzN4F/6Ofmc2U051I535fvnMtUJjp5ACzzP7fd+EW39mGAHWOC+wz
s2SQBNASMHCZvyWDG7OKTfj57FJ63Uh5+toaNeFaB01NHBmtefciU2oeQ+GP4RK0uuwdObFnuuaE
fKRgvdJx6jVaMkicCftgG2wcc+AIzj/vEGs7y3Ac7P+XkzmGSPcGKnFizOEfuB9FZUC3wARZ/RVB
/bjni4+fVBNoSxR6LRO7KoNORUuVWIclItDFtrFH9p8t+ViC+H8JindmczYnhjlY23jeUm0yfNNn
POHb9AICAewqoxnV4LcdjrFP+0VQhVx9X8SNd8Pb0rBicPFjd/+0givQWT7SUecA3+RZ/2MBFlgd
wCK8DS+dcAlDjSkVpOZLAbjCj1myr15vpkkzmGVD+0rjWOKmC9Y50MxirTkqC+n4iebi9cgullfq
L/zQOm/Gw6+I2c6HJidYWyz6Qbe0XYosIxCQSlBo9CHUJFOxdsBWB27f2gC/mh3s8GuxXmEGNixN
YZ4ylStmCcSe9xqrNH6OkusMHUKZ5hxO9IidmqueMOhZuym5kxnk6j787noFjc0fApteuSfogx6j
uv+ZtdbjJiip50QF5L07O6/xegruJuaKUHK/GKPEUn+WmFK3psHY+/PQtCpKJiuCIkhF61i+Wt0E
ROqbYPp/Bz9utcw+tNPh9Dfjanw/Jgodtt3r66DdpRG+ofZcUDrjIVjslTmyVNNQQ1oHYvRw2hIa
FvydqwV8NHX46d1I2CH6A6TgBKkfEXH03qxFNWWaRWU7DCLVxQZLbFDBICqKb4h0z3JaJW8glWFJ
xzFoY0UdEflTYd10t8gargeIcFn/kdxPWeVuOrGA9UtNTXJcjGDBN68NPg02cP+4TD6Yu4LpxjQ3
AD9qrG011J4TK6k8oC0F3TQnBRrWgwSsRqfNzYl8ZAM7YHyTIV+55+fJLiaFG+pd0QUtTKeLFm/d
xKrtPqtGJeL57ybRQ/wrhY3PRxtiVkQlF2SwKwZ4r/BMVXfCM/x2Porbl8SpCgTKa1mJLoqv2ezt
JfqHaVx8DqIDMGxewdUGXY20ADe72ghWa2DXUCmJkmHJOPZSgUzEkkgw6he4ArK3IHT+Cavce+Pw
/AIHIoCIkY3s8ooJttCiNkFA58xGpYiUebaaAq3fQcl3A5Jg+J1JDOzOjsFZyYG3x525CJYUeZlS
4T2yFXSXOJUovDIZMo4FVtTqwUF+FBdFkie8A9iDocjhkEDF3z+K75t0+VzgqrTTHWUvOnVAhpTr
Ke2/nGthDZ2ABPm48d6t4pizbVOthv89cKaxD/XbxauJm1+1KJlzNnCu9QXisMN6T4BS6l4CUa5K
LxV5naFya6jBBi9NhXGFUb8igUc1nprduaYoE2HwRyq6F1yhnm2IVgXiJNSRW/fzCLPfy0OEH8fz
rgSDxhOy93iX4JW+8r8M2HZSXIFqFK0Zbvroe24bVa6ecRg/OXx+YXASEDjfYGzokR4j+K+6rZz0
ybXibr5jr/beMNfOBHqPkwXqnNc6FveERjdL8enRp+ZyVzrn8Rwco9yfEK0N7kft66KuUv/1rt+E
0Q8+8pXN2HM0O8AgnwvOtMGFlAh67M+YdMFhDuO3W1okdf9Hh/jyItlSDtGidM0+Q5Sc5OR5IACV
GHjxbkNAxWA5lsC/DLpFmB68kh3Drlv2L9vyXS193MCAwQfutcQ68wZw2eNCZDveYEfHLJHKf5sV
N2sKpswa3+CzpYqMwTri9j5aPHE1LQFLZTFHSV83AZwxgEjzFi9NopZ678NlvvGw5ow/LQwq7EgC
3X4wTVcaRbwgGyn+MrTdr01ydkkZMz3zUjZ58/1ydxiJeIgyK/PzfifSR+FqajaHwMZWz4M41e+B
+fskuIkT6MqJIYijdabO7N7iGAS2kINkcKM+URgSC9mavfIMbBpv5szMp+GoZXkjAsk9ry/0Uejk
mpOSG+WTZX9pKJSeQFB7PoZGJYXwwLnYGjgCKDgBGf7U2jUqL2n5wS5Z29qZwy28Pmkh9i7Uaekw
mfV/JdnfJJBVcqpqdusOFxUf/OQdS3IbaZB7NnWBQ1fvPB9x+YI4yYi3ZCRO+vwFzXRIewkEFscR
3nBD4mh5vQ8xSlYJp5ri4w8Ck3KkP1whGcjuI7CHRMOavM9GH221KwdTo91dqkBOAmSLB9eYQyfp
fYlCxzOLkbuzlciMU8TmNTJysxGeMjR9aE1J3+ykWc5H3/hMUvJK1t9iQv6BBKWfPIIQ9b4y7brc
phtJoljgwsiSjRKtOTq4s7oj/hjVBA6ejKH7q4IPfD98dtf0e5uZ1X/Q8lE4BtrQsskfxg7et3dv
oTXrhCT0p6hz44k1r12ZJntqiobImjSJStAVk/jVxE3Bwawdnb4cd9OiMipyplv6RVzB6wMp6zTx
CMDuHR+AUm52OTB75IP9KL8pfxJ2G0CkFjSBUjy4WPws9K3A+u7S3KBW7uMZ9BwkP28EckArz38m
x8sZitjPGotLkM/srmbRUASvurm7oJqxeWFlg65uHT+5PWp04PCPqNjLoGsKc/8J7yWm2fmgpmEj
9ZzsSocEvdlMH/AetAt5euVGP6ZIUVrtEwqWZBoi+T2uU9tWTtTnG1qdWreRppcnkM8Ormq5lEdZ
iYwP4DDvQy5VEksOWbLzfJySKXWLnKCgcPzt7JyNnu6xdpZNRhDq2Y6LVPMrZhtHvMQnF9jFQnVu
rt8Rm27zoPriAdoEBix1JyDWMNq9jcwQ4htOeddwmsR083OZUp2oWvmVVtQvjaJYCBFpoFFcS7PY
vaS4m8cLyvA0GyuOusZ58PlD5UPazICLs+aq1Jk51Wj5zjT2WfhPPDzqhovqfKBzXVonb82b+Z7P
EG7DiLcpGq9gFvRB9NbHTYKeAP1lJT7EsG1QIB0zCcCUiA8WRU6p3RcYUyHp1IeQPryQ1jguU7P5
VcaLXJMS44vybK9Qlu4l5TycTkP/rYLON0c3xDff9XCAok0ht+a84Ndat4a9CpRz0QKUcDdMSLqy
94swWOx1ChMRHcyewURxJLNfNXWuOvunvMWsIht9K2Ug0HsRlNt9WjewqQycKEEaJshUxi+NBZRI
n9e7s9MVdKOTIWEiB7ZMuvvNIBzISvsUZqNyLiSnRcTIVUbqWIv8401G4YTHqojo/SApp7wKFR1G
CwX1ULMszajpvQZ3VmVqQHSEShInmyl/6sBV8VI789xnyE2fFAV30yoIaGAgaYMeUe6gO6YU7t52
Gsx0P2I16qa0IkIeWO4LBJWEv4tRIInkDoFyepw/Biqab5or1L5y5KGx16359nCBOxpNfsPnASLV
8c5e6271VP0fLgA/s/Mo4a0uV1yGLY9XN5S59+Gf+uz8teEoSqzjaj6AB6h4khzGVs7dW36tJOzs
NsPYIbULQ0NU7wKjyPwYNcDY027quvquryqkAoQfncFtiwIJ6jd0ClOR7ZLsPwwQ0zSj3UhMQeW+
Y7qWZISzpCFRKUENCdSf1x1MPDuldrOBaXXuM/Z1pZvJap3V2pSiun9GalS4MqozgSZyAw/81Gm1
aPUk179fyAkcwDINA/ltjaUCY12NMx4LbvwClpLNCHG54gM5Y3Q4P6ZS/FqjeuPGJcgwACx1/OgA
Ua2eL5dcv0XlmIBhbBRCRVqRILsjSbWuA/kXJ1deBbAyWV0v7XIHZcbt/xXxVxOWQnQdkq4mBo2A
TL/s8/XVuxH9GcKAsVRSjVOeBCDxWOgo0SXRL+KINdZ12wvZp3mAdVms1tIwRB2xDiHsM/FXFKwc
OJQYY4k7CXlfylAAesl+fTo1y5CrNMshbw/DJrehSKCrpUnt3EpAwNURnjwkHntNW2+vR4A/Htbt
FrqNKhG/QjVwW8hmJCEijqqJfyjZyH3KMhr4efb2xQlhuU5WDJYr4KKUwS4p+B+J9RQBijRUyOkB
KZ867nRJL3MJIqRKboTVd1rIErJFGrZub23N5FEtDQakwTdcwmjN+zLnZ28bdQ0bowt4onaWDqyo
2boE9MTyn4vLXjJ9xi391Xl02NT950Wo5s7SAnB9Yl620K3Vgy69ecCByF0j2t+DUWrM58iLM8RI
3PR667aJWoyeZLZ9MfyAxOIsU9HiWOSr9GwI6sJMKWRZD8IZPy+eLetXhS3VBZ+rEahsekjl9h+a
JdlLE/jN8pxHeXoVGKAGMWLOl3BueiYn7y0lpXVCkKMaXaa1UZ4+mBZaTHlKbTXqX3gWhvLTWCYp
wj0p5X1m3Br85IfJdYXWPGE//UdWLDqiuqldszyZX44xwTaQ5PpwDnJwED8d7owIhVIOV0Q6DGQw
ZZofDiRWzOlwWERX77C6qboDw3SK/B0b+OS1xeqtrjgEab6qaRI28NZWbD6cvUuYVavp2jmpZ8mK
XjaDVanDe++SbZ3oZgidCXmDeXuKs4MNEdjm8HtfUiL6lZXRZ1jLg8tMEJrKJF/1bjQG+lveesOx
w+Elsmeekoi/wQgAwTPVoXUN+/MKepU68KuNdy57KTeyCuBqWEQy6BHejc3ehOcjFHjn0sw95Ekm
xLtT1AMUUwiQA1iqpPtsHNLVO3s3ikSN3PalSo2DGDJZJWQuwilmL3LzJPZYIpLrjUvmmLrw15db
KT5kskY3XU9FseN6Ld5PDVvuqFaBhdgjwQZgXx/q/5j+K2vo2gR34++6tR+iLgp2Yf9ttuhssw8b
RHpnwgJTXvO0bOiV+moUkULy66zFA3CulKh5bIVgETj3sWWlNLT3gQ4/aWtJ4SixSvB7Plr4QbHZ
SmWLdTFqGNLDjSZEJext8Ry3ChrW/CP2cf2zWuWUdLdbHBYg4ioqcQREVLsYqHtzKgVQokiamKXX
unWHYpf3qhoSV8J/Y1vDmAit3iLtR4XCRs5aJJPeRy/NbqibljMARCwVCHQYhTlxYxf6mnM6BCb5
yqqoFixGC95+QlPc6EqzIWcDMWhP1WOL3Bfq6QVwR3l6r6Il7o9GRAl56Tat93XpoWmhyPnvU65s
FOJJJ5kS+yGZfZSVYthWm1RojExAUI0uIueju1wdO13+GbhKW98qH+PQ1CMtokO5gjKgbZ+GClgY
WRDDRw22QjTioaGk8hj1nvVc/x9g6IPNiO/VQagVAbF1OTwAphQGZnOBJ6bO77zPbR/gL0NXeu4z
BSUIvqUMS4MQzVwV8n5TYBcK5O3x90UFOF652LTb9dwIO4xZKZsXcfT7mVMVUJ7kosT3/viPeREU
dto62l81SIcqtzpy2Wkmb0qtIjUs1gMNqNc5SK0Khl5/o91+L69sAovm82fC83aVosYa5lAxDCKd
rx18atxk6Yx6adL0546NQowaTCv2N2KC92ptDMFamOwOffAZGeexA+6f1zpsOgkN4954rrXdTrf6
6ZQFeroF/DMcPB+YgIMGzWNVdWhw0ZwPsJG7cuWUu5J3rR5a83YGcdbtLLk52VtEXxglxdRivLyR
jnkAZZxvsMs4pbxAIn93sNcxD2QYTtWOZev3AgjIpLViCP024UN6UdnffOAJwlawEkqCdlW0gUKQ
kIHO1YxuOKm4QnLNzgDdK6SLRI7PS1YhBuHjJne6NRBONQ6+Zh9lu9QTeRIscrihZyHjiTdpocJ6
Aj5oJoL+sKUDxr2l0Ne7RIlv7/vHS9N4Ixd3KXI6gzsXga9klrzAyrDLVUPhWCZ1BfVB6kBjK468
mSvQaUb2y/bhCCAO6MQ5Z/bdXPmPSGBX1Cm52Tqa3IC9VGL1XKA9jBMkRxiokqWHMOyVJ3I+uX+q
rDrb6ULwxmZFZsCAnkGsSzpIlZChF4MN8cHdOCtPK6wRv1rDt5vPfWbVRC51WYq6dAeOF78VO5za
PFYEyeGc6761ivxa2r5hruJ3zPzKHboQcvHApTK81VfPDCh+1mbLyavrZkDw585l+tQfcCb5xjvM
N7RolEe28j0DNPle8I3CdKkoqdIwlcWOe5XpPpNXAqfcRysQKLLDfuJtY7MZL/sWJSVeJm8KB1Mc
5hUfeJGR7Vvv+jr7GWABjeCK2PROB4O4rjQJqfMlzjmvzc9ip2zKoygKrL34g9p5+trHiOW+MM+T
CAsqcRYa05qL8tk4x2o3XyIh1yU/jHrTYiwwOdFg0vS9mSOXVO5g7stjLnCsuCSG5jSOLqwzJMWj
j5fhTYeZ6W+d8nHkpiPha6TMYBOPxuAJbQoSpYzarMMdZKuE3v9gT+pAOAqYpPuBvz2dQttWUHrs
chRDiLBR8k0knzEkpgg5IIW1uNye4ca5s6I7nLa+GkBbWGojWaHSKqZAtAec2OhrMpfRtxtPB7lj
27x8Ez9QsBEmc94lrMcSfxxy9qihhhJ91AwoEvu2TUPsYZd91emBo3G831lCEChzRv06NE1G37JG
Ay2j/x5NYWfDi7Bk2iP11JaDv+hu85PxZLfkN4jPrH/e1roGiH/88L4zWTYJmJ3y/UkJhAvQq+nF
LujIuTIax2IFaCi+qXzkFJzFMST5iqrZbXiKimyvm8TWAPzJjdJc3iD7+lSmhL67vyljejoS7Ofu
WDUUs4O6hBoLRbJuFIsWCsBSERkAZMqpRN5nC29YzyaRQc2EkYmUDyLdDvMt1EqBzHs/haHbF7yN
THLpBlb6GbKtBZBPsmOv7SqcnK5BTRv0KsDuCrdOx3VnGeWg8wZDEVgAvnvhujaAzHHv7gnvx8mH
iKopp9Cog7RoB90ehdVyYj5b2FuZcjIe0vQFur6LmxtadC6qkVkszvjM1iLW09KKssNISjdzahDi
L64qxcOStxviIjY1SQC85nSIWmFEsdQpLdZBaHUpk0GCrn8bGY1jMGp/y+A9/+kHuoZi3R+9+HGG
40eXu732f06CkVgBoiMxq6152jPh0/g26/ntgsKIWhtpy2JpFp/k0X5xFtoQSyzUvuMhHeuT5dni
pUGvxyxqElhZZqtBipQNhpItyUr0qCLI+pAeU5xUOOhCGn3o3BQpXQlQH0O/xqQY76Y4LOVaRBUW
94ttnzxJu2Lmg3k1r1kVwaLu9SIggQ2w5JGJvB85noyu7BtxRCN3s2VxDOxEmN10kpaHXnrL2KKu
JkfNzvYXGyxNyIPsr1z7gz6NBbuVNXUHIoUoNaj3HN9HQ4vDdl/yaosJrzmixgfRnZs6k9NgsLDp
5IBRKJGLXw1nSEpHd9KExzlIcIyV7S4cwwjrDbBttTJ43MAxXyYYKiNW360Pxm9WiyQPsWKigTbo
8O//9Mc3fA9PSz2jIYzS2e9F/7O9bAe5x6gEaDDmSs34dynvqFrECt5yU6fkoSXdpK2VE6vjgc4A
+8BivLcAZCZkWh46TQHXDqo66NlK53SgqVsXLPguTbq6jmEeZDsqPcy1+XCXn9l5HGGQf8z5B5JR
5OqXHC84YnPYe6QYaLJgODl0jQekMk4QOgaTsAkz+XajnwN3vrwL6abmABvt5D1Zufxzyhb2u7Hl
dEtA9Uc2Ab8mXhCt9VppbRn+VNIjKXU2em2f15A8vbr55ZEXiTCxR6KN4tlqda1v2S/ENF9daJcG
iJ1E18XiPYZQcbtDM3g8asEkWmM2GhYpCUGfp/W35GIXaPchb2iG1gwoGZONESmCceg5wQwZ27ZU
Oky+4EixaEeDN/ErHcerHNTDxReM4sFS0TFbrvWLjocUDzy3doo/DAUYxr/CsY80y4/e+n1SGseU
FAPaxYbxxKXEHl2rrqEQ4LtqdC7GtW++pTBonDuQoAK3iJEBuefaDza89+4TdAI+lBEHoAyw7bTn
Oq7K63QoBThPXZhQPnp9f6JLoQ9v8MstYa7/M70LgGUQBrC5PkBOfYqsXzivpo1Ro0nIG4xAyOKA
sgNQ4eMaJyyYwDsy6t6sP7nvJfaz1t72s4mRsiO1FfoaZ+RKDRtbkUiFYJMFp6HJk8YXawAlXV8N
Ud7X5/5txULIoQhqIZKBgdIT+trVjdwPqgF1FthOfaWPrAzOHFCb0SQuVis+wBWVRnBmcFZjoJZI
RBL3zRkxsUPuSG4dMt+cEj2G0/8V4eaX/Qvyd8pnMVPVrTcI8+aJvZ5rDuh85gOXt4GKkCOSOF5U
bKN8lPxeWcoreDsXv7YPn33/his9qsikkVmBrlczHNc84NBsKpjV6/VHUPX+gwnBmSXxzMggDlyD
8iYP5UgEYyumxemPJRC/uJxqhHpbc4ntI1sXxDHnuREpNPnoeWgr09+SF+7fhbeGp1eGfrzfGQtq
mInbj4lBXna92S6Y4IQI2PUdQmPWH5qlgrq+JFpx94KEmhbz2nEu/o4xRlEs67HeroiEAzwtoCvP
S9RFNUOGSzRSvwZO38RHHPAwmIkpaUyef99dDftrCOmnEntljJ7+QO2sZdhU3wP22Y328biKwbMJ
c6maTELjntXqvOYjZ/CBgtMQbx1vIdQFf/VTVwD5T+HQh8yM+JEIVHmVURAXqII+zqDZU/i6ejUZ
SKAAh7zzA6KbhVprqKeWh1njElkTQGC8DDPmpRCXVzcmrNYrY0L0LbtQAMQc84jtpIGF8w+ZLnqg
4GERH6Rw4bGi/pz9zhExnfZX3lY5VxMtL5iP05Lx0CmUN6b+vfeOAPhg6GtNBM6H0qQHApk4vpzG
sF5hZHlEQKm2lJAqnYstmjhQngs6isVt2ikYMlRYshDgBB2VHPlsFrGNSZayNgzxvJTTdcIby7QF
BZmkB+4hH239oYBKSG4kI7FX9JeZYU8QZDKrt4L/7ePShLA+elaO0qa3ySCd91+s+a86qR/0dBYR
BrWyNl3MAqyU2VMhHSqZHM8UywYSH8J9Esjm+eZbNB51buNULSk0fLGuI/q3TQvbqsvj1diSmy/U
nH2Yo8uoa5lpvGFHgK36UaH1RnRYP86LM8XxZmT7FA72IRNv1Lwc2Vma8H1TCDLRHwK9ZXz0+PQT
BeNP6Mt2fTK+v3R33bIUbryv+yzqdiEMm7NBCa2GzNgjBkSIIH41DVvyRGWCBCdmI1yVRmLWj9hB
VIVoo1Jg0Js+8ckbyEiMs7F9W58sloARcJL4NMoBXOoCURYALvEpP6M07CA/3/vlwNZEQigyjK7t
1Lcmq9hZIrQhjrbGNdGT/rF04Isksn5aoKWDip4Zn1N7OXtFRjLMk/gC+hYHrDbBjFcQfDWo5hPE
S+YjrzBpEtOILR3jjx736RSZlxE1FJkdeGSOYLAGIqw+yo+FSoV048mFM4phALawGkLAhR0rftjK
aygOm2EfXVKQINBFYcoBBVMvwAGvWRycOEMgkFdMy3Yh72HST+LHA8zufEMLZrFBqS/A57WsyIF0
htdW3ZXlI2lOrjKpzQDfsAyyY2QDtFTBwj2u80zNDdg1Xq+WXmqjXvMEROHMrHmPqudgUszXkodE
8/XmqvdmROaYC2qiCrWT7NQJSwnSWarpQkP2MTVvdLXdOei4Vq98zw6Utd9kckENxzZoE1Q+MuDN
f6eCf8uCAurUjho1ERpyALlZ5xy2tLFJYRNEAWJNNMxVQdW6pKUY0aH+TGRFyXF4cMeQFq81AJ+l
tDRB/O1s1BMWWIn8yIYOhq9Rau13FInV9KglWq3TQ1yjqncT6aJcyZv5KjJ30+rbSJH67fpHK6dX
Wt1Z/0nJ8QwvT3eRFyNQHTzdGYlumAwpjuhKHFA06LOVBZYp+iN84wEKa5Pnp7LmHCqHWPNdnr4M
zS+nFPW9vDN4O/4hAOqqNwQN7YA+pEFQmnz7Qfe/9DmCg2/SKp+g/P02WY8ZVj1ryGTNslTcRuC3
IfOvORHvRPLREVuaZ1lDF/LTyzqJaemcRGBJAwHcPHSl35t9paEe5z74JV1eDGqri2OBKVkfHk5d
UBcfgrCHbvN2kqPbeyDmsijDAcmmFOMymAqdK5W/HYiebw7RJhp4Sdq3EdxgR8NISVsjj96qYQ3a
mlYEJHDQZMRqBG4x34fwAitKQPV1/+52E9yWFoocKslLJO07FMzWPTVderwiEUWiN/Zkgd9j359f
p0pT+2hswJw6DnE9e05I2fusqR8SnrEDMmk2//1Y0y5yTdwM4tiAVqyvUyPni/pWM0L2cthm94nh
UYs0yc2di/FK6R5VPMhF3CiW4hcOIJtFOBkT5FLKfH6mHWPBzgxoXKYHpphc0e4s97Z+/kthHKk/
Lm7x9MEt+lXIE0DlBjU75QvEFJ5jRXhIxbEg9DkkQZejiUJjschnZR1KsL1OTz4Blm+cNzq/5HD8
4reu3py7i45BtsuOPW4mLHuR/viO2TVnjyVVKxoLZMNYJbaELE96TOMZ+PytsWMwURzZId9erP4X
qVGJ0KgUUAiKX4fbHf33h4IqKOfTNnK+NBco+gLU9Vo66aifIeuLY1PpESrykw7TTqzfDGY65uig
HORTxivnufInZqee9qfSEF10LboWhCj8vFQbKyAMGW15OUA9A3XoyitaSs3GihaOnZYUH/r4VYvS
zBh7Zt32t0MYRep5iPLDhnZCI9F3llhze00fO1lY8Ka6vFb64h/WpB+VlPSAgDvgeI8H/w/MQbi9
dMFtmkDeytr9Pdkt52dbm2v5eWUAkedRo9GvpdfbSN9+E2gi6+Lk/THIHqv0yM64mjtpwT+QKogg
aBDxN4AcUSYm5mq/wcMOLXfPhtD8Ln5MaX525m8l+SpCGvUMZ1ELrA6FBffD0uZPZVXgoavY6o4S
HjZOZ3/52Hie8iq/qj322c2UdHj4IAtgk1Yx2kQDWjr4GJM+ZJxKVEAN7EUB0LWBGYLdlzB92ZsW
yD1I4IaIPyD1KRRQnCb4ROk8cT9IPMpQHIcmUsK/uPuhDx74yd4gDMUL7Ev6ropRlUTm9I4Jeqwi
KbJgI4XgUV7kk+zLfA7xJNpwSDu+uNWBSFvRhwbNahFOF5yJ9MG6L38ZX3TdDAipTx05muq6y9/8
KQNvDazmxMSeVYwUbzhgYRCDzwDc9KY/bsB39Bi5/uennBPuwamriZEK7XW2vnLu5aOOk25xUdAz
1aHce+6U9unnRBzfRzSD+XouUX+YTv+5KmkYEcRVOoKCAuPb7zS/6YYvpMGbxUmKd6ItCbJ7/cnc
uHIUF4xxVJDVPu7zh68Mb6uWD4mAWJM9BryXJxMDMmu5cvCHFBNfGPBjP1uPKgHKW6euZazXTn4s
46RG7atHTzzOTRnYcVP94QzgBVEybzWlY3VSx+DEn7fji/ZUA2KYuDQIwV98OEOjKVDygAa3y1xp
nKePJLunvFLIds3vafYGI3bsvwR614mSJRPDIWYx03Y+Ts31mRpVqwqxRw+sXx/UzCAO04ErS5Tf
cGGyID/JYyUmgt+kJ1m8/f9pS0Sl+5xRXfQPrcNH1XxeQqQYATfPppL2tAr7OxP07RJ1ZQzUGYh+
kVWoaIejzHkBVWf4+bQ+gD1dTA9phSJYDspQP6s6IKLDRodpOz5EJLnoYmrEIMrg/YjVVONNSqaS
XysA9bd7UwjXDlhIXSzaLOCBNqLA3zhXZkXR2arAFMJ+YMddqdbm+EJ2II3k5+AbPp0yQspB0ah0
yUQG3fBN4btsCm161VV7ow16tFVza5yvaq6PKyqabK0B1yT4biPYadlVBMlVUCqEiLHc94W42Krx
KTiHa7jhaZ6gzGt3K3z8XuO6dJ25KcL/R74TcS7ksXMZWjpcPyUBjNkAXrUhM3xzGKIL1uLerosp
MQlO1SqSDI4EjtgCWGvWj9Y4H5UK0A24s+RS33RZjeCHyyYF8VvVEvN5RbqatmkmmSO7tU8QLQR3
cP+qz+icKpdfFGDIhtAT0cFKczF/MzWuGCfba5FSbOlEHukb6fyHHO5qRKHxTqZ0SmLGPO0M+BlH
rIbTC+M8XnLLRxNl+ehsy+Dxv/+XDx0DUVbUIE81IVjafgTIprboOB1avBBwjyKVbR3tr0Hn1bHt
MMEDEuXeh28b9eRsvUySLAM2tjxWr3MDkiGBsJAOhd6LN5DJwEiGcgNLWqKn2GKdFIW2cTbdYT2j
eIR4Wwcuiftv+9kiHsyJpnniARRuT0sb3JB7IZX+3viZ5DiDjIoNWpA2+wgeGw3VrxG+JXij/9dS
txbEOO5z3rNY1J0YKoqqBscB9A0X4wOh9JesK3w5FPf7xun8w+BwOgvKMZRqcOBnkH2rhYWy1F5P
9DQFi8A8QS8bG+z6TctrUGh2Opy7tGjtYdiiQWfJVdRWiBiy5ezBabmhizjop2co3GyZDF4BYd4N
oCbw6kaMhSlhFm5x8bYdKQZp0UnqubWpQoQNZEr6hlLlbfWCEdrzjLzyq/dH/vTQwDKjB8Ys8gk7
iKpvVHCG0d+mOWSS0Mgn5njEweur4wXrUs+wt0Hiov5YoQviYx7mzPeiKhyQlWa4cI9b8F3cvs9A
kO29sHt8T3GDqlRXN05oq5VtBMmCjPmlPu0ngdnB9Fl3m872b06/iTIlGFninzZ7mx6gpqpFaR8n
X2rufvauJ8mpF0pkCczPNItzw1HlyG4p16s5O/Y33LO4+wGzW8ieNeLMFFRE1qQuZ5ZArqcJrY2p
pOkRL/+6yBUw0kdlUUQv4otnt7Tonb6qouWWff4lHTLNmTczNVfMgZz7pRcEGeQnfKCEyCEC72WM
rB6CmbGeu3uv/3J3ZwHaFJougwgp5l5VEeuoLK/wqyZ1LaRNvrlMAv8Z5PqHHt/S3yVS648K8FUU
PA/pMuk/IotanZYclljrRRwAnjAAe7IQMpuH/ICUqvUmBnpCXWHvIm7JUfT5PPSO20XZZ+Rl6/LK
L93CgjdCCPPapiWNx+nI//elYKA8VG3oi8L3fg42eaTE8b0CkUODzdN3GskeWqrJoGaviyrWwzWe
TU47BHxrJS8lvqBcmUJ9R+Yw1igx21oLwaMrnOQ/2mkTtu6gY0r7s57FZb2gpRSG640Y9z0I35Lf
Mt5OmReGo33ETflJr84v53fH+KRv0LTTDX4xaXjMxLfiLHpr3K/8B9WzdW2H/k8pEMUN/b3czgjP
9aPeBcKO8Knumc9WG+c/0KlGtvZ0ct/ygtTUQlUNQ+cf+v5RVk0QlItUbibD2yRR7+vh8zrFPX8B
oPlZLoVhIODXkIv1k7sxYRBfFLtlZ/m5xhEFKisGZh/B0meCf/Iegc6x57uEZARAlJ7ztsKQXfHn
7JXe4gkrya09g5mtc/eJE2hbVwwT4VdNz0PHcvY4veZp0n8WuAIkswYkSC8dFERmo2lnZeuWAPQP
k33Tn521Coy1GCTy8A5EPEzhAmOpGm+a1OOqgjclM/rokxeH4mu57KSLjuNdemJA5pnexxmio5uz
oK7a/b6bnCzoC9AbpniD4n1vSFYOH2wGI3xEz9tMtqfCGU6y74wG6lVLn0DvEVJqb/fCEvavhaBJ
mLQsyQaLY4h5yyON5cOvnGIhxK/LI9vtVZEx/4kK7RNjoajL+iuD3IEItn29/N4CCY1F4fd69iLM
RpYM8WEtLWEMPkS2+hLTZWA5AxmojaBjWbLc2pPvFRa8+Ee3C7Hr8Cu23p9Ri+GRpQKKE6dZyqaI
nt0a2dKXj/AeSD18oU3BnQE3oFWYuBANSgiyjTc0mPWP7Tjce4jR5vYGlM258VRMQRkorFiKeODG
0f+ICquRCNcTQTdr8aT/0EUcWfE013M7cRUt/TnvHoHtmEQvKRUQRxbP4UGXCmthQIPi65Rfoiv5
yayDLJ+Gr+va/8u1U4MkFDBQ5f9fz4nXVNlI30h9OHkU9L9I7Q6jXFsLNSskw9ZXWTX6MwsTephh
WYRKgGJiT2NirwGOIWHU4ISdP8GJkb3RhD8TVqVgcJ+T8hKnraucEVWx+Q77YDafuN+wxAIdFOpW
3VDuhw7FCSOedfyedtSh2OkBVlzWPjMqCWdAvJ6p18MJADx9lVnjmF/IJpVCy5e4+P8U1kuuxYGU
55cHftWLlNT53bWQ7NDuAueqpqQ9Iadd11hYShgzvEzsanebDa5pbluob3vJcPbirW0dfYBczM60
tVxtnlPg9k1Gryf8qmkDfMsRJD6YA6NLkpDzKZ5cEId0owcnz2LsbVszSNnYp5uF1ToXTfaI3Upk
KQS1Qpua9EtAm9GFdZfGgcfRgoxpxfqLbRKLnnKDVeWwailvCUlystwrqgUlvExO1Q8XRlvHCBQq
roeYe9LL9HmqpGg0qC9ElCgXC9QY2Mbf1uCiaNzbrOsPRoD4jjAy9vUXOakcl9r3a41P+zvwIIY7
fQkGynPaNu0SEZV5u93D78uN2rEM94jxi+VuhGjGewj3eOWRj9NIV5Qf1rSsMvMBsXNLTV0rYRTf
MKbIDb1uKgcm9UulYH9U696RQofqR4KI5ToykTZltoSTN+N7BrPOWrEwQyoAlfR2ziAceVG4fR+1
vE1w4x86OMv/R5on/x9kxZEB9ZSEvDjwuGy0qqLjszggYAq4YVfz3UhyBwAKzKzP9d80DIgBxTlX
dTUZaoDjtGxba61UcPDhwarGDxO6IAH4+d2tQbbNZvyxJLVXSQA1PtT9FC9/01HPkUWeTvruj0z3
ybmG35fLu/GPL1o8VxSjj1xVUM0OoVOfKf6UEy/GMzrPpwpfq3b73GW+ekP6yJXJ6gYy2JquMwvl
AWKnYBj/HQwm43QgusUFYB28Um89DdOoLo+lCU3Na4UOJj3TZU6fMMPALwxqHMQySv3HRCR0kkLJ
HbIwZOXwesXncVvQRly7Ky68Ui40CI5SrZwbvGPRPzZ/WzS4YVevEN0YmiCxVXnPD7GEP/xlkWIE
r1R87fMGd+2zqUH9tj7ZhrdUpOs9muro0aPRfLSe1C7rR2zo+vZ3EaFH6NxpeZXEWVgnDPIsk+Kj
lZOUszp8NZCnGlCOoWisf7h0166xgjUoDcT7vFA6Jv2mzpduUo0/kvQZKIqC/1x8G8dSi/nNVM86
UvSHhSgeol9wMesxkSjwyYiIz/79nBiP4jlSUUWrSiNlijJrA035L7DLzqNScQ+IiLWiobFxIouO
4Y1xqBU+QSJefguC0jRWPtzOS8YaQoOGMlFR3Y+MpMQ67ia0D4joEgvhoiNa9hED8gqkhDo52nih
JL/SeHHbWqGP1wgLfI+73ntK7lyFXPkD807vfZ2vfTHNDB8n2+Lqyv6+bSQNARWPAgZsQohnkSJw
M8fJvJ91rdzoiBaKwuCZanXc9OamQuuKEOasEWFWWxsyZOzn4HCl1KMaCLUZJF6MaUHE6CpF7A3I
MVl/mLTY+Iuk70SGPrNId0Fib56+OMcMzQAG/5EVEFhoFUqmfjYb0DMcxwHZJVyXBDKA+p+H3370
jqU3Tt8+RyjONaRWYj14/C91JafEcoG1beP0SF3OV6LzbdxSmgM5Kl1fh56qin1BFboOySOSRqxX
IPUTTTbpkWxhHLxKvMc5QeBiPgfNt+kaeQRDgDUIKXJlHtqH6iOPa2o4/+u90zBUbTYfhxu4buO5
tvOsTYDGM7V2yS2S8J92TYbV2DJfZr2RllCNtPlORYcNA6xPHC4+E74M/2+Fly1JzF8PdtMrLVwh
aL39vkQShRP1//n5GrPw/8jvNse36Ppln9iLXDn4FyE036Dzdyh20mFbtpVttFjFnXFaTEqr3q5g
pkrBd5vWC+s48Quy/xyL1GbUzj+QIxmmhaNs2OAGhwnoIaOVBGRm67OiGExwwBis9Sh1kTADLuwE
WHVxGcNKexa0mGJNxbPPx40eAqVQQpObbsUXMuP9Tq7k2RwIV8Yj1m4wkQMYNk2S8sC9AOg69WOK
FblqrAnYxCMOWQiJorJ2xZU9GlfQK9QGx92UF+hqk38BTd4SmDfapJJX798qUCBLLYTTKBXNVEnc
ftwErC/thmQdqjjLaCAvdLpMua9sXuavzHJpJhv3ZY4kSNiv3cAUpT93XvEbQrn8YDRFLbLyOQMj
uOl9Lp60YMwCdYjObbh8Jua7X62uRIWtSyVW/gFR+4L9EjtZIQAbJ2x56JIde5bk4/q6MH53pPNY
LQ1gzR/3g5qdzOaFyKn/BLZ2gqIJ6XlYsN7xTnW1rSVWNaSIbEUz6dztZAa4p/MoGbrCd7IwG3Si
u25111a1891jn8EFbHm5fmo5FlmaqjEOuBVRxeC0RQwH3uBWk+896ZSchUNpEUqCWWgoQoXWVz83
dQAfWrJJQ9qIwZZDjSf+rtULwIIrsUu388Ml4SH3N0VlhHyqCORy6EfXWaq8EZ7Df6a8QpOs3phg
ys7rAZFaLW8BIL82HkhJOuN650/6YJoITr6r+ylU0ffhUWgIvvB3gRfgg9p8Wb3C4cnknA27f25r
UL6C9cIep6Xv4KqN7Mo2Vnv8Ypz5Q9fuK8l5pHjU1bgaVvfgviLZRETZXq4+XhtISZRPiixSz9m6
Te/Z0TGGSDx0GHitRDtFtYpG4+7NXA1y2M3rq0YljZ1RPNpHUywcfkGfViYiVGzNg5ZoCNt+VoOE
cOoxENGgXR4xApZH3m0popcWqYYXmp84Rjrw3dP2DhG6xwxh45bBsjYwBUiP5njQZl7Qeui5HrPZ
n0xKL3bADdDHE0cVGPI8DqFA8Sh3OF8OPUYkpLOZQsRLdMsXfbaAU4806XLEoF4abRcyN8DwI/B2
envci3YwUAvcBeUOdFSQt4H03Xe4fpvcO5WP0p4nK1o3KPDczIwZVOZ3cznvZSfkDYCCS4D0yaXj
g/qlBJOfK2WK5dXcq6m6gGS7mpgPST3mSh0habAhUv8qj8V+IL95o2IsL7b4LJoCDwYWPNcEnmoK
lk1rCsJjnr2DLwSIpzO/2oqEdIHELL5Pwpz4eMC4XHogyGzUBPn095yBdB35pGa4lslROEiQk4g4
t2Z9+ZtpdnFCC0WGHOqm6BTmNNuTTj+JsQGP8XrvbbiB94/RkRCvOAbWjabvZwhurFspktlTWrVg
0XqL9E1mG+HDtTAHlqq1T6fI8ZN05iN41ZqRRf4N76hCyOO1NuoxPnj40GkE9CK5aQtSksAy+0At
EKQi7E0bLZqAaCCxQmU2yi1ELNvCuH/4HbHeWU+rGx+owuQ1LciXcfwSyxRPj9v0QovdTTu+yi2c
R2nY6XeFXN7FFYm7Q7Yc/EUWQ7XOU2Sj8Aj7kVLHxo12FvkoeAVAQ3X0TE2ErjoQfpkGJGF/p98U
f8H8Mg2HldXot6sttuhXiR3eAkDHtBF+j5qkOcx+bAydPtwIRwz0f/vbe20CDKd2q8iIxDoB+ell
s1ZE8TmaUcAgPbLrwYKJlFS2qj18iUmwK+8YWlmv4DijdHjaE4PeCj2jcSDtlTnpZpl9SRQ8xBw2
K5sMmCEgjZjDSi+EgqYccW1V6oaS2qNrqWViG7KLiASAKknbK6zKV/wCou7Wx9pqwFS0ZFeznv0C
4ZZNg/J9NyGBBTLq1PBGNOlMxOXGZGmbwHj79YgfptCI2bVfy0uDOKo8VDCR0EaZaxIKWuJ9qRGz
8kcqRGBCT7aEQ2y6BWS6lP4pzznNGqGoiW8SbLz+L7/2XTohj06yGMGN7GU4d+ishqlEdAoV0kpI
T7VuK0zDiRgQ0ouCtea/ECDKRGRTbdnIuZ/rEzKWXEzRMPEQ26QPvdNJIQ0L/ABT5Lo44FAyFnvt
H2KjH028wf9ZXyG880VYRgdPwxzYj10hwp1rvKP3J5QsYQNAk/oc0wcvpydGdR9fzuvqRaLHr/OT
AVjk+BkLta4/gXpZ2B0CZO2Dffy+9NYiYwFUmIjFiCdkIENirNXjwbq/twZ3yTJRyD0WwbaWt4Kx
IF3uaZO3sxJFnlc4giG+EzRg8MNYl51j8Ljo5laK9fEq23iOgW+Mze6DbOGJUOWiPEOLXEidQrts
jlvI8pMK4pAKbFrQvH7zMLAclp7E93+8lUMRSTXcxwX+HiDha1Ct5fJznhz01Sygh6TeMItuWsAa
542+D7G2POfbD49hXGfSeJCje9l+85c/7+3T/pUGGsP1k5daEXkUsS/1Ni/hNybHQm+dkegA2CKq
G/x1tCuBqy4BHJdgHKlU2NXlr6d8PFEfRvztmFCeNDMOusYKSzl6hDF+BbizyX31mqQGdiiSa3yT
E7z0ilPl7d+HaEuBYHnQ3ccZAFexXO9TA5//S23vISyuktFI2gA2KAapVwRbiLFgovtub65rslCP
GFUtKFx98jLVBbIRXz11zaiRT9bPUz7TXT/xuoaT2SJG5MqQCccUuuPSy5zayk4DbDjPax7Jtv5k
fR8aeuonEjMdW1Da50YgHJVSwgjmxULClBmmtQoP5OYhCB20aujwTrOQlQmsPlwP6HGu4/W99Pu3
C7Tk7GZ+7HIxd1z3RsKbwmNFDj8UIsBEaagz8mbdyqsfm9Yk7xZrox4ZGgTanb1TtMZdivGRcpWU
q3IOEdRKcSmx3MrRG8X+j47zEaAyMiqG5xpbnrUA3i5KgGZMwQU22XPoT17jpRJ6XjfCQ/LPqhu5
ubDDoeB/vfDuEzsQR9XsP/AI49+FvbbFqru1LDE8QS9fWz/OwpQW7JGX5h6alIPoPqKSiKKbVatr
BBqYE2ddTerJ4Fc1vqjhL6YsmWaZ5yyrHPghstiwL4gvL4loza2HDS3ARYw/hiWwPP4lzDMOzKhG
EQ6chd8eAYsZDoDGC4Z+Gv5K9fKZx3XnFzskTXN0bUzrxTJLbFeEDiKCauYupjXzXJUwAQEKKt74
n5EXpRdtqHtBCaFDq1NgTNFZB9ggziYYL+c0qFBtT1UkBez424nRWAy4aZqXJiRUf0tetZKN0xwl
gICParc/+9HEp/OmBeop/UHzH8vAylDBLpmJlb8lGUnasrdqdHPtBbuDRzPepBbKRr1HE+rgFx8k
hCsfRlGnlLzl4SapTbEDPPS7d6EndZj6c9TAcfR3bUqJlUiMKderbukeT3AzLTqa7ra0jpsm5hWK
gcyQTdrSIpikG9Um+DIDg2mXuhPJ4vAnSbI9oB8AMdkhWKQbK+zVT1J6JKhYMgwKDITV8XPlgBSp
4b9ye1QXqBzpk6V312hdjKbLzr7U6DUS+mY/0sSQwxv9aewSjfQpJmh6C5VGm8mme54nUf2UGpXT
Q+fkJcfmksZclmdvAEXFlwTCHxz3b/LNHFbXvRizXxOXOhr+e+rvgEBE2G2EX+sDmbaxaiu2eEo9
Nsru1oQVyvF2eGUoTIbmoCM8VLsArB43I8+8FKOO+QRpUsi4Bu6BpABeO6axNb7BdSgL+1v61ay/
drDtjYTqvx9cXGmGPQMleHp1vBfaCABtsCjxexjsE8VpcHfRTBT/RxFy1PKdoNHzABKkuisGyz0w
+EiR11Ti9P3KdY42NYRty1UL5TbiYVvZSE2SiU76YrRLJb0aeiYsAz+DkBXYc+fSqUZewvQ6NmBI
wEcqdrIZqZZqjnxqBBBPC10n5Fz16Pz5rfCcV3V849ZeOcov5caSf5BK1VyydlUbkqbwSjDsJJMY
Bz/CUKrh/rMBzVEhBUHM++LF51SIwsh8Bj8C8Am6ixrskq/XXMmUiiVoU0CqB3HyDD3scAujUZXo
d6hwVYyxOx0R8BziUmt1Jc2YfYyoGNXJnIVTHjX2rbIVs0x+9j8R1OahK9oJ7PCBtLEN9sYH4wM3
UU1S737hpyI5WhKXUa1S/gVkRQpUzXrRAzyZoBIq12zcFQ6LNSQ6/LL0IYlFfB+uS2BCFq1FV4zP
65yaalnAnhDts+A1NRkYbistRqNYIUyd6n9jDPhhmYWXE3cIXVNult5p1u9ysxW+RsipLxU32Kgb
WbtQF0a+t8mzEVqbk33xH3JnIu51Dsmf1vXNB93dV9r+Y1ahxcQ5b68sbDMM+vqQ3UnqpjTpCC3o
YnhENo8Wjry5voFHXD9i+yzhRTzSmRyiACCYBPsVqGixcJFK5n+1fkvR/QGtYxXUtp/Z2Y9ZQWzN
eG6G27pxvTB4saHB6wBX4Kghh/El3AckkOZ5TMbXvBVeyeJ9w40t6NX1rN+vp/KIr3r8Gh4+4Za3
TRECnSX47i7kwXC2cuUo8MNebAdJLpdra61yZEoiDSRh+hQU7ns7kqO9r5RLGhDSHmrUypzGNHn9
1z7TyEbx9BGapk7cvZeMcTZMDggv5EYcZe2VhCBiUnv46Tky2Y0xPPPdAt4fue2eyY3PaL7bm/i2
r3ijEyrH915nNdzpA8DJT0fk7LkKS2ITMoC4Qtg1t46vYOSbCai5OGUEAsncsv3q1WJYzl7pOA/y
nPesw0CIpWkH7aGW5IrOYFmPu7ReaEyufRCgOJZIUtMyLZgSotgodNR1k7THkePDKiA8oA2Oa11p
jL9SvrWDHdObgDRqvotF5rx2J7R0DD2ODio5Qi0mG8/4plLzTMcmpVMu4Xf0lnQ6Hl8u6lnWsfZs
YZ8Yy5NcWrCm1+GaSuTG2GwrmkG0TPJxOt5V8IynMhlEpQq290c8M/mlf3hSGyXwxqiGNPuwcmuy
5gucc982XoBlGITCy8TGDqMHKIQ/YKhef/EqKzQWhzsEovdHDe6hw/0LVyX4+s7WYUzMBD/ufPgh
kBHT5AtzluSzmM9qb0NhYGUnERnyuC2hAl/eubWJvX/qNYFh6Yf1dlf3occoG5m/3CtIwbkY5K2x
KgbHHzPYwZ91OMDuy6Am0UWvr7fQyPrzyfNCyy+OxIFoVLKp6eoT8QBXDdJTpSIdWCgiQtz37MXZ
4lGYQUGIJ+kGL7L6CVs+LdPPCZBlddWK3P+znU1VQtZpHa2cj4h6EpHIwhcYymV4Z8Q5N8Fhq1En
bDn7TKHt4Kq2PwDlMCtAMOczaDx+vDJ0fsWKiYQNFSLPT9xRd5vaLZObgTX76Sy2uWFfYUj0cyzO
C50Bs4RbkGendPAPfMPCBcXKkInEwmdEf8b3HMWRnWg1a7mupWOZsZjRhJMpMMQbLaLBWed5psDw
AgSQKUPDWSW4dROjia8w9h557EuzL9YB1uaRXLBYE/nr3jF+44tFXiehm/9I15dEA8pDPhTbF9gu
B0e0Gx8IgE9Q0PNsueHaPujO4cbI5ehhRt4sBAZpNRCj0Mtt6auyruorQ91tc1H7KeJS/bT+3HY1
/OSfNB50m2tBcyX3Ez4u87fRdhK5dXTxjG7CZApJRxASbeCgwBCqL4dH9kKvsIF5vjvFAmhxPepU
2gBv9E3Yt5bGVHfxQPXGjupbsnZjY/TqVdZkZzTGxRSfmvTe+VCk1KlUKSMJ3mgsY1dlbs2UWbDP
6bb9jbBwWMMMbwlIV4qJ9kYh0Zi6CgaC7w78aeKoA5YUCikSZccMLTRNOTBVb00hv1sc7P/afoCp
9f41xDVs+vzskGhJUiDfrXGLOJO4EKi+6qz1J5k1qZurYpMzOdkoDXfiDNOn01vUW8Qsw3YY5aQL
tTuHzXIdTYgVNesjf5NEEL6vgF1d+JUSWRo7jIpfbvBE/HUBlzNMDVKS1nEAoOFN4CYYrKH0ZuxQ
V2Xh5u65JXDHSpByWJ5UCBfmdwV4LqiTfOreYfvg6yv0WoCFT9vrt6AziVR5f8XGHoO3CyPf42cN
twb1FtiN1qXu4i+WYBOtW0HSXZYi0WMj84iuA5/jNilkKgmZ7pCriGLax7DWdYBW9BJUlZXYv9u4
WJ2V6Qr7gEleTteS+H3X8TLoJ9kq9dRm1z2eiC+iOiwBEhlhUaLJTpHcwxP+NrHxQRT7K02vTY1k
Us5YSJCtNkbrYzKhj7q1FvR+JlyqQVubxAoSU1+A9jmqlzSiE7rGFBM8myMs8bQRE36TtuHFv7To
6NFI+E1KcGQTsn4VguBo09Sdh7iBWuGF+txjYAnJ0PLTlJfTDxXZyodDa2U4JLMQ8iqe7MrNYaye
HV+RmGDwN0H6AVqjBp1b/DYg08Bsflbc31vlxUDxSeMViuYw9p5LamIfkATf/eksma1mpLJ3iwgD
WKTz3kS/DvyYFrYD/H3/7JFQulUW4g9mhCrvmrJboVloFnMFrpnva28tBj3r4Q7HHwusCcfwVqyz
eTmT63HVfOKAMibm/UfNc6iMNgNGPJFbkbQJkAt4IIZ53cY83oFOQisUY6whI17YDpOGRMomEWPY
ewBHQOquEZiibLspJe+Kc9tiW8Yga4faf4fKh1BFok+oyoaTlM41j66aCozAJZZStPqnDms+9T4a
AdxNLLakb9C+FQx8ZL3BZ6AidQNVbYFZwuc9YUG/+IQuKW/QDqayvZaoRqdkTE9pqHoCZSQ/Pfa8
++HbvG22KjDgPXODIuqdqrfTIq0lKhxobxbWePVyiTgcqulfmyXq6CMWQZbe4Ufb7pOObyNRI3KJ
P4ISUM29NateLVh4R4btISyeW8meXRugSyZcMBjBH1MKxPwwkJtyA1CM3vLg8eHdjkgikb1HrU+w
DeToPuSlk0oZJ+VsGB3XkA9UfMDNu7gihIpTGnT3OEeUCwMFuqbq1j/q7zRAJ2sLyAZwpM4p1iyy
KpD6JZ2x5qHCafYd/3PyBo8jTtXI9DsisOQRS1yksPnUCWXGD4hCWwar3MDWXvQ1M4YkDX1TbiT8
6m78m06W31iNhf5I3wsUmutERo28ZGY1yTE+MSw0aln0JwgCu2RIZf2WyMxcVcgJ0iRv7+hWilIJ
mGtBzlRS1SzCpABYcb3TDuhnP63cGWR4buTsLaBkQGuWm/gWVhM5rTBj+ohY7rfPOpKhxY+wQJcb
oPwrVkTpR8tAwyG6FvPN8DOTQrZl86Tn+LrsIN1pN9valnpi7254+HXEtuHaXCUUPI2SzzdMPG7M
qvJlAE0HTxtMSV78HQwPpdO0uyXbSRcJARJ5SfQ/1TZme7/qkTLgppzwuA1uOXzve+OIgXmU8n+M
nsNB13Yo/Z7b2D4UY0J/sBXqJuYOpRX1dfbqO/Y6ri4sJfstBjEn0Vt5fmde4rT/skfZp2Qemp5m
zPSBKeh7VP42yz/0NwEg73wrLcFfy9dG3OhI7bo6gs5rppZ/rldT6UxRRR0m7Bux32Y3fWyoQppH
WAAvqGZXsmgJMO61VuKtGiwVKszrp2hwkPGxvekSOt5HYOTDwpUtutEuC1/N4HzQBEYvVMsWssCk
mDBS8IiIrC3SPSYmfIEDMXW3vWx+xTf97/xghHOSMD4E0cTFVAqzGs6zzhm+5CfL5lau7dCWFYr9
aBXmSc6pHcgHnBmCgf/KKyJJsS2HuE44gbEowVufhFe8StvkDH9WezxFMr5IFa67W+H3TLjgqklk
FwNDAPfQaZpAt2rnvs2rbhPIrIX7xAyiN7ShhbRr7FN8Hyob+Uii1gLzjnr0+pTrUZ1extwrZnGB
6Hb7hYQOGvufRqkja4Sot3jlXj2HzGWuDn9RBahmphDKQjLVDIYw1YrcBerTlU7UiPO+PXyMaJ5n
/w6lVQ1hhDQ9hHyeF/xIbFJRcHrWfvbXaT4JLFvEZztaU13d3G/tovY2ZBrPEDLg1N8zD9hFJkQM
mW6gT9lRKec0s0mRluJ8pHIdK5QXdcWCxEmv66juQH+9hXCEmMtfucQeJyyi0uzNk0WY+XUEupst
ABDMsqfNY8A7toJO3sEn9bbfrOcfEWmE102HqLjJ4s/lCa4drZ8j7AjYj9VFZgvnFVLxUwnmCyzF
VmUDABBNPrqvkS0/9XJfATQblwi48mQUlUdqt50tvFxXJpGz2892dICTBxuuOiqRbLf/LNrWt5iL
gpoHs7MY86y27WMIK+Qmm5VWBe2QFKFAEUfRJ0Inh0l3C1mRvtNX92xTGuX4eC97x0+dME473eCE
rOkTNqamoB40Q7yCNZvayQNwgocKdG8TYzn/IbzA+jpM+VtPnp1ByP/VANkbz5y8DH1cf08xFqjn
TMdUZsPz6g12qhHUoJ22haAMJH5XyiGJgrUnfohq+PgA2D9i2HL3tpfo5j4gtJ8OkLYZHePRS3ik
oPSVPsaDXawRh2WsGJTs3FqkgSN9czENexbLZ4W60hbGVTEL2At/V3cvQelSAj/O3gu3cv52EM/D
HytOcYZwENffHSWK+zRffeSXX3+38Z8Dz6Am7JABpA/F3je8UwgwwLbDgsNOgRkDfHg1aQKv+r6l
oygg2IzR9ytSqBmdo+1Z4ugCKSLqMQSFPkgKxf5L0LchmcHSZJtcm9R6jHF0t6/nTQ26fSQ0g9II
nV0Emj6MBg1tKbKUUQaRRd/O/EDGcvJTPm6cDrmjde0ZSFB8lRNC/rQdwffNDPTLaDrRtfcnBipG
IYVFiJP8epSlR1X5MGWoKK56nao0468HuhJztYhkxGAN16aTQChpqcEhUdjQeEFDxNcS3VS+H6xo
00AzFGwGRQJX1KWBTxOP257oWXSOCE46esAS/LWMXLTRjgEZJwFRb9lPZ8jLFIqB2tp5miX7HcSx
ZzTV5bKx0OeKWBGPpsl+KHNQhEFvhpKQFgCOLz1D5oFMZAlj4Y9tlAD2BxhQzgKeBGzVcPga+CP7
sRy63Eu9eGaiFSlDylsYuTTv3bMlq5TjG9z0i/3vHBk4aQJL+kVOu+5M1NBlMO7JYt0OKDk51n/X
xPlQ7E67xar062IltCtxV59hoXUg25lK/j6Q/PmOJGqzFpRLk9jxR2R60W62T9ZIctfsL8miP+xW
dSAo1yGgLoL9MuBetJMFhkQadoLwkJMzdEnbSjoqm4no26UhlJnbW61H5LTOM1NCVNo1bxmxAiH6
n007RvPe8FQspiQomALIG9kfIvQ4Cnhf/NoCB9kb49aVZ9o+1eymQm+IkabRL3y86TlaIta6k0cC
qghZYwg0EQM+fyEoOCx3qqJzGChymTtewGOKTBl9xXFo1ePoXNBMohwua3JsfckjqUz1sDDdFYYO
Xo1rP/JSjuC9KmjPLo5S1pxQDGROWEJ2sPP7/547R97jrBISUgyZdn4f4lFLe36PfDhDsJWcIQJH
BWZjYmLIg1XZcfEBtL+ZxIiWeYUSL6OD+z+tjErXR22kRvlsiSvYHof5mf0/ZXcscvoQC3Byeapf
Kr0LLaGuCSxxGWlXdxOyjumyD3SQqe/a9iHpAtQRQxG/fKjhGuj/oTDFkSHWQ7JNYU/Nud4bqZLv
S+Gzxy9vJVrv/T0eBwKarwcCQBHetjxSkQ0eZjs9JirBNHf9VAOg7DwATmJR/tcywNq7X9K2FZJK
YjuerHNZ/0XjVyxNd0C5WSk0eJGRGA4lBislFQ+z0/BtisFrEYO34j+73gsePhi7nlOYea2tPuQs
hhCwjqoqlVnua7ZSYk+CkDW3BTXt3ZgW4VR0+ijDTHW8rcrMH0SljtjTKI6cN0z3Z7YyVkDck4HP
BpadeiVvXR4KwWfRlGvuZPWOsDdS1KVa/pOgZ1ducUkbe6iUy4cE9JtvQNapMOk9pfVp8RlxMi4/
ma1FZqwi5q487i/kgnl8xH0VOlyg/ytTwcDAofyF8qzCWi/OV0R7QA6E5I0HQgl9xkOph6goUN73
H+iKPE1LVT9E0bRly2X+gHAZ5/W/vkG77rGy0Tqfjq8Qz7fpKfRt5zZe1u7RqfM7ZFi9MUsiHUrY
epNdyUKB3h9gttzH1Swav1YpbmaoQCmx58UsIQO6sSojEmIxs601ZzXKYK23QdGBLKknRjw7/WPp
vGE+cG3hMOA8kxCZB/LpEXgDSB7vFEqHEEEx7niR2ZVKorXH6zXL+r34DGWtQIS18hFGzRQJuQHJ
xDY+ZoUvirO3vru8c/1+3top0SeHU+uqzEGlzbQCZQvq0Jz2XawKVZ89R9IFRFgBspo8IQEegEEe
Uuv3UUGa58Byn5K4ImKyPXbpCYEZZxMKCnOKN4jFZ/32+MQbyxErkAFBc5fcSwjaeI+yyuFQhb40
6j+v/OtDCptpqP7VevWrzDMOQNyUaQUBptW7udwansaJNOAQCcs8Wxg8d4rl3LGxy3j+mXCcL4Ou
d/mGOv0DZ0Di8Jih6aHGXOr0i8eCyGyUDBtDEkS1U40TMfJnyzN/H1Wmk/cT/kQ5gb0c9fEffdfL
pt+Oify0LZ3XCrWlQtmoG9sWUT6Q5z+C/6l3BVb/7gX1N/D+ckmdGMCtXYLahwttHoJYgqiPLpGo
r7R6Y3rve6M5fdoz48gcM7nUuv2VwAOrvi7ITBYWIr8ngvj6oKyiDR3yI0I7es2rtl1bS0XULD4i
HoZ+p/TL0FrEgTWXiC7mwvoyc5r11qu/JedrhKYtHVaYF5RYi9Du/gdRFScY3owqQhZD1rQN6qPW
Rec6kT6mnhOGg/IE6k1Yxb1H1N5LPpBzGn1ldKaAmZs0xplAdlyvbplwByN3a3kHgcxmV8KPSjpd
gPmepGCCocjZuyGB6Tc7EC50GsPJ50o71922t9wVzTecXwM2dLzCmp4FmwC3tvG2spx8VWGcaxQ1
4hAQIffBJEsEYe9uvjOTTO36hOMtQ2bDLXgqA+9vTNz4CIerISFLeOa4OoEWqn2FgTbzPtbCY+1K
W5zF28aPCmoHFXMTxN2DqEs2eFfOI5GzrCwUl+ti9zZKKwyva1euEyjw0zXYAL6GWuBucnVTxJPs
8e1ZTzk0oj55NqxhvSoQBjACqRsQRRxWdJvjLczYqJOX95CGhy4/JR+2RJlzZnW+ISm6U0Ffg6hq
DZUPft5S9dRkOs6rmPGqbcGGMOBrdp4qOT2nT8JOAlc3woTf8N95013qskzlejMoBpGhfaZJ8gVU
OUBo1SSqXMGSIbne6XEx454HwKyw7kHYZvxX+/u+5wzmz7DjyoFnYQSW7ocDyR3VF/nJIy6Jj0BR
Vjk1FnDVri3qUVBTEQBwrEgjtk9kHYazFDPjBcUcGm3jMgb+DpsCPX9oDF/RmkLHblOn7xge8xxz
k5scYQ0y0s56scFB3Zg/1/4Cosr5oeKD8VNolWiHbdEmgVi5L/xrfreXivxRZXyyDD4G9WetzX3W
I7kWA0MVSfhRQjVQLrmuNWnmVmL8V5xMh7EwjQ9ZS5uYGxznoA3YyOepSBaAJKDbhfqmAEyhKHal
S9hVHK6EHhDfetd30pdBcJBT6rFjVI2FC04/Eg+R6ppbaKMgZrsF0O2oRxAcpLVqJ5bbwKfkW5aC
fklXWc7zKTc+VBYINbdX7mlrMZzThYHJ/dqFXgsI3fre3vJLVFVKXl/gEHOMgBFDDNfP7hYAqxO6
JsmiQbHmYirT0IcJ2/J7nmy/Ah4Q4/NjZdaIBen+pJ1gr+bre1ILuj4YvRaRjvrHlynyzT9rKGNN
MK2d7Pk/H6/Qs1fhGOpJ5arIVW2qULGofxuzcjiwtDdRTsHnK8xFf0GjQkeJ8fe17SuISH3BBuAd
/g31uamJKvGMR5Nm2cj1EOHLfR1mKcHBeXTib81eU3TzJ/JCZ0iuntMQ61spTw9duZs6qfpd5jHI
ZbzKYGcuIZuzy2GfhXpM+aChZLdrDYYy6OPOY6y9bqWQ1S3OAbcdneBY3V8xsnVQBSGbQfs9oewE
fmw9IeixJZ0TgUogfpgnjdhTNVo5ZaB2P8Yf6ocqx6Pn8ihdShK2vOMFmr7NZQLKPs1PaFLJ7ebQ
om2uSd2/+JhiBdl7Ep7ddpEJValDXOzuGS5QzpaHhOqp2Us7mzhxMhqc42gpu35dRaC5ozpbMfM7
6sgkdm2h9V8RXEPsU4Pd+PUyy4xYBcK63+P9UWDgOfL5Jt4HEHxFeEoUZuVyba7PWnJdc3Nplskk
wfBxq28yTg3SqdHU5HmA4AsukIAUvIS98Rbb4XFibNVUmYmx03is0apRqKwQ+Z8zb3DfDolSfWQk
k8SXYL9HfB4haFBwa6lxpjx4FrdzvXBo3YEvUjRv9HjOfI8OdM8w5CYeWS96f/Ksna95uuDu4iwb
TaVQmeeUQzWlS3aWDPia+8mvheGWeHO+R7REAqhxhE0TF2QdH4wE4qdZAR1O1+mkv7u8Ud24R57g
n9Ss3orMMrdOvctvYJvSnOVlPL7tqwfSQXifjFD+dRIjrHRvIim4vXjEmLjcoZZDlmRmIcHk4bGU
fhWQy/e4nO9cG3m/IhLY6KNMg6KpBCONwNxYImU6cxeNu5nWaNlbmwG+5eqAGvR3Pm1Q5gisPFcO
hw6FMO505OmkcadIqxikKxkMi+I3gU1IDrRTChrBoG+3sbTED5vJuLyF01WUN/pLnHIuDgtH7Hz+
JpLRX+SPiQAsV/W5vYl+fd4FM8p2m3dl5u/oAjsKdXDqCOSGO+B6LYzCVKUwzN26hgkqXY4VFOKc
j3oYaeopUKh4VnoTXvOdMBOD7GEHZt8rPVyMcbj6ehZIYVmwJ2C5yeQ+uoOgu5Yn40RdAK7MvtJt
2qDUN0N6WNDkpCOEdcwUuPyzbKtu21VCoiAYg9/XuwEKzevbBsVrR5efiIumyDhTsoRVFX8EmN4Q
AcOH4mmUQd0kun563NuZ9BSQgw+8XF0dRdzIo5FQ2IWOUJq7xLIEx9Q/PXsShY01lScBdyc8uyJ6
3bQcz73tn2CV0eICitNg1Scu2XOK7AYUQKX7ix3OXj7xBrLx0S/JVSiMg22YL1VAF4OYlJQX3LFT
Ms+E16tM5sjlNXOOp26UTXMCyWVEsD6a/2GzBP1LmGpFcQvJWeUgVSjg0cwAdBBvOUcRXvUK/oGL
PEwRRmVaraKSgomxbyYS2cBPdofnIdlw8UDo1DgaBS1VxELG4iP0LDY+qwdN2nPesGHfKHC4Rrp9
Ow8O1QPSgsHXbNSmAEMSsWjvxKJU8x09knR+LyFXdEW4jmmlUyGW/N1CxuFWXN6zZlz/3HiohO2C
v+2xJvrAU+wzY4fD23jSTOXz7jbTo06kQM9kJfiLCPRt22iwLt0C0T+xaduY4u4sNcpPCHCNtCQy
3DC2MQPzAbIfy6XFxii+RRCpMkEJaNU7gbvrLDIZ+Y11XoAEHywqYp5aEkKCiK7FjMn7vDTfBWpw
ynCC5F8WsnJvj0PbmM+LHWOEYt0EEJzuZ3RDnCs7YYtPzIlsn6vF8rQ1BIyhDNWNFkpHCHIwGJlb
kU1fYlSa8rZf4L9YyQo8ZLt8pyMrFVZ4rLHCLiRAIP8rPm+J35dqLMnKYGYRIC9pMXS0HMWTPlPj
v1X/1QfksoreY+i/Vp1s/lk5sLJAjrOBPpe9B22aPBl33zb/Di6ce99VkCwgHnpheJx533up4UGR
7xOBlZvBFGch4yP21k0XDYxDkYeq+SY7mohmGhstHLyGoxOlGBeU3Z5eKzpRtzAqKg34jxlxsega
Qrb1RfN6DDYwml1B3ynA+V+fs0Q/MMqUuAaVPj7F7i7xBUgXCGbxG6RpeURqMxv2sRrSsqo8uvex
Vh6aJyQLRa9WkkLn5KKd+WX3kqZHQHwBUKkZZwFFRskWvbXyNpEjlSFmBvqlCzTNci6W5GKT3Zwv
r11MO/xtxW5mVaLaDumExAyE3xj2LMdTTesyzpzFIxwlBQMEEHPjIPL1TCEFf+v0+VeYee6zcV2P
yWPPkZoAOTlJPJRUSvco9l3Nvu5lnJfxlnVkWYCn87BRIyFkCS9ZLy6an2iQkPjpNRe1Qlkq3SSj
4p/X0oeObq/boEMWgGWFdsWUQaHOXtjSFxJZHpMibJ6tJWcpMxbOFshzxe7Rbv6dbH863gMdF+OW
sj3k+kPKJ9L9FtR9qearkM8tO41eFNOwCeTOokEsn2ibuA4PSj9S3C20pCkXqguglUakxSShhxJy
MfPLI1FoAx+pxS6H+3bBsZSGVH4vjeBaZ2aWadBjv3MZOp3fkJfI3HGupb9h4MBB4a+0JnIyGZ9m
MnSe0NlFPmpESdB63lCsdnDwaOP3M72Xfgw2QkC/MTWbWEBXVHmB4SfrKADMh2XrQNI1R7hx9jxZ
jqKx/BiRutYU37R/XeURdMwjS+f4s/hnDupKLYQMp56DeRu9UajXMLNQ7+GLZ4ARfz1seqSZ60pd
LYRyjRYYO2Pl04k0/iejeOK+IiFVkOhSfChEuSnYkvBKcSa/ZKqlNb3hXlFfGJkrhtkOl6X06Loj
Aw6C/Dpef6nsv2m6ji+Y48vE+ROolAg30IIc/772R/DynE2ichWJ6aaFaJwvaW90QLqbZt1SAyVM
uZZyYyIEM5eEdY7rLzxYtUdLE1TkxpW47Lp3qYIdb49JtiPKONPQ9aALDjzbCHPRWHm0SWnmt1/f
OVdn4uaTMRRa6+dGJWi7adI5HItbYdBixnsEny6ezGd1ZHKzlOrwIJOZHmgd0Lk9Is9mLfYfJrIA
zMPAITP9yBaGkC9ZUHn7i3TTRkLVqB2LooyCKkl+fdSw+Z8NDBmbHfJxFQdN/5pI45+fFtl6tIvU
O2pSMR09j/lL/c4vHtV8gw65sNd7jwD7USq7ymdzFLL+26p4IZlqLdHtAhDkPxcz0nKo2ncODxTM
Hm3xm+/wOqRNZNrasQcL0fc7ZR4HeobXt6o8D1i3miv85tbtKvgvc9Onwc2NS+3mQhRA1YLzy389
TLPLf6fTYAUuksvPmyp2GTsmywIctxs51GAvpRYHJjk8m4YYA2rxDnpJiMAVshisYXAZaabXAtiH
7eUWQ7eMcOipk35DIbB8HlxmuJybZfD1sRiK/Lw5CXjk6iQbaAsg4gqsQnp06L2Am2G8hCaQr/m2
28RrUYR4/p9OZt/cDRnONel1tCL0SvuwDjMo7KOHC+WNgJO6cI3dFxANjE4IF70rPVuxR8nHUj8i
+wm1VhuklfN55XklboNkYBpGaNrjVT0hJYQawQKMk+yCgNR0fn0b27ePFiv1qXQN/hk+aIYZdWm7
gW8SWGPUUOr/3/103hICmD0NtQICdhptq5RE/71rTqF/mEJpxGTbZ95W2kJ7hgXHye2j/2MMsKTn
WSTmTU6vBlK1ekpIN7qwnLmJTJSJxb/FGotesPsnzt2N7BZsxbyJAc4ddSQ/AQwyDV62whixTRwP
64lBvvCPhsGyAxRenYRbpsGs2plKl+t6IpkcUx1vfvjCKEj3Z2yEbbCPbXj6Rwxzq+nzqSHoXDn1
+LePgor4KWQ2RlrezJs8OLefpr0UBnr5DoRQOz62sFpbzW0Y//cJMrRFpIgHrk+CxvvYJHxuI4m5
fcL2/fRDy+ziRRdk386NjTaC6n4Sa54+3hb8QGq6np72+TmBbinUnLEnJ4Xx42ZieiL06Z6IZSBw
42pnYiCPLedW1Zt9se2BZre4g6xCtn+3z2NeesjqysNNz8HSrd+n7QJvV7D/jYwU+PZNqigGLI/N
ytIwfTI/6xs6u7KvinfsNb3q0bW0XyZHRWWdhheJUawBzCZUS5HhCWcGlhksFe4w/s2aMGy6KqQL
gVsqF3KaWduPlE+z8g3sNW23iVXoyy2UMSSoAcCC+ENZCxLhgmSZG+lGkcw+ZzYl5ZkTSWoP8RY6
l/4FSLpQEtA72cwdS0quGZQzE9U+MmUTQo9rB/ZWx43LQe5vCQda8hF9Mvp/n5H8vl4g1eEITIRj
1MA3x2G8RkW8MHjMN3b4A1iECiv7Amjgpzxc1hM0Oju9DAdxzr9gSh/q8/R/GxyQsyTW//U3OQ1J
xs+urRDmewx8S66BhbPUorcwY1NrFGClu7GP/wQWNS78p8UBppbtsVXH2YGP5nuO2Ecsf/odgzkk
aYWG4RgjLqBwrJL6t/CBQWbof6leUuCmxuqQXfwYgRyyti44IJxe9Xycux38mafqSa7U6aF5r8Hd
iFaFyoHtIOdjly1Olp2hbYqyswhSNsEwBo8MddgZ2x/hp5KjBZfnzed+JNGC0gJ/Rw3tzxl5UN/j
AUfzaYuHv7qbARGUEc2KhqRQYSjDhjPhwzoIxVhFPlbIqCLIXQSW7qvsnohdxC51TIJnkg7XIQbc
7obNp+mbbpQMvQN3EAboq+fr3vV3n+6lycRkT4AZjH4fCnnNI3aqwb7QpYrDNg+nm81EzlATxHbq
EHxIIUbKGELHW9Y6B5t0YuHIHCBth2ZVcteJwP4H2Pe7n6cTNVxRcR2wCA+KllRfJuk0jvFVHveD
IFSdQUjbRIXpZKZgV7jlcXqm6v/jGrYXaBtj61dStbH89wsoSrhqpI5a2hbXdBxc+0jc+rFW8jlw
Vg0mJdNIWjmNSJHsP8ZTqkpvMtQU5hdDo+CsNTLowDnmQdYdr0otc1PeXGN1p4G1/3ddXl28b51p
igElEjgJx9IUWMjygS1JfgNfgJ3c7QsghqG8LlHv1uL/kyJ3H8tWsHU+gq/9ct7gcYDcFN7u1ERR
x644oCe/NqKqrtYg1cpfk+qQyAN9Cx9T8YRfwpS1RHsN6P+/qqHMVSEmzKj4f+XSH392WBRUTXo8
xsv4Vpc9Rm8gZbP54ZxqLtokZYfmmMrPlv6psHESgn2tNJrhEI9Hg9A2AgLY3uoW67amYXOMCAch
iRcgJWhinneWCiXHv4Ke0Mu60+TQu6snNoTZ9e4ztsjPwr5DnBhHktBOm1BZDrsgkt7TYc0LVO0Y
tesipCOkmezt9kVO7O8/YCqmn2FQKE3nZTxdKd9WWjmZOA+8cHfUrLpvPmdvdn0IA4NVFBfNHvXJ
DEgrVW7XA2SgtBiEtOKxhm6bQVGiwOvZfsZX/JN0e10X0sp/qvr84BmxqAsh2WQv2kU/Vi+1oWoG
vdNbs7eo/6CDFNkUcEgPF7FYzK8/4+cN8o5Tgl8OZqLLeTUiN5puH1MU0s/LDstyKvpAEVortAsJ
1Mp1fv6AgSCH24Vngvn9iHFCV0FLai3uqN2WbdgBHRqqWgCGHoRBwqQzqpBJSQkehjBWHidM5yUG
Mo6wNSBXvNiwGkYJmX/K78nS7uvc1JSMxjCVF8HHmPBWRduCJWtlc95V04SaoSW1Hi8HJe+CNb18
cMNBiJL+Yv3c4fB21ryFMdHan34UfQYVRSE5glaQncVb9YECouzT+eKKdmjCS1gDD9qwBdP/F6B9
64aheTjBj8Xgh3D5SSzFpdfpDzqRvK1mXzo9iVsJbxZdQZpJLSuqvqA9/clyFem1UcuXOcTdxCGy
6whfW/DNl+kiyjazOPmLNoo2Ifmthm1/4Y5yhp9BMjmLzhUmp9EtEZicdMACMeBAzDz0kBs1l5R2
4Fy5rz0otzlfXP7OYYiMQojKJduhfhCz07BiwoneX0o8VzERglo4X/G7Ygbe0gCLmOb23gi9sdsc
hkMt4HlA8+AT4GbVCVIGWE4nfVxSzRPS0fKpBs4ee3Bc8IUXYIi2pgOzco3hS6E+VeGEh7N+b501
k2Q5pMUBqzTh3rxGcIJlB97f6MfdLD99nqAtNF2pM33fYuzQEcw+qsHSVaSkZdPe3AUuDrssxNWt
KFL6tjYW6sLcKV3+jbp6nOnd/dEG/5Xnl5wR6zlRKousWK+tqydmLi0z6L5n1gTlV1z0uknEn97o
ZbV5myzQfHl6PysiXNk6Q4yueAgsB0llTzw+MZEbgKbqwVCr5Uu7uV07eXVd+6/8n2f0f/2nUpgU
Yelv8f+Ky6owboUJ8v/FyzemsH6ABx/3b3Iw87ai33mARsBc1tUKdfw0Vl9KIVKDVwPGC1yyli35
BkxofSkVOj1uuZ+4RTZ3zmaReZL+eOCGWRDIJWSRybBwi0FAH6rAZIwI6jZe5LrB0W7twb6u+ov+
bspYp6Y3A1s2bRpS3fD3JD8/sWOroAAd3sEXonG2gxZ0lEahcDDtOqT2SuJY4YgJpZNz1XZZwEe2
8L/3G6IFFfERdtDrQNNvZhUhSYYA1AIQWBmjgG5cWpI1zIKkAn+/YW8YyiMaCcJ6aCudmewRR4Vg
yUaaEL3jOC9CcnknRpi0QYAeqq6BEL2yJfsQN+sflZnFARvcBHDss8KH4CHDXaBXuyV1CictpDeb
jY+zxOCNiUaoDnhePbzQxSG6TVVKfkf3XkptuhDGzfyJS9pkHeNMecxgag+oJ5ScyyfZHJmEeLW+
IrmfwHqE8rkAZuECKssVBnFWGV0WFuS4INplerKzjVTGgquh9h4uoZqGB6TRwIIjNwiB/uv8ft99
HAbY2q7bxAZG0fuuxUS7EQLYX+xT7ue1kHrOltb1I/rxvIWpteoS21aiiYHk7W7wQYBZExeBTDKx
vpKBPTvNRFEwT26ymH5Rewjk2yE0iJHtuDE2+HGfL0tjGSWHlyUEDyYGJtJWGoU8fDTA/3eW7dXa
EX4I21SK7w/NPLx3x4pFZG78dCmdvBcwYPj9g69NuxmEszQ8YNk6y0fJ0WYA0tGORkxgPsQU9ROa
KtXSBeiUtxsVzBvMOfaeSS2+gr9eS4oGhNTIze8Be2Awd7zfAPQvQ4IySzrFDTTAOCYfOj9l2FKk
d9yK8Q7rJjQwd4PjFiohU1K5RWnSGcQdV0WI5gFHFSoNJEeRGxF3nSeQIMPAA4aoxBe7riRdXmd9
MpNW0tpMY0Hw88cm7/QwJ7rUkJQ6FqKk0m9Kr+ojr5HrAdahsW/t4I3JUlccOeAIZG3FP2W8r5q5
Zcs7AktjJMs1TeFBHyOxQGFKJUQXgJipTy8/K1+onUMis0fIW9530ccTEXxTzBnNiDa3QiWIH0gi
aJvHlLLUSmFK4OK2N4KgaPAQJ41TiKIcyzWEcv6K5ajXzTpNJt9O3+axmh/8h14rqAbd3RFdIqVF
HEwlfCok7Tipx2aaS1oW8i/6BS8L4yiyWTXP2WUnl7wa8aYI99QPbTJrZwIYnUH9SdPhxJYdElpS
R32nDMb/AHSybzgfZ0rYHD+DvaIaTQZi8H+Nah3V5cmeABcfn4H5efHk/FspsXebaulYbmB8Q3WA
s5ldSMmDkyLKO8bCG+OzjYyfjK74z6KFjzfAgIEkBwhciyXYrpVtbAYekmsa0Zs9wDCfzCiXVCe+
doCma44YzO2uXSVLqphdk9U0SvS2+DXe/dWvkRWXabR03LNCTxWziafRAuyqedOHPJgUUv5fhtYF
GV7jIy9oqP++2HE9g/XDfFn2lb6pph5rnuL6lj+LQPSMNoEoVztAo/Iy83k2Nqgi/F5nnL+lE30c
sLg=
`protect end_protected
