`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
crsuNbGKr2+HGjsnrWAO3ApjaENLE5lmTkmDpqy6wXOqFQIJnrktoh4R9l/TVlY/BEwSOhFtvEbq
RKvf5np1ZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfoL36fNI5DjzIQX15YYPTK98uQI+Z0aMjl+hiAVWq0lzClrfpDjXWaPyQGiPvnYkkUnnCNmSyGP
qGrNm7GOsjezCGzMgQVr0792OKktWuV2kt0zVP1RUZuHk/37eznwh8N2o5rw+1YzW4dGzl1QbJom
tmB1UpBcp868gDBGaIo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nZKDyxkYA9uy2Xb3FwpEri9edMFM6SqsP4Aed0tRsVeeX445M1QANBu8GOl8sJ4QNxr6T3VU33/s
FK93SNbe96iXZq7rd0ZTftDGFn/wlb+m7r0WSjfp5pkNrLXaYMROFr5Y+cSF68dabG3s3COIhufS
z6LjxtxffkVZFl10/p5NYIyhVlCgj28/qTLowb5EYe1tZ0WPUAxBFuTyFKtX6X8Ha+x+nETiYK6i
PAhbV564AhzWOG1ohxDJJcn/sq1JfdeuDFdYSbNKycH1TqhYGY4rODz7EB10q4+UCVziUOr4Tv4R
NCotWnw5vu+fF2mIxu+vVyyYTSX+rhEfPs2iXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZ2XWhB75BM0Dt/9VMCHTjvBqUtECoyfIkFt8UyDN1IrerieLUkQavGMJnAyOgfgB2F9GkPnzVQV
7H9tsdZ87Y+A3ybRmsawN7gt2tqx/GGsvZlikuuSepi3sHN1vWxch8VpcI/SFn7CnlCh0jupM6VR
707+yLDj5AJkQVyH1LA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S4eCKuneguafnmn96ntdnponlGVTmyJu6zrxyF34ICbqsowM9Vhvgm6poU8XDQ/BrjS+RNPc37Fg
G4CZX64FNy0IB8M93ARmuOVvrGN2bYMf3jNRnVO/z1hOqr23u4iXXLcNjJcX+q+ntygTqDn+dkJa
tNf5JDJd7KcZbafDC5iOu1RcjafQnwlpqyaxuvNRdQkJM7f5tDyB/fmqWMaeSiYSf6cbwC2Jk6x0
7wUP2rAkEzcYQjkJqSGT74QQ9ZxpJuO1xNUbfsJDlmWbSmEyg55J46Q3XRBw9O4UV1TNB2XnSxvt
0rRnDIzS8sn75CDPR31VCmG8K+PwSCayofA3ZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12480)
`protect data_block
HGwVbJA7sypyD5yh/+WUmYczAUp9Ilw63ul2foAahIAqxWWNlG860q1IJCvcDi+ST5/TvxcuzPir
qt27wGW80Ur84JcU1ohvXeBLj7wUxE4SSH0YZIS2OeLGptmd6WoipbGBdDQqF0xVMMjgrKgcZErf
lwMei5al62lj0PDb+cw/LYrsWYwTZhEAh1QQr/aQVmVXX59BsDj9n1cBqUdrbtKzJF4iGjsn1KFy
IpTXkqC07+RbfwmuY1gtZL5gFNTUEmbshwCe5An75BA8XDF/ixRn3new5vA2QMpEc9jzrUs9VQjX
G3NwkT6Jrp0tH9X9Ci3PDiBu2Nt59+mPtjL8WWuVXJ5SnRA4FFDpXmnMDnzFiNHcuYFpm12rhIu1
2Dx7Cqj66JpzIn/pvq0apjYPvknsoYWVSZ9buI0fIE1eODqLhLJTiacql9p1J4xeZj6ikcOOEsM/
xsOzZgAKSYBkQ9cfAAwpvGnGUQUoEpEve06l/Jee4gCR59oqcpNaFk7awUmgg7Q/1h/ZGHuOk4m4
wYodU8wBf5YWkKYpL2Aq+ZoC/2e2soG4cbSDUTICLa92eYlK2Q3TZORaGeSjDLzLf+OyjZ7mRKxO
Wq2ZnOPLxlED5UqUvyNFYfVUyWC9ktHZ77PF2qlBSbL/MTUi0KI0AdJQ7p7YnRwKJnB/uGoEoDs8
AJfbaisVl0qjjej7tBX10auwAobsvdZc+MpeT2qbrhLVDoVD1aZ/mUO8PSszTcKXIpHU9XyMp38m
/bYmrhn9BhuQOKPx70XvyF+FKlCdq1+ZrBhm0sSXPCuuSu2DHXsR7KlL2JULPZ/WygMS3YbUI1zV
Lo2acO1o8wnIis/opw6BLBgBGI/nxxVtVVP7g3ISDTkyd3h7vBv03qyV2q8f0bu8CZesHx9PhAZf
UD5M+Y6dIWj9O5X4OglaOLQKnneSM3OeHlf+fkhk3ZUi47sz/1uHEbhp60TVhrUppoJhfS68U4Ii
cshkz6haEUb42OyQw2ufW2d2Kz3bc9iykcUkDyKBSr5HHfwF7r2PpeVsTtIl8K83j54sZVG8L220
KIwuveiXvuaHTD0cdzUDMb0xqX8RQfBWpSXwxp1Fll1WF1hvmsVmdfy8Ozz5pCDI1+FstTi+XL3+
T0opr5q3uekIuhDbd4oExxO0rctKeol65kOj+jfK4TjhkD4Zb8HtbkErvCPT/lCTAqB3tzZmmbq8
M8UKC18srv7p260omxmewaY78LGrnaD/SLanpKhDT0L5QkoeRewj/Ikz+e60rvsNMwOgYXQbhU8b
96fqfis08+wo3I+N3agwVvz9lazqVr5/qqajjwwNrAvyV1DtRB5sMC0g0gNrFpLJfOCS1+IG0tbn
QDy63/TpwwxpjcC045quOJ6kYs+Y07+GL0g0JS2oVuusjS6tMZ0MmHOiFU8BMCwT3Wgvm413RLt2
IUHH+t3G2X4XZnt9lZpkM5dEEX4fXqa4O5jDLJ10rNhlZmMilON/uebZxTG8LXWx+OqsUwEBfkNP
oxfyQf7+NzyalgoP+4q+7wybtPfTPvAdhO0hVGyFPmVeKIaJfmEVAtuJABfaHfEon8y/ncRhdOMn
gXXbrlgaVWC95YJ9emICdCRH0zv3NEVmxvHvwMWIE7dWthgB2+Y0+DNGs29z9JUJFGsI7dvFYiL5
kyXjfOp7ekLX6Bfqgr3BsMJWyyxztuWh02D8SZYF/n86ynuFuSFRJNo3Fgt6BmAHy1ZGE8RQmVe+
bFZZjQjuRxO5QWyPygRdcsEAO/ZoaZjQC+w5GgBLJvsR1v+ds7e2+JC8yxPWM2QB9WZMAOo/opqE
LwNhEhiRylgzws/x6/Po787skKmMYsCoq1crqBIOQmk8Qeew8EKeRIXidwuVFb6Rm/j8mjAbu65V
eF8LW0pUmfcL/bl11ep/z7/0ggzXf8Qd43x12C+7rjE644pvl2cPkNIqp5M+EPXu6EmYLjMRW7Z0
vMrCdIt74xCWptoh1b1K++082QXFbT2WeFzGpVshGE43tZzxrXfhCkuPQ0bHU/ttSyRMhk7BPBgG
b796aZsAqC69GQO11GEuRm/PE96m7lzWS3yv0TtAUXuhJo1Q3Be7iGdMgpY98NuhuizWET3nUMH2
EJvY3mAW9HgnHXlDas5DUeaT4iuWfj1y07A3ZkXLBRKc+Tt4qn1u3e/MR5ZihgXFrgDZxHUyAGhe
Jv1xraUIKOVPFEnc+kuDnpb7e7mZ5AodI5TZLNSuKRLmwjcgRXQ2A0il/Qc8B1D3EnH1Ec2sdMEH
CMdbfcSA6os0Ydo0uUsTuInmkq95cww38SZZwxGbVwSy5SBoELLm2DZgZfmx0W5Iuldie4SDqc3W
+FwRwvNYP5X0LcL2z9IdPI2Ou+2LUlHX9X47AIeUD95CABFK/ZRY2dqXHUTMX/NatcatvM21qrOZ
Ro6HLn7Rcw0xrdW43n06MFqFdiU2B/0pU3dJb/xtUX3AzcMt9N/91Us2cHMVny2qjbyCugVH6Zb1
ujnlgzH9PPs2smxkT8/ruZJ/nDHVlXT09GqsUyI6mVcw39G8yGXNcBuF00oBYwaZ2HYt5IU9zGri
OxHuMdrbsXc7BCS2Rbx0VX66g0Oqp4IsltD8yg/VrNjND0dPuM/ok8M0z4NIYodtu1B98N5e/wjT
85S4GKqo6okyJJm/o4TkEzKrg2mTBe/2E7qPv8EiSkdGP9na2herI3vwvvcdinUJFx1fxak2ICUn
jpCORb7iNPDFmCes1GiCMUIl8gbX0nj9tCbLg3zu7T/fSM+Nh583VeUxSHEjrabBOOpjuIvOGwwW
zaOo8c8Lk5x3wQVSAjQHkceMe7wzK2qGNjCHRenVj0HGHFcxF609Az7RdAJASduBwqgW/1KyCz2D
APn9ckzgigm3FMNpClANDuS2XFe7g/fn9xJm/8BOo7BdgsukBL4VSlH6VtXN2hPogPPGvo6Va3a9
KTYqYipApbaEPs8/CdAZ6BEtitmRWn1wPulaibuBfRZvkfuRpYlASPfSK0natBK0CZ+YVf+RX8xN
IExYWryrcjg9IgIbhFpqe+0gY5GmAHIgbxkatsLcJT9LOpxcYDvcRimu5OGldl7nQxW+RadCVuaS
rSBovqgi9hYnURgAwDz7R/IfibU2o1qRWF3LS8+esw5CfxOuLWYCLK5b5ixdbL+vWshL75xWl3T7
APM/dusTCIGZIgG5LacAO1FPKuSVhgOlVSNkuklKmQioREG1SNouZ60HWE51k15b/BQC+gE33jpL
45sHBGtSA4SkUZ3NiW0opl+80BNCvJmcnn84egBZsfpQqLTtIYz/xrHMdc6DEpNY8Qcf1zU9eB28
4QxlMQfXoWc6QAvAdQgMfmOGFOGjdRKa30DuitE8oLNUXojnz6DAJUpG1zch818pXcUORmUKlXfm
JwNuGoGVf3c95rI3WjjaXmNday4U+vQdi2D7aUaaUcL0EJLeCPfIuHY3lVSiUXDy2QnMOQZJa3/E
au7kDyZy+n6EOwGbHUFnfFdx/QXm12VUAHnU8k2ywIoQlQe4/QegK8wzNR1VNNh1FSzWEL9R973n
h7h3WIiQRaSCT7LSVybs2Oa/wzVXZ8jYxQGX63fV7HfrkqjF/I34Nlaa3DndkMvebfVel5bH5Uuf
utKOAPRkqM+1i+MvyHsDGxGQxNzuHHf6Y1I/c56bcuRBqFogzF1Ubhxy9N3Veg2iKyutjJGEcURI
L2O46SJ8CfgB1dKZsYthC01rB9Dhsn/0jL1j/F/2e7AEyV/OOpte2YXIAdznmB2N83nYEkxrRZhU
sZeYo3sjSkF4Kiq9np++uDNPmMLLRcLLZkku8NLHxCbMReafyiexKEx5hUI9K2IOcioztx2ZfTMg
HVT0y8c43+kIZrKIzBvouFZN/ebDtOTUYKjluiljrM0yMdMpyPIOwCTFuW1HJtygIUK2U+oPjwYZ
qXuW2YqIJZDOvADC4/lUs/TyyQvhbaN57lfPfPKjhYiQoQomoVp77HOYA3baLO7/uTVdJ0buLLh3
25kqz1sZILs8ZzjEj30PROXsq/nsGkiFU+IRyA9COKQJU7RawjxNa+KMcnsDx6AWUAxETiH4R9Ed
GmbH2ze3eKiq4D4e4YMuIwXo3uUmXr/nU7YNmjwGZw9X7pKCJMtdXQrS+usXTNOQvgCu9/V7zucc
oVthMWCSKEhy8m4RjRL3vz1rqO71Qgew0nf4CbV95b9NCwB1aWjHpp6bsXusnoYorzxZWlMROKUG
dzZewAoVRxDjg8AuYKHiYCWHTlpFaRNFsSUsCFYbYK2bwgbHuWOia5xijpY6/76/W+TNI/d1WCLU
0PIyK7E5kQMJJgfX3y3zOQJSzWdu+RJY8VIa154lxP67UvTIsR01VvL/9nVHfxCJaiqqF+gFQd49
55CVAL2TwgnzwTZQTfzw2BIvTH8EXM/pH3jQVcMj0H+NQodYrwlCGYh4TKxNpLyCszZpCU1Ypqyp
Zono0u1WKUjn8ZHts7etu3wIzdYhjpSZ/aNujV6tfnzytJzzjzfSE/wn7zKJxl/yDNO+NG3Heylu
u6KWU0QNHfPPF+S7vCk/SJg54UkTWikBGyNQ3+5T0WuP6OVRiaUFv2LAMfiosRJj8TPwAExtuWlM
U/WtaIl0SynXexquv4G+n99WOyQy7+5T0GxWDAKvLJ2CNPIun8grTzNz2OowVmnkN847wDE5ARdO
7phb8DneDSoRFE4NAR9pW+1kEUzA1Rqb08RchCiWZbsEGyGqzzO7Yj23Q4wpX/WTZWwoheW5rzRR
0b+/wJrFE+Y4mjmS3LDCoLYQDfq82YuqqDcKxKCNsfBlwhvXwmSLJkOkxeIdCn/zyd6iodOBV805
NInCo/xk2TaeS9CwSJco1FlUhfDWOQ3rBgJBuUMsxQq/VpRPpUxp0EyUEqtb8fUHNRjeXGK1/z13
DX65Wzsx93GTe/lA203urghDpczjJNJsLj9D/ewsm/H+hCwl93opwSH6jVUxY/hjRB6WfRqkneZ9
5FY+d9WYPgJtmgInzHJGYqGDTxzaQu4yp5q/OEKpvXjT0k0Gwkvc5RNo6Hg+AD6l0Kv7WVAHhfGx
WDa7CQzaNfoxAifOaekYBF3/nophNBctiW3C14NghK0qHwqvJ2c4Xh4txUNdPmEh1iNSFDvYXkyc
Gz4HxeCm1vmObgKqGFHfX2dhz/X8DC+fdLUbZnstamqESVmfAESBgihDDQSSKhQCvHnuNXZAQFBy
FLg6eH/JctZBP3yR3o30mHh9iALtZ5Fw4ljlVacnBbymcmYaw22QUnN1B6HxFnAdM/dxRdMvXybd
CBObk+azbIiCq345QnyikktL2X/CYT+qEAIPG4OpVi7S37+PSJUlJ0HtozfIOyKecNTAKIxi2a+b
AZc6HbB67M4tebwE6czNtiUINbadrg0E+Z9KDw3ivbU5xgRgUGweOqj3CL8OU9yii5ZjQoWB9rFb
YxYY4MdOF0+c4QE0e9qYLcbmZ1to4rOgnoZpyfcN984rTjU6VUU2lZRZyjrNni2AVU9QWzVJlKM0
dYMaidNQQBIzWHDF8BP+fT9Bb8Rq3EaxmhFSC+SKIBgollzf6vPd/cTdHOHohjXHh70oCBPdYTEV
7UCTn1qIOZDPD95si90vsEHrATUVZWhVKs0WS28uCK6HYn6YOJJBG/z3kE62uiBL6xO3sTv39rWf
iZ2wDVKYBbrbd2NJiqwWr+y4PJ0cPAMY/9Pfd5uzgVsk0SvQ2CCAMb5fs68RgvzhxShU25C074xH
+ddujqW7mezTljhNdFDGcQPOmAie6kHZdkNZNT6Xi1wOHrEAeUh6N2ZdqcLixTxHVOj7Oh9Wk3Cm
xCfePxFQjPHYAlb5/vf72sa525Gp1FXhXlNoOsalr+CEqQ2/jsY+t2d9arJ4QZN/iD75rd8pWtCx
vig7Bppr31wrUbk3sm4XGwzjZQt/HdFwdQqvxIplQSK2RoQ5yLa1zNjFf8GTHPV+5Yw2QIK4ahAI
lb2ET/pkvCNz3uPKqxeeenT7WthBVO+0ScAtqODBarPWipB7hRTciy0LLl1vWUyC9ImTuuQfOKKh
R3Njn6UAw+v0mjkfyIgg9kwPpLwmV/ZglLuiMOZnPuJ02LIe0aupgwAqU5Lu240J74/VjmqRQVeL
s0x9HaVDAH+aMTDR2EASmXsLTR7NbCMo3Q6b5PpwXDKGdm+g9YFcJ1w1gqLy6XTjigD3PkgE445i
hfG/VnSIJYGkM1X0SxQdxVtr5ZMTWAcQE/ro4n5XLaZCQ4I5xs0M3nZanyAod8Rr8IV2JbvWSQTj
LOukyQrV045AQPJhH4nyp2aGgs0/N+4pvxaGfvv7lmixk4fmBwKwleQnAyxr1e7NgSYZfi51+5XA
TtZlCTU8mzq19w/x9efimK2FxXPWc5ULIfQPei9SFF5alnlCmAeaDmhnBLQQPh94wg60Qlc/IQLC
CK+w6Olcryq7bvLqA/sw6EV2B7xtUd1uLCbObwSiGWWHDI1ykwrEZbuMIReHlEVdSGFXHNRLkJPJ
Nb84eTfeEUcEBLJBh7PUVSOXxexCOafObIYdH5xglbzG0U5INgnMFOMJGZKUP+rB0eFJC7E7+n2O
hwe5vnqVbW1WsG67TLs1EwxM+N92sJv2zq4KA34WA+KB95CAcXzeutTe4+MPMOsrfy6TxC0O1Uae
bDSa1yk+kZnfgkYFhytx30ApYsaELNdDF+NuI2tcjv/b6QtWfXQ1e8aoJ4yDNWcOGPN8W9tKLqJp
S4eMTwpb84WTNUi5rExYy+ngU+WCetgSxJrqlCDFOSw8AAqrHtw5q9O48oyrendCznX70EqCfnnT
VHBI7wYT/wXW9zfJKvUtwqcAy0Q0F8Af7C/BfviPxsVtU9gLuARHPQTwT45Z2mJCBnTu/RlYuOum
IvndDHCiof7cB53RpGX21/cKNR6SPhSr/Xynhd1mY9H5yYRA5vCM0hdBXTDbf4Pk3Iku11Sya2PL
DAkmBoatJY+HKdQYcFvw+UQ6PluZohnuuQhxbrc8OaBJSCqM4zcCyR9ncMLG3EpFPGm9kyEfS0me
YwF42VDlEsEIOz8r+HSkB0My4opf3xpMjhJgwunUATIt3jY4ezOIzfv571YIU1iRdtPfwpqxYudB
ifLdh+7pi5U44sNQBD3AJaFv0i2zBKQXAac4552rOCcwIuUzmPmoM2zcpbROdeNnSEI2K8DWAbL/
9zmnK7foeoL8KceuCwdxCDwVlxbyz2FcDu4En4HGXo3FuWAO+7wrnwZkTCCEa5RSIXirOhX9OsW5
c6o5bajLC7c3zjobeqJyBjHe70/TuSyclEwejfssnGz85nG97GdtGafq2N3EKDZMCjMRVT5VUI10
l/VBPdUHKSIhMjaYrZR0wGQz10b+Hfp5xs1iSLkGod5kJCHd8dTjz3HZRb4Lnk46y7dOu++xm8mR
WPeleZXj7yNdBWsySHK0u3ruVMP93cIE8JcSxmX9z5iJV7buEXHiQXfjt/4ikqIN7zZUL1KA9Oh5
dJ/ScWMt7o0GSVZO94pjppEPyW/IYZruw2x1l5MqVSK2e/f4tTndKtH/t6hou8zSHHQNjre/piWX
mZ2g1BzBtga918KmXz4sAVQ0d05FUj2nUAa2vnTS/BHX5T7PbtFtM7wM+Y5+NBLv17AXTHWMTSRt
8IFk1dbWdnx3ZqcMY5lRVPt1B33Jy3Iks2VrtsdmS1xR57mI+sLIyjLqOWTkoucO4hU2pYX4QLZs
YCOBLXeDtuyBLj8NSnVLkLQtUdBFyOf6vkjxAlJQNniGv+F6IB9TsGM4GK4HKHRMstJyh8f65x/U
D2hgIjakBQ2JX8Q1MLsgtVlBzWyDFOEjHEWiVr0iAjIPo7L/nT03fbJYRwtkwQIqbDyKenzeO0KS
DSmc70A8dHY+em0SjMHDOCmVULlt/HMOGwcC9kSZOosSDvQpKHxpo6RRSCi3Ul8q+sIqTH3JQVMv
1ah0QQQORSc2E75vrCwzYRHEcAWRjkda62QVYW205qlfkKjxO5Y6+Skvc7a6x3zdkHwRgEiQNieB
q8KmTSPZBA6CGFBMSl4aJfbCq7+LtLbVBtGL9G93yViZdNcxS0HVkzXrwDclFwgWrNmpxD8ZcMb8
ly4GgiKJSL+FSNC8fAnAPLaQnLVAPsCaTfokHlgBI/IbPkonE291WZEGwr4HjBHSMpDnjUbjqw/B
zRDNiE1JR/iZA0nwI9rsqKIJOxtU18S8P6eAvY+BU6FAIYeD69ujopGMJ6D9e3kbnSkaAgOQempw
okKlMB+913gRQDBIjXwt3lEKcSA8dgts7e+HUrAcjnYb4NKeCcz0F66n3+MlYhOf9a/f3Hkbx10s
e+VZv3NOs9KrtVcfVcF8ZAJTg7xaAxBsjFuWZI/A61TkEPnAiwfTXZ6wnOJQx19GYuwwr3xdqaxI
frEH43t4CHQ3jJTwykRlqUArZRnN9/YkOhmQqQnWhGLbUteH6yOV7jSc3eelmg1XQ2Cfl5NLpWUh
6jkRhKex2LlIVw/A3xYPWxe9iNTmGvmk04WvqM2TWDx8xKgCCqnNg47Q59hmVQ7e7O6PAxjdcDYg
WLXswkGxhILY+2riV0ggCbX4gsIdiMi13Q2Zd5bnMDm5WNCmF0hWbski6NMxLkjApfmbEFvNa/Qs
kpT6DGrDzUs40uNUuXIWM9s6l+aMF8Dm+fnexaTNQMlfLKjqxQIHF8MNkjOHbYyyJfG9ni7rQ3oU
j+bjSRwRaKorvsUHLj6AK0RaBFnYgMLAUAt430ZmeOX8iiuLa7Am6ZIsuyx+sfK0NLaiyIjRDPVj
FHCd6pOkcRTBYeMTSlOOOIgwNZvJt2bC0ln8Bu1xD8tS9I0d7VhyQDK9trFvnF2ZtL9FqOtLGNzy
acX2Dk5Ss90ZdccE9dM0dxnI7FpwOqmGFdNYr5qRr3nojGdVTTm7rBJiUgUcpSGZ99x5nJmAMbjO
w3hMg4WIKZqkOHxaPvrtVg0FJNgkJo0bLWE+wkn2GjSioWLYFvLQXX7Km9U2rqYE8n5V7M1D7Obx
ocSqV68aFiauG1Ja/8lHKYz14F5N5f9Yn/izK1UBBzpuPYB9VFLkK2+bPoK6L+UmQQKz5dAG7Vx6
f6Z2Q+jLp3N3gWvuaA/QOuv6EgiZafNRI7ouduiaaznLGy8de8rd1uGHUfOR2tyC1NyrtsGlERu6
hZvYCkTUKkg7dVB7ROR6Bqe/T7liCFUoJlCxi4FhB96jT6+xGVaFKdLS5O6KCc6OHhf7t0trKiAI
42dwKczDf6oUPunc13Ju8Skz7vLLFdi+O+hNR7GTb9k8H7SVx63/wmLe6m9ILWA4CH3tknOv7zxM
EyX96iJhH1Bq72Cj6dWemuA+zBKJ3Yo809wUr7c56ucP1O9XgFB7hfKUQR4sQDxq1X9fbSRqCKFG
1ANH1MFB2tVoEjQfuddwMHSPdbps+25YdWkCeaHUjf2VwIDggeQ7QiUZBAhRa8hxEdm/2cJrAhEH
SdMESuIDlkMSZQLsg5rNUucDASeWoRfedBdYotvmLrwkQz3tl/Xvi1lg0t/M7XBkMv2jNZ0L8L1a
vn6GIO42jylK39b4iyqoNKmivVv4wQptWMLMBpWd7x+g5o9i42JryM4IQgxsv/0zoVq2LRDjMzcY
upVB6zNKS/qwbZJCSrWynzm8sY9Gjr0SSWbtCRV3sg7zzKYWfBqMBX+Tz08wtIAlQHtCmtkxSRdt
0Qa3ao94fHtENpG7fcpGyUKMhPo9JjKWePPyR9qa9mudmz+T6jnHzLorQMs9nyw38TS2jT5eATVE
ahyLvA/tfomHFrORW68m4qlI27nJ/VU3o96O6ej4nnvh5IEzNW6PR6aBMfnoaD/swDgpGQs2Q5+G
ZLqWbMW8xdfdxMDj3SPToX2m41+Nd2tEPI+rH93Sfvaqpj5ZPY4uILH9ZncSuYl1HmU9p7EPB6GZ
q3v8txSM5UhlhkikiLaFp9D3Nvrdhxo+fxKIeb5MMuqo2/MX9eRyhY6NHlM2kUPhofd0OyNzNkaE
lOAzAexJnpQR4lNrFG6N4eaq2Vnq47Fvov7PKBHIeVQ9zzzpBiccNYvfHEWWLW8oHheUWbPagz2o
rIUKtWDp8z316JjelS8S60kRrKDcOX2qQPON0yzRqwUtHfQhoECvGvbJiV2rYjEWUTyYXt0AQWaj
fA7GgyMxxEYc46x9GgH5SX5QpuoNNw6swczquRbp6APmoiGBwx2dvSoVDg5aT5vWgBReydE+4Obp
PREUWI2ANFlINmZZbpKFKjDB6HJfsHDosoKwLb3oaBqnsow+Y+ctTLB7A8otESv+/x+z+l+Verid
ls+I+upXVeQjlgzijbMF+pgLCgVk1j64dwAXcmA+cyN848L+H5fFOJLiGbb9xjATcVQldOPC2pGt
sWpNm1mBDV121k2J0qqqoXs22mJlIc478R8QKO8KyzhGBkUVEnSomzisc1MQDL+VmKFy+EozOvNo
gY9GCE4N668zVAMtSGJl56EMknm+n+qkTJaT0dW2gCTDmxb4ODSwQYGMWIVnfbsc4EDAke6sGz2T
+g55kEKTekVuG4cOiQs/18ti4CUHKWlfMCAl/8VXizip/c8ien+iBZfpCDsuvFDCq9+ABRWhmSPt
rhMT8mU2iz1KIojO18VrMbhPLdO9qsSlxloDQqoT9lvNn0KPFlVaaOZO4kxtcXhyIKv+07zHCgDm
l1K3/naZMseh/Bc5Ckt2/YtwM4gvNdTKUlm6CFNnm9eGA+7SYQ8C2mbgY8XiSving2K/JAnYPlUT
hj6iIQ0ln0Wd3B9bHFbmrPjssE2R0Qg9Zre8Cr/RNT1bp7LZYsnKA0muPRF4skgryjiLxIGp1gPj
LHOQnsRNwTCsYhzFbuxamwQ4S++MBILRrSAc+KHI2UHaw7L4rGFz6zOAdA6HbqRRyBH8LNsyZGIN
SyEc6N5C5Ji0y0Kk/lrpXpDfTYxO3hRJRz0p9yNY8nc74jaCgCPqzlUW9Oj101UZS6/Gs4733QrF
y8jr8y931UdDHhkDUI4CBXIzvTmTeLjtQYiqHU6HSTT/3ccow9R+HnWNR8lKEfFND7ckudHK2FzC
Q1mkW9yCnafSwdB1rAYtCi2/CzfXUkEm2J65+EMPz4jialQVJDOu78n87oXFfmGnh8zdLhorxOua
I19mPo1yCra6o6KI+QULgqunLh3TRENqRxOajowGsz4rvrTtnlX6Aw1/qDkUR6uP2r/BgRNAL2LD
hzuicDYbEIvouRiDeNtD0IaP8uePT7ayEvLcPRaWv+lwXRKNxf1bphEDrFuB/plYX8jRtc3yiP04
cQlB+gLJuMp0s+R6fIHTABBE/li8j8pkL5UIMcuxAfESznbl6zfkdEIWt86dyO/RhiUDdj4mC1zd
O+nVFsND8eZFhyMHeeXEMW4HOORs4kkeAmyK7KdzaG5TbIQ4XztivA/6Cz+2G+4XSZO/y08IcpXk
ORAvEfcqyCTVAW7uarg36hyiNGFb3CEkcK1DjRO5XeENUxfi3S3lkMQbQu+2hHtJGk7BWN5WU2yp
gMyi+NmWB2B+Sl7iWSC19lvEPZzEdyBuUoQ4cvwlNmgMExrMTL+yWWYqYih0mKdkpdNMsLKFtAnq
yhHyWUfnKAynA9K4kodpRRAiZPMIVip0YFolTyoQBlkEKFJUomUKogBGtdXd7zRnf1yffwKmg2UT
OFGzHR0MwzY4deqqLQzrRoDBbM/ciMFEpUuAl3R+K0hZhXML9/6/CutpAsmL9nM9DoFeQekN3okn
zXU9EWutTSjhiXdc9fxilUBfcz6/S73SAUdTm408hFL2oIVMU3aJhN2abV9h4TBviZhCFRksyjww
vDo/dLC0Bv1q4vlIaRKUV3VsxXb9jQRkotH6JdduhCiI4HV5vpHsufVnsVBWah29m9PYOpRAWUQq
+s+IBmAcMpZ8cyQ+Io+bKnwWgdTTzAzz+kn2ny/q5Kvgf5JnrNHgCCJGMYXh+ausN2FsTZyCk15P
3xk2ton8vmZqQyTA7fRjB5UDml3cdvrilpEjLxKiMK5hwooBZFJlvygqoULlL5y9cr8rnNw90ImU
kNu98iPqR0oI+ifBBlKMiMp7QUfp4l6QA+GwFozXWvIvpnd6YqnLAZ6rVte2GKuXR1GIUn4tG7pT
a0/Zk0cJC7ZxN4ii4yQjBLk7dLkiLVUXaMsB5vWkjOrbuod7M2nFjFVhVT7zQUQzFmA3Ey8HNfRe
jnNhDrBs9CIF0WTr9YQqPKXM8BFuS4Txgz45YFFyhGpSHKvprtHBjBf075I7MEu41U2XLsP0H/qZ
95/u3f1nBQJGl/ndq75TCPGIcYctLj/Tz3DaZiRuaa6+rO4G4gklacD5yimH4iQYLqr6pQjMO3Io
HR70eWY80CUvXM7/l71pAqwVmvXvJFmqKHcvR2lx8K5Jy7nw6jJvkrIicllm9XOORj4dHjyh+tQA
WX/ggsOys5EsgkWrQgbd/DH9sur4CtF44O60UGj4Sv3+x/edYKc8XQFc0AHTsbKPSniWOXxTn33H
WaD1odgNmDCwsVHI9w7OcaV65UVeu48GHvhJq/ySc0bZOxEXEN3dwp8zKEsL/PMvE76i7I3BmNGQ
T+XcwYA8eSf9Xuod08xZJ6htWdKHQOxIDXu/fyWbzW8BDdt3AnpADiKTUcUlXYrdPY8M+SprOnoL
tjnxJSFHNceZMrqIiD3FJsReaz68lKzvMyCi/993QW/7f/UFlZUCW1Ep/AmkfV1jMVT3nJpPovtW
M2TxPkTBx0DLXilmo2Sy64c07ZrJinI/Sncs7t+4fr7ZJ6sdfnVoudaFxv1Wt94B8wNl5zYr9TGh
Yk8/ynDWxeGoREaE1EF6vUC5LMV7m7cYvQAiO+6e6tArw1uUUzU+CT72xk1+uOFn6/Vre1VkyPoQ
X5rpoDLfohFGbdaQvNbMgQxDgk75KkgPp7k7meomoPUSyst0JYx2+vx7MzqrRuO2uVt690MpmD/C
1FmokJ0Yfo//AY01VJRQ4Z3+QXshkDXfuxNwlcdvVFKFiTZKGq4nw5IMkrer+uz3yW2vygXOilW4
M/j5JUYPqCrSUf1XjzoihgTM/unWlE7ao3F3UmJV7aaGThL2pmhwqp/mHH0ncj3QWYtj0X5AlLgz
BUnUtmwHqRwNELxvopCzFlda001fbTCNvmfrizQW4Eg/mVbC50sZTuXdFZW+eW3cdHjqiowRMMBp
j20ZL++kHm1dXPRCy0V8fSYVvf9yqo0x5ZQDfPJfB+Qg8VX0Q43Zae5OxtdeKAVW+gj6aIii55+X
qAngEb8C2jrH1MpXZiCToufiR0kNRzz0xtOTW3wXNKssA42RrNYTDVlV0frbGdU1e2YkXK5OgfsR
0a6852c+VKt7V9vLG7DivPJCMH8uHV1dx/DHUyS8g3QUFsvDMQTLS7xreCxjAppy3cfpPtunXBYj
hkZhykaTE01Cex9SxrGD0L9H/uP+sjlgucHCqdnRneEv91iCQkiVFtKCkH85sPA0/L4A2mGd6HVS
96vmDfgYtUUX7anI9j2OtSwMsZgT5foWaDGgIiGr72iiL4f3ASTVYtPQAWVdpkRRYTE7195sv8Zy
unMaTJYQ/EB/wgq3pgPheNr0dENJXYbNgtaWekbyJaW8uJ4yJKxXBNs7fHapyUHdFuywhobh8u4z
ywK/ODxce1ejzPoofiIeDS6dc2okEuJauoED+HGgD0+ml2c3IJDn5dOa8voO8IN1nLV+z+2hLedc
8rgT1Ep4rqQNrlcU+ve6UD1qyJjOV2hhYWoMPaQUvyclbrCVxFOzmYMFoiBzWerqTreAStVrqVhv
VcGO50bpA/Nkw+yR5vBm6TgMjdALLcqwyH+J58qCZ6/9PZi2PRROZC+GicWY06kQXQSaYDcN2Zzi
o9iG8+A/B4WoBdIg97fDMX7x8ju9XC/xJONu6PjDqGod/jVAQEZMaj/B17waGTW7zil2Y6ovujOQ
Q6+hCvegDVMJdjg9TXOaN8kbQH2HC/n8i9TgrfKCn8GF1nhBTlSR/Fw4anE/NpKMReUQfEwA+qjv
DSEK3g+l2FMfurXiG0HKS/bwp4uETIfI+HDU+J3nkyNAcrrKSz/3ylKXPiCcJm3QJofpGwoBuojM
5HlYgaHa6Fjp3dNlu+jt8lBtQ9G1VEQAdStibu9X95H65nTb7j1T6W+qQLHyGM9/I+bAYjMM/Nu8
yY0dmHNAtxQGWtmma+ZtPUWRhlaPuvURY7hnBD+BWQeN3f8pXtF264DU39DGJK9XpRIqZZRxjPpM
F2ujJ/UfI+9wBe84OxfKGod2EpjzQTrVJ92aQHS5qamkKqoSqK01up7YFy+otmoEGDK+Wr6DgZQn
Y98dwrgb9g13GvH+/GAwVhf1cKI4p/S9gRNpBBfZ/NADgbB/j8qgeCdosXCZNZ5u+lfseSy7Z3Sc
6LnM8V7mGFYByQwSqfpAyHyPUP5sE92Y28aGk/bwppatN3WrxGdbjv1nxmsATs/M5yRqqb3wpa/8
6eBzZh7Xlgr5Ie/hGd6tefhL4fnKSvax1xlMPVtOYQnQ4O32l5ggMxE9dBwaGid/q6kvUEIoGd2r
Mv+FRYdKdheE1chQPvGg3t7aa+QFe2bVkZgIsurni65QiKPvbCMTMAFi4+8G7IWgGTCTq1uNq3nG
RRG4h6+9LAaiIvsDdQp558lS//fNid/cWBMyONeVhJbpnnXnLMyunFFDMq7oZQaJrlBWGjScF0pu
+H+jYzrJaiOnHglyHBGc8NhbEVM4Iv/E97RCG3PupxX61EWMxjP4ygnlcDYmj66V4pZifECA4A1d
i4C+9IcNxneoUdCSHy+24+3pAqxX6jFX0kcqRYJ76YZaIvpQYHjcZ5TKWK+NxZd/5tP4PgFldmta
lZfGXlQoE7me5PP1ceka4tfpRmUIo7rfFt0QZ9VRGr1UHlrTq15geVsvM54cw1oik0tt4EH9Iq1p
SnpwEsEFbzDXNFSCYMm7mtStAlkxmPQgXi/kcRPqQQJ27bNzlwgVizDwMFvEEbly+I+121wiS83A
7nx38ANyqBmgnucNv72dITB8h+LujyNfdtwqkUBYjjCbntG4E16W0QiOkxgfXQTNK9wDcKvxDIVS
EIqPsnfM2XR9MB32HmPJEfL3dGkuh0UGWy/0hS6nIx51SXa7dt9ncKl5elrYTRjyjj4+2mmtIPx+
yf8N3JRSWIgmQOhX4GjrClV5CS38vF6HcWqv/IWWvWHbsNrqY+KJYNeXBFwC0LQmCNai1aynRp6u
feDLFCeGVxOAXDEztw2TiBPYeVJsQ3QlQco6dpxkQMPyRm/9ksflPTDalxtxcEwA5yXIXyyiLwX3
7h0//LlvnP4nmNZwkMY/XRE7MnzMTGdv6PCDftnxEtUw7+Z8UIDbWcFrJ+7e8toSAtQXSDcJOSI8
Dy0kQ3w7xtQeTe+jQctEcuwID81OhFsDgV1GREWKGeCpWHWqWyNIlvyn1q0IrM4OspsDl6KtIf/W
deZ60jXZ66zUPWCOuq/3IaITZX/qZxt3iSMd/XPQ9qEH3n/3Xn1tHlV+5MBKw6E7O/McpKT2JHfG
2Lm9ncMEw3VBwNuQ4x5hCMhdsZIngxxJDaJG1fCtKBXNq7jYddA2IrU412Br6IBcBEVKxWqo0x9E
sWJ1DFtb6uamQeROq3y8IAPe5ijrsEzHI2FROZqqHjCwkKQ4Dfcw0XPe6eWY87F8opwWahqJRVek
Hac+kOnOuZSiyMFGGFCqNnXU2Gq2qm5hRDDcXozkyVvKd6FM4HaOI8MDSFuI4BgUmPdADd39JOgs
ALMb19XORS2wQ1PpJmEBuj3cLtL9d3TfU1ypjKKUVOwlCirSgT1lB9Fywi2f6cc7jzsUx9jSY+LF
PnaKJB9c8SIS1CUVCxGvsdxOAYJeTNczruLBsk1P98xlJC/LSxq20WT1a1SS03JPsKQfcT1PUKov
svFW5oWlgpG8x08oz3QrmUKuGrcuyV/XYifSYaXLTUShNu58tOfkyW2x4b92CdoUhhZJ4hdNHGQg
6GqPXeb8Y66zGi1GorbVbkI8sUby7gn6SrAX5DIkkjYoSiHIwmJWft/+za0S22rU7quWbbpynL4K
58bcqsxDEMzEOQhG7cCcAfq2xHHu/vru/xQjPqns+IxJ4Yag6JlTx/NihibQy3x42IM+jG0OIiB6
Us/HSEC6SdAniG52mhWAuUsvg35ForrJcGTLhgomvtM/BOeJ9euKEbPmEydZFRVEWiwg2q1CxplU
keICzaTRnfG3YJ6o2zf0cUhz2Ona/eUOlfBc/iDIS6x1rl5ynAVUyXvsquoOiYpXXzSPAMt5mdRf
TsEiw8nJ7GvoPRvr7rvC/d6JEXE+SlX+ZmpfVqKWNvDrl9Fei7xWFCRHILkYFumwu79N50n0QXfM
YvR8ugEKu83t1lVsNtMErCgknzfKmzkjrvOnajJENvk6iL7hwMxHhbx/OXWFO/yd7EZh0u/htbH/
rqm1tYLrQkKPTcB4nJCSRpDeSi0Zo018YhOdwJnZ09osvHX2k1irRW76pQXoJrimfB/TTOOC+TnM
tgWZxdEPryEWnN0WPMfGJ5eKFg4Gc1kG3srmbO577VKQHX5u7otvJ6Vj9rpDbBQA7DZk0lUz
`protect end_protected
