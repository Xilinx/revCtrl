`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
apc1CnSO4+T0xR0ZUVP5/vK9/mRe3Wp2sJuEVvW+2+GND5pkgI2H49+dTGseqdM9G6e2afbk47ka
VrCpABwiaQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f7SlyLV9nmSvqRCBSsFRHrw6gkFzGs6bg4K3McbZAPIQ/zJdiVM7Dc/Gm/Tv8lk3S3sKHgY2uf69
hQBxDm0KM11s10OJwjja3SYnKnNJZAaq6y7/9Afyyy/P7atSjGgcABH8nEyeQ+XCcIqEpYLT6o7h
EUvF9D/ONa7s0EJE6Mk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oM1ZoDb6aiWXXQy6a2GvOT4KOtd47FrXz/3g81u3MVP56zMR5GtLt7ryWgUn+rVf3VK7jzLiGQsM
w4MmQlFxy3MpvOd70DRf4eFrAO8knFaX8NelViGofkaaEwXl8NifzOmN4azyihdDxkszukClLEIK
SYUCXslR7lplKdOPsIjpOD1/Cpik+qHl5enPARNjAN5Tl6UL6EjV1qD68MYLhbUMb5jro2lgTNge
g+GoLkProEdkEeWXwqYRXcxxNpUVviYnaaqWEcPZAoei0kmDtX2PAvaYRs8sMIpXALSIz0GuW8DF
HyKVPa1XbYk6yBXiFqhGxRAcVAbrOv7Kgm6Pxg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RSIm5aPJ/tfv7oec9MY/ZsD+wv1orhtjRU7aQhwCXt118o42kowoxl328s/sJBbyFzCw0dXsDB21
6VgE9zya0iIr5nIEPfRr/74p+jO1YStFYlh+BHOPG4dIS/d2dZaZgN6dLkUeJV5xsJJx9zFq22iE
2CO8O9i5JJYI3lJQWyg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pnSKQgBiazZRJltZY1V4Fc87kxUj0Hht5jEcGbZ5u9DDWvUhOczLNM9CZh6kMav9h6qXXCSedMp5
IF7vxEfVCpdGdEBSwAZwRG5IPGkYiVUbYcuSJ48MlSe+d6AT5qAVDKhchsA9elGf+EDj3DMPaWs6
mNU4zA0B6EZ+0JAZlxeIr23YHgR0/H78dxw6+SVqdPMF8mcA05Pwu2ikVpqrc+RnkdtMILOREiOm
nWZexvCDDpkEv46NGoi+HeJTwqnDR2aWNi6ji+ox0k8C4qrjayUh8fW6DbZM+eykbm1KRK3XlUOV
zsKGT7nN0aVQAbFnRiaPXwpIdWN0hnIE0CdonQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3632)
`protect data_block
YvC8HV0/yF7t/AN7gkDr33trPB4ZC+dQ3hszQFD+s+3U8m7T6mHyVuvuuG+2f0pUwqx+lcmPbhqq
lEQDDXLA/F+uCJoPLT41crq+y/9caDcpP2t0NUOrLtpqoKVmO9CgDKc4N6XtxZbV84wBURAZLQWp
qumjNgUNnfyJKDcjf4D/1Si0Um/flZQpzSvP9HDppnzAdhASPBG1QWXRPi/pMjzx/ijcPWzkFX9I
V8KHQNQloJLI0VvZqLC4wWfTNzs4FWq9pdcMSz3i/RkvJwtaWwrKuBlF+18ulQhsdCfl00v1k3ip
clm/gUP6tL+gp7VUL5HtqN8A4Z04nmqihjkRoku4MbZuM2pZOth1CduNHb/lb0e3pjPJGrjw3Rxt
mTnKlmnT1pYSuek0B6o7gi2ZeTTPhPSj6fdwQqAe0NDjk+IhVqkusB74CfzV7bw0rNJJzv3Wlnlw
lainbdE7Xm/Rf7CHM92ZA+0Et4FF9w2TDUCXFfAOZl3blMWLfXlr3hXYTa2DjTTtl/TTwEYUyDDd
diRmdNw+Icpd5lSUCmduddEbxlSjBY0xMfTmro1VYNc558zJUsAz9CV/pKX3tKzCucXk4YnsEAHU
rhtxKGCjz+uDHXBVHojIU5Z2UJxAe+kRWL2pTXQQDDbL0vNewcDlsPvNlfd1BEVlHnNI1SJWG2TH
g1YwgQfxyf004N+SoC0pgmnas07Uvnz0XfPa9mPvomxUqDagnWcm8HxwDCKcZqPjKGqjhQoF2oKs
XfzxYu6jOU05ffxOGtDD6gjv3a7isB7oyBH8AWbIktuyGeNuGgsME/VtcLBjIpTvvMwqmsmwjWpK
rP0a8hIN+YT3Eo24NAUzZm58KVAunadKofJ0oCEtE4l4mRx7wRCeBsGyRC8DhHEjCfRQDErgrQiF
XVV8vYtbl96D4oT6V0VF97nH6etx7/BI3z/eqAAug4t2JtqmQUb8ukrIC7LrHhBARpkn1ZLxT/AG
0exCYgWgaFwzUcGiUUOlI1nfypJmAbsbGwg1y4drU0uUFcsfKitq4ktrStU2MNxlut47DyLI7Nl3
Zfdp8L7BfuQj/aMlAmeMTr5Nx2U6K8KvtZKOhK/yW5JKEpPQIfykk32ebxW/PJHLjIWgWL4AkQoz
BbKv2RbVoDMbRvr9tQDWON/q3VhndgKFM3CMMPZte0JC1T04TG2k4SZq/tv3FsDCN0NuX5xQPx0P
LzUuMgKJdleIw+dxA975GQkpqIq9WAKlLqYtu1tflqTyMpdzgvPekrw+kdlsgx53pl0AMh/2F8Xg
OSaKAVzCd+azMXLBmtHgZYBxGZwiBbX5ev/CCUb7nsdtEv1BJLc/Dd0a3tClVbxhl1pOp5eY19OJ
IAPLGjJWjQpOLkA+lhhDe1gwkf6IwJd1Je4ZxN31Es8t+oUQXCFT4IwKU2JwB17etOkr2dXZnDEB
mt2ZhmzaxDaTekImOUr2YAnz4W1H4Bb5yyp2TNr71yPu3QK5/Wn7JrWcEKP5nJFsq20W+S+oUDg7
a7l9CoGtRmBW73Pz3Ol0KNNmVDfguMxupHdII5FdM7DSmAT/9yJoxk6wFJsSgJ0wKGuXOvcClqh9
gxvYWvOtqMEKmWGLr1/9hEwRdQTkLFojhExoyhv76xu+fzEIszpnQisErRj1BAwhE/kTlczA/s/5
ZD4SdUKPs2jCc2mKg3bsyd+F7u1/FCcB2eZORGZeeqr6E5asMC3y2BiGxxddQUcdYSwU6PAft4Cr
s1prg4LpKtHcqJY2U3Ww6S0gHvQbTAB/1ROLHmWKHq7N786KPUV7F8Rk7OkR6Tdhh5la8Re3sWZc
rv7edjXqR7tlsXaiJoYbN+Qw2s6yJxjpt/bEEHQ2epM78mm1VgdZn0rYq8V+7d1Unb0m1hiPYdwt
A07wM/u+JzU4v24NHzN9qvyRCiLHH4LzB0/aHYmX/wfG6dLxoRIZR7VA2w8ZuGN656ANfVrbb2el
iZUiwHr29T1oayYm+3gJNIJBLxoFBULHYUQBybGmG7Kv6XHF8q+Y21r1yqnIAsdzWrGdxJ6ruryQ
5MONkEsQPNDiNTHKSQbqZK2l8HjUOzXN5H+z0FjLLhWT/borKNrRQUtXRwr40E6VVjZNuSYu/dvk
bLAgM4PfQds7Wk4joM/K2axL6F3qxbAgV2bheZBMeZT3m1EoNOvHIRpZvjK2MM+PNrFhiUnVTc1M
P4UYoBGW1HFVDHW/qft73C32zj2DsxAOZ9cIeNaZYYn1n3xSUIFHjpLFTFmVYDSBg3OIdhzW1ZPV
mddOJfS4SxJadHt9RPH4YJ9k0tdtxpil/1h+lpsyphBVzgR11ONHdH2FGNc0dl/qKdgFx8tcLHQV
VAU3whv6WPUK4YS3drxSHVEjyZIEWdnFWNYKF2CL6txN+kDgttJFi6wKBaENO6Bh6Tz0bmWxrKLy
A3vAXfEDbBd82oN28Tb8QArbJaQgz6gQDgnpwGyZCBNHe1OL6/pyLYpcntWhgfDxsbdu+KgYgKNB
ZEPtjpF/N+zL6hHGXg17wPF4RsNQfzVNxMtfbJxGzoqiGB/OidL4FUkbks3hak0j6oks3mE3ac2e
OlyDjdwpnhXOJ79N3pDbPH3fu+W6ojTrZhA1Vg7ULuZRoCd9N9xVlRNOcEEf2UWifQXcG0pVdEF0
j8EmCKsyfeJa0qrIq/b9B1ZhZ3wCwB48ljcga6tB5JXT77+lZhfVpNCFMeCIzjfznHUC5JTCjq2K
Lq66WVcqLIwjvHJDbth065iIrOElRVW41wpGh+yGmhKL+vsJYFHeg3AJF9LEi4SVPIU2+IBfKDDc
RkYLtnfqif3RRWxNgFybKhbqmAWqb4CPl/bjrXrYmYeqkTk/2Hk9dx/ccqnth3Vng5m21cwBq2KI
x0aMl36LFZKBRf7t1ZO/5QnmfekKxtR8Aax4LIZuL6bCJSRRQjMtGAyVxD1b80rIVHG746EOnPh3
lIaoCkh9RtC8Yl0UfjwIZBRvEtzXMHLF/BA4n7tM+ZlGjpImQp2Zc3WO8C9278SKAXv0mPmKTtAh
DNw1Jy9cx1hD6CjHuj8F8sEEc7sxGLX+L9fsBGP/KvLcR8FYkKJ2IBuPnbKZltxw7FsDRDX9Wre0
jF9/xNVhJEdJG9EJ/aLzd7Oj0kBzIX00yrTA68bHJp0ukjacSvJjiyFRbwcoBIdFanPMHPjXhzvM
ZwM5hIjg90umCLykk/iBnbK/9Un1dFGixIVVvTizeTEBrPbCIO5LQ3cE598iopIWiaTWatjI2hCF
G/NnQIdQxXr5YGDh2nkx1F7xVn3ulRu3UQU0mqRKs8b6eRd2y97CR4WvKhhRlzdpHTJUkrW1/YzR
wjBCcW3F2sMsIayW3r9b46S0RvaUPHZhnNoHkXQMsDX+ojxpnRb5filVc6TTmibUwiIe5wAHNyvJ
snhzr6v0DbPMcT5zOdBCtvuc09DONH29KhW3VsnzGvMIga8eh0RF8ym4DvWAUexlGYY4GFXgzDp/
8fMqz8pXrerx98k4cV8LiKsgRNG1Wg4r+HMW7iL/+tRNeOwDGlWVeqWAn+tn+alvUc6qo7LF90ow
rFY6g+19RcZQ0yJ43QdJAwC8ONFDARlLIrWT5wxgJLwY5vF/6TuloItNK9cM3ZpgFfWC49TuL2Uc
S8utq9/dyoKLeWIA3VbW1hA8kbH8zJ6wB4PbCHNMoRloGUlJAqi6FJtGpGrKMbvVo2ruQldEvDWv
tNvktVzeOBHOEfHxDFXNeQsGg181xYIlqSzrCJWvGwiIqhro5XC42UNE5ypAN31cqyikn7sT2qjZ
nAcMUJY9OfWVu2OcpG6uRy3rUxufNWnCV4W2Fv7D/UDhPoHXA5ekPdHP7tgnuReeRW0yuPehd+zi
Lj8RiDUGl0ocryvO8zNAEba0ja26K1XaMT9AReufOYLOkDP58XQ7R8UgI1cNavDHd/5ngPxrbm0H
fOewlmY6+2xRjZAwGwpBN+07emyxDIUW5jLyLNF1bkWxPXRlQhVfgYEbyi0SWRPnd2bEg1zXCEAM
TZzvzriXszHvJJfwceqW3RiDMdiEqjMIdsBXEDq6ulm793v6e0hkkIjAEnc23T7gd1aMSKlk96am
ys2SjXa7ZbeGui+6eB7k5D+cpZVYMIOCO1yhsklWp824ap8dquXZ+Noc2BA5MTyL+LuP1bGCpLHq
2VeF1LWb4o2MsvWtv+DeddlNj7lCe4pJqKifCUDP447TxzKs/2Qg6Xb4YZ8RPa6ABg4V9O+5BdH9
5oS2uugwYH1+HrasNu6DdpZJ8gTtuKzk4ZRn0ZsWtn2oqjQU9t7fWX3yJ8NH6dxg/6q4xjkdhzZ6
IXj9LH5O9/BrpDa7i8qwmj7wwrHMv5ykn0auxWthbG/DGamzSuIU2h9Hza9JZi9kcPBYmh6BTma9
GGx8sQ/l7Q698TxVyckzNDeBQRHIdV01PjWsaPS8PUsj66WEjM8J2l2HdSjC1YjxXLnmpwwNYyKP
4YL+rDImGTrBkfxY/H/hGjQy2Nfr4Saz8u9YP0wWd9GdT9/+wF8S2D1ZnMUsXC8RjGHmc2Q7vNkP
jCiCZVIhzoPHHS7lpDy6psXSg0wx/58MqkueZMHWCEBRvo34Ha8WmWrrc2N+rq9KMkKUijpX/9+L
4FjjwH8R2L6QBoqDFwyQw+rKzqCegVh7ellVS4TK1SSWkMDNiBaLVKNq5m3oLoNnXWaPdCoyFbD1
zY+91PbBXYjatSJanoHYIA8tPfryId7JtNGWqBkMuCKBxCCH728bxrUKEHRGB8PlYQI4VtlpTv8g
XZxQg2dYE93vSZVZpYT6ZvoBp27dDbS+Q+FOsqStF0s5+Il6G/YR9a4=
`protect end_protected
