`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px1erjyAP5O1QEY833iN+y9tZYCuy0pKG3XmEYRG4aOjgKV0uILLywAtgjb7K3DoVYUk+/qnYfpV
vmHxs8x0Zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1xUCzmV7ZIl5zGtPY07q3GXS92D0V0L10iIKk4ICSVMa0f8QHb+9R7N/nHAivy4EwnererRsZS+
Gjr9OwycLccWp/MR/2C1cGBs4uQcwOikro0ahCWMNof4qYVs+/ZM//8eTlsyVc0/9jR3v/vU6n5V
56v6TbwBw+Dfk/gqPas=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
habWysI1xS5TiJ6nfV4vEPL28kHCMXAs2Plm6sySPGwAMBgz5YGB3HQN+Vg4KFqH1UufCaDTLKo7
FJS0A2AJr8s8X31uqhFZM6Ud1Bhi7kduXtqVn7dyfpwR02JoNZ1yOJbN8VnHJ0JOHV/95TPnCD7K
tvKLu4HX2TU5nJvLxQQnGP5Hc3V54ybtGbW46SBRoY5U/Wop14wpvYS3hxGvee0WLquCRPcu7APJ
oiesbFkw7/aKUajVmAYfea3OJlhcXBFH4phZnzrahymSft+x8bzJ4AV2qjBCRiYbO76v3p57sHjk
x+YtSI/1TadF4YRHxnXv2rWGZ9Pmy8klOoXiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKv8c4Z1oQBru5wEsnL5NdDHIUoDkkU0V9jPweOqGUTqNZ37D4ZA1qE1rIwJk/Oo+4mpEHpoM9by
6x9QIqwdTWPyZJsuz1iQSFFG6H8OW1JxTkEuthYR7LpTg4NhTod26Irn/GHnVUTJmPP0gwIbeXua
XRTl8OMj3t0DKzwJEgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g1I7jc1tzmZDNp1aT/anUyMmIt+m3UwQ/3zLP/86625+2I6+SquMu9sTa8CtmiEetYPQZkanu7HD
hcCVknw8She52J7s+pbszGfxB7edYekr5pmTpIlrNPRCpkazz7s3QHCw63Euy4TbAbCDKvwC6qty
wvzuUuu5aQ6DCWJzHzqisQ76EUL8BhLYthDlNZPKSEUY7fGPrTP5af4yKZl68WyAapf3nZXUKe9h
SMfOfSvKl4fK60PPedYuLJqFpeYlIX+YMm3rqiaQjvJ0NwuimdPQbvQcJkQC1tb/p/5jpdc0MPZ8
fXTYqAmAFS8mkerbScmgZcfoV7z/hV9r65+J0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28672)
`protect data_block
hTX64IeLyHzfa3tJyS5DfnCGfI2VwUPJSF+Bc54ckFz+NzeZiFF5uvu2m2AY0CEoZr9/D7bPdcu8
4biucjkDKHi8OyYeR166g+neUnV7whLBBXiY/iPs5yF8+UExlLozbtdlZKRc63elUUwidCFznsCi
FdwKRRKr85hDOFynYtU89w95pH0jPcwZSkunj3hUU8bdMwHPOtgnPVUYUZ7mLWifjnUFLzrR2Sbc
icLuThSX412OqL+phUflb74Hd0pnuzPmWj+out3tDrAj0sdqTwTzXD5oRVJeLnYCYOVIyasV3O54
E6vcTED8jnLy51OwyF1fYBzoxRvViXsllO8OESfN5vY3Ta2NOKK6/xm5CFP7lJRqd12LmcQ2IUvc
uBkaFqfpfMC/V/DSi/3n5At2bzTy8ZJY+z4v0QiHDT+KgHKg/RJYo3YdSGpTZu6/8HTcdqdCViOE
4F7965ySL15G4p1Fxf1gwOHOiSpSXJXVRMzK33b8odGKa04ahBYDBlr6bBEG012J41+N6CkmwJ1n
p9VAf4I0hEWibNDkZVBuuSDulng9VVq54NH5U3606YATtfa4lMXTt5EJbrh/knYu2fow8ojzC1Dy
u2ntZthkm3pDvTdmRhJiKgTro8WF3n2e+pigbd6+m91EPzt8R3+qOMshZd81SYgYGsqtNiaygRjE
z9WyG+/TzwjBNSuPINf0qYAGod4GQf79Id8+/Zfk5r1DoNjMmD+q0mmuOayGBYo/Ln0qoj52IvKE
swzlkxSHzLYXJiQxrucFsSGQceO4ocKiUZXEixpiDIYZPIg33xCavh9Mve1730qGwJM26ZPE3DYp
lwkLhDDYqarKpfqbc99ucoBh9a4TRplKaZ1JSi2lGzZCVM6VQNvU0NcXdQN4MNQF1w9LfT92PTw7
ACT91MqkpM04eg/5EC3QM8sxX6jwc628JDnUoJeI+AmhDvXwroTCnd2lwWaOaroUZBBZmSTrf2Il
myN7I+2Ujv6BMGy35KAvsWIqRDF47iO7AF9gsbeQ5DOmDj2eLCDhLwKhhSzO+NHGYBaeSlt7EUx4
2FdPBaAczX13hCUctC6SzfGSFPEbrc3Mio40pNzsVVByvH1+xnuZypJzaeTThA0smIoCCCgBnNfa
H5FFD9HLxxpvhYJ033VOnMEtVjZmCKc1ZCsU9xehlg2Rt+xeq2fevBj8L0xQFaqPM2AJp+ORso1A
X4zTyHnAjQhScO8cU6/e8UvAse33skwOXYv4Kmc/RxFSNonl762K7xLzd0cjBtQPeSEOzUBel/EB
oGBbUh2YGdeGydWyKz82In+z769fgtfoU5gm0tyr4nVw2jyW6zPohrPZLSr7sWraMjl4OGiE/y4/
HDN/htHxttcldXi4XDpVE1Gokkiz3dywf2d+Uu/2oN2wnK4nyeLKIPaIPbYa7PC4H0DNsJtV1aUZ
GwbC6EWOier45nHAX4BpmH3PT5WgVeepNlOprxQ8zlWccvE7Azr5CZr6ZCoZzpcKu9RHhJmgtXDS
11LJ6JbyN315UW8yqMCQlMD4dCgLRNADwH7InkQKm2/4CMonkCVW/vO2G37N4fNSxdGR5j1rDHai
ZWjn5HP7cltq0tlv4wty8Pbs1OPbjkHCrawWDUn3gsLBocp/GgsktXdK52PsQyHpiasnU+8KL+D6
wBQb97J2mIHOTcqTICPyJ5pXH9Sfs7OLj6u6k3j0wqaMTqoLFA+BNzfk+MZQNoOAIESzvSDeHcIf
9Z+vHqpDUgGf302nTlv48cmw6UhyTe6XkxTr7d/3hxwBnwIkYQsqgfkRQBntYLc/KrVMv9bOL8Ap
sp8TwgvkcLO6P/Y8MQ0LesOqkMi/6l0faEbK2lsae8hpnueBCBjjoRwSXyS4xxNC8hxiwu5FprS2
mgzPaC9Zt1AvRUY5HmhAcpRCj9LiI9E/mf4s6vWWvPhUHVxdg5L2uoEvGiKN6qtHRdaZ/Rofx5f5
EHrsSYlMSTcIH5IWm5HuKoTONvrn06OoPUslCgZJh2txyrXBSwENLx7jR2pjMxuQmr1wVa+GM3R7
opfo6MlXO2H8FP/OkAw76QsiA5qCrgfrRLgrOHmEHcc5VUNr1W7NoG5L+KV/H7Q0o4iL8iBHSdbl
n8k8TsAEtbQC6Ie8EIl8kcFISnyeJoX7OeTJOrGkoWgtrSTc2EQuxe0uIoid/Xp2+6JUu6nA4067
YsSSkwcE1jCget37YYYgWw6naz8Q0gR/gdXOwpo62ucDmmeexQ5wsapDJKxK2TAJEKtCLsj+nxWk
hnyStDBA/EneUxGZNDHSC1Wp5MpoJI9M18erYqJJQ/Nh/c6NgrwU0eFGmJXo9fDThCioxjmVm3WW
bgPsdTkniwtrwapeo0FXW9vUhwJyU39VrzHT7vdEs94e1MtVP0UZV17haiZwjcz6Nvx8hkg/4sw0
8tTAxT+jFvGEUIDT9r2xASitu7H+yhoV+Uj5uCf7cDxQeQxE5q4Dixfs3TbLGRm5uOT9FRW9obSm
ynzaTH3p+EoHpl8D2OFzZykKn8JxGOKqIeMAI4VfEAkaOxdvwsIq5RJjMg7Lf2jgMMCwh07sVACF
v4YB2UWKJOr6+v/YZ2/CQJuybKbo6dQ7XmwVpLGFRVytspGH8NpOznGSydTZ8XZ+p037Nl4gK+y2
0DvFk1S8K6SJlymDBTR721sdJkfKhTYzPPi4cUUwimA+OWv3drqfzi97Md6p+UG6bRJ6a7WzuYTq
AbruUZBkk2tUFKdcvd2KijUqQbbDoaP2Fyit1mT+wEew5SiZ2j378oo60/gkZzd3A0J4lBZitZp+
F3+KKRnCnxP76NLFbTMs/24e+yB1N6WFunczw50Ptt9G47wl1RUxQhrwnoa8tBt/D7cQpY+O8zKA
7KEgPfa+b0Duv73oGDPV2q5fTvhLMVVou+n/fdavJCDCMunM+5IhJ+mQ7peO83MytzTPqlW2O7f4
vgYe7AtZ4nNxFwBBru+0KMehFTMbGY0rFP/Yfo0pLcmihGSBtSBOS703PYiaQ+8KkadLcuGymYqG
mgWT98k+zZX7gTAYonysO8Be/gD7i9AWlUQ7NchsUCjGQ0pQH4oFAO5cAioqY7OCDPuLwTNEU3Qh
hl6JiW7q4zgt3gLjotlGcwHxrfDAFiQdIylN277oahUm2veJScVV31JtoxV72urt8+wME/3UWFPr
eSZ22vFgG2f5CmoMaTdhmv+hDVZa2fapta+hZgvzGB6WKmdf7/hKAxKtx0hXa6ET/CFGdmjAD4ev
xvBBMKYKQ+sDCtEhMESUHWk0GyTSW+X/VFM2zkTyxW4GOoYfosz5BK6/9HfZoZPNPhmfR2dGqWaj
IBRsyiRt5Wh7e+tsYWFgdAgM+PpvEPzo/GKA8Z/aMRPYz2wCK+PqeSBvCfdVfuv5W1OZUL7VvEWv
s6+3WGXGusguSLFufqsZXvoEuzUThtrZVj2MTEI8gILtSaTncZs5YjrL48dSxuZ6OAXV8TRj3cnz
tUYhTTQoKCVbdNtyJexXUyzEXFmIMTtnDVYiVU4xghI+R+uSEfAGPvem4EZcs3qsnVpROtuQvd/O
FXawpHnavFGJszjXfbTpqhih6Msy2VKHVvrZGWqOfExYZT0FRaKu53QTtHgvLXOGJ6Kw3qzjoLEZ
p0nckAmJ/Ik6omfuQNKGc8JH3n1odNNvYFacNOeQ8h/3E8OHAfH7yfTZ6wBmnLU4R1DhFVCPoPqa
RviAmQYsCvrHThKG7vapstHQ/9yKb0XR3z7Fsd5juHrNpYCsYTubrOd1MpK5pMdz2SQBwYazSoub
o03I3L74X9FuhMQAfcTEszpO9s0qn20JqHAsT+3N59kPE15fuLbkSf6wdGRkd87nYn39yFf8RXay
/qYQs0WtHvLv7Pd2N70qO+bCTn4qdRc91ZB/N0LyBSaBic1QhoWHLJEfl8Mz5w2Ly/7Cb2pJNBei
bdiKdaV+VHId4VvW/+IHs2xdwNLmD36ajSYy0lZkwNQkio4mwlYxIdlcgBVvfUNXuAhqKiirfwvT
7kxwM6mZl7mgmGZfyorjSkYaU600WGeSUKNiHMhWv/AD6h/IaNTH7Pn4ZjMK7+dL55hcf2EsUGgM
EyJna8e+mmPLF83COJHXFu0Qz6BkmZS81mP6I+4UmzN55IHuTCvsSgZUw/7E0uw1W8CRuEE3vkaf
56gcBT+nVlHntwvPXt+9E7Va30AgFxeYxXu+aS3UGYbJdL5dPNfYbD7UuTCVZ9cF/SaInghyAWuC
OXKVWfr59H4nkDu0Tsu8jJyDtbsPKpA+Mdlrgj6WAc2/umJaGp4UDljekX/88ziDvVaq9s3Vw4oU
zGaMiAre7kuHR0jmzncESln32aeC3YWhKcE3qx5fRQBA7glF+/OlBugK7z5bIWBGw886YuqhkXNi
gSSfLWHXz043AzXwIhKFa3JFHdo7fsfB2LtmgqDyvzTaQuXhm2W5wa4k344i+UFYuZdDCJDWq/qb
gZFGiZNzmpeAondpVvbLBF74HfKg5EZ29ECkDRLnniG6koJELlk9zHpMQwVhbjFk5Ems8cqiZxGr
g+JuzqB2xpSBvBqFXJhdD5i0Qifw0agx6t5e/DNJIlvbUz2DC8ZJO+RnAkazhbLHAjj89mi/Lvmd
ip3uxF/OLRa/OaINFpnSUNcAq8zUbJ/DIcuZeQ91L1G9O9PmZS16CJITnSQr52gMT5NlOAq1gcaV
r9R4N7trIyGdADDG79XVkCd0HKy9GZ/qh1NPTZrnCtKfcT+OgHqu3UVFEDNGj+qnEts0cEv08Edh
MS4rUHjIWvD/AAs9rWJB3oYdwzJvvm/J70IEfznErHtrFYFBuiJmtrBPRDhS84Zb51Bt+Fcim6D2
5GmkrctraBPOTLGAOrOG2LBS5b0gP7WREFzmWzbC+36PLuFZU/USrjrP8OSaZslI7RubymLb5bIR
J2LkeATZ12ZEb0gHMvKEckhQxeVwE4shTjp5MgMRTNmB3IcVRMPLY92q/tJs1LzaXprcfzjd1X3s
aVQOo9zVzdB14BVhWp+iNK5kujfxHU3n+pmYcw0MF64K//DCsOcZ202oSu2VSwi1eCJysnePdvzk
iWmp6vRuBbDBc0xgTyvNiCx5SbCEKkbvq4GA7/Q8Hlk/WMR9YXEbNezww+ElNPtk8AbR5BhUa3bH
ne28sKXM4Sk4pXzsqeKQyEcEhSaAIEpW7GpfiZ/Pblx7VR/ryS7s2dLkgoCUDMBpe6f/L6YrGDg4
dkcxnWB/oSqPZN1FOQod91EohuDSaX0+iJXXcHWYfyMeVPhclwY4u5PZI8PyqMnrBgiurLawzKkk
zWwgoFwHlZxqN1GU8oyVQSpf/tTWnuEDsM2h6LIsJNTpmIKOXy3LzsA99GDQSigwt0016/PjCHw5
pEoMBEyrIpVtMiRlIfCpiHyICxFz83U04aA08UljUL1WpUsT+EQKVOtmSfGkF8cj5ccAv+mORFBw
Wkeas6rkDyZyKv7ci0y20p3hwXrjNFf9mvmTVT6NvmG+5vK8y/8DTsKW3tRTVS2NJ91xuH8tzYNj
8tzQl5jVFPqVes2hjep7ZE1lBm7G0N7NsCYL56MQ5echMU74tasoSXbsCGY5QBtR922mW4lW6DbN
0NzmMPhZGjPMZsZd34d+XolnXQvOQKyAHCij8dddKYqpsbVJ4QbbIX74dEcUJ31fnKSWRxJOSaDr
2uDoUdDwLwzQ/A/tGLP3/17KW8P8bsln4/VdnMlfCK7Frz/+vl80JDxwUp7EwcaAEC/DbZ9onf2s
BinZ9juxBkIChsr9wRtfoNoqhTZ9b9A1WPoGxArNtFGXx1gBm2pvA8F9b+OCE4BKgt4yYFvXGdif
yNdGiJdY3YRvSm0z68jtaAAAHeSMR66WvRiI9PQyUrV8pmkHJwr6AXQf9Z6FcOollJTEQ5Oldayt
PJnWXrJ36ORT+/UmG76bjcqtWkTMCu/4JdAV9rISYb11IZj+Cr9fDBSYMxi2Cdf7Iky0RabXZJwK
7V8FuLDa1sYXjYlMsPGpaY7lbE4WZmMaJx6R1bbHmlR2SagcIl0Zb+7+Hnwz1bwA0CQt4WqvbwYX
i/1M1/LjL3j400ht0q8/EeOK/4WruSpe/BKnQs3yukfbUWDoyQpQ0pFtLxwIZ9yyFWoF7T3/JKhu
hiPGjbMj6TU/SWEu0MRIJ5VGJEsHeZSk4WX7vtlGycNuz6asl5/6eKDoRsl4/lRUCcHy7u8FfQ1U
kDcrL47+uv4ioDFLDHKNi6VIffV9Yxyi9Mbo0Zfyd6ooqBWio4ZYoeQHD+snjtMRUzoOZ3Q7hkRE
wQeDZbqqlR6Wecrok5PCXZUNxwkVi3iHmevnNaEQSP7fVvCfvgWmMYHOmCS5QDxVJq86vYz9yugY
LtHhZpETSBJThpQ60gMyOjU0cuAmaqfs5KxCbPNL5JtPTKchE4QWc/ByfZM8xnmzERtmgsR5ED76
htSvQI2ByRMaxvcT1eX2W9JleoQjbKerGrY7HfxK0BmZuBYVwCpTjFMKnQpfUg3XvQhHgELfohEt
F0Nr5fzjz4Az3WR+8qtCVTN1tmAZHP0QzwwouMgsB9LOksJQ+YegmRqetZuKMRFLyFXGo6y9WfW9
q5UsZXQd4jt1/7clLRMyqGBmMJTWNTAgsXNIslFE1SmEyVtbkJrbD4JcjSmRHcvQj2FfA/SIQgmp
93DOqnLQFxY4etqyOEmchygM5YaCkH3V68fihEnQfbqZz2Q3yXXpUCosr5qDNfaB0wV9jtRJz7Ny
mpe5FRLAXW6+/e8b+e6sugHPtaP2lu49del9NsmgkEzjlf4bdPA9F+JNnNo8P815dzQguaDlEph/
lVaUfPOf5+lm696cbaJuVOHnfm5Au8fxs4AGXre0COsii3O/pQNFQ+Gvw2k8Uxz40oLqEkUj50+/
IeZFjgC4ND021Excnm1vm7HYWUFC2q+WS0VQs+UuwRXzjfE9lLgAwZDiM05QfSW9DQ7ih+2LHCpL
QsX9JUp88VZH4U8RVCwNuRnOolot2QzcJScPRBX3cNMNe9CrUB3TXDxrHcRV3diTFptbqtK7qQkW
QkqVJ6V3xlLnFT4derpOz/tZw2421mzOonLbVEqewZ6+1vSZ/l8rEZyW8I4vaw+zDtIKD/mF9tDI
bDn6WneEpChR4QeeV/6OyjByoY4kXF7Wd+QYtCmC4PJyC/n1rQZ9VgHBeflkioA/S4E+t9Afwh/z
E2Qcw97u8GsjvV8m4cy9992DgMkkX/EBJ2Z6fitxegM6J/YUkRpCiHB0uyaOM/vFlJFt3nxMQ1rv
mg+C2ue8aMk8nw2o1bkb8SOmCuAWBctdF/RpI4EKTR8O5KuMOeB2a40YFG3KdguvKDAL/02FJ4X0
9xwFhZvNFFdoVUZw6mnBHIl79ULf3vlVldGX85oMYChWCI5e1QvSnejHJZgCWlwfrF/077SpDsSy
EQ76Gn9r09EuRJ9zkrod9gsZhk735IUk8FuZySQNRjmv77OqNmGrm4O4L/ECJYjvuo02zgjbdEGb
/ELEridWk0fYCWrD0gzVZH0PAR5FYj12Geh/cOE0AzsPDfHLnvHXLICM/QsrgUL+R4+oSY0y31+s
p/+gMHHrhpDZ4hKVAumN4r/VoQbdD92pNL0+6LR4vppP+WokmU/Ko9xxEBGdAqU81lJiQKMXGgK/
k2G4ju6gDxN2D2SGDIwF1bCLAaV1aFL6TqLHRabDLvMEqO53Wm9ECxuihyg4OzBmRCm0dnag9ON/
pPsmhYpyx3aERB8pY1hO2zwrZM1avSfPG5Ppbo2QSaFBJ9pmgE6MYCZDkxEEOmiyOhEeT267FD9/
XUR5UMe8/mBMMPH3kLwKCQQ5N9zKbwpSTLGv//SFrtTN0oFtgH+1wQ7OSmGZkbwnpKZu2yuGeYof
i9uv0J0M2m2xGYUtxgX4B0Q0u24ZxcxuL1JHqpxVV942r2SEzeuU/jPe4VCKlvxKSyXzNe2skpZV
M6lPI84HqAOGrek+YL+mguUGKM+gfPm6+Mvq6sp2iZ4rjQ9zh3OmsmaAL3UjPcUcbwC2gA+w6Jfm
Sz5ku3XKX5QY97ckLn5E2uwZZA0G2e4g5v0E5jl4Ed5kOBgRkz4aS3rX7cDoOz3q73Vj0gBYc9Dy
Gf+6r38QqBCyV+DWwWIYeHzmBEpOtntgfScO6C1zj7dJCBP4Vw7lsgvKEDJdBNrk9z+a2Sc4JjZP
XxHK3RcWFDUgI2vQIe1MDq080IQY6oCpBRd+2eKpQy7XSDJRdsXpbsEM7lZqlIyFwCG1cekMiSp9
SByOoBcewgKkOszqptlglhRBnWBhnGIMP49En3V2L2Td5Wib96072h2uTkhbzpKAUeEM4HIxXO9T
h0zENtgxGh6ArzRe2cxkATBvukKabbaOLm73SgCxdVvuFwa/a336xkM8Zy3qtWhL2q64PyQQqJOo
8NXzYjOLnqouvAkpkAaO/fCCR9/0hQZuNbKQK+mpPThzor3j8sWU+c44v97aj9cfVPCDZDofkh4d
ZDzbKUb/lem5H0W4a2G5DYCSxG4OCaCnPTXoi3XYXoUf0PzC5K5HDNYVLL9q9qhq34kw4LK2zofu
V+shQq74T1luq5c+WHsmFRixxt/pxlMwIl0lYU/P0W4oRLg7aciB5oMWM4nRXi25VHDUYAQscMOu
1Uy0YAIAclMOGUEIOOZaltMruT8jnccWpVCSTD/2Lmx0F/3i2EAmODHL1DaQLW38ISRPT7EKbKkI
qtId+rlRKMP1JBQF3rxDNKkZmqo0L3T2ybCN1JrEOmEz4d1mn7IIEx52wieiMZdU+e0h7Y8sofg6
Hs3CEThnaqhE8tDdbUJeptF20C37UM9V3HhgaM0cn3/GMBdug88sgWHYTbkF27aD3U+5yxHCobef
rRCSu5z+SC5rGwVJeYgA/ET00nfplqVUgdyEhpnTwI3kmXa+zuToQ9JZK2d/RzmW42CRlk9OAO1L
SPbeyiiVyopy2J2pE3vlRzobrkNbzx+bvyLhRYScU6ZHXqVHBSfv/EbrRfMHouKWhpv8+m9rWhgk
fWbu/WDNAdqOAlOy+DtQ/utrzmOc3poKJAs8XYPMjgmmGeToPab60dJxv1Qt9MfU7p4umunIS0jF
5rvdg47YefeNgDHTmKw+5k24aqR/HOZ5x7mLkvEytpkgHc7fufhSzS0D2iNI3VZdpDXuKIhi0nX+
8BIJA74d61wdc0f1su/61FrWnhsnPFXjc1oz1ko2ypJAcCVp4qM3YKKi+swu4efUcqwwcJLbSTo/
ri3+P06j1Z4rxwPZSITYs8rhsYbVzHX6qrCVt86x3YWCI2FNoQJDHzwCsluIerLw3zAkTauJyagk
ilUXUS+b8z2hJdSDY13yKy9p5TIGPl1COM30mA3YHmPmCPums7CKAnyLJMbVP7OjsAkqKtrLKVDU
lDy7wXgVB7eH2VJ7NLGxOvHgEEbAP2Rg8xR2J8CrOoMb51FpLluy+rT8zBXSITgy2YMXCw3vduqN
6ibe6WSxGwH2mBEJ6iOV7yw3vMR8AhU6b/JiOnLCaAEcBF2DZWsMLRrOeDSua/Ft6ihm8rZoLvKo
W4CR3k+5iy4+vgHtelkJHIvmGfFMPMFIX+d6hjZEi14Y0oZ6+gpsy8IOduB+7xE4crphSa0j37EV
8GhcuSvZhvqNo1KBetbrY+lUQ1n1DzZk5lTp7HZP6T16qgGiVRItVgXi5UGynA2V199v80zgLhV9
hj91/ljk/XgbqIPry84xyZR+TsPu+N13MkfQDL8r1/SpPGTs2wGlKtsWmCIHQyBz3gFlFqnEQVu6
Y+8WSLPbI4GxbN5SDx0BHgsxTjf9jh42VYYOd+UoH9+bQ/+CuQJQlV3DB/gGi/6Nf2hD3trGpeb2
JoIpDsw9HaFUGGhtvE6qtldHjIxo63XxcnsfBwb3QyMNRwNjOb5ZAfeQMlDogTNBQJNlEQ3jyNDe
Am2BXAxxgYcHDPQfgB8Wi9Ps2dY/GMlGXtAmsvYplkTbGHgDFhmQhauWkZre8zoChYm+fvJMB0nu
6OlmWXCdRWbeQP4Z1SluKNvg0zkUHpA/zaOjT/gxZsRBzeHdUOuWyfZCfIv1OBBLfzqGe7R8iw78
z9fYjTgxmikjsC61f67MSF7hGA7opkJ8nMDqBA+7qykBRqtuVlxvCHjV+jvv9t9P5NbfqrCvXP4J
0tYeCzJ7suuKGqF8SnQbAbAe+azqBGNI2MXu+cZ+/0Pid7Hes2nEKZe7g9K55SZ4woEXjWCZt2b0
zzydwhXdw9FyPDUgWjkE+F/xGgmQKTxnvc+F3VzzcABkMcIcqS6EIeQFGZvgLNR0eWmaOPEnyFW8
6maPljefYTkysNdDGKNL4NHq4Fl4SXjvOlglemehjaNij3IbOIomPPuOYmcaIV1zX4rXtuvXexfq
bEAfeegHSpP+i3Fe0Gb9zMJDYXgF5vxTxBLZqG50TnG1J/RqbdxM6LOOQAsBLbFhx/bE/UOG4Jlu
0PfA1MjdfmgYOzkshiziaWZXCDskhIo9g96FiwEPzItQkAzxgR6wJtEYOMp87mgNoTya2ikoJOkY
kqOyp/WxzwkCNP80EDsz7st9T9xXm95N3oM5sdAQmtEQWCtd+PvXvT3treAA75sMvaosDtDh/kp4
ug4TF046y7TmUE/4Z2XyswlMT/ndvxbnCPC5Mpl2+gJK2gwSqM4sLa0+bFtgPI4A8pq85abjQX7b
DPu0RATDugEwHcdO6dYJOQBRVVejz2iFgZu30ZwO8BsCTLAaCAjAducRWhaDY/MLFdYEheKjiaFY
y+3DiCULHd4T9h10ASypGXdGKWvp8b+lVSK3GsXkvadVDt679UA45MijMRoPc2Ps6yO/DW4dXjpP
ld0TGKg8unSR2iJ/x2jv1IU8Dzp0IZA36ziasSjUYpXJMVxK+HW5RF5sz+pMhw2NU9dR8wml3olX
iyxfXRiT/c4AUGpbeEI5UF5QCi9AykBg32uip1TVvnEupmy8tJ6mslhT4Igpx+DweSdbAzpBydcj
TCdOWUYLy2ZEsrs/iBh3YWrDB8TzqRp4ENAO3rSXkAzxjgBzRCmLZK4iTJL6EFCM8mZ7XdmVlThy
aUdgoGIyeSj9uS+FDcTERKyrLPZ35HNO3k33dKRSiqiorZJ7eeQ3NwFTy/IMakw3rlxiMQoERCuW
GD3dUOHnfNDSfGLRn+NHJ2xpWcwR5aY+8EdADVW3xTyBfZaNESN57Q1tOCTMan9WUmFiE09V0MfE
9+V4be3z9sVGnOxH5+Fe4qVvMCTkOAlFk+MfbHhAXoKTvqPsND7Jkx+19JnNv+DeVu70iMvWkdDG
2Vg/vwv0EE/8jWCbQfBYf7DHvKWg2pabqDcKYwyFleneyBnPriSlZuq5TFOQeIKZBw5AgUBYJiMv
mUgnOQMwMXkusk6yNvwdgabjlanHGEnPlVcCM6DUWQOYj8jeRySgSQS1ANbkqSlar53hO8Oek3uK
FS0pxB8d5JO8Fm11skPkeCYjJDXw2GbynHHvvGfIC8+R+M9JPJaFY7MBBR9VVYBzwtKfWl76MD9G
hp4Z4tyaouch2ACzkVeYeu/6xhSIEg324ql32NVihvHoVrzT/vb5rZ3Sz8TLQyuZoVtSuJdBVyoA
NmuI8dWM/6jp7lGtfPUXOgB5Hocbu2Fg7VZyn3mhxuWg+gfPJDzBkX8D71uxNeMlcqdyhKdK0/88
mnvK/QofbRQiQsjqrzNcyF+LzIHG3iBzTOXFsiXu9/GRG9RKioLEMghNOz7puQycvLW6GkWT9xHP
SGpOEzl94O4v9ib2drp0kURaoAghGc83ITjXbLWmPxxil9/YBGEDlSfTbsiAKAp8GkZTxUDygYxt
b044gTiydOn9o/Z55Bdo0QlAYLaRNAYB9Bg64h1NaFdVowMhVU9XsR2XrKq+sYvugeH0GwrREeHh
Ph5W6M2+BHHXN28QLnB+oBQb+Dz9HAF90XjDWbHKoCKuuny2B8xSMgbMn8p1/isZAYZKMc/KN8j0
hrW59yxAcslYgtLiPUEK9cwIwS0KXtytgU8jFSA8eYlpyS33gqpyw+eqlRBJGP1vlOZiDySmLSgj
kLfwNRruJu/Y+PWOG1yX+lr/HfOp3i71QR4mca+VpcBUlCQo33mDNkguu5IGivsWpncpJnILJ/tA
gl+6+zKnK7dmfnqcq6iJ9u40ku2XEKjKYczhHy6Jjv0gq+nTZbMQvAYbVPoy19RnCNc4MLP0LGlA
zKRhwSBFzqs63+I5mzjuAKYd5FEU/oHRtETZV8KeRPMBWZ6qJ0X45Ih4MFXXv27ee3zhGYDPBvnM
Zc5nuRhuG7UeepBTJsuL6ICL/c5Zhiz6UL/oEzUTNOAW47y12KWowvR6wPZrnOb2qPJ4Xd/FFeyP
jcRcXSP9DdkwagbbnzgHMEaJSqZH0W7x147vZd1uMALfaS8iewQOp4hyikzy3xxsz1KLNCiET/ij
CO/k2VVEtLK+ulPqamSRaaupZSew5UsHdVGslZCfWdTGQ9XaGcUVvCOR7aSey5j9UCuo/wWyFKMC
d6ZpamTh76BbXFzy5flsrPdWSmh5u3jB5jVqAiSEg9rVwHmDi4d3Pqh7UUFSAQ9//4xncPlO+hsz
5z4Gmn1Ug3lgTgSveWy7663rbK/QfEkhfsS6sjFff63+gTtt7i1bEAUs4IIkpFt1moR468f+wxGr
C/aPT/zzvsfdaJ7p+e45MpciNZv/B9xFYp6p3usLf8/ZxUT+rHEU9HRILhS9DamD4NrUFyWPCeiA
7BPRgI8rokkCmeqtuqpPAALslzMMiOj5NglkzPM9g3ZerHxKwcE7N/02MSY7uRjHTHQUC0q7Ncy7
Vz2vSUTj5XYYti6Z3U2YMMK54cd7GaEOyAOPfENnnCDGqeA7l/pwoz2M7gQFl+UWzeYxKHgtalWt
OJ3wpqwlIA1DyhOPmuuq2O6OXR3qH7TH4vleYchtE+J6cIYt47Cn3lgzMz7LyNP3N+iKKfW0uLw7
xQ26Wais1M7rwsmmujbNrW1rinc/EMzpOoOUwS2ki5ORnDAW57Zb16iegVZtzwsLpHvzmhvAdKU7
okSj6CAUAsoWvbl1RC72o/NnHv+NUCq6YzKmGI6l96mGcAarzgwIOO3CqNfLYKH6mjDF+12DFQQO
UvmVLo3wP54AeJbhVPkqkbnpdLz7nKxv92zct2aDe1SZMUrmV6UwKSRtOsApY0iQWMT1BJ1uqmct
kPKSJ1kCKffVknw7RX3znAgmxHVhDI0YDe7tP/1PHcv0Yi3EkeUuTdaxap/EZwOe+F/ef1rshCxQ
BDiy4m89SHvU1U7/3N4a0vj+Hadw8wBSDoNSinXe45vHoOKxqNvc0WlKLnJcMUIujAfEVSlzRxha
SibyM4zFQmsb+5uTgrRjFM2xTg6L2Okw+tBvJjulR9EcCMgVHhJSHXc3lzH/XiFqwBnK/cYcMfk6
irzaHuygtHfhATG1Tuj6aCxfRWVpx4gu6PHGoPSQHv77cztA7UEuiRtqBLiDMKb+oORWmqooLNyn
hLqLl+AiBVAn4VZSA7XBqs0jQsa/RbUbArwiMBtujjO43vLV3CCEBxfiN+/xkdK20AazjMOZ+agq
n//O4ejhGGi1XT9RDCjpyPcCrrMmI62MHl4xea7xd/v/ux7QmFfxh4lU2OaNJv4jW/JJRRZCSY7p
Gia/9eqcW5meQIEeaxTfaTq3jcCkKz1qJYoPxWm4e0aYYSWwuhHW5WGMEStRQII6UbbcxINcuxyX
M1vw44XLAKGQeqgcbId0BSr81lcqIwej58IVAKR7+CA24QQD32FGhkQ+E+uI6qk8u9izfMkvuzKC
PfXVxntTjVcrdxn41bhqjdmxL7ocxlZbGF1i1tJiN4geN1+lD7JTAW8VsJbjPypx9iO8S6PZMiYe
/xirZoujStpaX3pETm+ij1p2pRf1QQVxBENOkhYp65u5yI0NSpr0DfCD86BWP/S1DeXeBf1rKTdO
oT3F/XTcOmVP2b/gWP+94uxEGY39/v1wLnD+gTvOf2Oy6mEXzZgyjweMkoY1d/K3kHip6i2wdOjj
tNO2+Z0368jWhG7kyD2fMrZEmK5F39s2E9BJBhnW1sGpujFadAnvVFlfOL4f68KUX9FPJHDUVplq
x8I2QBQwrt8Qhg8iGL5KbcSV60vyF5lbIVnqZyfIKvceSqiHIsD0mkUNNjxC6/D44NEw5ei1Ymqa
TL6VBDZ1k1jhxLMhszKF2hdmFGCXYaXRKpK4pXOrFdBxBKtp4Vf/nJax1adWKp+YunzkqXXdYrfW
LCgxJZkC8U7zeuJmD/vfCDXOOWz+o1LVdO5C/TXPFRYWnxMvoFX00NR2fy1d/df4/iOpxK+Zr2Y+
AP/qXbF9t3O2flv5msmAFsnjzDKBugPkfGndbeGA5CLP66DFGI1f9SoBuKE0Za72JBOse3ak+H8u
LAQ46vgTufJ6LtdhfnrZHLF0F5aA9qasVXBVR49HD4cEcJIcj+3b5fR4VcYSqUSVZUmti9KfYyGk
YfVx+FiORo6CsTey7Tc17dkcK/sOaGBp2OOl4PWxXs9jXEw8fEPy1sqQSuMkeEcUJFPoqfLp3vRv
/iMNI/ly0qp5rN/gAHKWi+BxdoQg7LLzRrfXqcIQPrH0GRR7GFxyiGA5fMMQDBzotOQc9kiaNlBq
MONIg7CGjl362u6iklZvTghVUTtNOJvVsThN/h7hRsZRibR9VR3S3oZcJMgAMpAPA+Woy1sNFbae
Vm2qqJObU4PH/YtevfKxlPDz+pHVlFm6DpACumiY13oPgbLrSY+z4GNNWwNwg3PiRDZl9OiMrCo6
eo90PHMgfO/AADPbv300xv1Y9C85cGGvM7gPxBRdY/GFH0rUpmlWw94UVhGthuKRseCTf6LTrOM8
BjXr1g0yfZLNf1OQ9d030uVrlgPJuncBtbKYJadgrskdM8fdeVKS8be0NvdoVb19bepLIwIuFIUr
rxmKSJBGCvzOwNgArgHwYCCgH0U0+p2KOdtg2Cnbo3MJu+ZuUGhsyY+PBIXqj7Z71F3WyAFXGMn/
7kRRuBtnzppfpP5OEKTeJ9NKUUN9iuZ9ul7ALFyJqmz/mXb3KKFnJbQ1vxwRDPZ9n05cYL36O9NM
NjrIvdJRigZP88pQIXQP8gNMKE62C0hajXFX/xtl7ww/KhBP6oVwX/FUTyATnSbbLtpG9cyrGqtg
/83bvN4sZIip382f91dLrdmpgTH7XSoTuX7Fr6hcWAuPbqw6wwZ7UmFhHcjlPUADgLN7rTvsKzy/
iHSh2PH3CDdIVHC6OxTe4qQHeu2RSz83+WK40hPH7g5bFA1xIURxlg1DHCk3IwOETG/3KY2Z3gmn
fxQ5sPfsfTgQUgd23cib1YHvrmmCUk39hA6wMFH+DaxG5VOT250jpuF1nCr2MOIhDeKU56Jbzlel
OAbI3UiEeDFRkvnXguc/7vSh9i28LfgQxFzyRTnAEvs+nRxiS5m//hvwIOukck+uMR/7VqysLD3J
myVXWu9PgD81k5B3fELUkKzR1p8bww6JD62gCOScnSfu0cAEyJLj3Vjgwpve6Kz4gdTCt88vcN5a
dQij5gZz26pbJDiseAKFoyS4gyooQwNdfGKFUGWyoBaiatGMycOtuNqP5ILfnrG6pG6Klg1oDKG3
RE4lAmu7rZHcPz0ZlBqIv4IYBj8cBY9bMpSQ7ceWmcveyuwY1E3wd8laG1ISdNB+0/ep/nXL9XvC
VsU2YrZXSxl4QpNkifiW9rjJygGTbBCmXxlIyK+rSuEpRbLyS1R6KNPx9WeQyDx6Eo1nMDVaon6Y
K2/LnbwwB4QG2cvNQTO8PpXmK7WqZSjc1j410EOP8R4g31009c4xFt/w9Xwc2rtY+0ATgbf1RZrH
1dtRZRY04lT++44KnDCE85PSTaW+1GdGhIa4dSB/HtX+HNBPyT/tk2ysZIGeQnk+EjI2784dzhVQ
ty+e0t+4UUJespNrtVLaKKs0hoeA3qR6OcZoYh20D3CibMLVsIaXeF0ZT1TMsQAPyHUiNZaum7GM
T1GRpLs2aSvU7Oi4CyTshH3/waXYxyMhPru4+uW6Bg9YJWP2I12sge1DaJSAmGeLx9CGoV6aOh86
9jyfmFB2l4CvdV3bCXzHzUEyVZ0EqjkZcwIuoGpc7S8kyaA8nuyQu7Xy3SouOvSPAJKsh/ngTVef
6AeTaVEgVMZ3wUeX0FU0GjPFy/IA0t4Oz/58Iv1jZJMEzF5MYo0+WftaFxCjWAQWHQ45kQdpMVQx
bem18SYV7eiohFQtsc5I7lfLniShtzZSUEZPJ+6wn2kktGwuC1ZOwjTJ7kSyk+YaUqs0MJIl09h/
d5aTeA2RcDNhzR0lqz43sVpjeZWNMiYmdQmNeZGHktVsLJMFOe3ZxoaUrHiTHIGs6cPDFXyoEsmV
Mmto1VIvoHnss1xGsDggj05zTFE5Q2QSswWXCISTR6CAephWduZo6OCl3vWMbFNkyZwJ+mkW2Kc+
GEO1t6i0roMGUs2FsHSjzc5ukd4J4n828Fll5tjYGWzB76VOrB9PjxE2I1cZvpj8st3ox0RSc442
nA34/JHpL2rWml7u2DcwzG5Hbo2mXgWjLpgHnGJp4zEYsks4ZppCOfB0g0Rasfa/zCNAnde0hV2w
i1LhRswZ9NHGqakT+8jMm0svRtpOvgsgGdsR5Nf14GoiV6b8ycEzzCwYOSCvHM+4kVyUcRwI2cBN
k+QKuGL5e7UKjkOtUf4JdHihB2MSlDGDw+jLa3InU1CJTUG3bYYJ1YkEG66TnOlsymBRYG8hJN4L
TIWgqg+6u8zxebqnk6d96hh54XkmyqDO8t4XRF3oAJ12sf3fSVztb+gIpqOo+5X1mIneTZFy/TF9
QYeP8HkkIl7sG98PFe7ooIXkGZAkxzEDJL15Hpzer6kneimbEsy11vdU88KucKx4iryhBQ+Sw6Az
aXbL5bYlcZM70wxhHslx9JOHmr23fJxPUkrBkmfvTi9Dpw2WoQDRh1K4cEXtX7rbPgVhXhl9Vtk0
O1yhTgfORCp74ygylHQDGkmxAjSKYRnrh4vYj8ERND1lu14jTTfucWl1fInvIRD21dLpFpIZUprj
1AvgPjUFnwI+CoHpAvSoB2NM+SWIotik74U+u/hU99c43OiYP0eWsjyCyq5fDbaCHiWHiF3jyioT
ANhEjOknz7fiZHjeVOSHBsi6N4HQr2YLdg5yDXCTqZnDrgkDi9/Mk0txrmGWEvHGatGQgNhHDLnM
iMOjeISTE3RFst+IU+L6tqwE+YZp/MnTsfE/HJ9aS0HuQ9rXfsuhVmeqiNaGTgs6vFlPDfI1wxpd
sa2bqDWcLKZ5TMbCD/UtgxxLMdlaAgK21lZrOteGfgcoC9FQg+anrN3ZJ0hCXLC8wtXyziEiE/2D
nbnx02CNrgU11KoygbmPUfpBJrHL6AbXA3IXqSokoNSJc8xHkpBglB2Mxsgw73Qy5z74R+IxU6uz
+X3uQGMM8+7+Y9Xhno4J/I744SLg3ZstooLVw7MGRGw75m5Mpymeb8yqGXNRreYoaJ70oyJ0a4T/
WlqT8Yv7GgxKZBv6RN5vBNdh8wVf6pfUgjIGU1PFC9qX7vV+sPjYqVTKjkuVk9/fIHhiVXR+N+40
a4EODY/VKXw/0OR4iE2YQljUv2sDPKrdClQc8v9op+bLTw8IjzPPsG0wlz3blSInr3AAatwDcRYj
WpsAC601dhPoeCJf7t6oGwOFs/iLwUWvntHSRl9Uef5GrwEdX5jiot/RynEvYNXUD1XK7zR8aXEu
x8kMrRrF+UrXXBo9fSsWPUWJl9TNn7bu4Z/I7jWRYQjvfdzFKpGHP7zRR+WyUbLndCmp6GEeGjC7
xwrMGYV1EjI8VFf9cdeYFJPCBs4KSDZJdsjG4ki1EUv0RHv2+6ljmqEf4niwpqZ0OwXX7MuaMSBy
ptmVxTSZuUXFpUXtst7Gz7lupLI4idiElu3Jj6zri9NdyWdgKxJNBG2tewcDcmcmy0Yue5SZveEw
K6T6YDWdIpjmQZgiU1UlTMug5YMSdmhIILWRgeVv5x9RsTfOXXuReg7f52cR0OKJYZxzXG+WtW9o
JUfOt86u5vPQ2hGpgd4lpMMujlEucLpzdYTmU+IKZQPRAlKRBEdEsxxb5bn1UvuKGxNRarezJn+f
ASdD1gkQiFooVb6wb9ZO+txpHsCtmy3ki1U4Pf2IJuAYUtJCLKwpcChOkb/0TKFqQG6w5z579XlB
EPXNz2J9PNZ3pWdAKyPp4gjCEmYVnEzLqvqWlsUkhryYCOgTroYOlsWQgfU3s4VoGpcm9hRBWy0H
j3JNDu+9gdrtKEcXMF4SZmGUU8U/auw75RqDamO0yrw+LbNsy8SXotywD9o4KzdPj7oODqOJfvzB
0RblUoMB4w528UUU9uwXETSsuhfLG8ePBZdI7VcGmCE7CB9ADpjPQ6OtcGlLUSTAuIX4OJ+5b1Ax
egUVlrNgnTKskhOS+Q7uYg3IH0n4tdVToH6aZHnmLklnyiwXSjcmciSpvxCCKpaboOMUFG5of+PW
0sndYQN0c3ELV4o950b6B5ltnsDibsahHRfoJKmZY+bAXVLlgoyiyD4uZCanUGyLJRdR9VfgWKJg
mUQkC1ToR4Cj08F+/OV1qoG11ga5dYmAAH2Sn0BhDVFM62gYXiVk6d2uJ1s2+ypUWykPAUvLC9tP
Q1Q1qqpob9vcucM+JN+NqwWKzjSu1h7Txqvxlq4NUV4zN2qa6uyIN9K62YRWFp+GlNaTExCImwnk
o1f32kOItawO85D5vC6zYfab45YzLtyRRS+VvGfXjaSxsg9fTNO3HXpNFhrTzBoL4RQ4QrFAS7a0
eJsvEom4gSYJaiNMnHxkNQ4qQ8FgW869hOcspVCM5naGl88Chf36Qmhf1R2YyZdTv0GRoW5ONT7e
HitoqPvrjdBHCo2+e0OtbNT6yxrN4rZYQ3LfZx+EAchDnEA9gqbihKRd6XDJ8jF512YL5efXuP+P
cXElT6sny2+v5fXvlnO7rjztaN4yKpyFDtYC5NZzR9ixdIOe1ybxLFv2d4wDn2j5CRXk9DYoTppo
iXYNY1tQtyMXwm85q56mDOinhs7G9nEGjipfhFKKAgZf+3BlDUK3zMWhQvyncbHzFJXPvRQrIPbS
ofX6riKTJQdTnlVzoOvrPJlspDmCzGNE3Ryo8tDrBXLMEsx8O2unT0cLf9RALQEAJ4B4+RhNMMSv
T2wWEyXjMrHZVQfcrMoxJLnuKm1qeFcUN7mEmJDdjVBXt229MFC9gvvTNII/HWb8rLgYLnkY9qIJ
vSVPEPQX1VNL2J2QXgacbq7qtL1g6PUvSbzJGNrMmNX8SHNdZk2Bvd161qCYTh+PYU7jbckNnV0T
qSetl2z+vNVKqPf/BxrA2Iu0UQLoaKlRdmpvi3ffaheMynUrq5rdgJS0o5rFAujm018QXI56xFfz
/KrsQZGECl4vQDqEkvxgZUcVKy8YLQxv06DbMkSeHYeY3gxWkt8wDd7bGAD7yQFJX7M80nqSD8tn
gX8wsLXxxLVlp9EF28sxYgMT5BTAQxV0FvZKh0ahH0cizp4Np1OKhgT4heXt7teO318IuROxv04e
mFkacCZsdP4e3N1Vn3G5cxIfZT9UGwhySeT/UpCxHQMDh526czaNxqIIj1FNa1odBsY6QPCiqiHy
c06J20W4THdyx+SwwuPb8GFd+1M3u9goZsATC1r5O1Zb4WpjUcLL17CN26m+z1c9H5UOHcRS7KjY
uYkNR6l9dByS+jxsRx1206mCCfTo5/Xw5RCv4Juud4blNM0n2X5uI+pv3d9T3IgO7/1rHIMkopQ+
cxAvwUyeSUepn9T13XHx8IgvMm7kMiU5AMR9ZCiXQLiFNkvtCT2J621glCWFJ0mXRqyTtmylP9jB
XQO2JwBCSIjvVDFNclpgU6c0P6s/Ii9jgLCJDRILU3DagvurjC0MvelJ52Evnm4OrqtQjI/uP3ux
4hZngVcM84exp6o3kd7qKw2XqSj58usAgGjVMz8eI4LhCa9KATsaT8MPP4BsNUWdJaBG0kYmR+Fu
VlYIzIwNeOvxzmv56IxJ5JaneKvE9qI3EJUeRXO3CefzTIbEiLDyJkG4BngzdAOgBq34qgS9zJYP
+f4ispRL5z4HiZUIm5QlENAZP938fS84DdTJSsg5iy44Ti87Hsr3cmE/lNKSoszJTfNEijXw4p1Q
oEvYsNt2xjOAtj2ZQJQfkmfBycjZGrPZc3/YTJCfoeBioJmi9z/qhGGpgZuDL8OohoFGdUF5BKvc
YKOUURxYB8ZiTxv2H8MUmOP1WpoMw/ZYkkV6k1QDC1XDRmZyHwsauTtnwI6uFDg5jrMl5w/DB2cQ
D5B9qVaCnFFuwajjqzWNrXYnU1ahoed0HeWNjUhhO1/p45+XNUMaamBINZVI+siV2nX+X96LMAlQ
KttAzI+OLxOlE7RQuj6jVoA9vKx6AQbyvan4nIPXI8c5psu1d8x2FraEkU9uYvKBobZfqIlUaGsR
HOLMD7bRuG11/yfkY7ulvz90x/SilT3C2JX2LFRvX7oxI4fokLb6mu99dBtR5fJChfmnWXq0I5aU
D1C8mQ+mBjiY5aKe2zJCyTserSHlgQy+lbUpdxlufp84UbXDSMs/uwomH4TEpuk3lxAvehF/b7je
U0wZZ1CLl3kYrofgybhcEiovPtC4Fios5T/I4nFDmU2/1HqDXSFaIEVqEiszqe6ylzL7wFQKf9Og
aVcJb7hnVJ8Dzoe72tNfp9Okdf2zs38tGq5PmfHZ39uMhdHDDMBofSZU6VGdyRM2RIiYHGzb6oSH
t1538gYdIpJ41KOiT+gGsfSDArGx5ORBSlv6NISPPqOz2a98DCxefAVp54YuEj25kekNNdtRGYPa
teoTyeW+Z+Zb5WGXryD2DlsMWmTrp5H4jEY7945LilG5eC2khnrFeqR/wCSvTT+1yJubEL/MW64P
3zu9i2Svru+ZCL3CwiGFmWLe9elwGvN4WDlKUB7kq+o+saOY3kBtyGjUSzQcv37c/lEb5l2eT/ui
G9vDNzKKwsqsqsAyzOW+BMOMYzSvs7EJ8mvtaMMbGUGKsSFlpnQZjFxNM4XjJDXSjUVaZlHd1Ikv
rEXWNXSzYEbmgV0a2ywd/SANrijkczDh3wZtuxu39YLvt3Sxp6UsYh9NU8dsZzHM0VY2RtrM1B/x
p+XQW/1nZXy1ijZ7KCNMF6QvlyEqYw6V7rzbdKCJywUmyV99/5rUiyieCetudNXfhgFrZYEmTjjt
Id9YWD4hylI8GzTEVQbLkRdX0tPxrIU5XReElqhiPUx+A5LrlO+epHk/gp+gf+FRwsxd94qthn9w
Cc06KscIvMEZm6QVnwc7zehWZi6Kxw/5tGmf6MRcwe5xub1dsP8Kwj5uOc702ydY/+DjpoVX/21c
k9EkXl32QYOdlIKzHzbZWL6NqN+3EfFUO4HrCrlh7eKWmt/1WorAmWzBEFdl7r5llcvVRahaqqh/
GlukyxFxfJxfMvgN/z05kayNjOxM+voCWP8fyoveAJW6kAIQgMRJrr5TRzYLBcHuLd3sd7jm42Sv
gaudKD1/WMJU7lT5SYLFapXdb3aFbppwtiK50q5zwbgK8K9i52ryKE6COmMJTBvcrqEQPZXKCOXp
g2YchbTW8QprQhYpO9Dcg4blOVyRwAOqXWP3+Ks2iImf9U+va1+gijjPEvv1vrxDdV3pbjWqZ3s8
W/AaQntPsxqRtyhncEmGXhsxsXyocQIEiRMFHz20S3eVgUENLcfwdvFjRhc6KyKBKzW/AdOPW+Zp
y0EdWbB8py9BuSp/lA64MNLAJTS3a9borvSZ7I0bGo08w52McJLUp9HYCKE84U4t8BSQznyQsL3S
eD8E4B4fQW1RNLHIlKyWt56BOdbc/BTsRQZYoCbQvuVgFbxwLfWF2dmBjpn10X+hdRtdbB30a61F
MtwOiv7nzQifdZJrLUbitUbCfz3Zv60eB+rpTrq5202y5VY3+T0X1mH6gsWc9Ycpdu7q90XFZI8A
VSb0PZKfU0Rx2pB4lDWXd+qhVvpZzaQrvGUatdJGymY+/cb/F/YSrmKxy+NZXeNJDDX7RFzTgHsV
IeFRINblAVmAUN2oFdSMQ4T1V8AC38j35tKqaMYau6h44MA4xBfJ+0/8QihGW8n7xs+C90u8FWxM
AfIvYUdCDkKk4qrdwx5StGb6F86Aok53CfYLfDvjy7aq8iyBuP8hDmVrsNunqUpaw/NVNLbO7DLK
peZLUC+ffjgj4yGpbutyiwwmizaoS+ZqsAEtD0hxMjolyiehB9QJsMMV4jCNpaS6LyY8LfGF/ZOo
5V8XKntg+C5Eqo1Ws7N2VyU131jmhsMQ+8qqoteM/chzSM3S0NNm1wIXS4X+GO9urT2wLwXeHbmF
2esBjLUidI6g0eZcQoEb/T0+aTpVS7HwQmyfVF26+CPcoQKxMt7w27xcIO2YeLuIw28pqHYtsKXM
VkqBNNOdHekf8Vvaw4t8W5vFmVlDLyw9yZUU4DKAyQQB4O3j6nlsoXNLQezl/dhWO7hufd49EYGQ
xIPdkaSLXni3UUHGEGlBC+LJjLnBwopHvjQgQXSZuewsQFy/05d0geDwIC52nly/EXLYsTA2SgQ1
TUU4WFhJ9pd+fw3eywip2I87A80f1qJlFJkG31a7WZfiqCixLD1ude6m9Y2VJadqtnvwZLRnHuZz
0eq31e6kxvA5R8+8N3H++woPvvsCqHnNzzM1QWmPx+qEyihPBOhwzwNm/QXDLjCCu5JSy0dzzfT5
BENDP8VKCFDSlXEXaHax1tDsI2RyHeXgYCUC6tewL3DvXlKqoHoCtpCSe0bpdL+X8HQvmNsfxXfR
RlehtzE1QbBs7CbBtDJR0HxJaqQFnVkv8MYJA/cYTgGHqhRX7blGYtxVLC6ZH96iyKm8YYmFjzLe
V+8GQqvqFpEefhKkgL4vBgFsfJ7i9SWNlDEaj5jqLR3g3cm34hNp5+loTt/v6VAgJeLbLpkMjBJD
ib7GP/cwELo+KFVuVmP+5wquJw7uYpbhHRoBdPIq+ZY2PDlJ2w/LZ2mD+gxdlc9OVWDllu0nRWgM
+IGhnFhAtdiGT938EgyxYGposHPNUXzNptyxrQKVGCVsGI1efuiIMIvLJIB9uDgDo4LAq1WRoK3t
2vzHhetG+YuGAL8FpGStK8zxDDMPVcZsHDQyJnPnJ1//WOlzR2vQE6EmZKmaowfhA6P14dP6Bc3l
v35FonQgTIpdjz8mZySj7NoCkuD8FjAgrB/R/L44Y/pfgLImaFbyc98RvnJ3Ezkk8GEjMTI40o+d
nkBVh9i7MSbXpqEL/WW7sc7tfFAqloqSMTRsuCT6bIUqOQtK9JD5Pwk4Kz1F8QD2y7FkP9e5wQpq
JmfgcEm1LrL6ddeuJ+ut3u2ub47j24hzekfux2FkPwU+hNeiV5El5Cu8ykXBUXX3xYiCzW37sB4M
wPcAYLhQd94/hpa6yMcPHQSp3iL6dXNnhFS98UBmklDOXZPVbyZ2usM8m7JsP79ftcA6TSNbuODA
37T8pqEzPrZ5pDlThyY+m/xDgDzD2XmyPTZCde2alziOLihk7Z01pvOq+MkFWAbgq6d8EID79W1V
gEbdmZ4Xkbzx5vfhWj5qfLEwSyaAcQxIezRrQHRQIoKh12kFa6s/M4hUTUVrrz+ThmSDICquMPXx
T84CrCO6c4AHsuFfJZnkyo5i5n09ZdO0X6IBTb4g0Heyjd+WEvsCFVFsWPTQ41/8PS7EAviQp+qf
qU01IaXgrLSOqy8l/OdqSCBHPa/+tpPW33dwYaY9BbRa95/RzbAYEn5soHlt93QdpOxCuYbalCn3
g8gUUeHiYzBBqjft4a4IiKgwvxbyj5mC3/3gbslAAyZoSAxXCCz8J9pwSArCkXtr6ks5yW9uwxWg
1+zn921zavrKwx4FHMfQkYvwpMBxKTzHxKMUK2RMjVBQsssW/MslqPVjiEN7RD749vRBkh+r1R6U
WlP5QadEl4IlLHlKMQX7/BPLsh8Hsxyxn82a8IlFfmMETO01ds2f+A3HO8VEhISshRV9DToIGycQ
a+VSuwkOM5P3FAAI515GGESaxOhQ5UdpaA8LcNDJvDFjepBdOzrti7kHF19/OXVzlFCYtvnRQ2UW
bcgoUJjy9njfh1gngxX2UGfCitMRs8FrAKsEQJWf0gqGdxyiUyqjhDRQBengU0kwuN0KLBQEHy2o
I0jSzxDx0F2tMPMzJCnI725yYKKi2QoIlCxDx/ehA42k3TL+/nBTj+fUPpy51drS6J53HoajsJvA
a8nOEavbfw65zkLzRcTowdnDjsM1YcpBvWUMR10vs3PyArFKAhVYTQMNG3M6GobLz0LSVDCjHGz1
INAslm21resBuQwt7eM7Ax27lAHcQZpgWpkJuohFz+im/1MTDPc54SgEFbOxKRMkZlnwyendLgC1
RZT2Y+Qqw3xIje3dLNDDyc/EoLvAYxN+lbkMPomZYJok5P0hMl4CxFhGDw6FY5AN8V1LyGkfinNE
X7YFWsEPp3sC8m7juK+3jbnzOado04GPcqO17c7wrxL6anW38Bc7Lq2oZWehE22tj1kfpSORELJy
xA8Y2W5Zt+C7g9IDOkdqms4Usuh54y3JFITT5jTk9PvhnxoZxcGAKTNZbJIAFVCGkXGXoOgiI5V9
MLO9JLzpaa4GFx2RfHe7QR+F7rEm9VvRAkG1lHQ9kIf+Q2TAWhO3uKQLeXr2OkuQWsngOOwb7OEY
u4OotxCS8hKiRvpWRVRf4lrhxHMyhQhmDkL6Sun+1xD07py14z83imHY3myQFf977pqiPgj9+arp
XlFnl6d2R2by3mPRSW0S3sc9G0degWGQ5O1dCQyoPZB2Q43AsgzmUkD+flY1rz3afLJzuDxCMdUl
6YpXnXgLudp1j8F/dUPtqbArnlIytxG2qMJpWSmXK+k3bBEZwWe8x2ndejgJu2w9Q4lCNei3YBH0
wv7Dy4c243GMkwMo1jLDtWqe9mbduMmWViQu7hWU8esnayMUmE+Zq3aOtKRjztPXMQFGux42WRcr
u2N34WWs8NaJnlz/h2qirHyqHm6pc46j8d9jcJ7KExDyr0K/AorW2DN2ZMfTBYz9CL88SWjnv4l4
qrkYMDPXdSKSD+NWNnzRTc+OrJYTxZjHW2/HVq+7KEkK0F4tmSFZkSDemoq36xGBHrKWrD4QMYPx
nmjnGYTlBR/G+8p4zGJKvd7+ar1t/nwuSGwcWoZ7DzcxfOsi8ANnu1O8SLQn/8e/Eo7dOWbqRQqG
OY7NRc7sruKGS9w9PRu3Egj7JVJGesSCj83Pz9NxKAo+icYm6jo3clAM7rv6aCiFan2HVAxxzb2u
XBz47QbDMKxgtf71kaOIjbp+ejRzhYIvG3tyyaMqPcHRD4bS3PSwUhe4GZh9JIB3DRe5pLxzI+gw
c3s3/NqtmfdQOt8zyccnTXEyHEk/oMzurG07YiF6VwqpXA3Wi7pbUQbqfYP64zCfqcPHu7iiJdVb
8COz5uUwTUN92rsNwtunYUSa94AtzYKAkfigP+//bq+PIctt9j4W/YVTH4TUUezHkUJ4lS7xZjzc
9Ps38SevXbX9bdqiedG6yhqfZxFisEBIOCblxaGV0iaprp/fOmjuAfEiXBPsC8E+ZDGG8p8AGCIt
BSDJfGHmxW68xNUQpv9SI5UKuZ2WCWPbqYLU1X00Q7fQMrdVE7/0A62dlUdp/ubUsk2R4tV/xbZ6
U7rpMho5R45ZI7ajZBBGLcGEjbFksMYDnBmzLTbe5yhvPrdrc46FCgile+pAKIwcEN38qH8XsQf3
VaEuuDmzUeKOmSjF2+e3OLN+M9p2Ocl6cOZt7cyTSxNH2N0nqZne+37ovwD75NYAhhhb5xaFzwiH
I9KlLzyKNhjTuRHcNntJKr4VfFKo8tA/06Z61NV34VuR1DCWuVAFiyT8/6qAl4D2qp5+LUV9w0OX
YDJPPFU4XKgDyWekVpVAbqnm08zyz6ZCj7s0nSFDsoKuv21kKSIR+XintbRMgrdmi/AonpLY4KMz
7NbrxdODnziYunkbxXFDm0gqD7THW8tjdUJJb+cuV90nQcwVWYcjqJNfSTlbzjOfOKpqXikXUla3
DDY6WxqlHXcdsiuEKE/ha/lK7XjEpyERBqP4DbnJ2Tr2XcDMGIAAVKfXN29JXMr1acuhXHsXMe8Q
k5VH63AL7NgJWUYt9i16HHbrJx8gQXsOrFLR0u9NnuEmRcQxT8AzsXh9yKq6rSnTwREuLK2yx6Z5
xj+N2fqBf7vnAvGE8Tb5s5cl2kv2eHbQueV59z+0NDQmuSTwQCF5zsny8PfYpfwIXgI40Kvbrc0C
zchr4rdwsgmj4DfLiGPD3N90AmD7E9RRn6h/t3QMIMlJgdTI03KTyM/qX3BUjnfrSGOWuWOcR8lz
rQTHYWALrrNN2eMyX1Yvh6+AR0VcVtHaLJQnwlsmnIXZRmdy/ckLNbBUOcYtvg0t8W024zJh9uVY
J0RudelFqiMWGg5Oj26+IaaqTY+GJNNKUQMQ9nFD6yJyusas7xE8nifMoi/WyFvOkdv3p4rR5Xp+
PVB/xVjlJ12xLo4c6W8SjiuQgMuzQvESOP8IhKPDvz9cNL15hUkRCSyzbaUUVqUptyltmp7uVycP
eViCt/fKal2QRC0AqqAglO/2U1SDKYA8f3KEKaw8FBuTiRLKA8M0WtSc3zPP1n7Bv3j4iSqyAlTP
GLX8Mh7nHtvKG4JXN1NJA2hVkZJaaBDDmidWzpBY6JNzJCKetns5LPOzqgvxI0rRrpFvJq24e3yo
rT5fC+z/p3ZJ2mRatI0h0yGDOI/gMhTa8+Cp6wUvHe0tWdu4EkDLFHqvyLm2LegZadkCLtTONj+f
cX9GWS1wPcB4CzbtAF9KsQBim9LeGx9NKkv/10J6QaMmT7GLPosFa4B2fsV/+I8mYV3Xm0ETmxeA
PBtGK9tDjKVqOSJZtQzcaafQ1xwi/DsDKH3gGK30KiDxy+/Uh+byTNlVRgrJvGIdQQONHCcCLJ/q
HsveBYvUgKKcC0oOUw9SWZ6yO2+dKfHy5mxySGj93fTiwJo1PFLKK/xTeZMLW6J9sN6KeaN76caq
zk/rVshPvygGHGUjvP+djEuj74QZbE/d9NaW9fREoR/lMQ+RJJYcafIIzE/qCj6J8eiYI0PDUjJ4
8u1ir4+39x4xCRGpV/fS9fqdPruiGewWILZKJJUjzz0f5t4SDqJLFxLsC2N1iCtbAPIw57yfFp89
G3TWi5HBrDxn7SI4CxtyTIGNNTIBwyizDMmbeTiOcHbL5QcjPLzzI4qFn87WXeRAGLQxs1dmR4sR
cW4KseeUfSvvMdAu0sboXlXHfHXk6FG3v/xpQrreIze4mO50H7KBIxABnwR2yR2IFHIcXg18Ex+t
I7onPnSd+Fr93+05W9WHZClthGHo0oKqvR/VNVCO+Z0OCRik1Rfgd4k5cjnp1Jy6Ot44Z+llinWG
iQPra/KW6kDQQez+Eg3L0+9g9MRaTzDf19FlrOdAiRR4+pRMqXDaiMgAePqYPI55gftr5IEURwxu
5MIrwXg8s7799WxHmxwkr3eqht6GWkwvnhcORaN/cjE7cc2n2Yha5cD8oliltsRGK7WryJNBMiuI
Xds5VFiBGTU3o7QKSqKjWCF7+uVu5NBRfsOsK68cDQ7U6wSv7rC4YXma+eWVO0J79gzfBzXaUoGE
jAS+1IVpFA7rWpb9Q5xF9ToO/H4QXKxtmudwymGnwHo/wG/K6oPT0pX58HdXVJAQY0TyK/arOMrm
aK9hcSq2Fcs7fXh0m3m1hWdmUlB0vVyfjIW7o78Z8pwkTvw8lML0FFJW3IfQpNpHVcyZyBIbG+K8
7rve3dQ1MiKL2eix3x/3Z2mK/NSY5NC7VNQothnyFzFqoHmPcZreVSy+0osXLksViBeqGjWuq0hF
Q+xe4WvXLK00iIjOBQFkCsdhGctVDl2iaoTVHSloe5WkNFn8J2im8bLRVdELA5CIJsRsZFnVvQDd
PAk1+TE+A8yZbE7QxQD50LosmG4c3fdL0f4ispmdDVBmshBo4UTjdox1tloBPvcjhKOfCnbsoo0R
jtPiY6ntFN3jka0vMsCYBM3OUkTaWW7IQ/vTa9KwneqDW1/d/eATjEAvDV7e7cF2qLdEooL5EyrW
fMg1fooWbkFtwyseG13GL0HgxhY/BqOhVpQBimuTEwTxmDdnGbSuV/YPyYXmKrOG7EQs/eVGph3c
yNODSl8xt3WJ3ah+JGQzuAeEOfc9hwHPFrcaTjhuJXiaerQP5pRzqnvbvv4Q1wmpXQ7Ere08v6nV
UwRgbV10TMnADYbkdRUn01V+abBRkebzXO9LWnMDViu4pwznQQjgfn2XEkKGgY9cIXFlMxrE1T9A
BgMblcwS6tLhgyaTmoreTv1eD2iWSdlOcxaOsPgyNXy0X8xq8INGPne6NpN4FW+cnMmJEO2zN25E
7O6/yEzbEfkH+1o3nfNX1JtJ++/CY5KZ7TLgljeu0/NwVuepnc2aUs921q22K9onCdhbIbgnTZ29
rJxKC8EEpGNqi1PgE1Dk4i/BgIMETlUGAMlp6m5Bpfdpf6HDXZW8VKAqb2oK9n0a0jlcbnazQl7A
6mKwBErGL9tp/qa8/5BC41kRJ3CX9PUKJXxMSDfVOlEV7BKiaUh1yNGKgE6ziHpU2zAGq4w2HZu7
Om7UaX4H1p6Bf521+0wxOCem7VReHr29+ZjPF8oh2OtSVVygQPvFI4RFTz7C5Fu3Fq1SQboRHvCm
3KBzDMPlInZC8cg3UXYG0R0cApOzqFSQ3OAmxzjpZbGhx8POqufuWhyN9Em5a7q0TlhbzEFa7OU9
wfaig+5AeE4wC8EftNE/K7lER3Pn3ZjZh6cp6lGYI/wu4/vBKujByJRlmbGz+DCaFStVOh1LvCDO
VsSlt9CJkab5bxAP5HY805a2DIuIu/w0tGMC6cniPz5Oz307K4cv+M7Fx1FxNV5sVzPje8e+SrHC
nfFqCx0WiXvlx1oQHUXfySLUY2mK2nvlim+2QGuIMy/myct4LahNi3chClcHgHYrBfG77nOwpI70
KtmHh5g/BWNOl6D4hN8mfc1A9xosruSO762fibMO6bltvr/RmPz40eAXCBmZ9OL6DPEG1ZmYDwmI
KRgydWYVu6NHwyyhD+RPtSzo8PlfKxTH1I7BOWiUYBL9dHEFxUyGJwY8MP7Q2AeDsS6IuF4VWLb+
yRp7pbMHcYKQtMXeRJlVBjpTCM7ix+QkPqPsfpqfn7+UzEC5sAAf3l4Gy55jRrqH7YMLCMzIRVe4
ujXN76MPmJ2tGXxqJ29lNRDK3lPt3YF8tLsvtHpy0qMAumYAlkvUUtsYKMuQjdKVu3TrohtyokEc
/NeN2TM3PdHYC01KxzU/IFpf/vjWhCCyZEf5/d487vORVY28V1lUJpUXomfkgqelbhFgaBHwVEyt
F/Fd2OTt44BNg/RyLzPFidgd/kPd/NWf+bK8fa4/2tjISM9xWxoInKtrVu8oXm4xpniDdXkLiDe3
STbclMj5k2xPD7+3KEbEuWGZCrH7p98+3N759hXIVdbnM6x4VM2E5ArYjsiz4JRlVN5dYpKwf6uW
6LuqoFe6we2dAEMjSzKK12QHXF3W5Bnmura5Y1P/ReWaMCeJqpJAWIwurpQUQhHC5KsgVKWLi9fI
acTE5/xbqrZc4YfykvthDzL5k6gUaaVz24ojoNdQJwNsQ9r1qfVD2f0ky1t3LJfdFXw1D6S/myqW
hWvSRfqvR9LImv6q7bHQgK+X25Vo5xGolQFB6GEpNs0cXw3VYCiwQHK2jJFC6dt+pw0HeI3eKeHV
WJ6KnxTjBBka4whIZxt3+6VWTlihX3M5cwYm3Dul7JF2r0A7I+smlbbMAv7r/jaZfUNYMsBhtwW7
Tgob9X5H9kgnT983LQMPYv2eoKVdKpcpKSQ+Z7r73iH6RD0Bx+2MFGjkzQqrRa3Z2bMSddI2IlV8
ltkpYZ9vYzhB9T/S4f7B3Q/nVyUu7EJKuTFQ8A8OOI3Vw2763g6VFxNjgRg/9OmFaASO3BdLjd8a
uGNfYrW9ovxdx7GrCT4D8bX+rs3wZ/43DPAOCAx+YjEuRXDBAIFb3MlIyO7D4r/AHxESI7kEglvJ
g54sdocfKiqBvckSIaAozyidYuwzLCDr1Mmpa8LRMTWjKyQkMDY7CciQtZv7Cy43mKek89CBrREi
H45/aYFdU5FuARQK1g5YBfWDYdRyMq7zSDg6tuO5MqUU4XzXtl6LS32GmxcuCtycHlKHQAdIJKP9
cnf/koQ+lTUgIfcU5soEc4zQYE1ap2Br1VK6qFIDe3s1nTtArMxSdPTcXC1+33l54gxYrPQts5w4
9eC2gJXaZQNo/zenJD2rjm5jKoRWr0I0habnN5oJNfREe1Azg8+lfoMx6cQPjJpFpsRc3A/F+Cnq
0BOC2VM7AqKxo6B09Ea2yLR3mxYywqaTs0WTgpJzt823xuDwRqs6qv/4q1j209rlMSdNH0HsaQPQ
6bHu0hnxnvZiDkhTcX9SgnrMMM7YDqCyQqYR/jk9JYWekT92f8RqvNH+Tsdh5bBnQ0GB8KZydzVE
15xMUVDjWd0yQfjfux9y/sZM7wUZLhi4MWZe+QaOuNRddvOQAw5z9kT2hLwXFPn2P5enV6BLxhZ+
UizGHN7fVPUpDLcF6+LuAQ7aZThchToJ1DwHr17R/YcwAodAbUVYiPHSBpGGhIgIFdmkmHdvBpbr
ENSSneRzr1jLriGIAy0gQRkvvfdYeMYcqxjdZuZ3cXAm/JFTmFq4RQiNCCwdgsjMqGPdFADBo3uy
ddcXPujPKztWdImfXpX1QcLqD0vjPYNIIVh6RYpOrnRK6rFoDp3HMw8+oJZ2t5X2EL0pSa352Ukw
wC2Q3wdAFY6aQsqk7HGSxURVC8ZwRo/GBqaxm2yazlBF7GNVsIHb/tND25PzpF+nhrGQc9du9SEy
V7XDjIHw8FoMxq6Dti80k6XNtB0y3BjRH3hvJ8gb7HuiZpm62oeMy3difyMK9cgKTKH52ahxF5RG
IYQ4WOWv9Tyjwjcadlek+Bt9YGnhNB7QfVuc847cH5R48zCQmAfgKMFX8n4ei2x24UgvOUL9N5BA
eau+huGhDUN4odMA21TenUvUiQcE9VWZ69abNQm1w5YZU8jmCAspHFMnWVKioyuAZIZXYq3LW8dM
kNnRqJuHqzBXaZuHZvyJssVJNSDaCatd+bxeAN+DsScNI/EnpMmiGSYJrnsuMbZqGOwBUjk/bqh5
ogelQqJWX7WTBKQ6jY/HiaeZyZpVTjle2ZWHPZ2USNYfOuKJRoYyGcnCeg9j17goPlCS8F71QB5c
EXT96kX6YFWNYlCu8wGRmBNjphEI72tp7Lc+6su5qRdCMKlL9SS+KHJDoU126Nisna+cSWy+ZKC2
nKUSNTNI1X+jV/d6x9JEd9MPK/0ZgApPTzj+HeA7ZiXQUdV/eqYM0LjxpRl9SedXAhr/TtCDN2vJ
vrEHM5AsnAd6/97T1+9mIbgDlwLLsqs6t1hb9+fHtv7EnxPc/feRCLx1EiS/OS6TIyX4QsH3BdUn
yRc8wMwW3ssFAHp+zZ4dRFntIa/F+kdUTCfCpZpH8L0bbWoii4DHvYXQ88FBTyVER7Ib1ZIbo9pl
JuQEl0240wlfge+v3oDINAp7gNYDd6UokemuPvrF0JiXBXiROMyjLDwaqrMx7vj6lhmMMX/weI6e
jp8FrBzIOM7in6g8COyZysaUei3V6bM4tuf8akdaWZ4CCIOkqVaJFx/Nb+KA6OEeuHDMAyPzcQCM
DQ3jhXoC5MowsdVGP5Dykqamp0DNIKnsW4WYumQc1aeWkffURB32G3qq5pgIkeZxm3FQvCnZeq8q
9ICOFJwklED0dueoLG+snOfaQ4yTOUkqvb6Aq2jVByjiEHhnzokeUGBfiLCKeAGoIpxWR38q5zyb
bDBMT4duum2FOkgBD86hbWPl0fNkLHrFNGvwKQlO4ZGitYZ/uMIQbCNxdVdrZuDSiKd7Zm2BHjL7
IQftwFOmQWnBsjyno8IAokpuNQVCjgF9tXZI3HtpcVYBJ7KXvLdPMhlUplOyyKBAMyeWvhFlWAQK
bHnHTPnbqf4KGjNcxC90YiXCNPrC690f0N1hwwh0iUmSo9E/s2Bc6TIszRZYMqzl4VmDzyra8hfX
8ZQKaza6pedlRSf2V9EZOwLHXybzJuWhd6djMKfoo8zkevY33178joK0byhKQ/j0UH4zFxslM8P8
4Pur91JUxzkHLs7WTAqyuWH/zk6ayZ8AOkStirvHTRSrQjOLWq/6Y1b0bNXuv2U9V8eH4z1PuYq8
teAAmFHxaviyr7U91hOyWNHhytxIelaYOmwb/nDAm/JTFTnnd8NPKh5ahZJ4z8TzFejJMmkL8Axa
tx9NyuzJgwKgy4IaYlr5ePogQMWxGvwfeSJTSxven3bzcsev82O/vs6CXeiBNDKUs6oe0Yb50vop
oTo/6HBKDFMzsmED82Vk/X9y2/sCN3w4HDPRkFiJyrpCni57eP4/mzk/EmrppLoHKVso3hzHdSKj
rNJjwPEvrWL7u/bAFzKo3lBwGuxx1XFpJANivNjiXY5c68oGs8+57+jHZj9hC7BmWrre9oGtjJ0f
x/qY5r+8d6GZI3yEEahgZQAJuxwaV94KRZOFDjhZ6CU9UqOvR5LnBT6KFJqeBMHGfXiG8wedJ2id
w0rM8mUwMY4lQ7HbDofb1hQVe6DcG1ChkEacMcZlonVEezxHjgk7LpixADxhfpv+L3SPtWY8bfRg
xSfAh9p/Zleb8PrB/1G12bhQm7Sb/7LMyVSvxehjX3gMu1n1rdd9ajM6L3MaFvcobkqfjrQn8k1n
+MBiZwECCT+4oivHv6kruZjkiqzZJHtqFuG5NNoF73UNZica2iNc//QFD2d57NtpCskTUYKWw/WF
7etAYIHqCmEjoZZn1CcDxKmIPX44w5r8HajQfgnnpVKMgchR7nsXFUbM0trSm3frTeCXK/eR7Pf5
t26IyaPA7Ww8x2mCE7yn3ynFhvWQ0cuOooLFyJ2PpjKMAA/ivOgwK7R5xm8nXG4PFGH86wMFvd3m
3qMcMCR1A5dUDDmMQVVxreZIBqhoPDWeTGl7HiNPIuTYi5Py1CXm//qj3m4WkROQ78oJ4dwUBaxG
uY6GWa3E6XGsJiFzBTM8PuExe3DK9NuohGgG8rJvWkjXKKvSzwGPjm5xS79tHRpK+NyFVhpoWY2e
xjPt/C0e3Roa/MhWcsEjba4k5FumuCVbERI1DW439t2io7mkVswCvfGJJPJYr/dZEyXt4uOCyE4k
MXpCB0LIDIeqS375Xx1qQZOb+cXiEuWl40s1Vss0RN693g5oEJwnWJHkbISjRAQLg4EQi0G3OYnJ
T+3d7ABHP7VjU+VMoK0tRSaJZzMe3u/dKdGuLsDJnEcAyf4mK1pdsn2WDuJnkulBMrfSW+jW3/mA
E8qpdfg/tZid0vjIWJJzVWSqPQZEd4aBy4JK/wXM4BNSTjMBTSvLq6kVS8l+W9dpsaR1YhxIV7Gu
V0CzsX7iy/JUuWi5FsKd+6KcVOjT/PBe+ifvSMr/Q+hY+yUnEjRGa3x1C9Y7FSBLmFD03pKL7ZrY
0FTGk8ER12eDErelINCTnY80nUWT7hN/RfQ11hZ9oqCgw3/FjqbKLMR0pItD2f3S9OnkU8rGcoq2
zx8d9QBobo904EiWGguU8WfSL6AB3sa8xWEFhuikdTTixiJ1HovuJ9lqn1sS9B2xDLgWbdNemmVQ
MNLpo5xo1N46v6auwsU9yerZ53mcKLOdfs1nlVo6hi7eAYxNBBzftpuswDKpdt4KRGVYwl1zvKUZ
2y6HAD/cnHSgHc9cSutOc+jhCK02ygbabZpmRXOdYCczCnwxxYKnZ0DG3g2s+WV1L+Uf/Z8D1s/F
7dPUR1W0Qj6vlD0N4MrggcClfaaHdaR9doBoWD1j2voOT/MgOiPEEO8Nd1ygyAv8tOzrHbNNT1qt
U7y6qakGSbesv7zu1NIvn8TLOCwBzZJRygJMkHnS650Lnp+y6ZK4to+sC8DbdvjdrEoBRCMu4Rp4
BpqaxZe2nIDesUHHywSYHsW7TjkIUMzoFKJ+2+dD51yj1a08Xi/Xy5LNHs026mI4kb2rc2uuU/p0
etrp00ZMOomDyRMo0W9tIm2hdxHQS1ox1cGGn9RjA16jwBGdG/GAu5DkZSTMa/BwgU4bUJRwSZBy
xoCcLvYswzOFzncrlTNmQnUPq3uBrJs4eG+O6ocxHyTSdweqW8fwAajfRR0+175XBv1ft5CLPexn
91z981GoeRMLzZbYwu5PW1MWAjYIf2hLKhu7fuvNvpOmeRgmT06LNFKzwSReiByTB2EHkN3f0T0a
kZAyn1tBl9rU3CiWR2V4sZkwyhs/aPdbGuM/DQJoWGn+vocZtyI6WYEIAm7/TWucfG9V3KbQluRB
OHzFHvPbX2ycbl0kmytL6NanWrKqQYR3OpFF6cZ+pRhB1QAyQdzs8wybkqEgLe525ysgk6MPuofG
CUBjSOjzLs9IreRgHMl4gomFiw8QdxaiCUbbEo/q66rjG18dD/uTLCq3a1SgCF1lXae7xpTgvDZi
zliK1+S/mZ15QALA4oQbbw2YItfnLhrZvtzgKHk6D9/K+SqC0MHdli+P9xCQ0ZKLfxalBQI0gwNR
CDIdzpuNx6Q0olQtOvAwid6DhZTH9JpLzH0X62UM2tpFvdDRu/ifAiVmOOOnpSeCcFFpjW9QPdW7
oinjGBzt/s6rK12pWsWru74MFwxpjUCtj53CYx7PL9g873W2oepZCuC21T1zfGQfK7tGk1NiI95O
LqPE86G7s9W0QzR42R0s2FgqMBbDuNwmonQ2uBXnV+ZiKZqhUEWh+p62xcn3dyTqInwPLr/9oTQy
iboX84jceGdiJyuUN/M9nMKxKyYv3Qz1hmg3eUftTq4MuYw4weYjsbTlrBRHtCUoOZVhjvB+qsKN
9S57V9KrfkqXNEfOHTSw6g50Y/P57wtKALpyDXZ+NU96h/MgQdmafuo5s09CgtyMwbo+svG3QKJ/
L1k0RFd6S5BEhwsFxWygd2huY8YbT26xDugj2/btn+0BRJFds6aFwPWTpEvxHzv2E9gviaE/dtpX
pdBzeTaEclTgIk8T3+tBtGh8P1wM/eflgsfpyCK8iCOyOzt5UacYDOvyB6TTfuEFSGn+Xx3xh6OA
LEJn1ixfln+IaddZheGFPGOqQI/xNz1N45ID0am4eljhQSNbgHr/v1pEB6ZoPbIMJKk8K55ayXkY
EIXxUxt1prjRKJK2REn/6tEXfXK1oRCuBspJr+cyoxU6LwXR8SF5g5DW3QUN+Yvs6tCeAOqqMxZr
DJLSUg9mPoU3suf/WuQs0gbJ5TyCwrWxcQ0AD1R/flt7FX8qULiTjS9sr3LKrjWK/wawKHqzl0zt
OkeBNquBQg6UfdJ2fsTMQKfzHowN+ddTfTtnp6ex0dXCnzJ8HIfvSuvVLLdcAD7teKD397wwqQ6d
hdFcbbLskPNPcqP4WmWwT/xMiZoW0WH6Co0i2+GjQqmTxArd4CxppWo1Od/2zbh0Qh1WgDRKpDGB
xyNh3+yomvMxSzJLPZC0tkDhkyiHkBBAgp8e9+pRdXM/bcMzhOKGqvQeZDvgNms2Gj7RN1UApPMp
b13X01SUg1RQPhhKqGSySqgMzFeNvNbPlf5DbwUdFW70uPnWyAnfMH3hzV8s8V8UnByxm4SUM+ya
pINcnqvRhj5/TdD9UUaJiUQ4aBUI/Xi5K2281O757jX/NFxjzOxRYmtU51Evg1782x7XJHwuDovz
eTmXfRqapZADuzs5VQnlvkIgD0Jb9P3mfXWExZP9T0pJbvN0hcklRsWkB5HWGtMjwMI1Ra7QcV9w
zWSDyxsHs9953aneIyCPt9VfKqjbZpUan0WNcepe5+TbPu5/JCtLAYxqhrgpVdraKE/19NtcEgVr
fARwffyqvXJaYFxr0HER/EN3xcczZNeBQ3diN9/PLoYx6ZosKDuMVRTvqbmjA5OGcqwo7t+kgjbv
sAPEsORwijsi3mIKwa99D02hNJ5TF96QgcTUu8/rCbUhG96p0pgW+hc1tLqNIYrsqvy6FBnojQFx
4YiJFyJQhYbVBSUIDlnQS71Wj1VuQQ/OEPrdu/3dYO0lo05C51Vurp3Og9Zf2rIiX+Co34wR1Ezy
Qnx2e+LZrOubszyg84jxzJ5KleJs18X/VfiuRo7NTB/AXjXW0D4/LlOAwHipEqDmWD4kU//jx19V
EXXKSxb2OeWSxm+Hmyu/1NtLHY0WzQpa2GsOIdLiY7ZSJKN4ocjoCuS/wxPkXwrStErMVhgtcZty
mXpeD7vER0r1erUm08t2sYjlauk7i7CFCfnIw8unMwAld6TseoxgnhOwN9Bt8uGXQMWuzkgeJkgJ
1ZMehXEoIZe83bT+rSbQgZlOcfce6/PzlOUtZWPh/xwJFrn75VybQIqhb6BetnKO2gMvUMZ124WR
O/qf1l3J8IZCZEZxxDZKwPOxgX7oztCOXuAMXUkCrYfQxWahei3Fa9b1xPxri/ibOUaTgEGAjvUM
v55BFyqXlHojaVkup61ds9udUMtdsUd894gMqf1/3mYQ7Y0qfekDXK8OoOF1otZQazShVY08BP+z
WGsVG8feCmMgBjghv5MLqYCxapnMci++4Hp5phu4O9oAQI42tdJ8JjwtqztdfvZnW70liEcTmcgI
WLHymwf0Z/Aoaxsj/tsTEXG3gBVaNAW6oWyjEDKu5njB+53IUhoByno9JKGJO1TKX/+bpVxfzrk5
QJUchmegTfM9cCUIBpsNuPsiOdol5VZxmOlluDs0UCeSi3bGQW4JLSYcEHV7gAANt0CSwXjxcVf0
PxCfmVTEWc93bFGPTcTVAx2lDhfHu00m5bbhMctpw059edvPmZ0Nqx5lgKJbR5NPG7mTbbpiUCn1
WFli0iuqq6ASIIMSLnfYOc/7yUrJBMBtzbEajmEUO+aK6v497o9d5lZE/+tEq0zgTk++bN9ZOJJr
chaYmalgwJH1AtHDfnYZ2glBit+bgNdOlfBnemmVlS+baWiyDmFyANfL7At4MQdjmBR2I6IWkdGw
PC6ycK+oDLsBMFPpUDo6C7B2PKkLzML9eCQv+NpzmChsjTWJe6e1ZmLuzCNKKh0//d44JbGtXRm+
rhpLDE9oH+66Fc2z7N1o5OWBo9m8u3IidxrokcWQ7AaVgqNCGNtYe2Hw835halMnnYvF0xGTYdH9
5URnAtKtHzQw6TbVafGXihHinxaRMrf1sBXEP7/AjJU60QPnhv8QRgP79qkx6zgnWUJlt2QNqpiU
c4i8D0h8GrBXv0zBFRMzOnzYGejMt2XoSrXWx/67qgoucmfQExPWKeQdx4XOqufN1Rl5D6H7VQLR
Y94m6k3RF15VUFZ6NC+Cm6DmDzJo0Q3nNtNgAtdre79Hg2Z52oaLIJzjWy0Lsy2Fins0WO7hok2D
BddmtBbF11A8rH0PZmNdhxPr0RZ7pTKQdFa22B2TFmdGjIy2/EI/jQ6vcq3nQrfmiEA2GOs2sEyS
CY/ZcnpQa+70QdNzMSjsVoFM7+TQCD/CnwS2LcvRVPGP3GWWzPlVjunJ9mWr5Lo9gougL2xa3UVL
wtTATclfIRVyfaUhKz1Mvi2RTgwYkaF/SGbeUgHuc+Lx8hXuCFrZEeJGX2BnM1zMeXR4KXyN//L0
wpRzaEiW0epayyMd0yQEW5schySJ/6j+o35CBUdUbjbCkRVPDz3qM7Gqja/80GjUzQf9thjJ61xb
Gmxq0qV2hFNe7QaSiaGKgO4h4x5rBSBUyKhBivZDvLwrz3F9K2JO+a872BBX7QTEl66D+Hnpctqz
Eg2pLpP7lRvZnEndWI4CqUlC+2qq+GYZhOMGvfTUFdRHSmH1z/hiLVNdm/hVKJfKoI3R1yOmoit7
njUdUXwsXpH0B2Fbs9kkRE2QwJV4Brgr67X+gOPUSunfCULZhXAFh98FD+qPF5GZ9pr+KB4pkduF
oz2CiyP0yfXMmjB4riihhSbJ4KVMlGrHyyFsSTSZN7bcOAFrHZc0HpkijWKnTVji2qd7UdwqZkZC
VvnXCHDWQqxURN1+Nbf83wVW6umWbHPvRX/jKVgIxoVAv8EsKENoCzJnlWHgiDDFNWIPMAskbuyK
pQ==
`protect end_protected
