`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ww1cFCaKpEaygJUT+P6Z2OD0uzJ4IJG8iyHDm5UNlVWbTWS9KXjZ9jEg11wJmlv8lA2AVebHxIas
7nZJsy/GjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gy0/aj7fr+HoqiF2MKC2DdMRffpsNgkz3LCA0LoXsy3oP+ExvEwYs55sO8KAxVdJaUPMOFr+w6Gi
VDRBmTTzMTTD1KvHQEhDppUtYnGyL/2qAWb6xHvmSHDtiAjlHews7qZ26fM0sYgNx48H6LSqgFd4
hai7P1C8/gEiLdaec30=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hi2M/LxF9qgAZzAUuc501Ws9I83yzxDz1ea90Q5QjM7jLsFrH4fLD2d0WWY2wDTdG0Ih+QNnE4S7
Oq9DybBH0zvBRUhAQoExlvdlIfU3Jr1YKpM3lLPQTLIhhCp1eQgIZljQtMN1p0u0HDYYsZO5DBeb
LZHGhmPHPWGqNQ/iLmQ+PQu0B5Cb+1VKyvK7Ipxjf6wKC/NZlztCmWzwV4WC+jY2wHB2IofyzZfo
xRBIRCIpTb+tTiKgZ9oAjPNYVjgXC51YW/c8ZhnzF0gIdh/tD6GDSX/DdrrBN7Oz/gtduYw5jR0b
WsJx7lVGCa/mgRPb2+p2mjuutW8gGGnh6+Yo4A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X16goI57idQ5Yk2jq4rj0BhsplRtdzoYr8oOU2lBTTonp1Nx4fK7AS7KgGuzY4UqvPTHmPTfD5ww
0YcXmh8hr2Hk6aIz+aWFV8C8XcReGDrBhi5Np0Vi5hozuTfEPpWuDV7kTmarku7FYKZbPt+lsAsd
f8+cIo7ySKaxPnzoHbw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RA9GWDJZOdw/NASVbYOgehelK35X4QCDpOGKLkbLHbvCU34C5eqCOlazH25KMTrAHxM2lx7+fAsw
HHb2ZWqK4pB4ww23gPcOsgxVCyXs7Dx/H6E84snPbj5EBFAp1p9GZJoguz0skOVQzCSeso4vwekP
kvLqf3Ypkz4/BbGmeIV5O3MvxWppwuIHCb+NDzDYU2x9uQ7mLUtu7pYCzPfN1FeLiv9ttZaXRuYJ
ADExpcAMpFzH3bwg6Tm6wL+J1DzA4jLGZxI9jxK+L6xNTv2NtONryX7sLla9heWPJCSHR4TT8ow3
t3QklA4V7oRFEhlMh0Nv7QVOAHjukKSZ99LumA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4864)
`protect data_block
2JEuFaTgqghMsv5lmjCzRKFTRu9v2Bd7cfnnEymmK1IpMPqqHVgKVztK8UcvkN/cLu6meLkuW+GH
jEF+IasLsTsQoEbARf7iGoWy/qxr/Wx8iI4qK11niwKvKRzj3E/VIfcoFWMI7lDjskoNrB5ON374
xdQdL472o5haNrGgEzQCs124gMoZrq6ZZftrvXJyyhHqGqmNNfQbG065CYcPsuRjXxzPltG3oMhc
7n7pQE9F5O4ObyVFgYrFINih1IyuB6ga3CPJSEZRwp7Gz0bxN4RD0DBaR3vYvY1rH6jZ2As9bin/
g6/KlClzLL3bvhOh9lV+NZ3eWmHbxrhNJBKH++Ph1mZwMT95zN7eoER7ysb5KV7rWbJdk27L1Pjp
J2AK+gNt7swd07+t+QM5FnqBfSQQ2y/64PfEyHTkNEdo4GM+mKi3AH8PslAcAFXIYE6fr+5XHFkf
I0vcZwAb4t17Xwwot+I+3SA55KPkc1jV16M274//n64FI5HGaz6z5RQz3eS/3YCXeImJ5+SCmlX2
ZaJ2hPuX1TEnI1Ktfyk/Fs8WuAphIKYyi2Nqrfqs9BKt2JtjpSq+6wf7tC+NZVW99sdxK/khYY5B
1LtU3OLzzfRSg3nQc0jpZazEojXeJh6sKdbQv0kD+Rn2s8esQSrFHC5HWniWqJ1DbvQHDVfepsmx
AHkh9NEOZeZvuxfjbHUvm00YBsADzr+Az3G6PtAn142pEMk7AE4+hNG/tACjIRA/Dq0C/GbMU+7W
5yf7zOmeZzfiMGYhoZSCDc0A3TujZxO/ej9MXgJl6+vKl9fKmtqMpAnHs4+01P6zhWfh6z5GR9/p
GiNO/IfutJNpOR8jYc4hWitEarSj3uoyIEKOtB417EqqwYbAdW68XdyBrNY1+ZJoNuYP5tRMRyGx
m4tS0rbFqhPwEvCYUwnSdI7wUw034fNi1JdCqycc7yOukkGEE3bo/CEFyL+a9ilZi7R8w9SqR4Wn
RgU4Mh5hH5Y+42e9wYYxA+Ylzq8gw8qW+Q/YU0/0u/83wEimNP7QeL756+ZGTjw1TDFTTxBzjUMM
/OxyJdpIIKrQmgBwbQD9u9W5WB52gcidObCqrRNaYiD5ZJbKMPODtWwKM+xBPReK5RECTIVAaR8g
/URa8PDmzE3+kE93orLssKBkVoKwi5GAWsH7pRvB8y3EmmOyldMeABfskoXsb0cH79OMV61GBKrO
ElPU4bcursnQOWwGLZog8r5+6oNOcdC6zk/5VdW7ZZmzPWZ3zgiVJKQl2mTCs78CL2O3ZmyUNUWI
Ms7ibMln/NcDSvvBPHe6XCPhd7jFvVW5B7eGni4odmjXmqFFzn7OUAjC2F3JkpjlhxtoewcBXIsp
JnjXXwP+C9iDMg5KWL/aKAReZMs6Z7jGJw6DsIMGKA14I0LqlwE5EXmNFOC5kuixCqA104lBly2c
xUfKfpr7zVxBSwijttB3WndO+MaIUxhAV6ZF0g5TEbTKZBxqeDuF8P2hlmd1Le4LtVjv1Lm/fOtl
M9LirFGY6w5ijydjJQmImquUjkFVzeTNYWFW/BHF9z3DgZvqJBlrw2shE4EKjei6025c1femgjCG
aSrwmiZzgYqnjWQZlTa1Yh3FRAz7L6BvmEe2Bn0D6luh/rML0w6vtsDv38Klid4y6JnmO6/OUqPr
LzF3F88EfVKFGpU51BU3DyFUQZmuAK05/lOeZUk2SR+R0QYi/bc2C3FqkeGH2idRVvwRG8miNXry
w3dxfC710bh6HbKkuhSogkN9A9pe1ISe3Tl2fhKA+XdF7j3YuWxJjfnTt4fHPGGFoq3cIGOxG/ef
nNyAWbnM31K1oKwqAfcVzXikSbbQmr51E2ufRQcPX5P0hw5QqwHKgU7Ka3PGOvC7hJIZpy+3QjCA
Q8EjbdslxHwYCuMdSiLij76F4flun1QuEvbuLTfzQK6+EzdsAvcrS0WYhM3R9dF3SLcfFlnVd0jT
FkeMu16FkJO1wC5nNLOKqDBkTfrUwUXlKVdbN/O3nHBfpnVOggyLpT5z6Lj2c2fexvMtDIGT4D+B
bH/JRHk2NlB3K9jDvDVOzruN+C1Zfz5yyGyQQ132DYuR+VIXJcJdg4/63C1gT72NnfAiwn3glPLU
t6ZUAQMDqsVVSwckicz/lrHMhhWg8Q6OBUplNK5+IvhNAgS2V5W3vDqzKQNTp1IhyuLXXM2LcwzC
OcHWoz1MB8Li2/6JzjIcpcq3ffLKaFIfjhrwoxELDh0qTcSDe3EtKWppIYb5VNLu0ycJSuwn5SBR
LZI8cwKVAd5311/InzJG4X6P/oNd35Cm3gS7jKvx2usq0+7n94ynIA7Jx9cajF3DXK18H3GrUXF1
nK519hZQiV43di4f420zM3oEac4f2yTdSzzA35G7dmKHH9BaUmAuRvZIZrMwXO/s2Rypb4N2Sn09
ToR6q78MItdQd9dgyf3budOZTyv3tuhDdBVAKxkiS0R4C7rSioYChcBQOoeGjdURMJWrzegldwDU
Kz0D34q+ZXzVG/QxrTbJbDlLNxLp8KD1juzeImE1FmUV5surZ/1d/GDLv96HFq1CkYc0V8+VVcCD
Qd138O4zHetoT5hievRVqmwB6ihTpaHx2U0Gdf5jGKk7d0uhbxWN+GdxQilLLIS4NntRQUJac3t4
HMKq190KJCIVnUFnRmnx3iO6oaVBNREGOO1bHh22osMvJYKrnXQgJIUoI/ORjFwdNM8yzdXkiY9i
UCC1CJ/70lx6OeGnOaPGyHOpfU/zN8qT3j6RR3jzmOKh2bZafICcRHHLHorCwntLphbi0+KR3LoO
lSJXXKv514XjmEBXC8ezIBpY+D01NDOtxmto1vr/KDwQDY9jOBJu0bOqM2GN3ouG53aomP/NP0VF
XpnyNMWtWGGJdNMrrmDd6bYM2Wk+Ai/CnE3fYle1w1jzes5WDvFiJFLuNJZwqnVVOjMBLS2yQB2f
tQhleRvQevR5KkpYE2YLi44ktOnMLJO39TwL1smV1k26t/hiVD0iwe6KUZfV/2idYRDizDxwAXm3
W/evPv4BP3KEdUP61Fe10hDutd5Sed2GFHcRy+bV3P2yHKd33ka4Z60MdQ4Az41rwL+qLKcP8Lb9
XyovU6rrELgA97WX5iTT1u9YiPmXNvz76VNkDxURb8eZIlLVzpwWBZubdW9+QyXfZ+3PjeS0df0M
ZYx6J45A4QMzyUTpe508imVTcD7g5GbvcuIZGLQLCbdCR4dKebN+1GC8A8/d5bGMfQorgGHLZ6Wz
vL17gRJjLEcsJxPbtEVJPVKKGLZvihE9aO2J8XERupmEa9agqnMe1b4+k8XN5SDg6RKnGiB8WmNm
dJ1+j7VYOh8PgDKXIUIodvfiDdqPQprXg6o080sfawKxPLHatwaJLISq7p89mX/YKGWVDbGX/J0Y
HPisNyhk29s3K6S8XBMNXfqNN6ZrkeM1bYA+R7orplm5gYhuNAp+svpNEfRhrgCEt8QqsC+3nAI2
ce/A9loVgLselftevBXZKBjBTfy4So1lGxVAYvBbag39nOZadgQ/Jfn9ztB/4xhvI/WEukUR0sdR
xfmRo4lMMvKrYIL6Wrj0bw8zbpy16IcZJkI6Kv7txuazyx6EaQ1O4b2Nb1DeF0eXQKKpkePtRPvP
2gJL+TtjSdVCP5a1j7eNV0F7YYigZ4ssne94W2tEvHZE5tR6kND2XB4PF9Bis54Z470y2rTmhRN8
jPhK/z1SdtKKlTRF1K8MroqluJc+/oEMAxIFDmFBQVNV+UqAeLX7ODHX6ruDTPcrxczCUKAadJw6
EGR10EuUEIv1swQ/n2/BChio7r98WUKJRXTrdsnYQ9jWDDtLjojHjSZwyJkTnmXbb1/EuuMTTq+i
4IfWRbfB61ZJ3J5SslP+1tGfhq7n/myFHbhTZY90SxUsLwsX0iiqd/Y1Ek4dOmNz037FyYFBBp6W
UjeFf+f1UfcTSb0/qtdO0k1GEtyV/eazfPNDDN22VxPx6Hch+TB0ZCqsqJ1yq99oLGiSdda8wJrc
tizrA/w+kYeB3i/jlKcCjWka3lQM/Zv2ft2GPC4Yloui0XkBpjb9tIwJIPFcWkJ4UAjXifJGBUtK
+cFb6/Lxgvp/+NiBBcDSLlCWDUEmQy40dA4tY0GvhpX1Jj9mapvOOc6u0GrakyTLD2toQVBl0KUJ
tQX4F2l+M46rDfDs00jsRQboH02/DAEFSn0SZal0Nbb9uamDmU29AaXxVE1etrdBq139sDcqE6cw
dvU73QQ0mM4kZve1vRlGf1b6FdGAM7kIIN5yGR8wSeXHY9RZsB5NfJTBwQFsYXbrJuqw4I08sUrs
355zhAiOL1SUCx+UbGhMz6pRDOWScJUuu+0R3wC7ghSX8Rx5IyYTnS4n2RgMXrcofU5GQ98Y0ZTj
FH6kyu8Ne7eJUrHFEuXyl+42jTToS2FLjZ0/h7AD38pKxwf0EDVpzdf+Eer7tAXfiX/Pl/lwwtR+
oe0y70dPKC58W6RohThT8kEs4XeMxpUOuE8DgEFNYFE/cA7RMuWjDH2xOZwHrkriSVXjW0MQ5v04
8etAGgFpgD4qcmjl+aMs2izHAAPkL152wr5fzD/LxurIEQ5ePDEwnAc+wN8TqzG0QnrfQ7yCAC5v
4qc2Ga7PXaF+wHjp9T1AN9s7s+foMXV23h/136Lgjf2aQWuWuve2NUBGx74co7ZwwBdUnEWEpW5m
xJIuItWeUOliNTzUQ04OQKIth9ddUK6pftfTESGlgd0PzVOkgdzOwTbqe/+F5Gu5yVqBLABBvOX+
zJDWe7h3djUL6ZQRonUjO9zMKGgU17rAkUYRFqIJGOImPD8Gu713Jl/vDWm5ijhmfpchkzvecU9i
3XA3gWSeSkm20qstOnb1jo8vEjjn/cYy2WwUryAWC3TohoXKFpCAmgW4mU9FWQdZuPVntrpXABMe
zxJ5C7Qu+trIaJQVy3wL8rh47CONF+ZUQ/LqlipfvCfJpfyYJO5ob00nb9XHgg8Ia60UwjrKaaaF
DWejGVXlQGCBfxmHhSZ8Kyiw58jmo+jystyO6UA7XnEg9FVHL6uCta1GGqCatnMVMmVGzS7ES/Dd
Jqhusf8ynHtgHLXiEML3g6uFG8iwGbcgUbNXQDL9ET0KKduD3DHP/jpKukcrbA6p0mHjUK+sg4Q6
qz4tgIzK94kPLOBGCmBac3vgoMYpOTrDud82S9e3feGH5DEeQjs3YljGGTTtPavIB3nb4kl2MJ4/
mBWu0F0h0RlAVP5XK8tk8Kp84ou+A0C/JZhhO6tL54leoEstVlMMdLG4kKYIwI1zeSA9wNNFfGhd
C0UjiqW2r/ffo8tg7l1i6UAJzYA5gy9zy4YVA8/a4hQeFX2jlZGuXipWXFbd35si2Uv/4DOc26+5
vTaKAKExDn7UigR1Zcn6xZVN5kcJPe+bASwiB8k19pGyW1CsCgF1PcnZcil1Wvbi/HppzigEcBZo
yGAGdbmFsm6qVDfIHSkFLubKXNBqRxVGVCXzpexaidk5zlQGiDEXFU6HPnCohryzWt/5MTi2xMwu
67TlRYyNYsucjOODe7Txb3UtyYHSf2HXNlPfKFOTPHjlpKmJht0CKR3R4nIp1ISLIIPeDYH/ZxFF
hETODertKSICkRPSrOD3TOseGCFULoQCiKdfhQnFnP57u1CJxDdeDdPs/ZrSaD74dEBnbsWWuDul
41xR0P/fBOAaA6dHc1eIAOfeebZHWOUypW+4O+um8owKCBI6fXx8GfZKLYLWjA1ERqFYZBTzzH81
JSH3LGR8iT3t6VzBfc2gqegiAEkM//AoaDMFfE9adFq04H1YjFUAd7yLYQtWT2NmFGcr5FNHOkfM
650YQqFzjFwpHOgmHNVnmnhqB360MKGjzauCWLCi8RbEbkJWe0KOi+zOp+5qbpeUcqCK2u+RrenV
OEmC8XF2t+0pZyaRV7PZRqF6yKeKWhMK9vuf8PGQhuzeAQkxIpUn4dIOttUCzKcuFy14OfMi1H3c
74fMWOB+zaoQ+izNNa2Lw6p1RZ3CwKXATROuXBW9A93DUzeYa2VzZIQmxz3xBxzBkdKMZyt2SR/Y
kPS0AYmNw8YuPQKUihAWisEM2hIFl6lsSwrATGXKfqjaUBVJJoNnRb8J2UqhodqbOt4z+KSZ/NSH
77fAsqIYs5PC9UNSsNORxCcG2v+vUdCjPtIF3Uh/7PXafiNCBUOeCzA6Vxn0tXjRTYGGk56kzBA5
VkDQmP2C7FdbtBNZjOyBbPHaaN4wHP1GBc4mn/RLjN2TMy1Y0AQen2s8THD/RNwF8GzeSC3Lve+u
r9y9evrC56WdrnMY3phdhtgSTSL3NtjvdyBjYfk/JmXUwGy9J5jl3z0Vt1tH90PYU41i8gMcbMuk
sKI24vImSNbMmKinWGeNcHFr9XBzlEM1kkvz/pIzaOlAvhq2oD5rl77hd1oqY1qtiAjI/ebQKt3A
WfLSt1T4acpUni8NOR4sICbhxQ==
`protect end_protected
