`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8336)
`protect data_block
wrovcHZ5qwQL2M/nAAAAALux/DExuqzw8KW6lLz8uZ6pvg6ZX1bbACzn1a9zUsNaRvNA2kkXgBPC
Ma2e3EkrLRAliFaJ0g+xc3B8vUQlqdnRAGv4r8CxkRu/vvRpGhp7XZGzypZx37qzMPeH70S8i45n
W0VPBsA+/tt6Znuqv85ffiGBjENggH6qBxk3uTvtf1KPN5ZjeSf4WWNXTt1KUOT/aDrx8+6ioJph
5xBxWjR9rt178PcQifdNi8yIzeWdAAnKzGCi80odXZ9mZ1W2l2QTU7w0EEw5jeg8SZdIggr9Hm/c
KmwrRnA3qm8nnYEWe8hoACrwwT/Fjr9tpVXT1eJrz7cnWcQzkAHr0jvQNJ7pqCiiSXhs0bjHlbOS
eE03Hu/ytYQpdg/OcZe425hwiq9NFEhEHqvo6jXK4uS9xRf73IMiHlga1QBe1ua4uDRNVXfehvvn
tN1TCTEGhve/kbAFLfJST0W8ICrMMh3Par6Ie2bTKJnQZOR1z2Jpv252nHlZKZGoXDW4riYGWovs
UQfLq62/my0ATSQPjlHywHJsr2kdJzXWUchfL/s4d9mKFsFB9NR3R4poacX9MDRoLM6JyjYan8P1
NawVURhCN6z+r4mL/XxAsgm0zxmxneS0f7vbfHLetMMr2Ig5pCkj7r5gGow86SXIBLywtPDVkOaB
QkM8BB+hrQ6VB/uvILk9lhySUOfL6dKmBx8EYElT+k58xkXI6kgbqY7IGLoMoJ815rFU0XiAwmhF
QSYqw4XaQ0nNBLO9ghTBj6pFKlYMozi3yDe6WzMM65+vlkJKzObZAecS6Tlg9YBXHhzN1i3EhXYF
2KjI0CWBGqgeCiK9kLMyXna9ciUXL2G/7c85m7mZb9RjDFUQzr6cQ6XHB40R7x/5rOzzuWPEnziW
5GSQwWNMfB3l7iGB9mKY6EZhvmjIGod3qxMs14bhV8yM7TwiMpbYlGevRPjSp7UwniGn7au+xYoS
GHBc6dINQ8tezCre9qYrlvN//oDzdWUjGFYj4SDryznWon7xhTTdZxZ3YS0XduZjNmBAZXUdHBKL
D0zQb6TXziXUSBjsCqRFuNh+r0oKIUsVMWfIFtki7i4HEm1z6Dm2Y39/wCy3IrClUn9P6yMabB/u
Uxm4AvNiYPoRjSIQS+IYvz4Q1KBbwuU4Lonl8uGzt1DSCB0HuZHcYb7hEZsVtgz+DClIKK+enjRX
dzR2+/0TATRSwNStJiT47BgjDMV/cLlLIpbJTUWZR0vCY2yAOdIQ71L+APm4IWTfUw0R8GaADieG
VaAodmGBGR1Eo9fS2/Xs5fG3O+NxXwzNRkRovAB+WIwH7jyDtdppMNc25fBaRvQ4/1gs3uxG1nMv
FgZ0uBFcEQi6RWdDZprXreBlS6aujy7T2qqvCitDMfBVrMPsJCGODY7fDejBPaFiO9LQL9buPXsR
zMvvADiKqJn2nTy48Hj7rFIX+/4MkevSajj2Jn7zkJ1vtHToZZ6tHsXJhttVw1JWuthcZ0lz9TZ5
ERdz+2tvpjSAE7GwVdeQ6I7BGPohnMYWS/lg3t3ZumAQXD/aFGmb7iD4E0N4Rdpe9pN507ZEeB9e
qcW/G5xd0mEmZ/1o+yngzz3WTViQSxX9yGAf/zLrHShdR/nAk9bM/JTEVoq9zmUQqQKSXqTUER6I
cya1MBIR96uEEk/prnwlJHLnIffYXCcjaUBQIqOOMrflbWl9WPD3itK+fLGjDabl4jY7UsWFhXXS
wI3fFgZB4dYssR1sWM/zaiQpaC2KsJNmot0B3ZFCj5O9edakDbfg5/i2PcWf7EiG1ePk3zCv34dj
fp6mWknebBtnXN5L/szhm0CeBhWbbwtWc0G2MkqjClU+LqQ6zVUm0THS+bXLzgUidO3XGvie6HSz
rDwO2F5FLZCHHYzBZZ1CF4vf5bLAtsC5IsowsQ4JtxNHoWR2ba2syJGUJ8x1sSJwk/bxJ0zg1yj4
9+z/mx1o5SQaOKqofhE4OWg++a8f/hIPG92xigSzmGcuiYJHJ+qJzxZaxjJGYEo4i0jFasXC0CKW
oRTb/OljgDF0c9z+70CHRgtO5Xabmp5pBXu/nPr2kv+jQataNRyPecrHBCeJ57Tfkt7t9jUe+2kS
DM1/TN/rCMOSw0Oqs66EBwikCDoydu5sqScu2bKKmTRKjP5Ag5NE7bOjySrYBl+hTJEsgHMPEPb1
dvq+lxTE4Y8S5HsROSW4f7GDXcqlKnoa0pGlE77O5pbY6Lk3goSD5q6xgfhOmMGm1bJ2CgwwRu6m
XW4aeeBNxOFE99Ky7HBmKEas8UtUZv0ZHPcSe6kCDDhHOanX6QJtwdZD93U1sGhjaRXkWx0NOofH
mQ6IqIgCxse3B7K4rd1uMBuh+OojZj3aeSXs5DveCOJRsbZ9gzGR6VEmyULGJa0lsntnZ7mJ6ZZ5
8RpElQXKDCG6R+OGXdJBa0XOv3l/FN8gaJ663j9aKml9OYpSlbrhLQ7JQ7vJeLZTZrbpFnhWccw7
XUVS9XUv4MiFLf8XS4qEbmBw7alqIWeAwtCv/wYCd2qCHgNrTlKG17G+m2y52lMG66BZH4jUPpy5
uPHo0JAu2hGeMzx7Y6tvGg+f0WCcDLVwdT/1k8FwUrEHPJY5tTptvY6VsSRLDCyDBtrJFJ9mxK1b
tmLnpGXgK7qgI4qrOP04yaaKafZaN9kqcKw17gQGEiA2yQvn4mO2ri4m2hTR1bznJf5brawYyfKn
ki04vigzOKOFFgTHQKyFcbX9aMamGS90ocCFVnGkbHRWGZjETe7Agz7+o0OJvifhFg37oP3zT2vZ
l6TguYMdtO97JgIh+7+AbLSjwSpROdazCalSU8ZkQ79Jr3fH47T6DWQIJW/c3osoQh1+TI8Nmh42
GOBekpUXqMYUhCtEBOHoYOZMH6siCRbTjyOkfAK2NKv+j5OmbUvtagWcfGWO7Fn1XMeHjOZGYGC/
srgp6vouMtBggAuB4mctYqsaKXmJ0Bu0uAjCjttq44YOcYrVf5GZ2b1kJUf11aVPn1+Wkq1qkBdL
tIReLnhLSJ4fXPKmlLPlI8H/+5x7W9XSXT+T+D9wwvfmp9dkw1CQSQyxfnCubziA53oHYoqjOFEX
30LvglQ9113E9zSsRXxhHU96UXu2ze8H8vn6uOJlDk/8WuA7PvyEmzbLQvsrpJSCBl7lpkdcBLbu
CYT1ZEHYZmZ786pESNuqcUJx3HTOLdTkIfTEbxuHBtKyI2ABQPPuJyL/9NCVK+UceVtpwFmY4hj4
VAUTTqA/lUocLR/n6L4J/CPnC/q0GXqegOo5oGN1lHeVJbMFtT5h0ZeYq1n4aVxek9Lu9PQqABWu
YWgA5UtrQvnQPyXCH/EIdu7vdAtkEDd7m5BQ+LQ5/KtIyxZuwNZcHSu7gmUcjJ+Yy3uya5N1tdrP
w5wxNpH8amSlCygYqWgr0dTJrBmEPh4ETuKt7eqSwyCOdSSS0C7q8eMsQD391X83A7mjluasTmX+
r35g2JNsI/tK2MMSt/vl1Okic7jW4UPklQVp8ul6F3elFeG7MYXptStLHbqbvDHDgSsQSWXxw+xM
2e8NsqRWnei0Wt8R75HQ0R1zkdgD9Wddo8QZWgAD2MVcWs1rdGCRLwVTzBnrAeFFW3x/JpVJthrf
+4SWyYeP2n3NDsAyKrc1z8Hru4rwvEGQ3wEVDGPx6djfJLTQ3dJjdMKi36Rj73K36Gf5lXtB/8TL
1WmcAaB0cjmXUvxd3K9G00UMONUi7hbo6RHVzeIejqnhseIZ3mG3zlPXxuOGbIy4J2YRqkzT63mM
BUL8xstmKUmD1HiUxxWMLs7eNOZSVJNnheNadmOWzP0CHZAY9tjLnoW8laii5lLr/uwWUrPK4scN
ZimOB+PHZ+CyYUtw8fHkCUjGFYUSXsJ+koER/ueFf/98Eltfp9RcBFClxzlwJVHmOiJxvUmFdxj9
u6SkqKf8wrU+11h/lTfo7ggWR40hN045uXxFDs+PD2JXyXoARwPu9WkGsPezT3XzFjUoPOHO8skT
Z07Kr9FTbDkDW+Vt23l2zS7v7YQl19JvuRdNlAgejUwKIKZSYQ6K84ouDkTOZ+ZQNFXfBZDU7dDt
YJNyQ0qQCsPQOPuSCtvBFPCnehCFlJbXuasI3z6IIbTM816LyeMg734Gh4QDSvNNBp4dO2pza9u2
WRBm0ggGVWm6kIayCYlrwOdt+xNwFvSzuRo7DFyxOHdXEjgUDpBA6EnTeJP+/EN6ho45jUyg39/I
jNAJqCHJPKjy88CIBfQrwxHRPuQoCu9OFZrKMdRD0TZRtYgsFd2LEBEv0rGFUGT9+i9dTMAf2EzL
5IAxGCSlMTtFbj27kF6DcdFSANUqthcVOqepxzG61MJCwv/qiWlz0ScEcaeRnsE1uGmdOEGyNMkO
ArfYq5Kqo7527lGbjdW8NpL7KSl5m7ey/qKBuxA5N23d/zVSWhcEfUXrty+0bFjKILAI5rGl39tP
oToW79mBKEh8Wkk1FxSGfRJ0WyBv4iNJMxm4BdFumWzOlTeT6PfFvG4pfHb+5kio9ebBAc9nS3BC
dM2Vx2Xf2tgiSgR8E4UaKYZxP/8S935x+cKk74lgHFyYNMmkx6wLxnVypmE6YEBgKYbzWLosZOKm
cd8zl61qFAEwcS3qW5MgawBd6zoRidoF7NlA7we4e0ljdkdpvZ2yJI7Qd77z+V3RuJYBR1xZzL/4
gUSsxCbyCtLViYvRGiDPchMW62GUyXZTbm+fhhso6F5G0MieCf7oo8ISAkJJZFPvRER7tj0FWIow
TOlsPpkFjSr/6QlSlxLthQiq4KRu//rIaUmdqiWo1p2zfkuWYG+j/oCFXCuxGmEjbH0b6pM3OIM5
4tk2M97jvm0NRb5VfX6lv97AJySMoI4R4wemFOVTyllL0tH7PzMazQNqqYoQi2FEtHrCYtu9YzC2
zDj50ogAPqyDufdGvxUh1u+8x3hida7MUxlt0ghPxoqAmhPQiWFmBtPcq4XjptfjFtbwhSaJe3I/
cFgxhbwbM/wpZqpJULzLDayqT543dLoNY+0Wjbssqr2Po9GUscNNYo4hQF+6Vk3pCNZ45l2a/kMd
YKKgRlhhgbFJ242lfMZBL5uOQxZVasPSebN+oh8BKphIj380hK0hQhhXcPXuoE8X5fgXKzRLusFa
12I0+4O+GaFD/idkP0mCS+ItGgIOqodSrVKewM8+VFlGEd8t0QhagDR/0Mor3cHRoyDZP8tPq+xm
Pt8CZBW9lYma8txaiuX3jQPp3fvS6QRXOdiStEMun5N7jzjo6FrvWY5/7EHjmwiyfAnYEl+pyYYR
wkDeaZBhrQ0fnffh1bPOKM7HHoK0UY3Dm5AIqJHXpR3t/5hklogguwlF7HyKt2D4OwQx1P2Xvoqr
NQHswYQBCQDO3S7nscOaf8SnjIEI91WYW0kT+jh/KNwxnmSsmjw16GWpiy+N0Lrdau6LGCK0xa58
/pxUCbL7+PG0BmoGa+IMs4qBWIJfn4qJgDCrqfe9FZ+aF3MgNaSG1mtFiDsVO5/QtPfslC2apDAV
3vKoM8qgfGBjOaQLWoMtKcBwm+y8SnSPzWRE/U6QIE+qRZYbdGCJhfqwQjIJhaGgPFTLFHIvA7sB
rAOes+Lpj81RoHCcUcpAXg+pBxfeKjQ7qAcz69opHGbInGrxawhkcPH/MGLemFs3aB9qKbsybi5V
TS5IqYKKRNxu1JnKKG3rBplWGw0qsh5vTgLwY9YzQHsaxL0qYgT6Sm3Yv/zRZ34me58sTu2n2lUx
AOdlntJ4ZzM+nvdCW2N17mP2XNtvYfeYhDYJ1E04kgzzA9TMXlv/8oxLKGS3TeswtxUkJDHAgMxI
tVvbKIkxUnkL6WFBeFw5TvAWIfoxm1XsuDN8pLVT/g2SJfeu7zq9I9xuF897+oPThNkf4SVZIVc+
VtgW+wEPNmIsXoiUkEK44+LjmwWOGdIg1vEp1+7VzIPYdoLNUYvjyQawBhbHLD3AskhzPVvZM4co
WT/HCI3Mgsu4ChdEP2FLI5OdeX7XQk5qhtqZsEW36FDcTitwLHHtsh7C0PcmpiBw+tU42A9GbP5C
Qlr1/YiBslVdGQP3MmE4fU59ZI/vWLqRgGZyiXtVe1j+SabUszsGXmGR/it0mSUDUnPJl2m5ZpYG
sfUuK7OvTSBvWWq/A3dWyj3tTE7iHTnl4RsASGXCXXOXSNyvAoFfac1Ixk2/CJ1f1mQm9oZGDRTD
1u/DsnCGGjz2bdRjS0hms65O7xh8XanHYdv1ghDPb4t9n4eJ6TCHMMnGH1itzwuP9Yrczw4hVMvQ
Fh5JMUJjMsNGgznMRlSBDTlD/+HLypjCWf6897z2lT8udxJ89j0vpuGCa/kiUGlid8A/0NNN94X6
GQL7Eu5MI6wLAXFe4qwAitFyrCu3m6GpZS2FQVjgwiMIPGsX5LpWbrXK0aRFQAo9zQJQ0rDivXyj
fOMd+TYrD/XsHy8FtrOK7D7NvTntMxtoisSHsvVAePlHamgPMF5j3OBbVxhS7DA8fjXxEGiUTd9e
O/swilBXrzv12Fyq3kP4hNMtDhzey2RoSlGDxqg6CiX957mv6xYANpyOI9NM+uCsVwNl5bFqWwZh
tYrly44mzB++TcGBR5kPSRPoe1W/4FVaA7ojCURf9DAhmuDooO9Ogqv3uFlRwy90VvFuK9ME+eJj
KnnLJ0H5/zoEL1Ub9KOMg9+ZH/2KON++hyYs4x2Sl3dXCRQELIQO4wNF+inaK6/1wz0PYpUJP9Xv
M40bIk2kvubntYz87vIHzEfWyrJ+KNcNF/ttaAiyOnbmpBkb4NfVsTXQwHNIHkvaCoGcbQNdM515
rQO9ptrK4CDXeumoU8mbo0Y4yHpBnvmVE+8XtMsOfGQ0eItn1wIlV+C/r6Pnuu163Hw4I1gxE9Dk
ffm4lbMY0wNKr/UkgGL6Pt32wKUGOuWcLvy/+OAqGGg2S7dAmkSDj3kZpznFiW1H4gtAFsEyzQXD
JeyzC6vGvgdg8TWmE1ZSiHHqiQWbASKmtEvgt9Fq7svcpoELdX/CcUGYyKBht0mZ0pUMBS/RWF/Z
IR7MQkC7bjdp2sxisP5iLJKIhrI4z8SeZImjHmMhiaHIGR9E5UNoERIjNWaj6kXmEBFeYVygbCNn
jGlEtFUlzZvx0zCoTDrk+hLrIuHra9tpPIx+zWHO68KQ22aN0lcBqC6e+HNGrT8Vc3/9gkgWtKY2
oRo1bUpAnG/s2ztNQHgrqAgo15HjzIc9o+CEc/cOh07ok/JCp76Orz2v56SyVH1B7zsskIIn7kTZ
TlLG13rbm3mdcjuqmFUQxNlZih6XRh85sB0rJSJYv7V7Zypum6n2e53WFFB3aCYEZoN5VuLZif+u
/Ijywxq2VDawLxIRitW/o9qB2jUgPEdJdsfD3AAk1AwUgwRMTnHb1KF/KrBFhEr7xvqVeMweP3UO
bn+oiS7U99+rOq8PsBoHLo7piMz7AHVb//U9z8/9b1wm9M9keWlSzmKLF8Gt7JM2lCDb/jFq2fQh
1RAp+FiSHSMUeegVW74BPhpNBSsf5UXHvyO9J//37pnwWbX9IJDvfd43Gq6zotUmIUWrH9kiuOUV
qTuxYm6AsmMIIkhholhtEeVfPRTSv4xZHP0/Bcyk4h/KJYb+Kid7OeO0MO25NzhkYPPt8ZHL9NTV
LLL4OhuZSS5hlMz3eSEPwr35tXDsIlJ1hnH0mPMgNJe5Pi5kutgwfIfTyOrBIAqJtOM0iopCcNnS
V6c/QijLFx2JSowy6ESrnHsBn33CvjJwlPeDDRBJa8V2TIjRNBffEgsxh7LMseaN6hEGKJnmuwOL
OAQ0o/FPN01w2Buuh5ItHo8n9G0cXVeULHnYXJLkvzeMZzNhcYnjyXdwh3bN2KyHKEKyPObXhzLX
hZ+TrxXdWVqW6LpTTj3VyGwQRCRByNiCmaHIcByiI0s9PHeqD17r8C/bksRc/hjGvlSCAoIevTCX
ARvOa205swebHvosiMTMlCrVK7uYo9HqB22/53HyVCokbintUUl+gFh+4COQ9juhQpe5alswYUTN
xuRLMtanzc7ubFGvSfOw+V/QXH5XeI3tbddF4n2mzGKVFnOzF5VZDn1hiHIJSBRUX0ua0EIoJ+gu
vYHkHrf3hIeS37mvAOwCl62cpJQho27dby8V3FbJYQ8mNvZzS6G1oqEeosZaX2jtI0+O+uKTT99q
CYhvIaTOTyXn06i5d3ssyxXxd6OHm9AGwWQuUwL9UEGN05Ihye5qxx3w5ICu4ATWwC4uGtusDQDF
1SoV5h29uewahpT2aOt3a6swOktPXNrwabmPiolWE3q/MBCf33HDjFGiB9ccgTBLc6PUy9sO/GTd
l5hhJCTg88mrAHOizIgJajQ5/y+4kJy0EFcYVmeNOY48qfjNNRGad/LMt2wkz3TnCTp+x65Psa8h
tlqPBV/3qykp5LpoVBzatn004o3gUk5jrJjASYYs4J1PaUC6lyjkB5GlaEY3w25Um8fff4i8QACi
VTOpdK6dpK3WzU3B7V5D+oJqM9SJDvCI1cED904kwaeAWdzsKTA+zCQ/5ZQjC+AqPPLQ8RCez5Ja
Qo58yh/iss9RGgfnP/tQDBQOeY8P0SvUVHm4Frn+9Y9sW7tqfHRKPRQ3XQQCRayvrLULBINxC/rz
7AMmKfOaOWtgVj60yceyVw4sgHjwDcULRTcphdbZ7cukExNhe271vMxMo8TBiowmo3kEMcb4+jvI
3ZpUkg8Hru0TfE8wEHRybOVxUn/CFIYFQoYka5MLkXhYD1A0GdIpLRltuAaUaXSbZ2U/47R/IRb/
5SC6W30A1T6Zm97NaLeIyxZdtHgS1QdVmIw5A6em67iIg+YOMeYoyAK0MLXibVh273eibsSYjvun
5UX7M1nXg6QSq+d6imCgkcTl/5vLQhXSr4FRqlCtxaCoGeEBpNf4ele0gkMdSFfqq9nLDAv2c78M
OW1oALSHR3ektei48UWSrsQgVIkPJ3Yo7/4ZM14ETnVPWB4aCFhnwO2ufhZUwpTZpFzPnehuXDUF
4ghcZ/iyXMo+B8QhsG9MdHlN7ZwFNcXbLe10knxJ6BGZcat/DK5ospro979Ayc9L7dQHOPELV5C/
LWYk897v85foItRExy/mUiuZxYRkJTve/p70X1t0zJG0RKBiZOVCbRQnV7P3n1dwmzfdN1lR1XHX
Eg77k2m0Ptj4cr77esyBThUQeT+lwZ3AcoFU8zMMB1XQlNTgH7n2zVj1eQnxBrHHeNwffJrsI3PP
zE7Th6vL5z6/AaDblG9sKExrXfgyVqR0Hr6o29MWTwxAP0lJ9Idah8PzMw+zLo5eCbY/deaToSlc
hIlxsDvnsV6O3q4pvoj8gYtmpEJaXHVqamc2Ls6Zez1QD7kquJPPdhfF98WwxxHDh0H+LIzY1G/S
IpJeG36/EswV6BCIdBiJ8kdJicnbgrnjVfJaCGplBSSie6SNVQ/sbY3bC5IFmxQosEYeIEjAkSvR
SaUF4YS7GboMqorODpEVjNM/GB7jzjZEGABftdhlDit2LgBPOEczqx+z4XyfuH1nBj5AEbj1rYn9
Nr+oeSO2zb24xO97eM38KGqefoRLsDlQDCIRv6wIDMFrm65Zx3bheHhWVhnWEhDq/SCnxtzOYDQy
Ny+TMX5eFsOyqZfH3bwvNqtm8lFn0IVb7uLQWwqWVD6FgpEOjZqlDKuvwvwhmGOgFbRVr6taW0J8
Ana2v7Yg5jnz+K8RKqmnJQoOGQjAPAX/oWeIpRPbb5z7qeWBix0jQWZdMggkvuEuYrkM76uzZwwT
dJ2G8w8E4Ad0YbHEuJK6T3ZA0V55pDHAhSB6kbAShJGQH+c9j/K59IuWYfBnwoXM6h1oUFZQlXao
xq775IuubNx+J/XyHRDIW7ZryuOLI3HkWjxPq98Fhp9zjTWYi9NWE4n2IueQorPp93g9A/Dnf9Sx
zOhxw5tUH4kKyo2A7xvWGb0OdTRioeXZquRTZdoa8P2P6FSCNUTDxOND4u8kBpPZHfZ+Q23Y/4Eo
lZkrbsFYlT24XRqs26vi2FOLqedDHrdv+z2bpkWLrvp8dvoNcs4VE+/zbyUfMuju3J4kcJrfWa/C
CPUIG4HUoGlEWjORyyU28s0K7hsH/ToWKpaB0jPXAd+Xf0QzqzjIJyUwdE3rjv2b8IZOA3Fb2PI6
n4MU+Jnb1JXe7OQM4UjGOJKx9jjqXcUzo6Ilp17tCEcxfM+piA4vAW69OnNLe5z7blIWsNBLvyBX
pOOIYgK1lq1TUxeOAYf2HyWHdwtn233swyOdDS3khHT9502HW/iF57pe2TLAUZjN9rJpVL2Psv/1
+1zU7km3v2jvBqg9TNgnCkPbeVbin2+MWUIG9nJOSLx7LRn94ah6djIEcgp1Kq09ogXZP/CGnuvu
YPe80jW9jjNSGKC2BqKeMmGDyMJZIRR53Qan9YcJaK0JY3HyEmcASSK0+Z1Z/GNqVQrJ+kMzrKQ7
LhFNPD63zQK10RBxW2ySlRUANhwk89dwtnhVNDp7vQDPS76Hgz/u5bBBDBU2WD++akwxNrjdebj1
MCSmSGhp3wlnfrOoqscqD3iNnxSe4lDO26GBvgAOgh6o0Uq/YBYlBTvGN2qrQ47J0AKd/lx2P0RG
2nbjhcXOyTw3/2T/GCJ8EmbjaSxaOYHSUPWvj7fTL5hqoeNwOVuDQ/iKxAkbW2Ww3iVXh3sHPpiH
OMMs6rmUgRRl7TIWwIqCamOevVAGpd/gBOnVK0dzHwAOlQLXgd7kTgya55VhSzmrGIZ5QSsNiovP
kSwNZJHvLPjiJLoMELW5fwZCuGzVp11V7hx3px2z7cjDvsuISdEAHC86pnATz5489DzBe2jok0da
LmANU99ZoAfvUJwS03Q057Eagej7AdT8dPLWX6WYn4k5tQQZTyZZ+BKvJeuKIXtN9QU4NsB/HcaK
dQ6lZY97yEKqsy7rEaw2ez1NKsh93gFIRzEadJl+zOcR35ekunqxlQRTvIP3vlTtxlt23MgC64xy
CgFN4PxsSKOvACwWjeGieE+WSQKF8+hCIjBOJt1aZOnMJqLkI10cEW9wR1zuG2K6OZb2Tj1RiXZN
Qn+qeAh8/WJlTLuorN0=
`protect end_protected
