`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZT7+RCzMGpoBYSuObDu7GHIWP4wbG2z0+NZPy5ctMvSzcpDtYTeVa9Rt2jwWGft47o5EJP3ckUaz
ga/PA8jA7w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nez6Bl347nb6+rwYEAGUgNCAGAzNmFU5MeAC9+3K2UzYt8qxPFrJ/SFJLhvmq05ak2WdPG0DC6DY
KQm2he2dsLt5QsRiFYmj2xAL1KdqCGiHsVFY+u/PuU8GEcfn2GTMt2pBI+06udHlKRy3Gt2+icT+
Rzwp56VKG96Z/MuGTf4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bJ23shOZkE3PVggRHLeGJ2PbG8xrPMkBPZCJ8ZYfdCaWhZ4ZYd1C1zb43X+ojqULL2oHyUgAMgSj
ecIJtiACC+HQhYS9ZAedcNObDtyg4oslk+vfdk+TM2FZF2Etrw/yAEbq1f/PH0Kn+mbNEo33Zwe5
Rm8FZ1wDWOyOXh016tcp0RwCvdj2XR1Kw/zAigz9XUFsy0aJtcUXIJIlKcvvsjSATgFtlJhxEDo0
pnsWRjWP0UYdXkfmSQNXFz8qVRQRGSAtue/7tEuKBK7i+2io/Fn8ReAkkGJiWskeE9nOr9dx+4DE
9tfPWFjj0ZgyCy6JPKhTrEZyje87nH/0x9mcFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dilSTjuujT5h2DrLDbS/v0rUBHgSqc1odhqH2k0dTfIZcb7N2jGBdTrXFekiehlmoGDjU9sGGdlh
yFg/bT9j8pTdVb3lIkuOyMiLP0CoFYVl1z2IegKN7b9yFR+7EZbxn0N/B1ycLjS4ssnQq+SGbWl2
k2N7LLrQtkLu5td7xjU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pVPXt9t5C8qS/9IP6M6Y37REfDMW0SGfG45oP1DNSuCggimX25Htte0JNMgNJo8ar+6qTjWsopD4
IXOQzxTzbzczkdAIs6+pl9RpNOeJpa0bvybm+uwfWb8+Rcnz3NLflVxnmjLM1ayKKYARNVh7gQb9
C4SQt1FdooQ2JWlTXbp3V2aZpvw5F49u06L9Z5ayEEDdOQE/HQgnVfIryQKYB8stQTSh++L7A6Hi
fnnwsPjJQ2SynIHMSopYLmrhF02KU9HJ3WVKZ+nUrhCKV9djJvyWE9gZFn3X/nfyIkmo23lpYTgC
rYvCI0W4K/uiiwV05xGsCFhMYz37LiZv5/YMUw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3744)
`protect data_block
6Wo5rjfCVuPcU2g0iGcqP34p7s/KuW0ZmynWdo0NUbOe4m5I6UBm71JQObfl/N6HjzN68KxyjRys
HLuzYukGLpkMzdpygtvUx0ING9I8cRbga/kBx3gm4ajD7CDe8uBpZJmMIkf98X3xHjPVuFLDj5vW
Gyh1I5hDgVdW5g0vmw1vlS//OyH5EN7cv18RAjXDk5tyr4CfRyZt06pVFcd0ydv936WOBvbhwRmn
3BmOo41fMDKxSSLky1ZxloW1b690QHCyvR6nMUcloD3b+PaeTvYKZhMy3tboEahOFXPwS1S3eDem
dz6iwEGoy5dNLpkwMZqLWNgi3nlGZdA6yqzjrMyLPaZylFRrG1PSDGKFqGltggT/VIfFlhj+O7ie
b0mW+jpmTkyOS/V4vge7OcluHvT8WxKhMVQTZkkB+BrvS7CYqCkoNDvERplImtaeDXmMztDxkXg9
fv5nWlM6jLbTzMjndjwuhKWyhIi+8UpumJETl91zRZdC9CDeJDt82NqcBcYBqKxaECvcAS2NxgV+
kGs4gZiCbW/Q4oTZjRUlnCLGia9cjLTGDjHGoUHrOPUoJee+nNtfqbQYkxPPu9mvHpQ+t87hd4um
Pk2lzEEtLiGrXXtR1vAVsgU2E1tmo8z5vPcpZozc+TDyA8bcycU3Qz4yRFCr1woAYQObgJvPUQly
lPupuKk5Td7IoBTzkMjANFgBHlF2kZgqZJ/JM+K3R0iybVjSN34RSEuTbTBtx440qqMXPKvfLeKl
brL7O1L5+FGvzwdV0YJ0WE7vcfOIZcYd0Ub8IxkEDd7L8C+2vEUkgGXnUqhogSX77XsIMSIS4lNW
5ZtPmXFXJx/KhCOJMnf6C3mRVn6ksDCIXSNLb4sXkMgjJ7U9f8BLFBV1t3cqLq1Cqg+qC/SRC8sb
wMc+VsgqMJA9D+mjDdJoDh1lk1304XkftVkiTtSv1yDMsooQs2gyJrIMz0HcAeufGJ3/c65klX+p
AVXu08dR0u0E/f0ZKKcnX4hrkRJL7AiN449HvkTV0vlADPcjz5bl1aI6F8xRuVnyEdxcJZ0sSSjH
M8t47g4jQOVaC6GJ5bv/Rj7t+XqV+Iu3X+rMWy8q/z5wHRqkSdKPx2SeyxLek6if8z5tCMASpWiq
HrtZ5yxD57vpmPysHJ0SzdDRCb1mavbGbGM1KWS4M6nuEhQ6yXm7MasG0guI80uWznvfhu0Uruga
yhee4m94456vkXcrITmGnZRoEE7SJnWWn6o8gARP1Hw+JtQOQB8gvVPfCNJoVqpTWKB5bsTfoaa8
5cydzfFoUtyj7ERkUDAKglvBeneunLkdWG5j4pXOZYpOjLk+sfBeiI8i2YnGz7S/xllcuDIune4b
/tCVn7dtE1w5RxEJ7gxnv4CcgncRDDPGyiv5jLwV2bc7PIaf3CZBakPyQKDBvyVslU9uicPnfl29
mtlB1rRw8jSrATs1mV2s+Axff1tHEscEj2X3r5oXXVPZQZ9LXh/4m7pMcBLKQF18gNEnyWV4W9Yb
Mf+kAyGRhF19X2MqM5yBZAQ5TBC4pI/wcn1RXIwNaHDfizJPavANU9JqVUEyDqKWDrj7T7ucefay
VF1lcfhy3ncR/PkyFXc8bZWS1sNQKpSVHm3qlQB5co0BQzhpSfplXfXh+KTP7P12rw5SE3xIK2HJ
W+ZpNJsPlTF9PrTuS1qvnOJpCw4e1WNT8uvU8jFsIKxcAulJN0i+X1cDWsdd136kp5QFqjkgsMN8
DBupNOVBXKJo3VVuWOkxw3SYicYX+GyWH/mIQPPBneEaxz7WRX2srtMgQpTycbsPjUSNSDZHIfQR
kAPUWzRETvseb+G6GjbxnWoWWcLCDvEi172nvsrxxMlo8FziK1aTILxUaQZXE+PFbmEyzsc61H44
OT9RH4zFXEgb3ziplsiomrK3iZu685ZCyWThhewGz9bzkMCSKq/41Ysud17zXBNUaPMjMfMQhDjQ
w3QwHqFvLeCWS5GiT7k41IpLwzqH59xKqcfVDZVuCWbmwHxo1v+bu86x37NeUSCiAKSDMO0OUwgV
/Ru5cXWQ2uW+KTcYlOKtC8vmEauSrJcdbFKMhJsODjNOaxfgZk36xCEwsECKrW2yENQhwDJOb6kh
AtOjuhVQc+dGgSI12iTQPfB8M598xAsk9HH6Q78PnBeNoFk44ZS0UcO/wRv0cYVB+/3G79nwe2xx
GTTxxrpj8WnGpveFbhGPGA8NkUHg22JtDHqQOfrTljO8NyURreH9hj1QLe/dhyMLNUe+A1Zy9RBy
jumJWl4j77xOOXBm+Lp09Q3pHUAyOa4w+Su5bFoHBud9l4T2zzM/rhvVwHt4qFLvXjRPLSC45zQt
92/eGDRmi0WbBXxKWhTmFnJv3qebVSlIoC+ojZkKOSBVR68aPktvut1QhttfrtYhaHt96QzlQ6oU
rkyWoScfLC0csbjf1/TV1bT6IHK5/4ouejgEt7BE331sHVkVlu9vHw1AoktYL3hKk27t7w3HBFvf
B1APfhAzIxKYoi4IITjPhxB2EgKFFbnwQfr119Cll8U4mkrbt9+H1bLtfS8R2yWR/frsn4IZRg2M
7s0/Gpa/WUnSSzOB6vzj228ybl3qpFjrya0cFooX2F742V2YSILNPoieoO7BwzY+7PA8M76I0gkY
QOeb/vYMc2CwkEfOEAOzlVIQyEK+fe7nFJtwt43DKNt3atjRxbcVuZcuq0Vkqv+oHatSDRTfcSs4
1OL1QZLH+8Fd6OzSo3V1inQIhkxxyexFHf9e5cYHbveivxZe7bzXIK75YW2rQE9qny/EfCka1vYs
Qwi6a9QMvsMvyZx+LE6AlcwN+gXZRfhud8ojMxEocl0PAeP7cf02sKd3y6km3HgJybdvOl+v96y6
UQClVDQKSNLO/gDA6ossGSQuSfPnBXrDGeGk3QTNdrgc+ztMur2sSX5/oaYvpMCimLEfx8EDyrEC
xhsuOtL/KgkRighGYgD9nLHY3kCA70vbAVepLc5YqLpEEF1I8YmMd/Z6+kOcfJkJTtRnYNbny/YR
o/A2qTgv8Y8N5GzREzOyBLAe2mUPribH+xvIrus18rLcn0cNb7fJOVBqKdyz73L+gUQzR0L1Tzjc
m/HSNXt374++7Tpb3tl7P69BYd/0qo5+VcaRU/XdHLWvfoUTVPN3drFx6F5yX4RWHDPlTTWmFaa1
QSauzPRKFVAv43AQTg8pXZmxDnyYvMR8rtA8lQYOeGJNOpJ2yUlb5rFOpHnugWkzvid9fzbTE19m
yK6XUAi72DDZB36pfjlx+SQ/sG2UOqI/sbDKWY5Lh08XOr+mt1xbrYSdORrQwh4wATmd5qzS1nqV
f2XtLtq3fgm0nPI7D+FekavV3/nbMb6dxqVePD0cuqgLFZgKN58tAu+ulxOGBlCpMrruHA+/oAqV
b7iWbajlQ+6gdzjB9aF/R+0FeIwjTfxH0b/DVLUbAxUWTnxtMG2kbI1S7J4UbAgYzAV0aP0v3l4g
yTtdBOicy3OUhAKtJeayRo+AeYTTkud+6eYINQYqxfaP9THYTe4vcaHsnJaFDJ1G65j9ld0oSMMg
BQ760lX8aZM14gOhv3w0LJymYbesphHAqVvVHk3JXHa5LPi5VS2mmhxkeVyxjkb9MjKROV+Afbs2
EbY8yuGVpyZk5jbxlkF4D4aev7C8VSMAoI/+fvJAw3FZsoUa5ezrE2GwgBLcsOr5wqR20rK2CqdR
7SuISiKqRfIM3M9c+FKU4V4AliaGvQpiGI4SqHDvmyrW1d1Vs3ZSykW4mSQARu/dMuE3ovBKRxtM
fqbLnOZkJ1ONnu6xriL1SIRRCTNTwP2lfjjMhorMgvmGmKbYoC4br5wsPgSvLa7QKbmeF07lo87m
CCyRnt/dO51sMM6Klv4B2NLpo7lSbodNJVvkHRP2U+FMeU/MGfpCQBVr6UnIf/tQO0V4PiVqsfj0
d3NTr0EP8n4QFtWX1VFy+F6frkW9FTI6hLXJ0EUj6VafcJdwPfhbu5tLFDDdfH6W+ytX39r4DpFu
fJdJWQapmtAxHjVQKbMnRmBbbT3xkh69zSEdp42/SJ3rsbe86JvLpvQroBXxije08Y1Yhm4tuqOF
fL7OsikGXC44APSD6c6XIqf2QbG1LYIO1X70nhof5EmQY49VwDZJujF6oX33IgRqn4N5B0mX20v9
U8ERx66QOwzETGpN0rF49GlXwX4T1bfKiKjC4RkqCR6nqImAQ+CYXCzjbcczqre2G2iy50z550HD
aw6xkD8CO+iVivXvZ3+DwoU5bZ12/Ze8r5aj6Xj2x9g/qCmk5VZdaqdBEMr8pp2LUvl4dJ+aXVa0
PThZJleDXIWDoG8rp998IWs6qGDikiKDoRQzhnLoXgd2wudw5AHj6B+UoPm7Mbx7y/QtQm1kJ8xS
cx8lqdWySiqdJfq3pbe8L1RwITTqlqd7lCQMKEOTCsptoS0BqR+sI6CPirlh2EOdOmz14D/B41Ty
mNXDQOxMSzms8UNFeLFboeFWbximq1zO+xvJZlgZZm5bY0Li74uLVB1JgE6E6AbqfXc34/ZlAc5W
JgUGetwe4c5/jXBX9wnHHB/okuIs1kSKi3e3kecBAns8L0vf9o1RmXxbfjM4Hqigk0UF3yuNtT7R
n1m08EyfJIIc9OSwggW1rd6Ht2JGgOu0xOWmvNSEzjLrngSc4bQRzF0q7O/BPBzzR+ouWPtfKvdD
mZJ4ZTMuo5Fw7yuS4M5zO+/NaPyiWe9Hsixs6Va/XtBwWNqfpWszInIKNOVZn+y+0H3fVgnhB9wM
rcxsachA2I6v5n5BQm8sxl+3VqiOgZV9FXqR9bXaCoXMofMwXbx2F1PJIZojm6Nt5zjvgj8uP15s
mIwrSWKALWIu6zZJ//RCQLAWdPfl9B6dgTyV4nggubJp5s1s+HpgqGvbAILF6PFEnvlMZ0C4cBef
UJt0lC64jgO91Blyi/+XkoLOuBqzLmSa0o1rr/p9QNfqBa5R3KE5
`protect end_protected
