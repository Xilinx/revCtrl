`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EPdxM3QhbgUN6r8Dgx0n5NBf81Fy0ZBWeZo3Ul/S8oly6CAR1aMUAG3u0HqY/GcYye3r33iDCZGM
zMAJNvvEUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MNeexIWnSmsqqVBUWqYuAxFn1Qgpwlhl+uUjsZlepkzjRg+A4F18S/FvjRGgVbyIyv6Z9xHpJa3a
tlIRultIsdXbKfruxy8+PjIVNeLneCp7igD4bmraD6wRcpRC9QZujV5t539qBv/U+hA45lD6NQie
9hZyMey0axlwfdLia3Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qVjFC8ZO/8qo1YHZMnOkJDD0DZWqL4+t/rbLKxncvRJbBjDhoHF4Gw1ihBQRt+h5YQqw5L5232Ep
H8+Dcn6h4TNoBTlOgTlhS47eBIcgJ7e8l7YMYaSr0KIsCFP01BIB6MJ3jwQ8MV0V5kIO5UhXU56U
6VHYQ02kDgWAFWD5ThTnxYK807VmI56AxUAZY5iGzdBWIowqIWh4B4YtQuPVuU3O4upkPiHO+Qk2
R0GsmMEO38DB6pGo4u9p8S6ETs3bQ3EiiatJBzD4tEILiSGduOPXdVRoEf61ZhjQ/uxo2mhqcQlK
EmaGfhML8dP1l75ebPKN5cY1OKpe/taOhWlDsA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZGvh9vUPHsWNwCKG3TRwMskTk3+hCaHjiqHio21vlP3wCoLJRi1iTTrS/Y0WZWhS3KwhhXZ42XVV
XaHp4U1FmSMk1hVV/Menu4JBOy7kXHLso2bdsfOD//GxhmDvH8TnBk6d/LggoztJdGy/x2CGnkIC
7j2kXohQf/FHKGT8YT8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OHc/Hnhw5G/Ft4Id460f7HViWwiW2C7RsAsbUFzYNpqrIOr+DMMx6euq02Iz2BQkRa+DxdLbZojE
I3s3is5JFUKOYxcHAml7Cn0nQU1445lBTtvQAUdGtADKIeJDOTvwx7zrC2jKhr/qsDzIP3b5t6TA
pInI+gHlsjH46XiGZIFF1MaIt3qPwnWT6Ydq/AUsryp4TNueTJmlU9oZQdIKMn+b30eZQwrsRwRA
UC5Y+zA3eVYdw+2QOU1g2521OFxuC7VaqzOB+3wW9e3HBdEp/EfHj2taeE8UReX2Rn3iZ0B3rf+9
csxMMNr/KsiEOted8iwjbQTSaPBD3lW/EgGXBQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`protect data_block
wrovcHZ5qwQL2M/nAAAAAPTTJL3DAs4mYGP4bETAu4/EzXErvrmLIJJbdiDdU79+/mH9o8cD5wRC
nC/kIqCFEtx0g5ouK5H7vPIw6cpSeFPUAB5WGYyDf3/Rd6VyCFZll4Gn3T3qd3VxMSFI1zW89/AO
7ZdX/BgO2fOvzI0PEQTcVOpnasg+bLIIVoLX1arqL5Dz86V0zTRpeJh8dx4LKqGEx1ZSa5ijA8uk
krzHWFJHgAQr6ICkw530oQmQe+4JLDMBQA1AZThQH1hvCAP+MspDc0rMnrlum+RlotvVo7HsRsu8
EFrlN/9Y40CK7gb8f9a44XboThOg+yXb4QPg5hNZCD5QK/G84OFjU0LqhaIU4pPiJRT4hHYJxOUx
Ua5pARoqJluSBt3NDOJYGVyFu0ay0O1jnAtUow91Dl/67Y7qo0xT8jroEpRXiMVVrbS7igZUg2IV
LFjbXGe+x9ub5u4Kf7QL01ZtSV1wdHkTuTm1Ni+0cBzQpu3cXBJRE/jY5WscTOHmuCotKGc+qhSk
Jyc7CngSEFL10R8W3aZHIYfC5MnDgKE1MfvcHZUyT+AqndBkuECiKll5TJ9cP7pZd1k0Vwcnlb55
rDG3x985WDTTn6u9jLHWCq3V1L0VPTJG67y9vS06uGrBLOrKxS0Mpu0Xlp4SjFZ618lxaJ2XhP1W
Pwd/tTCZMWlP/167S8+voZl6SPgVc1H7zcObFSuRiwEamXU0fiIpxJW9LBU1w17briM8spvx6P+6
AMsCJHiXNA0FcDCglw75D2tYddduDU4lyKyh5upVDBYZmpzye6ozjrfgMaxblaxVlfwL/OFtjsOw
GLdLZIv4RMYZWd6mRjmrgvUQ3lxlZBUrqY2jvu37Y4tOwYUEVnALMnXyH/jxUBog3C2jyaXeA7GX
Ued+uE7dpPJRdajQDrRIbULMyFvWN5B3xM3zAwQRMJqXI8EOscgmLaMdb+ORuILkb69hFqiOUwGC
q1j9nJOv3IEKubG97OgpR8WwJ1sovIsAmOptuUUP2VPG55DX+8ufeoFY1pA3tszwm2T6cW5Bc+TA
nZqEFCG6gzRuPDm0mqmU26RSNTZh5GoFSm9y++3RHI/C6i980IjWCc3u8SDD2ym4VN4S9nBMUgEa
B2/tFBs2MCUlXUg3QpvrLskc8tyWM9Cn4hvuKPOnUmQ2nn9lQRbOzNzb87vR91MHK5odgApGMK25
aRQkzMUJvh+CUdIQ74+fQdc/hli9UCD57IfmZXZdLxq5X3/n9m1j6lvCUWAUncJCy6muoWqw8WPq
mG4jtMjHxF+aeW5wdnIqeCWjJWfID8fpmX7hwHc1RJ6142s1sCEM0YeEWXT0X0qzE1eRrY168bmF
A7AfvabhNZaiZWLuvv/Ar2B/vTjWtoX0NUX7HMjeFa8DB+b9BSwCq/oJRgWNRsw7+AHKS84w1wzy
XpdJID2hj3Y4wVFk5bjqQCfLXTYVrY+NRPu1G0CSeTMUZ0TgKNQDfZl26ZPnsGOXLxNYWT9fQnme
ye8FzLt4IxDouLxRMZ6WWEbFpdpn0QQNzLNVlliSDaeWYiExW4Q3DnkG6t9Xoiv6YHMktXAY4xz3
JYbzt/NOFiR93/Tn4c+FcxPHktfZXR1P67pS+/hpvQ5SpgY7SDMxkpKREpEw0JhcBLm6Yu3+Qy5m
jUwraIlFNLJbShXwGtJSVrC1twgUQIpQHzcHziDdDG5Ixg5fiZlNu/Ol6ngKB07AkFQFErqiaGhh
K13Q24DQnx7BcSqUUQmDrqGYPe/Y+EXiJ9M3wjDTXTIk1rKn/J1B31joqSYZZHoshp6bW5R/bmEF
OEypiqn95HhDWML27dyjsUjBPo3Z22hX17pUBj4M+X29ZsEl0V4FL99twSv+Nz+NiT1D9We1Mrhw
wEOoAWcgP9QWzkfCffioZ42MI/aEolJWG15jgXGTHFtryugZxxo4n1/9PCqmy2KwJLT9bO+7K0+M
iLCUWJo7rEk289cQKzQpFN4SM6vgxT+1t8AlkDYUJ4ADPSg9DqinuCfklbv9g498LpK5yGvNu+ux
2HoWwiODu050U4bjAt1ohH4JLdxOfuZOeetsvnYL7ewSkYD2TsROvXNwmhUlgJGe5TU7C/gtKh21
6IskZDSpCYTy51MOIGC9C86AfJM9qkHGUvmLBWCA+XtM+zoXsjERKkouCSgxIfwvuEof7bn22aWs
thDx2OxF4w+G8Kl8EOL2HwRQFLqjP5JQ/1OTL1EhFo0BqtCo3rcXUVDzDxDSiW5JGQgW+LWT1rn6
Fj5P6JBjME5MZVMflQSLYQpKa5H5ynXFhvxZz69jsiIRfbv4TRt4ppYAK9wFcH8uzSHmGCCbRGc0
g8ow2shlsKsPmyOTBq/pzoSJ3T9H8foD6gWBMqCly1uY/ZP4Ls+YF5+ZCflqe94GQYjqfJEikpz1
xpesdWqyEMcc/S7ueiqboTAd/00ZIKbQ4kPqufIq3+McOmBtWjp1gXdvFuPTo2icSXI3hPm2qyfp
WyP6i7HNfHMtX76HraM9Mn/WxGPiVgtqQngoE9Csnb5gvtVTmqahgoXzlC6gRFHMaCvrpCfLATG1
z4wDRDqJvz1vdGAH2kJ4Iam0chocdkYy18n75jkQkVL3h9dJYDjBG+pAL0ODGppNeYWcZi9dxeuK
6tUlBCBQZC3FZjCOtto3ZaqGT7Kv8LAaAgEVcoJh7pT67s++YLqmdxv+Aom05pMAInj2mRKhYS3Z
RqosVqlB3rDoxsdfBQhdPZhqJQzRk4LAw3h6Rh5Ezks5j6FPhI+rmq229MeoxuBE0C5XYjjzWwQj
KbDtuNInUnUIZkvNLYzVaYq7NTnoHtrAdiNwyRIZTt3Y98mQsJCcupLzLcyyRCbizGMLe+3vpIcf
fAkVgbCVPtrTuhwY6jA9T59tRfR27UNxoJ8xYLfL2+L+yGqbxqlQapOF0HE+wAuCPGwd0beECZ3D
KmcgaEWrKKpsqBBugei8avyTGzy09LvsqVV0Eb/8giBicjA///EKecWMfi6wSSKwgp62YoIb3fZ8
KJpnj/kxLKLLj49/jjGZCsr4yO6phO1ubXoct7AkL2XY715EELRSkpBhYmTfCfjcMtlH+MxsW5R9
R17AR7mt08PjlbT/j8VMVMFU87hIV4vQvQRfgujjLSdTYchy1dCg2cfQV1/Q0Ad1OuAjv2roEZJE
lEWfwRBSTDASON1SEI7tTCP5cWQl9fC//jOg6/RlY8fZYMheIhgcOcL8K/1lRctvDj9J1pFCABVt
Wftbccd81EGOriXuOL8ojoYa6/DGUmFp8inZKnxYQvzRdsW1zNKqbowGSgv3rUb1zZfjfBz1VDRO
uqNf2Ssgvn4rkR9D9t2px5m4VTXGzk+X1vfEcx3Gf33CkXEcryvRGbnT+b85NXTYPs2GPsqRiJGT
E2+DFF0hmpMUVV59vXnvDQApuk4gTUkkZXFSbkOhuEStboC+xhtxmETkDygKcPkoUKQs0Tq3K6pw
mMHV78nW4jBsTHM7h9z2nrUTBtT7ACkNTOos04MOqb9AqAf5CrjrpdSRh+nONe/bOOViZeazNmnc
mcjUJwVKJrpsrozxqsCnyGU1I7UPkiElJY66SfaxF8Z+Uax3eQuVEWfuuB0h7DFSSdTfc4NsjHQM
xPw2Y6dpEpNmt0zPil45I+y7kQ989NyaazMxyPvkDimrHekuA/pYkX0BApmUkxWnh67grNeveRi4
LsA94HsFBUydQ3ArdZqywPvxexNAESGgTx5yR85pbO+HjSrTqLkgDIUIvA7WD8wA23HfuXWbGacC
IQlVC0P6Xi1iT84CVt8vrBwVEYuBeF5ptdoR7VBtJn9mf/lBXbYiGEuKD2oGjki81xRUXp2x/nvg
Ho9C0r1gRNIxqfSTHfc34XsL9FH7kc2h1kMZSI4si6xInlwMTAQoL9creToemYwkxbd2b7JRWxt2
VKILCjCZ8mrI1WBKKdp/f+tAnr5w5b0tjSh2JuHb90Sffe2RxjpGqqOD9uCHD3LWqRiSpcgcgZdH
KUSGw6N0PyAuozh36ZRnXfB1pt8T2sO6JileoixFzBU2nfN9UGTwZr8tRk+XcfNVEzMoYWjvokXa
Un5OjZdvn0BKQ5RQHDJZxDMoN7dch1vl19l5/8IFCrgozyYjGHl1Fb7W2pxQKpcX6a/YM0R6ytgl
gbbUndvdQjX2HJ9f2TLbMM+REdJ2CYaEvIwe2MFTfZjiBkYTlhX2Vr2g1F6m1K8nk5828gwVCxEy
Ng23XByzsxh3bG2VXODS/2Eh+HxFsV8CiAUqBulCnvWra2+d8X+453ZDUQcMs4mYf/wfo1alKYFT
qfjLZesyDYiUBhcQhhx1CbYBv9x9mYSZN7htNeFiA9eTxUjB/8hYr/5B5/jwAg1e2SEUTR8JZgPy
yK0S7Xc52guaWRwY9Id2joWXkJdolINgfEwu0mkOIBTfRVCgudb3+SDbPxhrF5hmjYyHFc8KeVQ+
PGHCTelw3tgkFBOkbFO4YNfWtF1XEn5lCDX3cKcprPqw7LM2KbosE1FqJmyAdJ5YAuPHlElIXmMP
PZl/TtehCXLzE7weTcBzZPrZIYxaqa+ZKP4BexuIfcmYgCsvKDMHv7KTdjU5R071oo7Occ1c8Gj/
ZFq0/pwtobOqVOwPI9QhfgfTvBivHjnW3/gBTzJ676gVILsKEZXmi2q8b3oGDUZOTTz55gFr0BgS
qpVxpzPHYvxA8//wQHKSYBY7lEyTj76Rxu+7qSZjY33F50tFCAkonS9w5VR4aM411qklcycx4ZaU
4YfYaZhnHTnXHjilyddl80yzEQjvetv5ViiL25WjF5mnfdzaMFOm/dsgczT1ueuZLlEqgbLp/S5G
AbKwNzSb37IHE9a/W4WiC+C9PrOju9MD1DetfH3wQw/nFC+rpqygHMhRpYFa2aU8sPkbn5HTX2s9
2fVOJgcsQ08l0ZVak3hdA/HHABfN6A8P9JRKkEH9OOSVTTyhtNs83Nmib3EPrLMmvfDIYVT2Hxg+
tvFkZarf1uU8MS1KoY7bCMgArSj+GLSzJivXoG3ZWQrFUIkcisA/hBg1HD4DC+Q5QQVmGUcvKIYU
ohOYrCaGw9hO1904jCXXJNBrUKZNOYUE4cyReczq78FZMweMaMV4p1cwxIHkFEIPqK0wCAUtoPeA
5zrNxSZH3kd5XyrHd++9VGLfSG1f+GVGH8Cq+kQgGyNxuWonR64EHhVoAWsSNJqC9iP/ACHd5Te1
nA/sEhpv/oD7KeqcSUJLszcZ0I7YhzxIPzN0vyOltsMpCUDYOhqqgkgK6pqMv8LBfoObaTv0CVeM
xHUXMwguOrLWDgcFhT1I9LwzTtQzhg+fMxdLcuiv0BsBtQXNS1bhIFdht9+wsrtY637He1/91iLO
FOop5er7DkljlOTb3SgoLOe60GTfFCx0Fe+uTOWf+zc3LE7TXiFnUUv+Gl+2uS5Ui0Qe1NmZgcdu
qACmufDZyTIt1d01LqJb15M4zQnPA/Vt+5K+Dmp+6KE7Y9F0y8I1C5irajs1DSvfBdPd32oWxrX7
p8GwWZlhgXNqfXmFrpaCySNMToYOCVaDrzo+MXXoJ9ZUWy5DRu5FCfLyLbEu9ArdhO3VLldH3V32
1icmAWK04d50dbT7iECImvXGe9dKnA4muYrhHh2ntZnzqxhfLJo6aX0VVUMhgyEsZJwA/KlDhtCq
wtetUkXIXYYR7IVTIK/jwJR4jArF9IQAk331NXpdbzQ8fvk3Bgw8IdRJu1WShEyHlaQHWIkfrcva
+VhLSpbe5VtqkXgR07DTvhnBCX78lxLYiqiPYuWWwXK3wGJ/unGwjH2C5LFjSPjRN1SNQL1b0vT8
e/ajga2Dg7JPbzA5Gv35ewnvlcDL881v6ozjgC9X+ox1lY/6zHPXAiJfsaDkzVko8VDtwlwX7ill
PoqW1jnezQ7zy0zpVA+c4NKDGsCUbkyUQL2HqFBoDmEV0kv16EcVbguaC8i/KEF9Zo9bprT2sbWT
Qs+m3sz7+eiKehiaXU6CEu/ZPNRYaqelTMGJXIwbVkH6FGlH1XpFVOoDmp9BHwIgHfcrnAqkLfeF
YDH01e1qYTYLCyQ5SJBsHSHVL4p3vPl7UH2tq1qvJri0JHuaHkqQNmnBQH447UL7+OlBm6y/vHO8
hS8Tbg6jXcjaZSVZ3k1wJSKJxsZQq2V3NMJk9wwO9H9u7BCoqXVdae2GtvAWo40nZ5G7B71fahcC
cwhB5zVeKItuP/royyh2lv91pQdRJSHwexUqtbDyOlOGhvMqHMbuflPohUGqB8cFd2OT+ZnJjRUB
TbmzbLgGrWaVIxDNMyZ0EsdJ9J9P9o72gHpRSIz+cwRRHLhVdTqspAk9XeMZOy1ujtZrkoY9Dblg
axMBtavG5ldop2YJ/OESLEODfj2MYNJiONxdOZ6nLGkP9vlMCFg+lP+Pd7XY4EXYmu432CLWHdKN
eWqbh055BonlRw9WFNr7O5cpc8P68tdR9UbACLuM/Z3rNs4B15U7+t1mQ/M6rVmAgmOtK2IRXGN9
od+6/gS+2kSx0frWuYRm6phULg+JUschD2pei593Zah2YXl5mKbOE48yllmQI1iPPWxM4xV+p2+6
Q0iP0DsK1n2i2hTWb1+JUu7C2vbaBNVy+PbgVJxAr+h1K3pmDN85O1gODNv/LHyLvZVp14T0To4V
sSxDF2HLFsrKaBJ7taCGEF5KcRzPdLUyEbPEc5aXHboJeRnc7SE2tyeAZtbu//YulJR3nTTT3jbj
UaOdPwuKLlBSeOu/20GJyTaoHIaqmyYOFCJZe5AJzccCUTd6WPIYIn8lL7LMHSlvm7Mb7YRIPQQ5
k8Dhw6RCX5h628bVoeJiYs7at9jAFEZJlO29i7DtwWH49n9d5TWAT5DTCES1dU193r488lj8u66L
1/D+x4cMZCW4BRRjPYFsrnCP6iWkMR4Oy4xMfIO7SCqOamsXHJfTLE+XeoWFJz6BOg20qpwROEro
0mY9oA==
`protect end_protected
