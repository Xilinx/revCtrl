`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ww1cFCaKpEaygJUT+P6Z2OD0uzJ4IJG8iyHDm5UNlVWbTWS9KXjZ9jEg11wJmlv8lA2AVebHxIas
7nZJsy/GjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gy0/aj7fr+HoqiF2MKC2DdMRffpsNgkz3LCA0LoXsy3oP+ExvEwYs55sO8KAxVdJaUPMOFr+w6Gi
VDRBmTTzMTTD1KvHQEhDppUtYnGyL/2qAWb6xHvmSHDtiAjlHews7qZ26fM0sYgNx48H6LSqgFd4
hai7P1C8/gEiLdaec30=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hi2M/LxF9qgAZzAUuc501Ws9I83yzxDz1ea90Q5QjM7jLsFrH4fLD2d0WWY2wDTdG0Ih+QNnE4S7
Oq9DybBH0zvBRUhAQoExlvdlIfU3Jr1YKpM3lLPQTLIhhCp1eQgIZljQtMN1p0u0HDYYsZO5DBeb
LZHGhmPHPWGqNQ/iLmQ+PQu0B5Cb+1VKyvK7Ipxjf6wKC/NZlztCmWzwV4WC+jY2wHB2IofyzZfo
xRBIRCIpTb+tTiKgZ9oAjPNYVjgXC51YW/c8ZhnzF0gIdh/tD6GDSX/DdrrBN7Oz/gtduYw5jR0b
WsJx7lVGCa/mgRPb2+p2mjuutW8gGGnh6+Yo4A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X16goI57idQ5Yk2jq4rj0BhsplRtdzoYr8oOU2lBTTonp1Nx4fK7AS7KgGuzY4UqvPTHmPTfD5ww
0YcXmh8hr2Hk6aIz+aWFV8C8XcReGDrBhi5Np0Vi5hozuTfEPpWuDV7kTmarku7FYKZbPt+lsAsd
f8+cIo7ySKaxPnzoHbw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RA9GWDJZOdw/NASVbYOgehelK35X4QCDpOGKLkbLHbvCU34C5eqCOlazH25KMTrAHxM2lx7+fAsw
HHb2ZWqK4pB4ww23gPcOsgxVCyXs7Dx/H6E84snPbj5EBFAp1p9GZJoguz0skOVQzCSeso4vwekP
kvLqf3Ypkz4/BbGmeIV5O3MvxWppwuIHCb+NDzDYU2x9uQ7mLUtu7pYCzPfN1FeLiv9ttZaXRuYJ
ADExpcAMpFzH3bwg6Tm6wL+J1DzA4jLGZxI9jxK+L6xNTv2NtONryX7sLla9heWPJCSHR4TT8ow3
t3QklA4V7oRFEhlMh0Nv7QVOAHjukKSZ99LumA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15200)
`protect data_block
2JEuFaTgqghMsv5lmjCzRKFTRu9v2Bd7cfnnEymmK1IpMPqqHVgKVztK8UcvkN/cLu6meLkuW+GH
jEF+IasLsTsQoEbARf7iGoWy/qxr/Wx8iI4qK11niwKvKRzj3E/VIfcoFWMI7lDjskoNrB5ON374
xdQdL472o5haNrGgEzQCs124gMoZrq6ZZftrvXJyyhHqGqmNNfQbG065CYcPsuRjXxzPltG3oMhc
7n7pQE9F5O4ObyVFgYrFINih1IyuB6ga3CPJSEZRwp7Gz0bxN4RD0DBaR3vYvY1rH6jZ2As9bin/
g6/KlClzLL3bvhOhbtjv1RatU87XN/IDxll7fS7a6mxwPnreBchXZdZeSVFJoUuxMvWbt3k3R1rd
B9CvCxo59dW1xnCS5XechQ3z+loSZT+XAB6bgElF1vNiQhQ7+3FhiU1vghuePbB1lF1EME717a3W
lR7is8iMzVt4i6CAFM/ak25Cz13n7Lim4rIQv+29vAPUjo6Js34mFrwFNI3sA5s7vuMTa37UMCtg
yXuYGXLv4X102Eg8ZA4mxr2nhAQAEulmX9O/n55/bFxHqebXDbOa2NsSCrcZrxrKTpFMDrNs87iP
Uk0ayFDxNOEVKOgMGPx6q/guu1O0dKrZpPsQZKa+Av0gFD8aC9QTanCthuHe/7c3WUeurt4ZY5+z
0pGgd+5Ce3kcYAfXPPtApct+1NUh/7LlLdp5FZ9j1t7Ub1XiqffB/0q0nQ1en4x+h26VyzprAlWR
3scBEBJifrobgdGE1mxf3wHE9l3B1ShvvX75UpBOiN7vrUnzYb2wuEYx5hbHroeopq1uhhOmYoGy
eQ3cFZUSf+OwSNq4UZzs79Bzdu6LMLzqogJiwqFgNk7WLx40RHuKspJuflqyIbu2jFP7yWJvPIcl
4S7sk67ZTK81UYIJiDjs/HBnQsNIFvL7cXWybaKPE/oJFdKxM8bZ4rwc+6n7KWvHKdrCc0H8B+3N
X5cT660ZX2hkH0mJgQzLMv2fNitvEaOIbbAo0J6wRjk2czalj7kb00MGlgwTYkgioM5E6g0YDzhY
nUqkFP2cGPhxQVLgMEWjgAwd6Y86Dw13gb7Svj2c0jRL2zb/SjoGGFmI3Q0S5BTKgrItxV5zHJo/
8WPp3xzZvrP+poAsm8s1/YxyzsQtdwWkqE/jC3u6RQa9foWb3oYWqn6kcMUePsne7Jmq78LRIfDg
WLDUGIHzOCxPvJUF6GnHMfi12Y1p8B++LN2geJoIyBWbjusxENGUlr1mbYIEi86OPls6PsLhpFGZ
rl4WSyOq/zZ267s1s/MK77IhTLYHd0ak+pM4UpcL5h6P6woBPduUN92Vji3TIEvS2FFRZ90DIukV
UiV8e8CMhL4NVEBgAi0yGriph9hUMoVBXECco0RuYspTe/jqKBF/TFm1Z+RIqaWAWBi3vZ4o9rWQ
JkWneD5BIrREJHhNEa7uWlHdrrJzPcqxn71MiDaGu9Bn+3yPgl+KopwXQTT2A7dk7bABW/Atm0Y5
MzD0kyHhfYtsDlO+gemcpumvYI+e00PKC2MYyz61Z6209Z1T1kGbTFYiRfBrVqGopE56kpSN/Xdt
Jagkh81haf12WOv1gvfMLiGHGrBSMH24gzGN9MvlUJZRDxSoJ1X5oqOOnINQ1zoO9DFtfaJMPjhE
3dWhc9E3BOUjesf8jFLvqHLyx6pn660hYxU41ja8W2VLhz023k0J+6x3UwRl/SAbsmm7Egfz96+z
DPL+V8QgrQ7O92+nI97kLhVgJ+WGfRtvZujruzMii+RVvtVOyhS1pFGxjpyIJHcAG3GBrFhCIGw/
ALJJvQDZgr3A8QNf49eTGxbmJHijh1DjjJiAEnUyIaOc0sjQ/TEmyc45guPXeMWrv/tftIiipjMs
Nq6MXKfChnOXy/XoBSq3p4/WVBwOOxup5HdrSXeGhM09QaI9t4ON6UTAaM89OPAsqx32EdtTYTHU
r3YaSWklJhY+UfHpvH2v+6Nw/ZsXtrNdFvItUg7SBlkjdT+cQuXjuHoy0XbuxvSwPONKz1SvgnIV
7DMHV9R/keVEmzkpWxhPKEWY+w0JY/YlqgYYlyPraGEuCxQOl4FQT/mTtEL19ocvC9IjgY732tA3
t9SXlB4pBPklFoGtr4NQHjeB6ke2a1lrKBw1ycBqRAD+0P11h40xOI1C2eSINmSFaNVEtPkClyLw
BSY8Hpuw2kAIx4IfNXiAGoRN3EsRgYVj7ZbFeNJ8ZRH7TYNMirLgM0pbu/t8nhK9mX7UoTM/XFBj
SbeAPw3uKevtgWcYM6L30rEsTBiyf5oyrOM/TujWwMC3NJSk3rpt3OBQ9y1ALmLo+/wRgnZ8zAm2
1W4/q0UigF/95/Iei8n9htMLyrzh6uzJodp5gETDcfOhz1uS+qj2MKHFQ5ICtGw0J6FYvCmaPYIT
FInGicSA26dEXXMcU7uECuyBP31PnZNQZ+wVNUcUkSILTHiJXirRwOlENbJy2TQd258Q+6tybye1
aNJc+qAXcRkDFkGddojOcdFPnpwsA/Ocyxo4+e03/DwQw0IePUOSWTNUjERVfm+rhDghkLdobZCT
cIz1izlsOkjqBImJDyrH16/LCXZGwDLaOfil15wZguyPzS9nCbVupDmqael8cq/1uEvI9WxUQmb/
FmwfUY2mK/mmf7DFDLd2U60GVU62uzP1MJny08RkThFjg84CnAAckg0X7v6Tuin/QP0RnOstqRib
ftVBNa31tCE4xi1MFL51QblHD7FdG+004NuGCiznYObZKM2FNWWU+VjMBsCgffYDXt4Q9KjFmqk3
xOJ1xtBXsLrmpjS3u2nDuy7T1kltzJaIJp5NcQMEsxtkt874Fp0BlNsPifFu0hA7bL9c5E3omnbv
I99dHshflytsZatBSEL/bSBUZJA7CZa7Dg7ul0qwKQ3umpxntKN3acXp5DYvSFtf6FRJmX6A9Ud6
YXD2OrGOI1+HaTcNQ9H7saDkNFyivJwvfHIZ+NU5zR04RVSMqWDNAAPMUvKehVUsdLULHPfNglqw
x2pyOawGAoxIFasYE39lF4lEsD32kEkZMqsqKsybCbPA9FJzQeYaPO2eh2Xz7T3gBS9XGQUdh91V
ozxszqAKz8olo6w4AG90gED49McA/js4mw5NgVJuNfVZmEJjTVtllqGXnFlGuu9piCfsypK8M+26
yJWQld6zrQO3dY3n28XxIQIXtk+ncYCmr7Xdfgf8tlHED/njLGw7gRngRLTGpGzMCYVgRJTwSBLZ
fUd4qFp6KXfjoJNCSoYWr3wpcCbUYQ9+MQZ/G38nrhEUxLn/sydvY+f8Df2VPsHJKPIUh7lEILnr
j5jahYx88uAW3BWjInqMPtAKEuydQC1jB0/k6iNma7PKDVcRQGbNSRrO1MTKyolMknRmyOcFE0ch
cw7MpDLSM6DmoZPEJ9prYB0W9CENxuzIgPq5WaMi74LWj5aEiT6Ncq7gVyE/ATchYId8urwEsGGV
b1GmG0kcLaVzYeWC5J5uD6EnQgtV96AM0/ZTamqyCqsUoz06NBfq3dvrM7urkBeBelRi6ziuWnPS
M7pvp47cbFhkVGZEbsf0GJDI0fUXtVbQaoypK2cshK/3vCjBYrV6KnuG/EPqUlpasOkbVxON4Gw9
DYBOJSLY1Ji9KmHhVs/s3fhgUmPQheHQGUjELRrDuJr+TbUl4gp8OANr3lNrPzCCQmoyCTJ3lAEp
PbIesc1EvMcuqze16fEKzpCAJstThqQz0fcxRRNC911pyazizAJhTdgIGVM6uFheZpDO1YSrRX8R
wLC71/dNkwUEJWHeJxH488bA118Jj59tdzdZiDGnftKZGbx71oT9scKOpc2d0YheBl842dekSqyU
88s5qMEdwu9IhBLsryVPb28HwfhTDug/mL9F/Rcm4tNIsaOFf2xRVYROoFHG3209Scc4/sW/4oBo
ZIYQ4TaAER/6KDQ5Z6XblHpU04ZwDIopmkBDOSxcPLASJTHeUqtLelY3+GLAPw2NbNsba27sBskH
oPpdhVNpId3f6i3xDq7z8YuJiBHaVO8inhazu8xq8OVNeDaLKEBHWWSim9QE2DWGuC/JocNHrwUp
Kan9p4bltC4ckvUjou7/DoT7iFd2OWW1KUpfkmHX3zn2kkMtat7r8UXyJRqYWnBsaP7zUZ+bP8mV
RbNTmFQpR17d0980hACtr0uDxPq/Bw6Kcp3W0PKG38ZOyDcjGkSaQkVtKS/XsCvEO8W0YCnetlVJ
upIoNch5d6eNW01hzFdl5y1yKNQN9wZqw1FsAcCh6qds90TfoXd08cgfqYmTHzVl3mocarK2vrun
7J2NezeeyeOwvHn5E4Ms3KAikzz5VQakLhSAiYtOHdSe9J3i0IsRn2qQLtdpW+pSXBaZlrc1yuVV
8fRokvZxfHXz0z+gwp4vGiSr/2PVhTiqJRE3/MT2j2tuBYN1mbH+ag+iqKbwp428/jxc6gRbdTyM
TepebTNi796iOc9xA0bJO2G3dKgdXeAnbut9GWLULKmtwr1YdOBvOh9lWismln8g5mFk6SN6r4lE
3crGvroJ+8xmhRrpAPgU7zHYeG29zWeUqFIgoxGONCJITGnYC80oBwFj9PH3Y1QqIC7isVAiiell
uCVm66XggkxarHqcMuTJzLhFe2ureafGI/dLq/KEH8NXkZUYzr4kq1W6jY9Gkj/8AjUjLm5jqMAa
IZ34xtIejOq31JDCIAxxpuR54R4+KSbiPdlHSA8QTxzssWBL3W5tMITFxMF+0KgmcT/r6Qvj9Tsk
HFaUyWIpPVtZ3z+/WgGB31KwHN6Tm+CMcP8ST3WEX+Lstz5CchUPnl+xSthhgTJGXK0PK5lQngMB
r4OiGGT2J1/1OEBo8JYs0z6fGsaazGLXE43tdRiETEPLJkfTkGu3K/mICZ3hiMyxiouN9KekTL9A
xwFHCkzJppKxXdLl3jqK/1BmU/tP27WOleLOQe40q7A7cFjG+UyTBwukFPx/SorSTvdUibN3s+Jt
+C/pxcfOEIbvvUbolT2RahpbrIjv9xnEpNfKQwt76QLD4ZjRYfOkGGsyT7OxJ6xFdQYhlQxeLLwp
9CDS5+GyLMCGL2ezWt+YXjw9o5uat9v0YSddKnh5yDxqhTWB9f9A0zV2PfmZxE9+uhDLJf7nFHDm
ZUQQYolYngmh2KC/lT+c0Kfv3DbOt6hIn5Z13E+2NZI8bq9GwL8IBLktcQ5z0wdqAHFuUufPu6yP
zoRY1CmLB3eL0V3ArV44SR1rxrQgBPXJ5WUYXjc3kbkS5OOMv6MeIWFRhO4C5kkiT3sLPZkaR+vr
yjmnOJ6M8qFGCURrJfy1SCJO+3pJq49rg3AGgKu99o0nY3xcu+LnaRRsvmHIJC00ydanrf/cOI5F
/ladtDtIZMaEGFJ4uA34K12mQUna4FFMaKNsjAflNFMH2dc40CMbuadIxCiM+8/yHbuGpaCtMXXH
/olbLTXVHe8uP90vA6KDvZrDXQZJaKTT4IdbHjj12f0tAEk2ekONuqhofWtfukqT3V2fgPXYJhFb
+/FYq1T6xpAiC1yuawE9G/zWfj615HoSC+n1hEk5qpVOayW75ufiuAapK+5HFnypzuICEwYjUyPT
YTqckVvXyak44j/P/iVBOIggjD/kYngFhTKJGzog/CX9hSzuFA7SHhXWDIFLUiAFc23KDN1KQ1ct
+0Y9rOfig15+CeJViE9VolHZ7zE5/Ms6HeO7taPV2DwlCWZKbquwEjwtK6Ksg/wBWZT9v/RuwA3K
RJJiGvi8yC4pXjWZDCkBMkB92CmAGSs4/LmcjWcOwVui4rzFoQZV/l2nnF06d9wtEQ99ay3Nxg9p
BMCb4tKungTYu2JKeY8ValQWC/TR21xEySzpti8dAec82Edt2K1sCvg/ogBWrGYbbU4rtwWKhqo8
DHYQi6mMW3imPIbEKNVm/NSO8zvyJjX6di5jF6ml2T3wyvBrWMR/fBnlURxNi/d1zrzCnXsXUw8a
iOtTX9JYv/iNYGgUXL3F4UfRbLk3QM7G8zU4/2EKzsK/m8nnepiLJBl8S11WC9pAZOmYxBG7KiF7
IiIIqBZ9nrE8VikMBaTxCVLsgEFOPr6NjWbeRWBQwHzIi4NEnZXtsb4H7eQolBMRauRNkGS+ypAQ
FkOPYRIVGCMfZ6FBxZrhLJRpQk3oh52tkKG9FTymF0btUw9Re6pGofB2SAEZwiPK04Ou6Sudl+FL
E+CiJJ4+JTfjzVeQ0BuNTCKGKSNkeFlI6zfiOtJoHUcVVdLdM5mf8VtVK+GmPUYOzKq8qMxBVLZZ
uaylLeAiuoUSAH8mgiEv3qoHxvzEdXcauQqpbiYTN/qKfTQiVD6D8C2urOT2FFoyvZ+mNn2siR/u
+8VEGZnRJ0KJgbfYYK6BhFXh51lT0bsVd9bkhubpdYdcWkJuLdLqU8IqlQHTVItqA4T/ssYUNOz2
9l8EJyOjv7nph9/KZHD7LDf0LkB0WZpcsEEnaSxQtM2eeiLavAdW2d86eYaWHBTewmU/4c/Wiq6P
yu/GpeK3eiIZz8XP0er0dyEdhRLohWkwVI/gorQY3fD/MR/duHMuiTggwrkZ+G5wAEjTaBdFDwvP
C6qR/riYxGfoq7jKq/IP/hhRurMg45A+P2/MIgm8E2zuPKl6G4M1/363Tt4XtzDZJ5pmfp3LidFH
UFWS4sqhUQKESTbHOVZCv2RItwXBhIr/8Gc9VyT0HhCQn3n7oz/mIQCA4DBeWyT3a6WPetoQz1fn
abfcgYhiW1aHEqBPGfgY+BteTaf2r1cZXGuvdY/0ZTGs/kl9fwiMWWwTgtnyfN1JWWuaBBUifk5P
He7ySIZjar00s79nRFQMGhp08xM5ZYDdjJfzAgDKS4eJoR5278o7LU+VyXW+vbVoFcc8YF6JYa3O
/Efft/6OMWRt+yDlWQKGjpU2wE4fgLyBRACTPkKpfnt8ci1vmj+i1p1A1N1nS0Tb2E3bChxTkOI2
r+qB1TJ/E9SsvhbxqtrZVerzcWxoeF4btCpZjKCI3Ul1qEgvEP9WNEtqzbSidMMQg2v4c+gA/tv+
giM3ZP40tMCdyGGuWSKbR/uAY76vHi8CAd3dluXxeYnYfZuF0l08U56lvkf9R0oRbVeVVryp7uXv
Rzt0oz0CUh2D3aFj00e66AWdOgJOkH6oNcvjMBAYeB3tr7w4pGmOgED17fGt5pz46A7AqYiaApP8
CbPL3OHUuj+O/LPa9+dv7KFK1Bzo+EhQorXwG51DJlhraXS5ZU+Xji3pq6FjGi263j9D2ElysyyC
34v7nC5A5ZU6k7oQiQ92UnIOAtgxELlmtdwj73hVS6fyroyTtfoCeAJqGfZZGmnOOo1B+bxJte1X
d4gE9dVPdgvMA9bSv89NF3x37eGUMYiFS6YGw30VVr3Bgvdbb0/gmyEI84LjHCCmUyqUhrlQHMA/
p7VtUeWQiDGhQ3snlNcF3LCFWEVlmWN4LcUEwNsPKgNkXkxnZs23NS1vOg1I/TiNifNYDgCdy6JB
kFIKZgMK49N8y2BidVfW8qv6YGYycSaFIlcjb0cplad8kwI282KIqeY7t5lwzpQYlEbNB+f152qN
7qITMzj4NGAUNN7xHo1PbEmA+NtSbZxmwNNVHlJfhgdOuM7+FZw9G3X8jcNZTHdJ/qPTT9j72+Al
t2Az3pp2GYxjJVrdbj1zNuA4ayi2yuIPcWqmOlie7ERCdvWjE+eDGQ+ie8XB//Xt9d/nxwr0maBH
RLAUkT8j1ojpsIClQw63T95K+sQINkO/t1qr8Daq5FukPZBk0pBGaAfWvlwwx/A3tL5o1CbxTYsh
FGmT1AaK1IqLCz+0+QOK4t7bt8TcVjNEFEO9r9yzKVphQUORE5L8wyeMIdmUlatZCHvxNqk4toxS
+atpIVh8jHs0b0fCySj8l6WbPfdZPKY1iFvIkDa9W/VPksTNXMiuEKyARu249S1Ef56Pn19yIIHn
LmoJEbhpOIlqkI4/ypKiM8xD/5a1F43aQ2E+oQIxi8J6ak7xW6HhOEBQMV87XuAvckcSKxUAoIsi
uX3xcbqsBaRTcvIP/EO7bNKVlvty34Ksz1TArWCNy8gTk3UH8jBySMrtqYBein7EifFeCXNEKGbC
0Fa+DMg8qo8LIeL+P9wvA7dEXFAcS4E98xvEZrngFVZO5z8Ru9DySUEuus9aOqnLKyBYvN+c9dS7
mlFeyoMytqkWaEoGreHoVDTiynxAj1uzMQOLkoTLPph4LbSAWS62NduXznFrrnZx+fllbfBvY80b
D9zTLe7Ao4RB6pAUP9efcgg/hYntObhJ7kXjRQzX/IGnO6/rExY/QIC+rEwZfblFoOfihI3t77sT
RcuuNufAgixVodRlWK7+cE0VcPi46NkpSZnz9gpaOi3ZvX2HXPIFuz+slN0JR1+yEApCkXF1fkMf
gXfaox2/baUMwpAm9+q89m4ktjYhZxPRXuju9TuuKQqyRfIly2eVm+gEjzhLG1A2BjUgv0qwZKRG
cBjWk2EIYCpVcyzIsAnsS3nkXjKRf2actBjmp1PyvlF92CTSlS0g09/rufWegNPO0kmU2FjX4t88
Shf/SuCsoNokUN/X4VROIPhU8Nrjn0hfLAi24H9B2BUiofPuNgELcdFyqEAzi+F0hZlMerpJ5IJO
z969yOqpIxnZsYnepqaXigjOqwGiijf0EYW07igfGinAybXmojBdTN/CETc+n9hhEPQx43YZlS35
ODA0f+0NNkpI2j0JWuMZFBzt2DGCKbNEcZqZyY+1UDViJWUkFuqwqKnkiooH7Of9NaAYKL+1gucS
ebnFQjkX52TDonJmALDYLoDvVedOqQTro9aP4GsdI+s+GqLwXFkD16CDVQPBdDranyYSegSHJ7sg
ZRFJEAfh5BeSXtAlxENLwVZif1pN9TeUkW5AcjbxFbbAqIHPgPvmH52yc8bKAelCFuOsKHtT8JGw
fhhnDuo6EfEv++fTL93ueSo4+TgsodTrjX2dGsZESZHm+JdavDGckuVlqD/9yT7gXkRgMDSDgsGK
FX32PAZWuMZF8grA7gm6Xd8gO5AkxqpVsv3bTXtunU/TomOoXMo8jfCme7/yU39cA+dAFBy2aOG9
D02gbGnpIWk+JeaoDPsktiMRBXl/C4kdbQ9/a7CWyFzhh4FUQ36JIvbJ5Vy1yqjHnteHP7DK9n8+
HKdyChCpPfgu9DoWLzFUV82/20EcL7d+wCiQrtD5R2UJu9O2IQcbMeKgrfOVji1vYWjEKsXVb9BQ
UY8KqDtrfa0Z5EgBZJO27KNtUUJ9EVkEM8aErl+lbgiO8HCSUtC6O+RXGWU8caXXI1eAjy/7NktH
MJJjbrXduI7raZ2d+B2oJq/4TVV8Bo53LQll7MB9MYfgK21sG0PzxOP1ndzt0z3hJEVmgtATsfww
EV68L9ZgXp9Kv/JsPfTXfP/waCObi9ED69C6tvXxYCIXEzft3lOvv1Bl85UifcSmDQe5BWlnh90m
QHSlh/oFqRC0TJKCYJQ37lGkdDot0gRYR6l04f+tHaW7AAQxVlhtBQo7sHua15TwBHcFYrytPOZB
0fwG72PKi3n4JJ302qwgOF7CUa81Xo4BQ9k5+2P0JITE3uElyxiqk64Aq5e4D91Rv9yoSdY1jmIv
6S/DhOE8HxMVwI9oqeSyMSKrCQA9lYEmTRgEO2WcpLj6+aWNTzBS4hBqeQvoYCFBDMP3Fqk8AJ4D
dwtTqkZigiTOzP43IcUsZXI1NbP2x/ceD8JBe/kb886fCS1tG+7DOHLJEdJwyxL5fJImALTe1ZtO
ScB3pTHBO8XHnLpdlFzhwE0SMInnmqk8y73c8n7yOdjD+TX1TEp5uOR4gjMwnXPKSSb8QNrB8LPK
AeJhnrIFXfXgCZ4uuYAtRTCGzy6Q7SGN33x/AtwvHkPOEgaxKLxImhO2nIb4TgQR3fnZ53PI7rGx
9ziTIoY9IDnok1LvHmsD8NcfYlXK46EZW3L58NK2Yo0eLlAimQHiFx6+eJsBwuNRnl1K859FGKtk
Z+28AyDK9pQl72dPJ1UoW+tOkSEj0zwgLXKfgxhxTvKsTDc/v1X7hliaP9jp8uGamUSS3QMYfXux
uVKK7A9/KBX9p1JwR55fIevBVduO1mq01rPvwYWpYFRE49qtretlT3eRcC64PuEHyQ9Oy8eubbaC
GM4AtZlHqaOXsqRoY13knKAfbkAEjNLwYYKUu1qNo73EHp9w0mbb00NS/3Ob3K3G8iFN//2QCMt+
It1vhpSvs4fD1zcTvRALV2OXjmldN2oKJeCi9j9CeQZA8SLlBS7x2Eg39fcz3eoVu0yhkAp734rx
OyjXoJ+67Ps2Mnlu9+C70KMTi8X4XPacREyT8qovLaIDq29CSevVv7/cLVkdcEakN0O1b2fXRMid
GTfu2+8OEiUmujypQnmXf0QrqM9Tl0E4oFRUbrKwlkPU4P28FUPfpUDZGfKjeT6bjs7G6xhKuLLd
man8/WGwMPRVR57ZPZ+1lLq6ArxwNDaDKwQnzR4uNbBDGBv1oI6Sqhl0gI47owmZo5vQDxVNL1Hg
f8UcO/3skiueZEa6amqeIwHj1HtbDhnZZwtyNDB1y8ODVKnfUEHscEDu/haTtGuo0vg2ydtGc9Bh
BmLeo0uX+9HJD/u+UrIhT/syCmqLIQC7V+TIi2ka8X+csa08Uiw/VaTqge0HYigpG9XK7Y4asNEr
XcVwWI+dHEbibhcd22EkmE1ukMMWPBPRIANOsdCktX5tPofYBP5u5+xhARhNVXtSvoO0pnrNQUO2
yGhpH741J+L7UV/wXOD1aKdTp0OTSr6sIc/pU7b6Jh8a0xz8A7kjphW2TRrtNcnmnHX7dU1BzzEj
BBt3wr72nLFeTmrL/LPHmOOX0ceSMUsJ50Vur25rq4wUYk3srvqQ2k9UnFFCm4+vcg2KLH8V0fJo
vXuiybIoRMUSwurle18xpIjewb4SOaAB2GfqCELbgOxDcQOYkWffwPPndsWUlKO9AP1Nl3RMrosW
INjKZYQeXiR5edy33atgwqtIRMWcBcSpbugK9x7tE5uJUkXcH97vOuORbR6GWqBfW/Bdqvd4UWM1
gRD/iT3kkMirjbpfYl6OKO4sXe9ZIGmI+/jId620PlWss/sGb6agM3DBc4Gu3qDmYT6mNM9K6a18
k9jXI4U33PZ0zdcq4ZxCagGDwESZZVsURBj/Hh312cPzdCIXvdz/fWiSNy4q0AyEhGVu77ZUYfP7
n7v+s/CkMIhBB3505/i/EmfbuKa/VlTUbOEujJwVrCzmv0oCLBYIFZ0AdIsOlfabPrWiYi0zGd9b
B0m/UbUxVRHn0CnqQ2jGQVGVlrsV0kyKY0DNfd5/nB8AtrjaC5RPpjoQFN4UZzbdC1LD0y/0KPu7
3vLStX4566O1g35+8YWIYPhYawoSUAQvfvrJCMBvpLjfZkaejuG2x63Pijo9ZaD6oNWUfoIfpexi
hEtBSElI4esLx9pa1whSWUm7Wbp271/z0QBECXZgoiEM+LGWLn1AgzCI2c+qTTEMKE2roJoQUjs/
P8idJwJHIsduiOfwB7XfMp1me0niSQymSSd9g4Ekrh5U4+jLHBhKeCnoduahxuJlG3n1FmyiP8C1
tU+Jhf2iJYqgZKtc5+aMASo0tcbkTVnd13migNXq/jLxxM3wrTXIsrKvnVEpjYzRqKMCE/2fyXI8
ShYpN7qej/9QYbr0g9rSZKrejoFlzRR0ghyCrv+66WevqmXQftwUcu1czU4Po4hrg/9p2rXj8PMn
i2/CAFw7ZlfHskvNZC5mBqkXna1S2QUFQ3vS6rbbR3n5x/09RBzMNwJnV+WK+N4ERYw7h1tVDQe6
WDsSfyqxhiQQ1shH9sKUQdwjkbRRffWx0k46I0VPkzFKRkc6gSwzvvNUu/ZY0nc0UnRxhNIgMhac
0x2Ba5JzZz5qEkjwc1WlO9+FMngPJHQJlKnax/r+OZi+CfO6xgirxxbMbs9x+AI9aA0lInZXNV2M
g6+GuKkUnWUy4ydiPxDXZ3kCggIJxP6+S99F9D67WO02xeBIQPTksN6oP3/V0bIrdVSkq9kTA+P3
OQEhSjT1kO6XcQBZcQuNVkv2H1GwKGu1jSAyb7ODmlmaXeJVa1FiLOXIAqV6etNqxL2WC4e5W3+6
XA9gtSOwIBvGBkXL1jmJFFHclq352DvlNO2R2zGPM/cT6Qgctlo6TxLXFSBavd3rZQZUye3MbLUW
RUwhlMz/Ld/Rfz33AH+rY8okq2wfOejIrcKtAIg8OMp+fZ4h1jCXP3+HQSHXw14B0LFWWC6urkZk
PniCC0fhUY86av8POY8U9VbFYTjI+hjuDLlNLUB+NKVc35jXLz84Z8KS/V5GynMp24XvaIH0TSMu
oo/tteiSPJdzfYiv4QeTaB0gElM+effmx6DfQgwNlJm5Sd+YRNI5elOPzUJ9ChAfSIotToh9sCsx
pJYLLl2ChnhQgw/nNkqrbx0OvtcWWyl5oEQU7JpsA3P5hZimkptwyLLGFfg65eXX2pyulTPfqs9e
80Yefx5VSTZrH7e4iiTEIsXyW4C1tJzEx1dB01iriht65avyTrGtdFfd9kEJCEqR2D8U1hUlB51g
+N6tZNAOsl3XkuMKuC4jpnag4lH4Y0Z2V0EgliAc+uSYEBpfUzXnW5VuhUSmHXjfBwkcfGkg474v
9iMbigQMgaY8hHvK+j/29lBGHaijCkSpvuQ2fyiXdsPgnHg3nnbvRPLhZmWNNSzAi+sVHPe/+DKq
7kHUURqcloomeflTWYa+GDk3zXHirS3oLShZJYQzbzjFC/cszi5kG1P/FG/trIFI5wUIUzn5tZZd
XiyiMzRFEIoOW3RyJfQBbrPydcQu0kD4beyp+BV5uniGLxFDxo5mh5EKP5ixMSuPZ6NRMu61r0wS
qEJLXmI8v5pFxTSIeeQVzjm7L+ekjCmsNCjiNNaGf3luHzx+2j7DoqTWbrdDHik2pjbTvmkLIa2q
8sP26AEb8+41fEa1xgxYT/9u5MYfkhEUBVtfBdu4hyThAjVpWleXbERDH1q8qsFzw8EE0qnTRis7
PFsEgzPiZbL5B8WNZJJna1otWIz1kgKjc3jb3Q+jdLGoOm5O1A/vUr5Ju10izt6VhWDJzW5QyVrf
fJeCO/tkbq1V6NIk/BmSHbTymZ4TMQA++CuIwEuskLZV2ZWcl0FZONOLIaAkJjI2W1W+o8qZEoI2
a5L49wsI4mOC3+QnMvQsXPSr9KVkAH8jzLmMtKcRN0gWyW3Xy4VPyX4wzh1t6C3VQ4F/llYsz+wA
VEV7pAxO/2ovdtuZGhXuwteyQziE2w8iGyEtr6Jv4+bvg0kDhIGsMevR2mxMnvnELCmXZhMrzpDr
33JFZygd8svAmfvE36D3Qc//HOF9yx4Z4nzv2rx+QHiIdP5uB+mZO2cR/q6ANYd0fTKsf9jrk103
NRRhkbKDbP/L2WaMcFWj22WbwiIkOR0ci89mq598OQ857LaW+nRv4YKdkmnDDEUlsbk8bdWkZ4Tv
jgqPPnkAzVdtDb6bl+ZtoSO7eGHlPn2x+tfXSPUPGMsVh0HpvrOlSCbl3L3F/LZpN/s539aLZKOi
x/lFw6cnv7rBCN6L4O07uHPfmGrYaTUiI7MUKJUQmh22xLWUC7ny3htJ50beqIY7FDUitF7P8lh2
te3Xa7w1MaYcSSeeEOm/JQp+Ply8BFlOKF920d8UBLZtlCyUxHmu4Hg8gZ7/21D3rASt8IYlqETI
pQNstNlfceV8h+L4IHaJ7aEqfvMZzSgXJx98dKsaJXRt71wRQtN7/rl7EnZpcRz5pG6LK/cHwNih
K6LKb2YtE7MMJhK0Hlc+kU/o7zu2iQ4pgdvY6l/7IUQbFuVxEVfzZQ/Lb+0I3+3ayLBGvHR+819K
eMrxTCdAkCt1J8MPmzMMOTg3O70434R2hJss/lW/NGnaoP69zV5aqnPyQLUwHLIUhjaY9ioif+5J
FA+LbqgWvI+t5aCV347tdlZ3DUOksZZMTYFEsS485vrKAlF1pQcwh+0mIgEhTN6Ig8LHK2lmt/J5
JnzEM7ktCX4ajV8gsxkwC7M/YUjHtwu+yt2RkAWPcZd3XWAubk5hd/jfEtu2YSYdnptEXbDssQJW
yjRlqZLcmDIrAnYRMnNevhsMQwXwrujzdMy/PpGtgPJVGoMZyTNtKEbMR3qeVWTMn05YGQ1Pk7YF
u0D/ikFIiyqvTEcYokwM9+Pws5P80Ad/xx6e6xDEX8h1eDN3cUATpqP7e6Ofaetr1zKviW7DUfYm
7YzIMJ6IJbz8Jqxa0ZAuFOXffXouRAQhhu0eTztPplx1stF0B3E6B5rWPXu6cK5fybp3E3Y6bDSY
hCHVwuBqSTXVZYFNORvX7DQaHhb+0nT642kr5VC/CmX3gyjAS3uRYygfdpoVt5B8EaV+6PnRc6uL
JgFVNTNp6bQSZx8/y9orItE9K33zrjGDVG1R3FqXEO/TIq0JYtzo2Yw16fn9Bv7BTppLkO7vbPV1
2odqzjM8yVRwnErJV2eLgoQcSYLAZG87Up+ATqRMw7m3DYuRDT/B98BQYylWp6eWcvvSdy1bv36a
Ke5eQUzynUZFNNmyEchDN3whszG696onCxHjc12v6LhkeaGYqan7z7/SsmVTV5jdUbQzkZZCzuOm
1XYR8fVIcW4AA70YXRmCXe+C1rlFggV9vPuuLIoS9zTu9Q8LSC28Gg6Xp3sR/4zSsUjdqUH7VQcj
RNBorlcYY/dC5J7lQyL6Mef9CXc3ml2bw3VxbU9g0es0hrqpBa8aeMYx1uQveJiadRqjfiRci0YP
gal86AKeByD3ARU0EoUhBTF3CY9qgNdCZuCunTsSsNWETh8UQ9lpK+XkbuFhKjQLYoNrMqvHpeG1
Fh6M8duNSfYwqq/7uqACAdW3ka6CbBhY4YCRkhh/mTfnCrW/n4Z+aP5QgUrJ2UZTRYYofHZZ+dJD
b0ZK/0GB3fow7/yDGB1Bkz63xKT38WfDXIy2wLdY3R6iCKj2pSG+0WWFHScRTl8ao3QXpTW9pUQk
TmYHYR7O+x1u+sTctKWC4aMdG0Q+7eeJNhTk/4vzMrHJI0woumTaYNjxeW+HKTuT3O5Zq2YtmK42
GgIRUKzlmNC7VcrKTtn3yhLGWVy8dQK6ThfCFtmRvwxNJMqu6umLjlQNPC9MKUkLd8LqF/3hwU4I
+JKlUM/hbqDx4XxuUhTkUU5agPF812mX81xLr8L1uKXGDj+zaZcIULBU2HkaJw2DNy7DPQN647GZ
m6FCTNeO/HxCYu/Y5od3OJgjHTCP+E9p/2rRZmKECLxBAogBArOzRx5S+40n3j58XnW+lxd3Zltt
4XSoKYDMYD3NMtVAUewZgYMas68vtjPdTqyiVPeRnfrmhuJrG+I5qsMWYwcjcudakJG5B1cHnK+e
yl3qfHVK41seOuopM06F6bNddbIXcjESPaWffnweBdokwdMQmKOATJr1g5V3FKosSx2qkxQMt7Jz
8rg7gTKeTwdYcf48WHbjKe907DO+XaZyRmdqvw9ISIun127/QnkQfyXBwYnl7jat+le3gTBELpy1
XYzg8JytuvBYGwBAsTIW1kXrNNZPNoOeOA6WWf2kfWt9A0UOehke3kAWaPlbMcZysE5653/DjhLg
Ueh6Kzs9uv/mNIvGmSi4Jlj2oJS833HxskLHO9LmTULLv501p5F4ktAfwIjXZckDw6YT5WSsL7+s
SrxEJF+e4wPQePT5C4mSg/J1as3P/cAFpI3NL5e1NjK7P9sa7mMbppKSaauHDsF91oldffAmSgdl
KW5j6LETpZJGuhllEKYDiReOkXdUbOU9/WttcAGEtiuwsAMFQZoD7EzBghKF1p6WBr+LSHiAMfKz
y0/MNJBwSrNdk95vYCjHH0aLJTVXoZUmYo8xJh2C8r0HhpZ9H5Rw+ubbwKzb/BlJueckcK8+fv+Z
A1gxcucbxTsL41gDfPUOOhvcy/OLqR9bNnCHxNnL9cK7L9QHNzv0RN9g5by06occb1+eo58PHCbO
j/h5hPS5IhDDTOZvQzrbu0RJjiygNca7h8kTkfCdJojo5w6J7gIsrtx02Y5qG9YnzxlgoR1dJr6C
olBHzuVPCzCsuP+Wgw6tUByltrHSmClVE1ey/dUhRe5tPy1YN7Lsh5bohMDSe5HkhpwpcGh/6eJ9
Iy2CuW7zRvnBR7hab7f1oJvvegtsuOxZZe5OrVa0h2ZqY5vAPCv8y70P+/F24K8LO2anrV62NHQa
+EQVgXeICA6LRBvFJRtcfzpPuDp6XAl2xec9hgLiABwhmZ8O4ZIGeXAHvkB+NCmPR5KLcFXB6mDs
UihzxPc00iBRC+5F2RwdChPQsLLLr9r2W5ZPLw5LcdziJdldTs8mfTgqNbwV1ndf7y0wJIRohdQx
c1N9EOLgE82lLKQ51SI+ecgMEJm5FmE6TRL4f0fqsEfUazcxks0J3DSp+MXieykuP9sbPQBc7UyW
4EQ5VVK/S/O3QR4koS5IPItn83Y/aSmlqg2Hpd1nh/ba7kw1XQulMHAwPfHqGRY6CJSxJnZEZydu
lZdI4LW3cF5KlTZaju1305YomWABnfQYPoT1pnS5bSYa3vd7Un3hbNN+dFiz4hwB7GckGT03oqYH
l0roGIezIEhhBciwqdSzzEbq8RT6UFJg3lWBLQUMo6CPbs22Wjj2RVWyNSTT7CFZ0M3rGmH9LBsL
1IQGOutDpMRJuOJh0FI5QnWynkH2y0o9LJMgDc/2Lh41z28gXyokog2uvlkrfP0u1pVf2hxjbiRM
S5sVd1+uiM610UwNkGMoAkxbS8yTiysPu6Us2Mt+qXqxdVErTm6vlnuYbXplSGCbI4XF1FCHfzMo
lHimiU3RdksM2xFwejHt6Ok+//jgClPIlfHHrxmuQgk0X50jUFvTwXhHL2z7QOcXNDjUZ5H8rm1j
fnNql1pjhZ4pnskKzTKbA3EW43JeN1tfQvwQ9Iafcgu4nEbLGYddhajSNwNL8MWRQoByBDN3zB6w
tTXSTH8cdaJJQdmD1OR/3mbDY6+fVT+R3E1m+6bLbN8IHplZA6li3lVLrBHlXoJ81PjmeltPRANo
cdC3ksEUG+E91LsuWKjINgkb0LDrMqRjM7IFXUs75NYrUHu7KqjSqeiLSKCRh2Bk0kisW+NpL56+
maOCXea9jI3NEIjz4+TLWGPp+K6Oe8SNm3sfjG7mKvfgJneG3y0ZBdFItDocRUwxUxZmDSSVmxkH
TvDgjRZpTymtMzGVfntg9OVGmV32/4KOKyWXAcqDodc5dfJ8r09p8h9J7ydIDXwtHTtYJXflr3/4
GTP+5Zf2RFxW03CD5CcAOk0wk2DY/4CtzySSCmy7cMKU1heBzkJ182GtT5Wn05EwLf016/QAIxZY
cJE1JPyrkmH1zQ9iChtWiBhDG+2MifAfhLJddaJ1AGS/haX72S5X7HEAr3DmUvdC9r3toiBjfhwL
zUoxY3h5A0+vaYoRZdyx4RGRUuPh2QMWTF0EOIpZTyhT7zWMXQP3HegYUIpKElPbxVDhRSoDxpcc
HVSkCBBY8DhBke228JcyTUjFkKygXJS+XPiTesq9qZH0P5DsDZnb6qEHQoCpwJVvJenKOqLWRHmw
gWN5tK10pg0k3hk0WDvVxJy6UjwgtP+ZTvHFCTgXd/Vaf+xcjRaXf7m5qYZY6w2tYDEhNnW3ZkWO
s+G1M30BGcv00HaGpYxnp2Ct0xmovh7Cx/f5m3Fstyd0gOrzMGQMUSUCHgF2/RDfjnKu3rNsR9qB
yU2R2hRLvYymG/PFM5XEQ6/roUt0oJvbnjQH2awuqZP+kUE4KEW7f0U7C2GzlGDFroJ00eE/7dr4
rhIiyZTWxTIQ0R7ehX7xkW3/BN27OT0nWcKB+LVPeE9KNF6w6mpcGb5zc4WbWfrvcInOfuPzUSAC
ARf1wrBzLnklIO1lluPb1pcf65hLu2NlXNEnuKsYmWRFOk28lWxvFoL2a1Va3gVuB2MtIehCp6Nl
gVBHNACuCV8gmWDON/B50OXa1dMf12C+gubHZaOvtFEtfKXPRQMCxf8xxgfZaYWLXAhCM5IMztLj
f61p5GPwg4LgSNPCEUyEB51olf7oA/zYG9YqbYPbwTwgWkAZMrA3GVgNhratUQvkgANLC7pCOww6
PIRQ3QMhOnBmJlkH5n80+S/lLfi8dv4SO6HVTMrjJxLNHD8hdoXP98P3RCVT3NT6kjaqqFBz3pNC
XMZnYtAYqLn04jFKWO3VXqnTpblj1GkelmvzIiJgWEh/IQWLWbf3xF4PRpajHR3gr9IOxlJ01I/8
6ZL9oNsnGmKr61kT/NqLtY4G5dVZl9CnWb1pw/g8m+uTdv+9gTZhqU+csnO0JHW+0oK2sYCNAdYf
sfQabZXxGR1UWVcFEnD/wOkbIxPq8tWsuXRS07tjNXdVKyrb+wd0f1ZyKBAFtLjj7wUAhQTwEwtz
+0rA5TD24HisM8pSMnWF7rbG+X8T7ZXRUNsBO0lyjKKYd9ycn0wey71zmq0qsJ57eXcpIF/x0Ouh
3vCjDj3G/CdAxJwG41ejZMYX8/8T7VkxJmsVFC366qIdSUY8tIIPT+AcCFscgh5zskTfn2RpRzVA
hB7svtpvkOAMw+jbeY63+qHiXhurQfk4AzGEFuGzdKQjl5zqznHWCXMsQ195OEABrn0pR2ivmlth
UUSirDIFKPnNaM9zfUmzm1SSgWXispaw8RkZ1i+p2GyGknOwRKKQBdBpReby2YZazR6wvCWeU4Cr
CpC0SbR2llLChVuNNV+LPAj94lzNvTU1uyTmKif2ETPFrUN9e9b3IzrCH2DOqd7asX4z3OiXvXYI
UNZAW6c7i9CjwOGo8BvAx73NJNjHx1M5FQS836G4+qkEIVIBo0CNYBAoN8A8k3YXma5mlD80y2eF
jEHgd3KAbFS7wxDTYcOax9qzlPFiaHkmp0SmFaXaJ2vl55oBCzA0xL1g79deFdrReupY80eSxVTU
HTG0oMyRYB2GgVEluupohJwxSbQ0+XT4XQo2km2n6kwbk2/yQfQcJobAqzcN4ZOb0T+WQgjZGdk8
YMlBMQ7UGk3VFJ/LQVvCTBOMda8nIM3sNfyjjoSi2F00Re2N5Qre8U6l5vTD6yq1K4RV5LCgJjUI
UYPCUmOGokZWWTTbDZiH3lc5WrvLcRMlq/0RuTdIOgG8k702QWkOE/CLeHC6jGmm44GOlAVgtYl2
Dv9Ej46a48t1G+7fSMmUdOoAEmF7uTaqEWWHcdX+8GwKmacyf5uDJHisQnmN5kHAjydHPjVuPSkp
me+PZhg7XinORUGnw8Q6KCGwEWUvYwSZM+jTOkb1c4Y4hidpoZMnSRmOH93VSPLbuZKcmkvd5usy
XzpFzZWmoAf0Ghzjdm34xAwcBapFey+gEulV9d1OK4vjOipqdytUF2ff8l4t7sXF/zFp0yqpVbKy
alAWmnoYmtmVJzR5M80b9f00nF2GU0Dj0bQcO0nBi/hsWh/DZQ1Y/s8u7il1WZTFoUwVwaEnmWLx
rFEKBKKcWO5AjxSgDCuJ3okLplUkRWH/0K6ppaiMbRoCbYqvBNw2XMNYt7g3NA7bn9zSJxrWDlZI
nOJ7WJ00tMY2fsx3xriZaPu1UQztWqICdjr1N0WYuEa0oktWwoiE1e+FGdXQNc9JCkLNNY8pi94/
LtNhs2wE6ZquG0XNj/Oq4HEePuC5EcmymbTGX4PnQ745itFCAQTq63i1f5WmKdBKB50HE8yvklW2
bSiLJV2z6DX0Ak8EeROGYaaIQKapAWOKsLHYfCcnY/lq4RaZRrlfWWKieL+OxEbaqEHn1Z7yd4s7
EfAmEs1AmffJssLYY41KeBC+jfLWeaIJ9YnAp2Qq9s3B2NUQTULuf9iR0VT3G6NAykAG3cclwQOy
Hl9vO8EGHuTiJ01ak2nwiwthY927wZ5e1A2kajEdvKb//gwr81urw5RiUYFhMe3d0w0kZ/YKNgHJ
UctAzgh+Mwy1TIjbnq8EzOc1EU5ujPZax1kl+FZliEQaQy1/O9PUcCXRWwt94iwAMwJZtk89OzWj
Xwhk/RMKYObVvwwGmDFzeA7OMzuODDQufQxATSaUvvKXqsN7WLYvr1jGlfJvzRnIHPHC4LF2jhEU
+sbelY15NFe/R6fuqfs9AKx3xFU5KOhg6/Ue6hmp83aHwQLHAw0XXnz0NZdLriV+TdzaKwPe68KP
YAPFcB04aoqU2hE9g6+riu7HZlImT7KPFbYtfVrankp9//VdqK8=
`protect end_protected
