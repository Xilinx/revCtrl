`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 280992)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/oC
C7fe1Xyz7PPjJRef766UC2pssNmd+h6jWR2MDwb+9PAG72uT4E/pH0PsFMx6PL3sMYBjTdFG68hH
Y0UUSY7uDSZnPp5llv1mKdFKHpXiW6OQucBNJ82kdsh/FrEfoqTel8ydcp6VAhCv1ybUvnZHC4lF
tLUTeUEXyaLgeC67roPOdhA7vFirHDnlDuij6kgIO+l0sJ4vnT17sXGaTlvTPH11rQD+hPOnAE8d
3IqFBA79G6M2pFD+vqHpX8iTtM5VOLUiBjsHbnuYvJ9cA+xdvzQbTk9gsuq5oLPzxNI15tJ7bvx4
Vp/GZ+lV3/QQ8v1T16iysSsDA+WzJcbdkwB4axtg3MJrZvaJod9yLOxrKM2GUsa0XN3VQxOHqgUb
e8UwzEJBPOapz4PebUxAnXm4tZc1cbs/uC20QmfCSCb6NF81kwCvDA81s4NHfw1oxPZfwQfucig9
ktgxWwo/3byVIoUPuH0maNqxKejBpHSZtgRjcv3GVPAugbwgQ/2a2g4ZRvPgHogv3hbsE1bT6jJr
FshHwiEhN3bQIVMQqwAnvwdtczjXdFYhi/uqmM4lN06WkieptjmSKrWnPL4pq1oRy+/YpZukVhCR
C8u6DREA6pP5VLmJ0hoyLcOZ2vNotOEmNybRwY6vEzfkwSGm3RaqNrjt2WgfI/g0SrmrPhbhQd+Z
Or8UJa8WZWs98vSfOgXzBA26w6maxjTH1l2mAYhxFs3SB1L0S8OOuKnwGZUCq3QbUDwL6w5MCss3
098QDlnAfcux9RQfYzLf2NQRMuH3CtjjYELAp0PnXwnP2nkJkcagexpDUcVCTagatIqjDPxg1D2P
MulerlyrsVhf6bnOc/wi6ok0d+c9999VhzcBEKL/1iFc8LpznLF68ZgemTcEzm0l1RwWpAxatFI5
AvvEzNFlaoZOakPbKMD2f+QVQN3vKbQKDMfL531Eel+WC5Oco7j0c31LEYslB0XIg1T30pE0MgDa
A11ZyPlibqC38umWeXDIKzKrSjqO9BC0e81BDJDAZfRO4W8dAsAVQj8mC94FZrLW5sTXROlrIc+J
jlsgn73xIKWd+Vw23hTmpVygEZdgOiYnq2AJVojBW2fG21VGNKz49Z68jIejQ4uqQeOeuerrELNU
HfBMwfiN91Eofubxq+vVEgOfWVxtbGbb6aTvz9H8YK7lA9mUxx2RXc3OdwlyOSjfltxU74u/+iv0
D22018qB1JIlm1nS4eNbhnkR6cDm9atgPsaCs4pSYqIpbWrLlWzAb1ws4tdBgewi0JgXXB9M4u7y
5HfTvZodTABGCC79E2+SDXNRSQhxXGppp6tcbTnXHWa5a5SAJsKCIk8rCpZuUGZZgzb+Q15gly/K
WQoTzgt1GHdw8LTvaDyh6cKZVD8g/Z0LDMtMfDC5mJQusAqIUmWOAkDV7Vp9RgB9q7dcDK/CIABQ
rvhyWWu7oLrbf7VtjDNpTRWYNyh1uhxchOrQdPwtauxFrADG0xoGi1D4ESIxIvm20U6mzRqUrIRy
gT+fioICxD+Stc1LM0U32maA0dN2UeWxdHpSXdpaKaSbuIiiI8tKtCchMn3duGzEP3nz92K4x1Gr
tsjuU/749HouDBPhjPPfg2a4FwB+AvBFQ6K19gQ1Y1v6N2IFdSxrO7LokD4B3ZHe25307LNqFh7q
zTQIeneur8QuFExdOW37DgKA5s01tsIAHni43+F0YqJ82/QpfHw0tLGxtgYumr/A79ej86Qx0137
ex9Y6D8OSjRZZEWrBgSb8kvWV2svcGk9Uw+/iZP6EhNXLSVYkaFPocMbHoEEr4mXARHlXTiAjmmy
jwVW1qMvebu1F2UmvR2x3wF2fXs4J4scku3QtevVYp0fsG4TB6YW1iEtVH1HXbabsKY1AtN4nlQ5
e2m+z2XAXHJnDNdQl0eu4Er/TTIcbLv+PiDcO4/ydh5XjnhNThsxr6qAxHR+DSIw5jevIirHf7UE
XnNaSPeaJ5jC8PTfeUz9LFPapws7DJ/adPfaPmV46iwM/al7v6YVgthwJldMzZFgJMevKRDYsa+s
U6W/8C2wSq1kLhvtY7eNPY0fIKC4girenF1dLTj9n4c5wJAFyavdRbFCn3de7Zt4Kg19epgcPNJY
LATXnHlvYK2fmex/pvwNgdJvxzekqVDkOe9mxjNRvkG2Mwia8fNorNOhiNvpX0FLH2q7bvSlCG5u
t62/MYuPAUOSRaxy4oT0pjnOM5H69LE3YlCM7dfgzExZnrngzUuuChpDxM2TKnzcDJQodYEPNkvg
KKDRo/HPYkVi4pOASX+4Vspughbo+V5ndzGluOf38Kgam/mPSWQ+2vk8DUZ+hLvPgbVy7sbJNuPs
IHT89m0EnwtuQoaAK/aAWvfAlupmxNu61q3CJfJhZfngHy6A7Gb6MHPUCk9jol5HJs+Y+MnC2FFi
PeO/6v5iergQYSSM/tjLscPhoaPN2SL6uLHejw75JQ5Ts0RJbogQSJhXCXr0/ZJGtlVuusZPXjEP
Exbd82VJJZxgDfrBuH3LRPl5nD5llxRn4ll2FpHDAKgofsnTSfz2HJxAiy2QMU5Si4in2tbyFdqf
1pjTSzEY5L+nsl09zbONfynGhKveeVinWO4dBhBxoAxIacZvXPNQNsWeyd/QgfOMgJsnc88rpvcR
EgfptSuPBJxtpT1c7OaUJyAc+MlMijonvhANcCD6WUQD05N/dYEIg3kxYLcVblNXW/mAkuPkBTrS
//BUiB4PNuZ1oMGHB7y3ZfMJX81FbfFJ3ILWucnf5tF8x134TuhjBZuJCd/rGw05bjFn1JEza04b
nCZkM2CyVgyxRgIOCTOt9eJhOkYUvNZ/fqLzJ5E2SKWJl8/B3/lEV2ou8QBK/Sjr/skKJwQe6qwc
2965Pe1n4kOhCY5OaFhyAf1OVXaF2INBHbkOrpGV6kctrDSuEM0gh16I15YDSvOCdAr6u+EuR6vC
ipFVOpP23uILMI5djlm+dG53gcvoSANTwYpQ4J/12XLx3rw+0myiXhqGapV4dwdD6VLWWsZ8Hr/A
Cf1GGKULgoPsgzbTP9c+fykHhT+U7z6KmH5s4dmYMnHusAuLe9QNs2AX52yfLbOdK2OyN2epk2ql
zshItoCeIAzKS/wuCImLcyP4q2VfnqQYOFMAd0XSmhUga8SNg9JNyAEwXbPSBFVsGvFBUepsuQNZ
bqb1uoY11bdDUjvQy3yzi7i6+qg9B45SkTfYocftD8wmtosbB/zJnlY9bLi0AUFrGn2gHL2x2kzl
0IsX27FVgcMWfMmmyn4xpi+utfLsyFMd1KwCfJBOdbugUN2f+GEWiiTJdLFkn0YcOqnY9osb2Wgc
h100Nt+P2we6WZqm2cZ8zBOv7A3rR/y2lk/Q5clUHd9VOj69gmCQrCfsIMxRRUqGR+CTz7XUuRTR
KIz+euHJ6X1ZfjKX5AURV8mGrZ1omH/KngLu7bsKP+QDEFcjA3jjzNIcGeEtGTiSlHEwYhtdEu6+
Gac5RNJXjPFLN6opyFpCgQy0RTMlrmlP/2odY1PYmLXiPv7mui59s4wEdnCcmdTc8HLHE9mxLZRk
RCRqGnAuHaI3FSNrpIRZqNMnciQ6zafPxlUqeOSpiJPHP4NFfDqQSGGYT3FMX86tR48WgmGUZFtE
uVDX8CH+O8zrE5dxuLeM9PSWPoaZlYkUK6Hl6L1Z1bLwR64HnutiJBGOtRQqCNJQiDi/DDHShAyX
f/A0rr8P/I/1bWTbAgVreJEW10UVI1KhOsofM7wLo3B38GMiZvaYdOCPbNollWm6g5V9hcdOgztv
9spl+Y9pASMtaz7sCbz2nDN2fUJNu8bEc0+QvLuyahWg0LzC5pm4I5+5ZoVjaKEWhG3KipdCXIBS
6K3JJ152xf0o3NlyhJf62uyxBTcmeqMhTELt28sPm+4odPj7lxhJEtnP3fEz/Zf4JFzeNaYdYw2g
AkZErbIdJEqlWfLpgpP2b9pBZ0WE3Sx6FKomKqF6dAL9CHASmE3AX+clRxh/kF3ch2oJd6J7uPfn
OE7LGBAgoELR8LKHZOtmMBcks0JpUW84Tku98QtEZD3waEDNXJ8ucEMKoLjtA0/r3lvLalPh853p
ZI4z4bwJkqPJ3JmSSnIz8Tu55sH9j60DYBLskfn6FdHGUa0A10YqF5X7GkxcuKNgb1Smxrlx8n5N
r00oUdF35wIxVmvadqUIWg89US4PYX224KozheKdXaCj+dTuXVRWQ6kEZHQ/GKWY5JdvWqC/r03p
9xnYd+zZCaVArXEUIr5G2h1igp+irImxvMyFEXY+RfgtkmvgvdnaG6A09mB9yPQC4cyFi7TJ9jsm
NfkrHsQLq0UPEOe0iX4nMS9sVL14mEyw+Ka3ftZhQsPvjYfpv2WbVz9L2Qp8uRIQywBJwBeGnKM+
VtTkC3cWQWm7PAx0qFe7fj0EkSZ+8KeHKSkdUuH45wfv5EwzNMMPiX70L2TRB8G2W0rwXY/a8k9c
aFSliq7rZDCpIrPj2601r7YKW6Phc9D135gecSn8llL8pFQ+Cl28XL9H19KPBCbyp7CKL2YsWc/u
5ahyKa3xsmWditpGnFWXHqBGBwrNPzxX8y3uytH612mmsTc5F1tFsn37tdXY9rnJPxeMGpoGuW5f
Xg6QJYLeMgDu6bVnB8Gvs6aZdGgvL8NZqYnn2ckKbOLHZ+sSsVB74QjQnCLnoazs/TzI/6TWpE8E
OvejhpuyLPsEMpEcvaSl9cX5t1twHR810ROhcU+ZiEj0UQcHzxm1s8p8kwtEF47ynFBJGtQHcpO9
naHvDk8yla79oYCwGg1kICzYllJzxVgw1O9sFqS1fE67YEZAgruqhXNdtN+8V3QMuiZWqBNoVyHi
OpsRuQvfM3VLWwicm3S00/Ke51uT4QwNOpt4OL7EyPZaaF5tHjQV14hY9Mdw+rRHMfpGSc0nPU4m
uhS8tjQUm09iFludzYdkkiRVH+gPd0Q8TkQkErcliqtYNpWg5XWBRXM1qysPilXrFv/6+/ga7hcY
gaHamKMzKixabicqGCBNwGl3imLjCnNu6rqI3S3l7WQ3oNahs30VQD3OUydYW8ky/vnkDOBe6Gsl
GNTM74w5+d88gt2R13mxw49ggiWC2KgFxR5XEvoXpce02sG5dosgVrXgMFXgRLwuWENvkj6hHqfB
fS4r3vgU0nFR1j6mAfdJoZvK+h1dwe3X0wbo4riUpFkd5rJxZcAwBzVvYWrxdfGGqBBqDWYf1gAt
9y0JY9ItYq5HvUbeEJjgeYNhyIDT989c9dcVlQbjFkSTZml9++19LNTwkpNrrtz8EK/EDFqqzvQn
H4u8zgQdZDL/ET3yvtaSjZb3rIdt/7ZfCb2kr2ppxsMleB4i/EkfHThQI4k1PTM4fiAkr53F3hL3
2CRJQTrOs0FuRAk4CkM44D026kMdG8fdDW/qDD7Gl4jMJXtFHWt1xwM7hu2gZNNb/+823ZrIjZ9X
aMjBlJn/YpsEWwfSalNF8JiZ9AZ9h+HhZpDQr8eBYAO6k6lKuTNMBFAkLdv5eGbM4JA2xOFpTv46
ksXuRBQCmkcJkWIygAKIzcRhM7pwqwv/9GqjZF+7nP4hF8mKjrM5vsgqq6JIanVt5SnjukZjAb+m
jRFacQ4IpAaQcHCOeJW9S6JoUwr1D8BGbmCu8CrX//MlNmXPr+LqLcJngFRXO7GJIpcdOIS7tqII
CyBmTI9O2ADpQbqCUx/UlrmPuxDLgei2ShSu8LEca7MiiptF+ht9k7jwmDWyEbLyG31ZwqO6Tsmk
anOwDP8cXX8UQqnSq06dzjs5GGm8uyoE721jVkZOF0+ZCZXjPyeJCm4SsXPB2sGe0sQbQKP80eqp
qgS3awg4xI7xoXzyXGdURr8yhG2WdfvT02RbFXvtJy5Wil1lyKgN0hOPGoWm1AmsTvWYYbK58uw0
+BdJnximNpJxoEndUX35jp45/QcvlJrLde0zPTjo16yWikdjJU5bw9LaIsrBtltSKUCh51xYpLPw
v1fUAGzuU675Ve09dygK1U29gkQM//o2S6D6VHo8//MufiMtzldVbYJdtZ+0v5S2XWWsUi7CYTiM
mSRjnXwGWOb3CaB6qf9BT7SX3iWN4yrHOCXHfzko0EXmrU7/T6GFHQTQmvHnQZD0gRM/ncgUbEH3
Pr91GCpKe4y1oN/M6uHStvfenMJDJyzjHKtCizlJ0cpd32+bwwgBy6XVWyW7pM+0a6gGwYe8j3Kl
n0rpj1GRaj+4CMJ0hZjEqXbbRjyq3GYtu2WgV0qF+HdpTNI4DqONPr0SpuyzcRfJ8eFRQFIQo+Zw
pvL+DxrNWRdc4z5s5FeXvtd3mR9RYnS2aY2XyNFL/H26+ePe07iscnrIuhBKpvzfD/BiEb0aRFcV
79OLZAh5oIEzg0pmUCx2DaLqEuvt8lFSJxVOSoGLlXeMssoWUFzFGRA1ilsMldpgB7CX9re84pir
eJNC4MF8CcjmKeKQVN2WMvQYz+Ohz4SrCLlBjFV0y0qvolp6yyeJkPmeLV8dKuwRoTPFlO98gere
19TWZGsqduHVdsSMIEZSyWfdndsSvBiax3otPCpomNwVpm6IKdtC5SYa3SsWN1Kvxenv9NEsQbf7
Rt1imZtgBELXvUb4BoOv8lamRc0Y91q3ba4k/dz2kOhMslACo3aAM4bMDimDYaxSaA9nR8lmdWt9
Was75siotqYD4Dey0eLeoZ4MlIpL+881rfaME7J9uTYoYcmWBr5CNZSl2j6lR75YvdP/5mQ5aQpz
bSbUnSxNa2mZ6H6tqkNRS+JcWXIECdtRVWht/Tv7kYKYsBe2zAqUBw0WkP9cmeaqi4mh2uuErL5J
9hGXl+Hqj1ahiinsLi4Jko8F3yPP0RjKXgw9d3B3MHQGod3hzDBZtXyytHhUUp/MnucZF4gQIw16
4FFVKXF6rFyFqmEwLYS/OdlizQ3L7yp1OsQFY+yCOgoTwlWVNLenQxbz2Kg1yxfdymt1bWcaKHN3
YKTQPcA2W0cJRNMxDRRxKf1vKQYX+QeZFKPFsTDTBPQEgtVRGESSgmuTCpl2LT3avzLQby7n2lYs
8ZOVGzrs9bc5y+dsMP6kVc6nOu27qgsmVmZWO/+IxOjTzIoznq4yRAYnAKqWkiiSsKae1FBRR5J/
WuIY5CLQoH7Hfj9PRQWycb54R1NMZaRMqNu9ljhHmkD0BfQK4v3EJZP8QPDvMVgFzxAqu7bGkZYi
Q7lsn+rNrthOehMCdRzr0nKFsukaBh2iT+nWKnBhYxHTAPNZqT/zUZw2vtHQne9IDxoHhdbi40B1
3sAg7ZVMQPO0ymre2R0VKfHLGSyrmn2YJo/PEs9pR/Bwft87nkGfFHiAdb4SrCouOLOxNbOU0iww
eVzzegBNRu/WiKOaYEb6btaLrGM3cHs13ztsrU2GNp/VhwZyulPFZxFVmxfo7W6bFsZpts3k3hr8
PT9CxYXd7kuq69P1016fmWkc1DUUnV9nsHiuNCJMM7SXP3hGSxeHLQAzw6QDJgmXKCslLWg7+Ipu
0FfMifl0WyIZO5LOMZrV2xfCOMf5plzqU8UHqR9CtXrZyf/XmJlddoEht6ABSc02O/FDTNXwecp/
4SmevvL6eajvNDOOq9tfBy7FT+EMzENFbn230Bkhe4/1qwC8L4iO+sxMdnmLN1jaAVTBdLZ0UtZ9
VjMJbkG/KMxOo314HoRpP4xg713hHIS+cfHBJP8zuen+SkD6Kt7HVyUO9FGEi+IUuuELZazAISJm
O0Tep9jdGz0oH2bHkDPciu7oyi2ZcOMnrw+c1LH1wWsbfE1khAy3CfUkhCpme4XjB0gD7AQ/36co
g1cVVJTQfA1hsj534ItiqBrcN9y93eJNBwY40g6wWKlptrs57ZzrTidTSgkfngnvpWGbGwNPPy4r
5g0lCqDgQVQoj9u21M3B1Rrjl6xH4woXbwgHCREYGj06hEVeSCG3qUkVen8fybXcskwpBkg4NocV
V7ILXvnNqnGYJ7qkObzUh1DfSpDUC0f0HgvJ3YiHcOM+MO1jQxwXFtfD77roRUZVjADnJ+eHSYDa
IpM15th6UYpY7TDlsZxN8K+/53VtxzktGQsjRUmKBmsfqV1colT0pcCClaRV4kF/bWHNkmstLOpM
Ju4d9hyG1o5PY6ijasIj5cyFt8fAfVz6xvlGPTn9fsboVntToiVs3B+Jsh4+b/rHmN8JBd7pTEyr
KpHkQ7z799xInZnCWwzdwWSpk2vuAh/IWW2GpmO/oGdp8L6s3jV3jHB7M499gf8edvRTxwxdM71k
KolLtGCPAg0SdoLPJLQVxRQtoCQcQdcL6Nda2czdZ7U4FTaWMw+WNh1OQyEtQ5aG4btv8Wc70Hyn
/rGvldhaRtwvCYHtwAogZclh8ZFZbqr9LJ4RpelllifhBMEZhnqVfep+nJI/srcZ4atbVOAj5rac
KIGX7HkHncyXVKfOcbumTwGn4nHvm5N8EgsGLhIBrnxoN0oXd2bXSU5Uryqxjcim1oCZpEsALrG9
bH5iPHUhr72Er9GMBem8V295Tzys0YXNhquK8NPlczkoL2k+ptc8r5IuKCy2vRC3rpHiz96KuE98
lsH3VTqKA+nWmQkI/TAqRbWIP7qdp+rIimvjiGcnyvnfAKELKStKEd2qZuIMbEOguMb4MuH6Hhzf
UzvC9/tc39l4RpJ4J44thZUpjOMJk+BOXk685e9yeMv5r++t5d0z4u/+wmsvRbmuJOhDSLQqq/bj
6rzzIf70Pn1vY30nqLGNMkvhhGHUJE6dXxd000OVeUxUugOHyVFmVelUT4w1hyh33HsUoUoxQK0y
Rr9W4O3oQ5lc9W8AKnX0vsRgpOK5EeRaSIrXdvytf27+JY+pnV5v2MG2kU19XrUbtgDuKwlrkcsX
lj/E2y1sy7BJZb8ADfYy0xmKB33zZ0qihD1dOr7EeR1TnGhxVG8UMEU7vfFjU7DvJwhCN+NnbZWL
0rTCWeBhX0Q2/yo804nHva6/jWsznxkOrebZcFDR61d+sB74JzDJHuDN3QTkmkN8pNcymuTaHLFo
F20rjrpwhlODfpNsKyqetbAvzL6nATSPIp5QSPz0M1+qltUkGZI4Ya2Smq0L9E7B/hO4Q8nGnk13
NfORSHE6if+HYFgZHhzrd0a5eKG+r/9FNmuoQBJBwPEpHuWdKXpHqXplsWWUn09TazrP+xwen/5E
Lq9URhIp4O10xVw6F+yD882d75kipcQYxeLxE9xnOW3HSru2gddKym2mkUL6ZpNkXuRYCIUUbEEO
xyk1mpI9qpDDuvQ7YYVGuJM2HpMAP9exWB3bDjMWgyoCtsYkEP+nMcURWanMx5ChL5L/Pvgk5LNq
LeNu4QOrg7nw8Kml48n4jjV0da00AQ3bmsax1dcNvnDMF179SH2fZlaRvrg6bsa77zRlnRtCGOaE
Gw1ukhd6+ZFhj1jnBrGaGIyodkGNfpJSzCRp8LFC4t2+Up+aPGxcQdWPcX8wpjXZTq9E+hoEdc6J
xl1BsRPKsbJ+JssD0UkRVyp27GNJX+okcIP7I5MhcjNYsKW9jGI/VPFMsSvASv9rANSEc/qXjOzM
Jx5exdOI2nT+9YRJ7hLRaEXGDfxD0cnNxpuYRctaOYRR6KNxpDMbOXpWpIUvOqhvQzeb+jQfbsUY
8jt/dHsal975SUqN91tJcaaC7YSqPSgd8y2NOIFohUZlBUK51YPb26FqwMNVpFfs6Df2NogteGjG
3Z/0nGLfTu/gHTWoRsxYwV0QRhfy5DGtejmQpFALDZ65G2JHeZqcrUkCWtklfq67irrTWFFv8Vtu
VhZXWgSo/ajKCwiUiR8cJbxbZi39FXAxfCUQdkWS4tmBTrNpLDCSj822wz3U5jo0viRWyqKZcx//
OiWaxmHFmbWLm9JKUimcaQwbBBfdzv/5V+YMNNfcXdBHdViokBNTn7PlvPhHSUpaRUfnSdMq1Q6z
DWQjsMBruACBfo6u8QwWpBFqLAagkmJAZbwm52flICfb/nlqYO77M4bZQnBF/i1QBU9wilLDTk94
Sha8p3esbRM8t7qZOH5MKfeSXNbubT39llP/H2VmFpJYuqrHDS/vQer395fvLr3p6dnuKkOiCxKu
xswDnxTrjitXbamQQrow5h1hSYk+nHMcuVlb6Pu2Z0f5wrrTvIGihvSr9+hIJypNybqZRHrSiXAt
2qF9UK4nBopmyNpedTQb2hYgYw2qorvGVX9/4miRF5lVi4/66y2j6lD1cjAMSZhFKnFxS3CLjzUF
+7yo9aXtAvpagPV31rysB9TOXslqrLR8l4QSeHNmibD3RMpt5+BkvZidUZzeMj1nk28rWWDiB/Uc
nTzhfQhMkIHMKasc39CqCo/BIF7/a5CHHsXwWbj4IPAP+vdhWykN5KBltiiEPAepnMv4cgHQpA0/
P5B1xs2qtDLPoOrM2ahDNMb7Vcyy4nEeHX5y6IM/j5D8fetPQ+hFD43+hyMhgVZcjPAmX0+rGflp
EYV8qV4FJ/9J6UTy101iLinhyV4iv/eTMuWq+M/01Ombsz43/kOeiBmHkJMc58kpQQShwWAwPfgc
N3vdRQK+CyzVoX6eAgYzKmKK+LbJ9SEjBm0jzlSqae8FkfxYdyl8iS+6t1T7ePS2zZSxGc3l2hsC
93U3bdXMlY89ZUPaqy6rNfXfizCCPpd4Jow3KU8EVkhh5/S9160C/ArH+vUAN0+yz+il98wNJOX0
4sSWBuqDp4VjSZxldXwLrvxS1vjdaqver3bBd/7RdtWnp920JUohnYQ65bEy3MLmgrj5nrS14BI7
sFXVUhc9AHS+Ow5S7EcDMdZ5m/62PmrTJKAym8+ItDorMYIoDgL4e44OJ+ElMZogVxrzassYpV0c
7zQcAAmGOLKnjEd1ehHsWLDoSCX6DrazpVoLJhmb9uTjJ22WScvSWC7bJVMP0hTOrodfeKQnJ9IJ
by3Q19DbZit5OzYgnbC/+TPmiQuaYoaPva6/wdGKjIt6d8utG+pB70/y6XjJUiWUI0kpaYESUpFe
fCIJjJv9sBM7JDHC+mHHdVSTa59QkyfTHYMQofoFnRtriUp/zitryc/vj0PibvbLlBbJSV5Y/2Ry
ypAQ0SIwqFekxffQfAxtul0D1q/MeDHEdsYxqcyyM2qadZ5ZHgE/18rkNmlM8Dqa/kvO/L2qoX3x
YjOFqkFh0QO04+1LoVySw27xLyOixKd5SbhpIX66u/GwOmEPwQLzuWDFB7kO5ZIGH82wM1wsOEkY
gLuwbrkgnieWT+EQ0zTLm9roUDxq8SNKq6Qm9wpSwMggSth8Ju6PUCmjQNjFZuTTRilBueMAP3bO
M2pzZGmRlhq6iq4rz0FNnZPrd4PRQ0mYRM8qR4Kgx8svOkBOHirlyqv6dMtRY+3fbD/72LQkmDvB
CgkQBT4ynlrjhkga6hoN6botw9oihiSnVmQ2xFzvkP5DLjkXjxoVGtTd5gXRMFK4vvbnSaXo9hiB
oepCSlsNU9LeVeHBkginUpVJVX7GChIF9z/6Pt9SGJaCE1YrfVzQONcSS9vjGfL/jo9ClRCLwQJJ
GJXIz6XhTHWuZufucvg6W46ycWU5kpumRs4Yihf9ESfWLeB2+4Vx1APRYO+oYnOBs0saSUCKI7S5
kNmS2nnL7KQEe5l/tHAp2ypcUfLWteyWpJ5FQd1wCTiqLmbOBv0ArAtaV7XkEUP+XNKJhj73Ckf9
Jj24ZCGaW+sJN2qFL/giMD1wt3PUl1SqYRbY9b6tVBc88GNyCg7h3gPmT9pjgueDDcRg3QAoRgOF
wii4UTIL5fqdLY874Ao2a6kHFRDwcQUmvhirNdkfbBevNBmw56NWEmjedWfy6cerwFFVg3/TcXlU
wVj04R+Rf+XMi//57r1u2OFXjJ+HFuVgpZ3sAWL0Kt19U+LNgdSoXKIZKx/3uckQblrbwkcscFAY
HNZ8EHO6eb55+JpucDm7wIqESkCn+Uy1Xp7Xkao8rFU8HeNqYLqx+EzI6PyITh4I7d4SmvuHM34Q
515gQr7hRdXtH5kvCE2yrWOqg3VPDadcZLUhTr+zkNmGLqlZuyLbryi213AyCbppfcLfWO19FsME
gXLVnM1WgTHOiipMOTIg0PvRhoFq+Rg//g4IqUOP40j7lZXEIdtpnq7cvbL69+or2LDu1gbXIy1W
c4donbtYb7vKBT3n+jaWpss9nUUR/U6i8eRj7Zvll74zW113yO4u4YxTqbcqFGMdWfY4Fuoaljb1
FaAb+Wi6ydtFg23/Mw1U6vfvuAZ0583keJOkqBgYqHbVdly8ZnOpLAyHcXkJC1MT/JAf50ZXxZja
OE3cKcKKsRfQhj6lpFVDvN2zBfzJlXk8C0t9QS9jVsndVAP+3fpDTa78Dr9Kdsad6tgV3epFQdDJ
aAYe/qJukXnbLJwdaQ0sxcDULwHTPQG0JnLRPfbJ/NIw/JBV+GrVVwVq0W4pGZ+Rom0r7bHuRLhi
UF2WofhplMcOkysWVoN5hssReXz08jnrUXd61OWFngvcIE8w2WWk/OnB+u4pbbuoscOKK3tv5mWX
qQshANb4J+SmTBuILKFOBbqBS3YkQCQk9WNeYwhx/Ay9wmJPYAry/RiXjNFNvalj0yj5Akvoy96g
VL75w99rf7/gY0SklccRZUycvAhFNOUankvx9+Lrw7mu6HK2z7xsD5kpCGkDAofZO1NPejd3ZboD
JEGEg/zad2kEv2CGioYpSOuJ8Q//El1KUl3WN/qAtAgoqX4fKXy6R/zr6hN6pVd6H15biflnuvFM
sG2t0m1LA0j7K7849vr3971uTSZeNsakUE9TBfuqBSIqas6bPOqzNi5j894MxO9LQRnnbHFP8/Z2
h9uSA6eI0NYceVou1j70IXIOZem0L6H4kfMmkLO9wLpPw983adRhjnoynKiHi3i0hJlYmiRh7TDJ
ZK1y/IvJsHW2USF4CIKsCQGBE9A642fv/RXjIhMl/ECKOpLcRpx5H/ynWmaPq72dHwCSYv6PprNc
C5awjKhLskAMgKHyT9F+r7eoDD4cuJuLkT8lp+ihhebs7TIQoewVmvwmaLvYMC1hJaLbjUhh641M
vuHkkxSHWVjzSkomRe2g6PzPShDjH5JO/uQS/9Vza2+Gw2uZ51abZ9gewdsbSNa99GjN5tnfKkFR
rdCd7JWO23j6sBxjrJND2W9ov2huqZhH3/5pUSLt9za2JsGEBqE06aj2MjyTQeJfJX//j50hpaTg
r/Hv8TRyBSn3370OzziNr2So1WOnGg+/hz47106C2061GWeqtc/CR/QtfHxdoZLsBtydOlGtTbdz
z19UvawQbOFNQwp3c97aViQaMr2MOS4UsyDivZ55BMedLKFNMB7eBWskoC4ABV5Q2nwnnl2iVB8U
w3GVlG+c0TDpRkIoaPQ0p2rXZRsBl3fuzwAWR+rp1nuKEeeTheNqgv0bsQlQPehqjllBvDcZGdYn
xVTqEFwdbMcveBpxfhCF6bq8SLI8f2NeXsVQVXqVQH+V4H7KTr4CTbhlqyfUy+IUlZvmg9Mrz/iH
a6qRwwjQBycEihe0s/f4CcMsNkhkcYHwRHX8fpPKNHYuLrBISGZyvqG5yMsyyUQDcCThu2v4pOfq
e/v8qhLRoIhEQbQHhol+urF/unABivz6tGrEN9QrFm6F5zyb8ONMYZnvHshPpgwM1eoV2PKlhL68
iVpEneihepUD5sWrNZR488EJDaLCRnI5MeR4dvO/QUbt2FZAQAVvQ6oz1nZhOgv0wdNOAuPdbvSY
5udsTFMMjc4AtEoUr3MkiCHBNSvhh0S3N97UkUzo9JasY8ztQScd5YFK+x/5YWNOIl2tCkN5i8AC
a/9rpV+wiHjVI1fSHz/UuqQLWZvr1fo1Dbqjl0WD6GnM7ZrsKm8Lz6sFWkJuiXcxAMyTc9ihJqYQ
znbiuZocBd2mAd5me8kNTeENhgcLFzu/gX6NSbmrek18USUcm5FqaIOAsvqq4FvX8B41WpkuPaZS
ERf7zluRS7jlH06YjuN4FEP+SxM9bmtsqIzEkDKkLoJ7ghpIkRtyEjjiSZHBfH9D9kmjTacW/SzH
Y+m21/PgdXyfccFIq5d0+ackh34kr/BbWV0Jq13KxUc0OVI7gxO/Gfd36u3qkrPwpq0MhSgDWzj7
1FtNXbgjXxCkSuUQu+PibCaayg0Dsnvz5t/ogGpJKRY9eEvhU450bG1xrw0HzeDPdxAzBSip4XqK
CWHFh32wvDwNA0G09ZsVzf/PIVURB6Vadxhqgonyg3iD8+EBjJdunYwjbTagjmdYRznUM9HAsXEG
NWWeivnYmaYxfjMPlNe2wjtP0X4wBmS5nZX3j9qNlzUAI3ya3Q9cwkVjPLQqAc/VdMX5QthGrxAu
DYgiGmgIDhZABaivWkGxtEqTuaevX+gHbKEYRjPJjSepXzmNtaMhmgdLL9Lyu+ML/+29waVL818c
fqJ18xqecCEa5BtS8JEiZ0Jbfv/y6vJ+8JJoc2i3wjJ3GafOhyNRgCuJ2lzl+Jo51388QKx5bs8p
VdKEHT6+ckDDWEpjubYPbpYhDbyQ78eAP8rNq6G6fWSGmCf9PYjOFIxQKRxS6pgpBBhHK9bJhHDe
8zVDJHRO4IBFrrEHG+ZsnSEaJRB3J4wVJ+7+9dezDf5Hpu8kQ7EK6LJ4FaoGbhXsnrUBWmVyHBz5
QWBKlYWW0GohOadkIHajxIGHKhwcfLCa3ORqkChztoDuRXv/Zh8jt5RY2npxPFfYJ52dFZsg4oO4
9bJSk+ONFOpgFfTduSYFJsPnFj0o0rSD698vfDts/NNiBafKuZJwttHSnBrl4xIKPeuepMszke72
KXn9Xr2mQPyg/tpum1TwRdILScrIZxCgVrqnFsYpRXmGK3w9uBthThkBTgJnfN7gXczOzCmZsy41
TAangHyijdNNqtiyPjUqlUFKYs2AixEofI6mUGE8EDHnvoaTYIaygCZmZ2fx6pYyX63/+wveDmOC
2F79tVp4Rzs77Qp4LD6fVMqObT7IE75z/qXGo0XXnhxkD9dI7QtFbBSyjgrKZs4K3+sZxFVf6U3Y
+jtROdqcOig8sUKTCZiSzvLWlI6Okw4kGszeS9ILK38sq5bOZiaubyDnahCQOkhiNKWbTzsJ/HO1
bN468RFlrid90tXTtFGmJHm0d1g5lw83QB2BM5XAFF6gdCR2CcpIzrPRwAWLPCIPTApoL8My58Sr
g2krfcjBAidWuLVMarU54ZiG/b3nVS1ngNVSglV8fyZQQWI/aXD5fa5II5XbTyCNVY7hD7Xsibtd
77xwhabWwa3WeKdQdzwBHjesuXLuovAO3C0d4WAiGytIsv9lkmoJAWy/gGdmEaATkDOAMxRxIjlt
Xk/oEWTWhYRaP7165VaiqV2WB6nzQgMH3SMTCvdAjFl6By+qV7YfqQsGfjURoflx1Mr66oUCYlER
JHZ6Fq2CAy0gWkcisF1uKjjEHg31AZpkwlXdtIDTEG/Esw6RKOcYkj3cVKFJSHF3mMThHe0mg/OK
lZgHAQdTyt/gL2hkNCuGMU5AJP0vKS401lDNKyDk7eMwjXzCM7CFuQX1D8u9f8HrH0VwPzpT+2i4
Jbz31mTu0S3ziK4cSn0NYS1SiOmHlQSxllc0KjbhznqqcEvzFT56CavzI35pnH5s9HPN7V7DU2iD
nWquYT4CTm4jnum0V0TsLCdg53T9QCTZr0SerO0JDR04f++qs9wBHDPv3n0yLUG/hbOx1gky+5iY
qkk7JrAlgJ/tj+oLDHy5VVaRQDzQ1yiryukxHj5jOckRfZhFt2LB9ju96TNjICJjdkKUj9GifQ05
AOGXNzRcbxEVLLZErXiWmq56YAQI5nqe7tWMmSslVNsHeX39LyWs/QRiemiPEDHGVsAtS7ZcBATY
Z2oQvgRt/KjAW2objZaTSpHHaZqOGfpfZIw9eEjUp7HWCYedhzS9Zu0d8wa3cRHnWKDQnSYqe90n
Vv09c2HQ7fkkYa4+Jp1t+OqvTPAZ7CiSCr3/B0Gh2e/+bOeYlpbW9Pir3lM86kIfDOe6lRIjLAUi
dHIxSe+5mftDDxFw3iBAbMN9Z5l07CuiuHtR9gU3zVyxhyNeo+YPiSfoO1GknSUSIuMCzQkRfSJ/
n3X7NNDa/i8OM/RcwdHgoUEVJp4uKevoH0mqAT10XXeH+9HWKb2fFDN5UkOU4vTLN7EZYxGz5Kks
KQf7zKstTA/hn4zkTvlnSL9oyDuhsgzKn2gIwIHF4MLC8+rfjFoNLDwEoxmMp5FTWHhp9YP7IX56
amm+GLF1LNzKHLaNaJO9xgkgyXQeODUuZ1Pn/bZ81bwxt1Q+j86CFe4TZTPlWL+5ftiF+ucRZEy7
QWx3Pw8OQ7izkoZcNa9eel3ZVSxrcikceMGfvFolQsLVLvQkgjYzPsaRW21+gbVdSSIk3pZMpwjM
st4sD9srtXu/SpXciYvOYqPyw2syqlmeeBrbraNYi1A8AoRICyNGv65QHe43uB/BXwccyhgmsA+j
t1JA4Fh9yEmLlY220MGg+YWEIpgz2zgdAtdzSaEqcKiij+uw8cN+/zRBQIQ1L2Ysu1JQBUpSt2ak
1pgEefHupj/G+46QXiUWOHzEjao+rW+xcxvL7KEBlP69Nt1tRqE08PJCon4CMfyzcogqdDzw8MNh
73eRqeWgGJ2nDpDTBaELBKwFVqW/abd4psN07nz2XOxySYWX5vJPc1kDTnaYqVi909+7UEV+s0ap
8t3cjToLUEsC9XcG1tB6Mac730KS7l4jORtHXOpXDp/KAC0aT/ccnRmXhFAo1vsGrHIzPEzjUwfv
O5i9G36UChzIRtU5fotklVoZuZEuF9XC3TxDn6aFE+jUQN8wij84/xEC9udKE9JwzUeN3WsUdYg2
AkLp3RXommtIwYTxssuhjfTaohcagnQxWHtfDLZiQSzCaZMwzHBm9XiJfuoQJpock7MmBSLUdjBB
rg57FRmWTateOWLx0KYYSvUHWddcGOEBLnA2S1iKRj4dcJ20ZdfSfjAF8FxzK1VzBGcyzK2WmugU
M63rLrmpmAORpCiIvhoQ9pCumMiuTqPVz45+ItBOV4B3ce+dhOWIC20HndGq8uwx8UCIJxgu3d9p
D3VjWcFsdFFrwfyxfANEITx+xMYVTOAyy8UH2EEw5jyrlNSwTx1T4pJ6cR2aSfZb6+JLyWWOcDMh
gqHTzWpFM3Cx4cqm2fiEynkznzMQF4fK+1X1+jU8AtexFCpmzYBsP5YmVq5YU69k46q9reqb/DGp
URapQSpZpkErzDKf2KqcrEKqa1Pu9DbLtVmQRitkAPuuLeJFHbdloUtRg5Gx0HFnJHcko+SHy5hL
CZRnj43M6Xe77IfMINd5FetZ9bw90/pkZ1jB86Iu7poRZ2Wvioq4D/nPVraWBBudWRw3onWXfVDG
d7Cy490F4V6mf8irzMdqJNshUVIF2VgX05lza3ZU6AGlR3PiichdxuzJIfMAvnLNzNebtFfECwp9
ged+HwoAakgJYP5OgZIgJFyxJR2vXhbMcAPrbqONv5W3zvM68iiyB6UO8ONIWBelhbfWGrSOkNn0
u1mA8YTCQRup2M2c9TZZ1bdC7eeehuPWL/oJWbP7FuJw7yCy7hZAgEQSyXqkELxKYNv9RW3K5iaS
abWISG2sLFnGNgzt9XzgUrnMeiwDFnvp39QiIOeolYRvQjZayLwjFMfPdcZ9pXapIZEBmAy0L3QT
GaOcXNxSyv3xrz0yMtp4x1PpBoyG8ADY8SrucEEz0AIc9BnftPKbZtzn2M3foFj3351VAbuYsC10
rieyW4331JYleii4u9eH/LnYIxjWG7MmM2TENklMk8/W4zUVMrPXcylH0z3KxBCBvs2DXlhfRu+z
xJn04CmoIHyBL9+V4fdqfj7G57YvQdhsTA724rV4MoEXaV0Q9JsMM0kkLf9g+mDePnmet6aU69JW
ztMtUSyc+pz7JFAWTy6k3kecA70jPgkOgaDob0i6xm/u4YUYSnfZpnvlFz0qHmHp6/mwngGcgETi
S7LkyKlwF45idA7mQB8SSF1Di3IuTuUy7siPxoiWVGGNieCh1+8YEUYk6QsYJLU6Ezvo4OBdi6RK
pjF/Ynwq/xSbcvwu2jrqmzVOkqrVs2el/XxQHP3CPR/IoKeUARwhGYKzw1SnAUAl+6XNMX4sj4WV
bV/zp0MMEfR0Gcvcv7RmiW//LakajdwVjnZ68aKud3/w+7XvVkd4ishW4cSVjQ86pXGIC/QaNope
sSgSLs7bNL6gCDDApIS5B9KTLglCAK10+zQfHggLG35R6g8d5iAFEy6c5V0aggzxKSjY9dho7/ZX
mv9WE/upbv/RwJISsv+R7qp4xfZr0GtqhnjRMsYXBW5Z2JbXxS8hvADQfnDiZybt88hSZn4ccPGr
gXZ+myfwuMUgYuBCw3zaM3F02KJv3WPzQoU9TTNaBALzDvFqqdy5uM1C0PpjeDZeWZMUCmtI9eFv
xoxqDGhMfxLipWON9aO26iCdiblXzbY+XhG+R7A8B+boDbJgZ+GD+Pxqmn05xCpJJKsH8zViyy58
gCIZBGnsmVfAchVBn0gIZSJdAnFV0zKrOVbgjbIZ6PdRm4T4hZj6xROTW7/hF39atRyOBK6TqTHK
ygHL5PtKVSrkxghVlPAHtB8hLeME462waZw+BUMm6EAGtSz2VQwP5N9rFogCq5a7Wh3aCs9z3ary
bY72W2yGPWgUt+Hc1+DL0hgDcWWTWXFv+r+sty3QwGYgx6HxIVpWKLZnGR79zRxT6Ep+J6BAiyRO
yUB5EYsDykThYGT8hwbYLg6YN5PV+XwePcQMRK6ARIzJLVp8/qm4FTE4HbJK9m9QjOfonCMZXl/Y
E5AmpqNWHG5Q+tox0lNMKMarZcypZFKYV8udmt5t5hVgVv2jOKz+82i7AhJ4n+pEKGepVuXw8sRG
meH9k2jLdfgJWvjQDZbydlQ3rnnUWnMJVhbmtRK5W0drfyS2R/LpowoZjG0qsui3AewD/KTZ2sf2
wNFM7em4w2I2BQVVAx55Q8Dfi1btOx5dPpSwpFw3MMlJmH3dAFIHxWZcRlxImQnRfSNgbscB65Au
Kdx+H6XCk/5LQza0lw87AZXWP6Qj3k7mabIb5ihDIiGrkg5O3qDd3PjdSrvnJpv3pjP1SLEZ/s30
9+NPLG6ggTJiNoBbeBTZ0Iy2Pzhxt12cs2Ve6UgTr1njmX0j/6/IRh/hGR8NdMVWnBELeKzdYhnq
V/0/ZMYPOqtVNiK/15mdNWH+FcPiFfbo9APm6bft8epn0ACrk2ZX4btHgUvHXkYyn2rybmOWByQr
0uCcSxaSbuC1tfi6SKNFC8rxQyOm2d02xYAc99VfiUYX6NhI+ewThQh8uk/GsQPaxDjQ8wPBdEmo
8EqoPtSpHdORuC79MfRmpDsnUr596+et6k/EonJxdT1qWW/H+vhvy98MpjUvnjcUDSI9KeGntbOL
vh4kRzjR7P9Ar4LQ/5oM2DNIs+eAEYSAcBaQB/7ON58TakhN5/yWnxjIcIE8nFWN+Qog4oL3GgRh
blXkUWmyGiloxk9hra07WioLcJNCyvWukUB+414P30b+ycdemwY+k6XeS81fPFVRRVCukxRGwU2E
uwZPGZj0Diw/xGYrLynmgWBcFC5HtjJ6BNNPA8T4y+IjBJuIhAN1ACT60K6H37sHhSph6b832Ahb
3TiJF034f2Jto1O8V2sspwZuEqHDTh7peEtb5AmQlkwICxjqdnQ4cmbu8Nse/rRKmtajkeWVSE7N
g5yp406HrvjNcN+TnAsy5vc1bunE6h3+ixJkn6zwLwd25Xk1KCyEVJ/fQ/yOdKPKaUp1rlFUutuQ
R4Mxvao83TtyU6RNzU1BxCDkiF0ANYyReLFKL/rugSlaoTfggGAxP90P95I3C4pwaWodeg0yf9RD
QzaTGo/rdCIBroe8CY+I5ToD66A4WbcKMradcQu8YbtOGKqA1LTokAiHcWAVkP9sbHsV34ayjDKG
pQOnGUsZ8r/63YsY2JenkJiBROQglY2lqtil63StbT8fayPYDh1yNRdBKc/xD3WRCbIF9bYIclUp
4pRwzDVV2TcjdtPtfQluu4LFflL1ZTmfBWp0UmRph0WpKkMJjhjQAyn4COv7CT922PN7hENiv5Bn
A3jtZ2ITU2j6ir+fKwJGixMKLFhwyws9tx6YDxIAg76TGkmkNWBHXti1LR13fmBJJmQnuNWvWHmT
hwtBlCG6iRiFU7L6dUNuI4BEqNuuDCmYo/RVAevkpfBgcNnzppakwypnstEZwEIMPOQfJ7oIj/bt
n5leBQg0OPqoO8fDDdDsrNQoFWcptHKf1VigMGehhJw73J4yLMbXVmouMJVCq5NRlQ/98waC+4J4
bR8S1dhwMAzToNnMDgv3Z1pbaJioFiKCcR3X6dzPcRsAcw8eNUg20TBgv+MLOho1wCpavyR1RwPG
XtgntdcnAQxEEdnr2notacLYqwttJz6YDMGL6kBjKlyZ+Ud6CsDFsllThX+sJlO41x1l8e7nkuyq
unEW30wyJX5P2dvNV1dIlm5ne+6oYgtJFdFSnArlP7apv1TvGiwf7JhHEuJzJkoDGNcPpF3vjvJV
fN8hOfqlMGK/T+Xw+TsZny8iN6EzZ6d0mQadvqovmAttwM6p1kI8R9e30g4X4rJB7hkMLRNZK5Nt
wkuoU5O+N7P82rAHfRTn0cycWwqRCeo4sf7vAAbRxyNIev4zfPUsBES74f45rOC4739LfDld6cVh
OhHAJAbgbKEOZwwN6tJrQvobN7ys4NUrLrE/pp2VfC1WC9W2NqAEtf3kr/iNYwOkFGD3bdMlScwe
wVNGa+YiRdEeNV8GCtx4ZACVh1HdE3kjQij5l9p3ukyxSSWid8jkGDrL3WtZXllDVrg4kZ6kcjZa
yy2CwTMQ8Ad+tLo28Y+ucXqgjPL6z6orDzoOx2Et/XrXR2dT0MmhBUkdZPj0OECO4Z2FfZXH/JiN
tcn/Dw5sD1mSsNgnXiYNFl/rHMBVrvrmpD5CiMV4Up3P4Vx/NEy+6L78Jf4zPAsMtVrhfroAr5cB
UyP2DuCG6nkYuXv467fvmVyM1b/AX6vdZkoDbekiNWqsOcMl6ilnsk1LpAH0JhznG+dpElK8H4ST
5XI8qKHZAaDzn4DNNloxMBdul1wRJlYT76fa6ICmPZjSN9J2ZPp4ls5aX25UM3R2XzZp2ROuTQsk
wtHRwOonJCZRwpemaq0LW4n6DES4nVessWthZGRTOETewnUCj4Rwjkb7LiqtzHzs9MS+Y27NVEDA
2LPOywB+81gVmYqXzKj6THzWn6nIrm8LL8Kce1H4yR/v6fTm9LMkBs77oskj6tMHSXMQPyfN/sf6
Z8Zs/NdNlc/VYgIOzneqqmCfAAhI20mf2Y7xr/e1zhajk7JBRT5vOov/LRSN8iovitZ68WxWTPZj
SegaWkrQU6afH76UE9GYvjAHgdGCU0SRaNFPOOHK+VIP6kHaO6lTlpiXkCb7wrnaBTe8G7/bKiEA
Z/bSNIEqmA3q0jSQkY0JKhI/s0TkBOvjghU0T7dSAagjgGkWv+kB3kZ7fZ6Oq0lZlA5aR3VFijZv
666evdWPgxF0PcTjKQUnBA5sbZaX3gihKqrbuojZ8jIaK+aDjUFhvjbrkujJaU2esQFz7cYgsJ1M
yhGCYwt3ClAvN7XVjHdrJKlSWgpTujVyZoRYR8JWS9BfgAn+b28y4kh3mn2NAi4Wrcg0q/o/Hc6I
k8+8kDq7craZgO38j5s3c1s28OjiBbqOnecibZSIqujJciKUVriZf+zayF2sPOxyOGHLfZbiRK+s
yKjOphtrPmhj8a/Mu6aCzVuj6HpxXBIEeWGwYmbcLmun8RUsB5H1NFmqExE/5GW7YA9zfo0/hsIB
iUjR59yYkqMdHYMVuxKciJbkG85rIyW6Q3jrPh+owJCAkAPjRXJiLxf3R2Jpglffs0rfeI4wtEyG
kEooGp2mRO5JCthDFnrsmfmbtX5x7cUKKqWXivaGLAkggqUFl6nbpfrFrqFzI4f/p/l4nqGNudDN
M9vTgAgR61jxXazk8WDlAxmuOrXI8XswIaiMDttihCdtRqQPh3Rt/bTf0oeXfCW3Z35KCl18Xxml
GTTGY1Q3UfUzgCVNvJp+iLr+pOb0qAtxMIbk0bqtrTvsWUEWCzsxpAE4XX0DVJfYSfDvEb6U/6nq
TUx7jeNkhm0jDvCdUcypeeMLcIsGL13USvdnlApeQPO1Z7SWPHAWx4KYDpDcuYAtVeURnBBxsfFU
M7V/cAq4fDc49D65mO5sfMTE/ZuTLLkgD8e65gzXEmsyJrtOr/e7qfN8tyoEDU70Gm8n+bbx2hjq
/TVyT7P+5muHj/YfBOmkpQge9SMZo+fAH/h3MRrfU4dyUebpfWPsE3n1Ip1SugSbyyEqCBIKIshh
gzpRTjj5gyZ3O6LkEn9oCtKtjdXU8q1lG/66OyBCLdpzf4Si/gc9NA3Hoj2w4l8BL+dVc6x864+Y
kZh/h5fMjxoAVNFn8zyijr1qdWTu+7SqOrjCHsY0ICSTK1xMyJUaY4vQYiWW7T5xXbRzD0Wq2XH8
k3dmJhMNyuJbPumTrw/eymlNZKtF01kpsd3h69I4pYpO3qS6PoEBgQYNtsvYNr/e0g8CgtUcKViV
Vwiawdpt7Qd2QhJ39uffWqpKpE8c8mRGM/eQug1XZJMZxpqs0IuUkwD9bK1aNGHNYJVYIR1hIxVu
SCVMd7WEahZnVAW2+N7mMzhpfLqhEp2K9Il15KENAnsZ+IqF93gTZg8Bm+LhlqYKm0cWUP9Y/dt0
03o/NtvCAW4EiQPxM+CTAcbqR0sY1ktAueTFb6Ff/jBEJ5bLU6ArugBC5+MxfJjB33Mmqw3uAoqh
G7BpePgv4GCyx1xL3z4HLY7Qf2K6n5N1EChs9UJFZ/EHKC5vLucsqvzcqWXkLozP4kaSO81dviLo
EYjYkx4cLh4Gjz1OSVQd/u2wXE1j4be/L4ee0bgcr+/uAE/m7hEYsk5iE2VlukevTE4+6gjqVUNy
bxUrO6/McakSCgzgfZSqMYfNrl+64vWPM38O39jN/6Gitb7UnBBSDzQk3XOtW3UR3lY0QPox5wef
p/JLPnw0V8Ca50pgza+oocDMlYPra7RAzXu+Bx+3ZZWiToBG5CBG65cCzAid0L7iXNygRwtNQJw7
qVvKBmwmMYdV+NeUcwcz++FfzHohvUCpWUzRgn7Tkku6sRhXFA/Hr941y3xOFm02lVeBR4Wgctd9
P6l+S+ZV3zpsY2CcfqnNQQsQ1sh5zvvp3/e0tWQ8JcFRKuGUEtNZ5ZM2t0TiW60r4EPa5OX83Vkr
qJOXePrlHTbPddyLvHpGquSenwhhD161/A3fg7K+TMyhA7g+ibdr7pjcqNqL7Q18J05LznJPOBlP
70Gm1J57F7LyI8YigV+6dAvsUVVVuti2cc8qwSWBB4h151riNiWQdduzpZfsBtg8KIs1V9E/2UGy
iy9mrwImN9e6wIzHgJtcWb9ImnS2Tdly5CLY1TwzEyu4g9NCfEvxTsPUrBtlHIMZTBUv2U3pl+oh
fIo2LdXg0d/7tU+lXLgouMi6tJAHea/cV3agxsgG7Heu/HiAzaB/HhUSPcV1h7UN02IFOuKumaLb
DtlRWnqLLT++4T+gnDhgv9EyDrla+c+F5Hj9Hvo/UKE0gbMAiDbBmG4A6rPaHReI0RjA+k8FRnM5
pZO/Ye8LIHwlGx8qWfvEMsaHED0jmdkum+GHazv51lU0JqaTEwT1CkU/f2qF8Aj2wIzuebk+d1VV
IietRYoiR5qOdSdMacDL1XL8KBREFc7SzCuZios4gjRa6KuKKu8a3AcP/it20G8tCjQjTGmWruZD
zct24wYEJCgPuqRoaoOYkAUeOpVaRxAl2YSQoV99rWKpI1olmAaYX7pvkSpD1IJqT3hpTKh1zpT6
vMZjVkVJUDiuxJHnVDQKXDZjk1b7yRZyVHd3Jw1HsBTtT62nHLeyQVupYNXU7u+PfkDfcA0RiETv
CKvlsKbqyCaSlmnM1TytsrO6h2P3s844+3SA/aJHqDbYQ9KA4RumPR4hGcbAk+e2rQ0+GXDvrfAK
J2b2Lu07wltEhnrFUrDJ7MiaF3QTCC48jwRgw+l/efIL5VZaI1QNbAHNlauhDH5Q/l0M2VdpzMt4
+j4z0VAs8A7c77O1qqgTP8ZbTZzZ1twI0T+YZzMA+LVPyUpvDs9kfcfoKndzF26aN1OPwxMlNys/
kJbA/LCsvQi7SrEsrUmoY4RwMJvXEvKw8JcOFsnvtPXgDyPo66duQSVcCayG/mB0hFeAewxoTlZ3
KNcE046Z4gVy2q6x3xNC/GlYc9RwRfPS6EetnZJ+4Br+J4LYkWG5VfO5YiWJq35UvMIOSoHhT+gh
FM2CzuFmfli96y1HjxAq3hTCbL2JIgulk5bvH5IheNVS997ac2BylYXU5xEC0oV0Kj/vVWpwZujC
t5XC1Aj3XsX9O5QwKd3h+P2/nsVRkTOwouvcCexalXp3uwggrTITTBlg5ZGnUTbJZRLy3kDJtGAL
/W75THABN+mi9n1oeyl98hGVpil+xdMnrcUSePOJBJm3mq66vz2llSX3Czdg5Qn8UG56gZOu7bj1
6DpxnsBEUEVDp31J/V0YaKPYDZ7anAcAsajAnP4yxgaE0QbvQYoQ6mw7kfOg1dHrqrRCq/v7c7T6
PeztJF5PQkBb+/TjjHrdiMEeOykZM84kWJLI/yuVEJPvKhNRaoUA6MFOy4iv1xb1UQHrKyMwrH5K
Bo127IiaMBYTOw/4spcvYvSS8lIMiEyoG3HAkDeTQaVfKLYQbFqMkx1mzqkyk68E+WwHQfAjrot3
OOPdMMnmvoAL9bktH0TvlAQG62V+qjoqRygRkMXy5xkmshZDl6Mpt+RQdCaueT0rul9vMkyhPSHr
syFw/KgJDsmw1V3eSkP5RA7Z2SM2ViW0BatQk/u80NyTpSe/IqIGogA81n8xtpunC5y47j/EtFh/
QtbjZJkpS5rjQmL1Elms3UZN7D3gAftGhzLO1gXN2lqeluKiPIphP4IG3PWhmB4HkNm32DqodBuy
YhVol3KawZ7YnlhxtKvDknYw+Byw866W/MG1TBTLyPnSLmAZ/6Ws1sj6JUSZ9GLc2RiEOMMpTuap
qyd+RIkzK/4Qno+iEOsdBB09QPn+27blwS1x+Gnxhtz1FavFrKU2wLwMbL3K623NzIXx1bxFjlNT
eoDjtcopfWtz1WshA+vpU/04Qe8SrWKr8k7Qlmz4o1OghJlyMthJMNQCF3DJ3VL5B9qp06JAw6d5
IvP2+Y2m2oc5jovDllKbju3YoQ4xGxGJAZpqibv928aAt9VBON+2JKfsWRzkWUAQbjMaEEh82kJX
93rsgeDbf0WshPaYBaWlwLgC66SjW4PUctm/kyZTrBeEUVHT8ZMuSCa0H2YYHjXIg/RcwNK2QArl
tI9sCwLpK0e9EH9AqQqhDEJ5/AJ/QnHcSlnhmxClUkR8ZWsSJ0vVd5bp1Ii0jZd3fjEbtkJP7/W+
WQPS48+ns65rrekCEpe7pWcgJxww9lhAyr0YiwUNB4igtiHBXfr44P0AFcGiqPfekGLvTcJ3hxS7
wROSq9DYzSALWEsRS6VHhCXNLZD81VeropngA/oWuFcBA5SEUTUqmPFvS1RhGlqgAo6uGxoK9JjP
tpPd5X3Ze6dsig+QQzhIh1j7Pnt0v2nAtOaMIZcKGZtqCwQzvN+TFX5dCbkEuNh1oD9UcAnQ7D/x
aR8AxTF5elzXo9Fz3ut66/jOE3XLNdZdk5fSAplH6vpAiHmxGyC9Xc9vAGOgsPx5uCQZ/cyk/VZZ
XzOZZqrK2gl4HhUaoCEhcdMQQ6jTMFzsOksRdOf1L1NpgaaLRqNKNM0NsmnIk3OYeHIG6p0XVpw4
wL13YE0xDRm3jpZHQMCniLrx04ZG4ZY+XUOhYc2QGv92TB1+kj2dPgKZBEpCbSElL6I2B5xgCcGc
7jB+Cx1y+Adk3XD+4L1oxjnx3bNYTr1uSKGbSCgYqBkcIMs8I4y+YKavxria8Relur2qETRf3mo9
vN6vr1NkwaBdUpQWbIc1erQ87+8cXIsTseuNlBjJCXUzm+uUrlasXIQtPTcPpWq1IXtu8gu3BGRr
BB2TR7naTf3EH6tXYhWe06GcLdKK+NKrwq0S8vcP+9bPprvNBWoOFuCcYhaIVOBeZ9jP/Uk5epcm
Y6N2Hw3zcNOK/AY+qnxznCr1n2eQOgudCZjm86BAnKl6NCf8NnhYe7J8EczAnoZkbdx5uYH4dyjM
/imFMypRlu4S38pI5OjElzUSOgbs+1CTmwdbp+Hbl7PqMpFwTJCEU8Z5MOODKuGQIcTqZFFf/QGk
n+XSccQ+d7853ZjdHg+KGBCjxxjGDdGOibcuud8Cfv+bCSCWCi1w/JtL2+0orkYwZKWR3hNrrDke
n/m0mqWwoc+/w7BE2hqqsMqYNvAgip2sTkOv2AbyhxHQa2+C2scgz3Oyjz+4f3p5bfW7vAlkFqIi
vKMePEltfkFjMqynh6bbHASyZTAuwYaMzhclsYu5ZgRa7StOrEANAeRa7XLNedlfh+inP+X6yLZz
uh59G81/kwZIIGg5K/Hc/jg7SCnnY6JNCjMgx3TLg+PYz2OciT/D0NxPXKfDt+RDE7iJAAexsUzS
uk+UWS9Ixl0Rqd5JG2eiF+epiFOtgsuPM/PNcoY+oFVR1HJ0ge34fyKMR4RwSdvpMROIz+x+GaPG
RiCrUMzvjcniHvRKcWRuEIw/CpgjttAV87LEBT95IJYyAtUOjP6lmfTVYwUFToSpNV/II8fJ6FbP
u+gE65ZsD31Kt1uCya4x5iNArDmc4gNW4bWSR0r2YyVfsTEQlsGbzTQBQgezTuJ1lenL/8rSD3ZG
nJLSeuAcC1kAuNa8ei3vwSv0za9Zdieg67GLQZ62ZRRoDctTmOELlgqBuNOyPbriuYDZ6V3B8EER
zOPUtoECXELWewHjyv34X9reIsnyyj73l2gG4fZv4HIdHfAsvXrgwLG/yoqbwaoYg8aljYlDu9jh
CpDPE7vC7IU7xfczpl8ZfuTprJe26GvHiO5YziQtjn3EH6pQDikOCB3l8moyPyd1ZDnSRMD8vltd
Kdkv7CgFS623aELfzaicJ4WHDyQUkB5BgzdKQRTCl/ZGBSxckMkKRPMHyI338KLp3MBvUhK9M6Va
pfCaFNw0N2aU8bxZFhNP1gaeARdBOSRzdMT56hOQKcKeQNzuMt74dbugrvR58yaS2EQkhAVI6Jp2
gnd7JMEC91aajmKgcta6oH4FIF0p3dVqsQF5uR01isyIU45/Dm+1Srcm/3mlkWXL5q8jnlbYTVGY
M+yPGyKmQNE8frz8whAa3NSKIsUEANOyma4Mqc4qv6ZyAwAgTmA85fud25nErYiPZVxP6yD1iIX1
uw/lGXWw/B7iFgTG9ni3KrMs8Vx8Mzfip2orvagvdLJUbi8aLEiyw56JhEnHmBsOzYvkhOqz/qmr
DmI1deiJPzHa3HTiYswfOzxRvGZpZdlr4YvHDAdarVF9ZWm9thxS15Qx58qU9KQowiREEI2dqDsV
Cf0DRAPbYeqVs0eBLCQFCc5NL//u2CN1KRoHB4wyJOinsSa6vH+GmehqaskGiCAeg3D42LT1Xw40
eSOTkCnLSF3avUx+qsTy1/hFGmzmcwnjkSsG9+W8LuekHWv6pMxok3DZXCgM2/tT/vxVdqMNAIsy
k0b0TCEri6TTag4OUuiEnZ01iBxnhmldwuJo9f5L8Kuab/+CDv4NnFfseMBJMsm5VSXjkCrrxxE9
DU8MQ6lviqQ7NHMajvyBCPP/rJ2rg1s2ABxuyWQ2Iw8vbCP2S/6K+kmWSjdkt9K4Yb/2SbtdzSuj
HLl2cUNcN4E/OJ0erImBl0jJy9fCyHmjhoqbSC+L3gyDZLCZuLZ1W0RoQPpHf0Ny/YakiapeEH6F
LJ0wUVNUzM4fV7RjyEEo8tvyz/mSU6gochom2ElZD32DTJP48LDNx67+L+BmgDeYUN9eKjZQ8guV
GP1sgXP8jEBW2JGKypmoS6Ub/ype2pCZHyHk/fTGCbCRomwmbdPZ1CO1PQhDhWnldRHiLWOEUOPb
/GvldTxN3BUX8xdY0GIqb9/vIuqDOmQPiT2XNziusPiX568GRLrNgv0yR6sE4ww3X2ydQscXDObm
VwUZhmFTwtN9HvGbBn+Zh4efv2lWFJQsGsxdn8w/DHE+7xLjGivNoTqPME7lO2UVua5cEjsxo4S2
gFAsrGgiLlHLr/sqg7/C7QAC2yR53Ezxgx8IJ98nus3K3dIsJ8H3AUsvqIj51VLL31ANezggfdxk
dZ+e4BzyYtYjxlH4UAY43N5vAO0EnzX1aJPsNegeKSMLOzae2BTgtJJbts1vWRcCQfNblmHtAHeT
LCGJwwKRvUxCcXVOPXmofzPJiRxRr4LUUTGHHiy02x6G9OmiCmFE4dzQvuqqVQabpccoqqEDgyxp
TsBtsimcyRBovuwsbWL2FkB661FcbOq1S9psCclIo5qiTiIF5NTi5y+uzX4ULVB+jn3t83KSebwk
m0Jzl+q4qBxoz01/yeoPf+F3NF2nSacqZ/wCCZVhgjQaQQVwn2zie+nnLWaeTzihp5YYH2DXt7zU
VaYAapH9dukS/yWd19ZEGbIxxmMrTU83eWZkK4hZ4QS0/BK7XVRG6+gIhjMNyNja+AdnZmKZJOYU
OauKC0A88JCcNgM7jU6VWVMrUFyY3vnx2HqkZqD9SIusVTU4iH74c/qCIL6QbxywjVbsNdSsDtRg
8hxvO6H/wJdV5fXVXgz91Ty+2Q0aBuvOV4QFq+VA6yRWdtNJ2Gl0qlgGdVYsybwJVMCc8QhWD4C1
0uE3WCBcsNjVj6L5NCYh2Mkn7iqrVQlJ6FLijMTXMOFFLbSUfSF7H7vATj0Tl0oGZlHcK8ao15O8
tKTcP4VnMRgdhhnbf4qS5dyyz88k0hz5JdRZYSXasbwQhzkNH1CfZ/Iiw7MrwMUCVcoDZSpnqAFi
hQx3+NOl5hqvfyU4xgM6ML/hZE+NkQYBiqJGjbr04t1HkFYePxWJGIXFh2TUGMVxdnmYiYdlEyLz
sOkARpJqtOiJNFuSd6fWLjj518NK51a9rEPjiDNnBdYRGlF8Xw9cCcJeHyUJIjkNad5ipop5Kt49
cS05gGoBaG4Xbkm3tRPj2wUXlDCUUIZV1joygk3nCuxNJzKpSrIFjdqJEKIVxnpxlDrp13OYwuGu
S78fLw3BzbYp3NW5WzPE1F6MFg6sCVOgE9EnNbXrrPO6jv5b53Xt30fbvdJKaWnRvoxt7ALSD02K
DiOEwGVtf4Z5peOSQYczsBHTxCCsKY5VwMnJdhwI9WHG2xQbmoxt/ozS2+U459TYAt8ZoCI32+Vt
Wi5ciPhjcQeZZCIw9q3dROwbMbPkeiLKYHuBhFwPqd2Gq0nq06N6arf5biVnAi4mN9jdY2en1aEF
0b6DOa/WLfy/b/DTCyaby6CbruRv9j5OO0Q9quQYB/oPFWrl7vr1g15GSunleNwb3+wUAFiNJR9O
9tudbeDrsYQLhBWGeZEoXScWh5AOoISMFDEJ4MbEYepWJ8KgS4zCQiQdi/f43/FzKBT0/vm9z0/7
QZ6lk/ttPPB6JvEFDF9qi1gNfYwJykawGzZhqQaXztTg3Oozw3WSXCfC6OtIz7cMkZKT8IzoKekJ
H2EENnqOah6IV29Yd0e3UA0JE3i0CgFmkqBMzA4MXogJAwUJiyVyJazpEahs6YrpDsJ15NVwsnAK
kM8eU2UvPVUy72W7Iu46DaGvWA9oeV0n81Ksg99Xte8vZmpZqOUcz1xIKfVpzSdjRxBzZWMmUM+P
B9zv30BOMr8EpFaxRy5EvREQK6UW7GvF7vB90grE+rgUw93fkq2wZe03w4cEZKS4JqXA2pxG9TMv
XixM/s0t+OPlJ6WGLd4AFviz4Y93fdtdeaebVYWLiS8eX6ewfFbXBOFB1cWgOofH2QU4MufcsX9L
ppel8aBCqEGCW+MZVhcw5CRwEigo6ijTvgx+SIr1mSjjDbze8YN/9SaXGUMcVsXlWRbNx2FEdqsD
JJ/wkUTizEnfU/1N+zQYnZ85/Wf5xa5QWRiOf8KJhu9/7Ztaurmlu4EenahLjt44SrdtUIqII8wc
1tdHk3M+Hv306R7l++ILPxBcM6hxDW+57qr3301CytGaV8PzptxdPJxPA076p0TxVbCI8xY8bJ8Y
Z/hBonwSIRj9jve4lWDUzWJPjT+SL5HPkfMMQPmzmY8UaV9uWYd0DvuiysrKrOfROzjG/XAL62He
Umah+8symjNMx+97nIIwb6VRQdU9l3VQyt7PKPGsYhy+H6eU5Qg6lUVE4E5wYDqvyG59Kk3WPzI1
K2iasJrBrOdmRPCbfaIlcGHIUShabQz2hq0Pk2ttuwmlwyHLEdK/Oe2RuY00AreStTwfiyZ/IKC5
/MXulwkwXsGlG05GVMCQR/Z4PSDv6aDXxh28CnVx3y9UFllXzsocdnQPc7MME5RdTbUhX1q+1fva
L/t2c1QLWzzVxvjSF1c2nboZl/junHwFPFMvxg0PnV0FzWxytlWKqI6JT0iWhlQgoX9wUZnpRqPL
MAp3gxlkXuELkbxHqBlmMoVQrn6Fw7cAm8eeBPcSbNSfi98vhDwfayI4YgAj9JskHe3/1K+PYABp
oe4qEu1Wi/bbnuTYsJoXTuSvpJOI2PkWuGjSxYh9ml7ZaJ0e8BoYHHwsiEQU1oZEUuClFf1NFvJ8
rf6R0Cj25GvdDbjFPxRDN6LtyDirHpLMuI4id2Arf/sb7pcQsbK0sMA7OgkwXLulwqLKc09+HQe1
uIqryMlsKGtTUkyP/uKc6BSlK/3h+uVmAhOJn+H6jpCemrbT/vj1k1+IL99b0dwwISBPzCEYVX8K
gP0aZi9+r9l8LNCTy4Mkco4cmAHOb7X6AOeTAHB7+g6rTMM+iq3JM/SsBz1xnPdFGCSqK9CDg/QY
6gq0RSq3tXqz+o8dMnmDp3H5wEQjZO7O4TrpJNnWw24N2KYqJfhZscaXX/PyxPVUySfrKZYz7xGY
IasbMgwIGC7QOPww0YtXapdwO007LqQ6bo2tLfkiOWUwaj5NPql01jcOxT3ZhbDVcNM0BFL2Kuqx
jzwo859zPBaWZ9wfZ1XPse65q6pq5kf85+e462EYq0FF9MLpdhzUXgtbdYs2lEStR8Y08g3rz880
xDVDDs2/qKSm9/a1rVArXIN1RUxEFn+o3K3uGvxqYiFtpOqsl4hsocTFMUqPgWGQuOWeNRWGHWQu
5f8NkErxD6wwm4JMRzC/WyPRGUM3yVHlvC6Y9wplGC/2YTTieSdVd1Lr1A92yov3k3kPO67hh/sp
IuyVe5414PPX3ME83pinlS4v+pZnz359a6PiOYcLkmhDSpp2qlo69UizUt0KeY6GoLoYk3HTxNei
xS63xbAqoBWmT2QbJhUx5R2buLs7Oe9Rt6FQnhmDWzpH6gFG8mdJIZeEE78ZYFLiQIh+XpfVWr3Z
7Qr0xX4+U52bGL+GFc25tNJ1rCgfqOfPhqdhsZOt8D/x8ntKw64rMHq7Wtge9oB+Xa/O25l/Rjy1
y5F7bSFj6NAfLSlT+EWziXkpjX74UCr4JY+YwbVqelakL9d7NTRhLL8BAo2qG8dtyQG8KcFCKH8Z
RQRFRFmS3QAhapTFDmcGnxHAAjH28xJnMJGH/RC8wdTKUJPur0MlZRxt3SOPUY7XZwzr8BSZd1I/
J1JdqfXDbh9NuGClCDj5G4vIrI0uuCCpvzTIhU33S+oAaqoU1p6saxrDEsGlJ9cPvBxA0Pd8K8bl
WGPgZpCyPkf99pdex8lQXWFsX2hBM/xq9VwU/MIKa5DCCZYTS0dWd/fAcKc0hIhwLYyiiYW+Z+Sp
CnMTEzaw4WTRkNxFmki3iZxnKN9tJmNhxATqMFTMuCIdS/X1gRVAG/HH+JxPe8TLj1NX3sEXwBkf
4ndegD48GhWYjm2KQ7cXwXfRTTY6DjtdUVVQ8GSB5cfoi25H3AUtrCh4vqUTO+T7QjF0ipjPrg83
6wIYvmr8yDTc3l8fEBrsY/w3ERIQNOpr+4YT0f7FcZL7648bwOnFTTzjbz5FVd9tCi/r/7S3ThA9
uilL4hkCEAj+QgCJa1jVx58WMbmNdVvH1Z/VPHJgs4FVOs0jflZZL2Fqn0QKv0R6vLsNRdtlTeMP
4bELM8bvXI6K4nBeu/DoV+N2/jnos19cco8t9zI81B0qO0PqXc17NOtl4nkvzHQ1dROPOFT6Bb1t
wviozUntHJo10e8KbZBa1jHLlF1ZhgiPQqJLQgXLnjL5DeemS7IMKEyfNwiKLeij683VuimDua9F
JRL87jgJGtDL5dQC1clQbZ+VXeP79qEnxiaFyGyXNQlVVywR+PFsEv8c+Br6TrRf3EzmXM5mp3mE
YXABt6GqctwIohHXVghUpi2HS3wOJalq3K0Hq0SL5I2e2GUHaZ1uYbOS6MixIketpIxSOO/+F20u
YZbdKkb7nQWHGDZtqwQ6wcxliGwiupS9uVR8bSy4pp11WQ1ibzxa0zl+LqxfFWoi19fvFK6W9Fcp
Lz3Y2E14WQlF71th4kQhc4Vmmgwh16HWqw2UYSwABO0O9NP/a1Ni7zOEn5I2nNTYRiAExnAaE9PF
+n8jWB7T7ih1PnCEeCr8nt051heqQ7CdkHCMwFp1qkMnlQwdJEzOAOGxB1+gw1ViE9Jd5eTs7jQB
ixBFVdoeyHWOoB99P6dNOQLB5eN+SG60rHQD0IZeFhGqHtcWtkqRFDDbd6ywBq5rsxznBbRorkWx
UoVaieyRLg61GfgkqMDyVZdFoZcJsCxyo4f2JkaLkTgh72gLV5xPY6oAfw4CnzWZiRsaowgu9wLR
fT3gl9HlQ85VcZW6FxsPTJsy5yWuwB7Ger+PCed/Ump6EIrPzoJZL4t/DuX1scLSheG6+yCeK2WQ
Mlp0lZ4vPZSHEJtzKfxC4xn+AHuun2jeHM2khnQzoL52Vm6wI6jemVxQTRZlS3mvrf2MQzCZ2Vfr
rqSR9CeA/RAvf3q0fqeyUUpH9+3qAk7F8ozoIwxjdKd3cLDYswDC6DRdket9yjLkDR7fnPDunpGe
lazsCdBaob2Z8MbcVZcQy+bP6HBtC7VGJIX+VOpOT4B7L1WQ99BgBlL5tV5S+W5XI/i+2Jz9lFuA
m3PXyxQuyMMFPcJe8eB5BFblgkG+XcunRNR1nDNo5t9iRkpuHi2HJHtZ5MQyYabfwvVFciKTcgmG
jD5tth+BMkmbkpP9NrQEqE6CPp+H9TVpIvEQkkYuujXkPyLWxqFPcId2AEvktK9PhuhdztMRkoW8
Cg1+yd4InTre/TOTXTaNuQO64kAQEoHthrtcgfahVJOOfZBgndVJtOU1Xy2xeYnw7Fo2T/N8t+zd
EG/GWXNh3e0cwGu3iKYI9zh1UrxkL5cFeIIPdtn6kwj+M6xMhv89Sa77yBP2rKAv36clb9QhAG1v
Eh2bF8CJ8Y0qrHW8aTarZA5lA7HhFqWPbpgodB914t4mNDcvSAFyEEHiwEDGwiW+LCiY/QYlsgci
cABrGQSV18l3pd385DgXF57S+VsYTtlfj4wK9ykPj/BEPd2OQyRZDCj9ErolWQRFtEZc2kKHQS20
jJRkqufTwlCJJcLHdezUT2dxjV5lDjcxUTROiNxDcwtefbzbxSuV6nS4D5jqCt5TkqZ4+0K9jofC
qEDvcQFSg3bYkRYJhHjWeQoCyGcxJL7W+WFJfTnBgYysj+NMW586mtQ7p/hheh3G379TN7W4lnSY
FPUqUMai9zeAy6mV3o7pFD9m6sbWD67r0bTJ8a010q0gdz6C7TLcbPqbh2PofS0XIJ5/x9s9PcyF
UZboJ9mpDB2/diTvSP3ekhU0Jk5N3a4CnywzHMKjOovfuhKWJ4XOQ8T433lqmyWfUd80BFD9QaZM
p9Wit5+WBEavKXhTUvZL/gaqJ707rOAfrFlbQfm3h3+RsBgZAzpn57zrDQu7FKqRhBlUgAFChemy
aFPGA34mg3mK+D3N8PkIu/Ra1hZNd+jWR6+ADn84hZQoTnO3grK2LlxYAICpoFeeXENp4cpaTn4P
rzfi0JmT7nFjkaMpHWZR8c1iRi7LhkTvzsJMBBVglpVEhpUoGr75bcW21fuWOlmLwZvGKLzMpmCH
VwM2g7GeLZ5i9qteOvouSAOq8T6122FZ5mARay7fU6OY8GsjrYrYeIWPDnutTQPd8BhKtyuKEZqD
ukKgYq5tY8vONz2jCSYnO+xfPpd4qE2JDfewkZwY1L6QYncoTpz/2Xjo+B2g+fUw3r5kraePidYd
WGI8HQ6SI2wCxEd69K9MKP8urPu1M0UOv0c4RoJZM8qK80tzcuZ2k5sQKirWP0queo4fZsraxTOt
Jq3rujshQgEHECQY1KhLuOHKJXgkRcGkXoiaBFjSWBsrWb/DI+9X67CZNUZmZW3/zSp/obYvd2Mp
d8nJttbVmCCLuEPN8+PK/QO/7cOquVg7ZOCxNqR+s/E2MfcNXf7Dt4fH3YhQHW9YTkFlxJ2R+a+j
RFJfeqkx2i92t6LaUxmneQKgfakuLrW6KsVIuk2RtrgxC8NalgeOyoeL+/VgrCPVTLAKykDWvMBy
qyzAwa0oTtqRhjZ3ODflPE1WvOjnSxRl9SFrq/3K8YO4yIN+XT084dC5o8PNcwOqoNDRuXrEC0Ng
ofa7Qm58dB3KlIYL6VRby/64+223SuJlRiq1pbUU68xtps9Hp1BcxvAE5jdItotqoXRF1MQ+uAcm
QAEVxdBh/j70P53vaZp0EBp7mhq93aGRjkVpYuh7uo1NAD526ZZieCjtKDr0hFtKhZHSSZiyBxQO
2WLKLPkGw9qNPq+29paX7p4t1xg5hhc+GZLJI2gtNumZdTQp8/027x5veKlBmftGKSVMvSX2B8DA
08XaM8VtVf1bfLkfGwhMnQOfpyylmE0E+P07qcly8vf8Xo4L9yCMEXaLc4UKZuXkui7t2vHMLswe
cRrzU9DyJinPYO9drOTohIM7eUWGTblTEm4mPBAPqGnO5719j39VHef1o3M7zjcTaThK86xcqg6+
AQOZjFuNRsAAbIKzSGPwSw3di0XFR4nGllGRA1D6BQbjIIr7ZmFZPCQJwTQ0hWJ9WyfYJ2l5YdlK
b4GBZhvvZBMd8/f90vcd1yIVRBxyDJDRYZ/9iaSS4tW1d0GaDIb2CGlIiN6hWnsvUPtBSugFuAUB
5mhSXkIjDyCUWmrj9Mr0T4bR1Cq8MEu+EL5iTG1a4OzhQ0rWUV4/4iaCrPBqq7ndJgubwF4THLhK
CP7+4jHJh9V/zqGU57LiHG1pgjCT5CtDB8npnQD0jhcaAyLfkNDWuWwvw0pCUo/poKhlK4GDTeUd
kR4sQKV40/BH704AMygNNUtpZbLlMo4HcOjfyQttnxGdyJjNRycdRG0d7Xb3tPyaAPWFhmlfIm+y
DP5sAPnPW4RPqzPuhCvRzDVqsZvU/0oIxJd6K5o08rSVUZ/2Zpy2nOjFlbnDUX1FHWOG9Kc9/5bp
pqx1FjWFs9Tq/YBTb5T9rbzPK7niM7I88dVk4La7IWRJ+wW6KStAFqbNh+SNyXPOltPSJjlC8Z1l
i+o70NDm53rFX32d5v8ykU5fq9ufwjSQcP++Ku1bABw0xZSz8wp8sJh13bWj4cGt1lPFPmehXq09
0fJp3o4SZiYFkrqW+mhYPPvQ0+NIZdmm021OUa3hmEEkLYWAbB1ec1xXS0hpAQqR931vW5MVusqT
7twmWbNjs0I3m385ha9v+U4H3h+BApKz6acSrF9u/gLm8B1toMftKpn16Hd8qHwVfXrDiMAIghlZ
mbj6aPDPa689hBpvwXB7bhlYxbBHv466tseT69+8Oecy6KddaHOMIUnhGXyFW0GGgSicyqvMlJJD
th9/23OKey4I/lkVKhewijRp5ZPBJ8v7KDlv8CksIIhwsaBbhviqczf/E2vUtfqYstbE00+x2cTQ
MTB8TKJB483jfENnVKBE3umWUsHHHILRNAuCIuK3cs+xBtEiCFnPJd9eVwnDuLWgXGeRoG8ACnr7
dqKa15zCBLW1+0nSa3rfMIthuPpcMVEViv3qZZ7yDiDC3dxNnS5/NA7YucS9l/CcCEy7tkOZKrq5
0x8Alg3BiSf9bArfw/B4wWs7tOD1C1Zh49Ehy4jCH9hlkxrAdWe7aYM3SPrJe+fA8BRutESi6uDy
krs1J5UoOePwCyyv5Yx02N0pupB8J7eT3xYk3aLVL4Wx+5tJgZRFKr0pxm+jHfeiEDUSGINZo5Bf
vEwWX7/xubyZ2PtdIeY2AW5+ahJWBrUdPFuRG5TJ+2vJOdnsx95MqBIlO/VO9yeTSS3hVFseDE/X
MeUbBZhzz/b0Rpaw8M/YjiJQCdOI+rEmdGTgx9jJ55mJxXcCuSP6Paie/y6dOpsiu2i41KPgoGPO
4XY20wDg91NPGSdIIeUUUjeq20xsSpMhtiL7QI3LddkPd0KmYsSiYAiIpg0XzqDSJ9ooZzWun0JA
1N8EHMowxxv+xKowL8gmcTpS3N4hoBTiJc/ZlbGcJxNeFYpA7A2G0v9igOQ9wcJ9Fp6fgU9nrWRu
upE4Uy/m+Kgw6L//LKf1R7FeDIT6wYaW/xLVVgzmuqhKx4Eaz0WQEEJoBd6EB1h1V9w0HbFMZzxQ
nr+ge3xhLmj4/nqx9n1sWc8/m1G1fscXmGdrji5K3YUGZNmJqVVvlcJ9uNY0H/BVt5eYsnitiI5N
W3ZR7DjcfIbkygvGE+8dsuHbN6GAg3TlLUBOo9LLzuRu13B8czGq9z+mR4hia/ucLuis6Tj3vhBT
ZENH4I5xSMRRrGqRxOSGnHseyVtzoI7hj8rBjNVePjbSFy/1l+8gR1krGpgBZpMIhqKeZ1Cqe5Oy
LhV+hNEt3Xus/Ig1DPK1pJVF5+OLw/haSPK2jWAr5/34neu4vRafnMNgvr960oBQkyGbN0kxJNUt
27o1CYcraaDRVqngZk71TQERQT4SF3Oa4Bpk1KjbX1eSV1HLgH58rSQ5DRVWmZkV4DJhjvtrjU4W
+rCQaEFaY2q6uyXQlMJBOIaD3zPM1icwA8BufdlIRxAuJ2wR7Ywv4g57aLBZwcJetHMaesc/UKRC
e+rLWiyQ5I9C8djx9nI2N9MYksPprXbpr82v74YkE0R6zpFz6D0gQ/U7ch58bY6IE/gXdUDbrM8G
tHh1/Fo5Gas8O1JWzYjFoS9iuIsxLuJS/ewxoofKqfAHPvfXM58IeqLMBXxOxfRqGYuXOVwngK8S
GF6eNr0ALbNqrbtp9u7aS6CyTK4OUrUfWiZ6ebNyBYQKD7+A8RptHvyCuLiymR3tVU1/JPwzy7FG
8DkFPmu/hYY9GZZfR47aHph1eSGo2qdlwfCCJQYf+q+68uCRMxDIa1Oq3N7rLEDyTKYJZSnIOaPv
ie+90+LDc20M+8Jv0N3n8nTdP5K3V0ZiY0YJaYUQgfJDHhZ5MFQV1KUnL/UKCXxeBzTGeVmCQ1ar
gGLHmZiodZvFYiW1jimppJP2JL+mox3sR7Vkziv1/Cs5dxdy5pDdrITncZM+TtxBZgBrbQT5Tuf0
dY3+7ina9zEjF6eX2Tn+7DlhdfDzBx9icYsJjLpb1UuwsCKuQqcO3XzzBmTdXRk7P34pxUsOyJzO
E2SavRZGlxjErDZ3jSbXzRDmykM0FgFzRTDx8AT+kCk8ODPPXn6RpyzcuRgMLnP4SsQptPDJcJss
wZu+R98CFu4q9S92C1I0THnbuo9pyTWw8BdK3Ui4YFlC5RU6ZMKIItcag8Kw3r21IhezlruTJCYY
IjCcyKlWzNuMCZ1UG6dJOQNvhRtPL8BIQGYk1dP/iJUpsBOn/Zd2GfjJKowI6RQoCCIvH/tjgTJL
VgAZvn5OXM1oThs4TLJD7K7TbHt4WxYu2Wo4XzMGoUz6gUJTXZiW3IkEWLgy9XzHWruyqmGrV3d2
Zhyeq36+ZwyF4Ze+if6MRHt+5+GVjRM1JWtwfrFAM9hT/XNxtWipL6rsq4b2JvXMRgxckdlBHDHF
j+HnTkIRO/EURprtxEvKl3bJC3uWShoI2UvSdk7azRAecTcueS1t2Gm0MDr6Xp8RiClz0hNdfJJp
H0ghaV+UI5l5YGj6X5H55Ta26oMJiqSo7BQLC3QIk5I32aQSYDbxh+gXou/vos6IIy5qH9cjlBMj
MdJssWwNdMdDed+jFbB+Cj5bALniBb9roOAb5rhFDzQFNlx1qZL2gKZQ+rnlpdCBMOKX/skc5fmH
oWVsUpyceIoHGx4EizAnGkbV0elANbfHzTJVoJ+x9qur90mwSgp3iGNmSCOz/0uNKyDKaN6IAEoq
wUQJpgZcknE3V79vUq4CsFt0RI43VJe30m8dggLYW4NOWANbChZfnRHocBBtDnGufuwSvsP9Sjem
jGUbCxk0YZW0hcSYedm2LQvLrtRyJiWKE/+/dvB3Wob38oayb9B66ZdTY45Mp8TLWli7KZFrEJ1a
DAoSrqtLRgsyhXgIQeWueBYS5eiiegw1gzC5ybQPi+eAZ40U3T6a0Ky3QDISlP02MnePnRmMsPLk
k57/XtTHnROrGNhpFypWvFTuPGsF568DZI/O2pc2duvIMhBb19+5PIlzerqtSKKblpmF+HnHznE4
6WnUaazA/8uH0aOu9PLDORE3UaA1cnZ0pzMUGB4N10n7YysO8sDtChAHoYg9DCUbabfxNHNF0RO9
Uhhcof3R+M7WqmL5TOLuLVjRQgoT/xfgW/l8sX8HsVeP4kbB1RV4z2LMLG41XqxajFIqOC7cJGaV
aLIh4gXaJpEo8TRAvv+y2pJiV9YiBQtwRXZKnUqhSKgI11uV5UM3jTRKZj8NC6a7C4tZZ7dTZHQH
z/GT0MTWyYT8sEBCQB0ix0Yi1crNBtiXyFvDuWUWhjo0ISzyh+jYzR09PMNucvPUqKxc3w8uHsoi
0op/JevnYWtI6BlMWNijOKMOVrkWZMKmyhDjZGY1YPFkumbHrXmYwiInCBxJurf4LY+S+VVedFZO
U0i3f5MLTHjDazWcbclibaK4YiZ+f7WyLy5sT2X0K9yqCMk7xJvN8CVvF3w14EBz6i/KH79WYz3f
fbUnsQc0m/0MXAqhphK9NHDm7Vtzgbp/Al19p7XY7s3ZjCTQ0fzeNaSeyAq+ophHHG4b4NY9kYZz
IxiEuQroEE+otsiIZ0xWi0JwicoSw69ZWiQjLrNrRKPJVl9T1MQLsy2B9aGrSNifgrl7yynQClv0
+FRPjIxwCTXGlRZMQo2dUN5o02ZA6l2j4g0UY0wIkYoumifwxZuM7hw2cV1Ncgg4htmzI5EXxjBj
No5Rr3//V58na3RSwbfX6DeoSLfj8rfuwgiEWyVbmw1hcHZsZc1/wYs+9uAePza2w/gnNRI42IUA
StVeYqno5k5+yt0TIgmkPcY+sdX66vqwk6r+2up0l3RWUHY+Px/noPzwXE7vjuZmHRhGo+A39y8g
0t14FuOMi82C/idSqimijglrwV+/GjUhCeGfmDetCxPIpKIKRLdE+jxlLrira0WDQI/SlL/e6e9w
9TnTch31Str+pvVjXUP2mCFqL6NdfILt7+vCSQih8p0sKmcofsV3P1B5j2+ouuC2Oo74re+kNZD1
Pu7VO7toTWhIjau6/zkRkIr6GqUy8FuOQzYaq0uy0+o6mobPSptMlIBm1mDafwcTIIsI1xix9VsC
zXrTLbhZqjERPSYayz5/Gp9w0siFjbHGHqEoxgPmFovznMKgQvGKWSTGfCJZv44KcmXBOxIcDy44
5uuUNDg+O/N2vO1k8cB/e9L/tFodfXWgNY4GVb28bO+p4PdtO72BkPcboM5YObEq1FdbRG7DNQLf
xqqm4vQexu/1ze1lEMw5uR5Nu4HVhoJ0b1Swe3pkFTYFxlO5bQ4lhoLxu+TZW7J9av9lzIbne2ZI
rbPq59NOcb9qqSEcCFSAeb+uUxoT5cb65yqMZSbbSPYUq3WcmSz3DKokkej5DaNtUP/8BGZJ8b1t
GoubGCYnQtCRt9ejNEz3HytLx/duS6cuO/A2DtvC/2qrjSZ9hwKsbV5dLImRXyqTNPm1ngixN1o8
WH1E30FxyhqdDjWWm8X1itJBqoo9zZSYTLBsn1JlnZ1StNx34OGxMKPpseW9yKEEzAJFBVig8Jqr
6Sveh/ozqQWGH+jcnNTmpA9M3ZSPfU3oqBA5k63eNsQxMq5zQ4n7ARZyMEydPLMLfjK/HGUifZxL
i0hqqutPa0N4reet1A5FVM0tLjo51rpfH3yWoqzfM0F9n9eEeBUnLrpbl+aLD1JIx4LyEJW4KiNG
WHgZf9OutRFiG6mT8DFSxX0NnNbGPDH0bgaGZNmcelTTcYtsRtpRnxFWWLPE+s2lg9aY/SYu3uQi
c36Kg3GpRIS6huk3CMKUvH9/vgTQqfUM3uQ2k+nSnRMuewGs1iU4OdGez1Sj/E70bhatS9z71M1F
w60ek602DrTL/BbCXy4gxnoj8pnzMu0rhhemUxDigvje50qYdB7F5UAJzTlKQ+Q8v34/PR4mMB+z
oUaTIpQgydV58n5JRvS7VZZRp1J46AM0eXRKrMvxEJsOfLY46Zc3BMoB/rEczoq33hMDQZ5CMAWV
YrmsEFcsKvJrr1PMGCW0C5Hp0F+rSpJsiRJYyDIFprkE5XbuYK8SW551pkDaI7gzEu6aGQs2uvEg
FKU4/18YtofjIRqkQ/T6h4XbHdpQ5VOxUNT646E1QNE/ocxU91wJHurhCGPpS8M1HjiCu00PumZR
YNfZ9IRZlXTV5RLwpTyQCtqJGLTA5lton+MOH628RqADX936jXFfkCMkqd/WitQXXEkxHgxgcbB9
sHq/0RyOQ9ma1KavSkMHgqBHj3YcQGke06LL+JVUr0nJOHBWTv7dDvjuUe5X253KC4sTJ7Y9Yjkv
OA2ZxZLUmItxFsY7uvB9ItZ88bOKMkOjCoKPn0u2VN75helQgPeMvIryXV5iUZdGRUoYHjbmN+Xy
xCsw6GTSI+q3syvfhWrZtZXeSkHecs777kQXel16xD/74lRNAGa6l3lkOhtVb7ujAp6C77y1uNxj
VWP+b1yKbY/OKGm5q2IEmr0fadzQlL+Ig1hBGZqe5gD7sTnX3JoB0D/XzDudt9VmmNMzLPeVWSWD
0ErvZvAnw1ADgMAHKwD+S/D/ofn/hwr3Wk/0maAXgYGxPPoZwNZ7z7V9Z0+kIRNE9Zo8APwCmsYy
Yd7l7DqTibWIcdclIgH8RfDlUdjrJ1nn7bndeamXIFBdNG4AqfobCoYGzeFDkqn9Ro0+pNyxbZ0z
9fzqdMLeAFgsM0cFPyQ5D7szVZuz4HNt5Bgphp/+7Jak9wgnVVeOFnT/iBnuV0vYZ932nlT8kwkI
UyEvq7kIO+OsuOujMmK3ofSNTc2ZbSRWXiAqOucYDcj4JQUz/zNa0MjXUXpicuADmfQPJkIsZxvD
yztICNicEb/rrnbpJEiOVijjOIrDUt6aavGXcZ0Du211Bhdz4lloAU6sZeLD4WEr4UyaqGj8LyN2
7cYJy7FqhzPAVxkn/w0ZkHkKMTMli8yZQtcTcLAxHl028oD3Bf2VMnd6Fb3iTquaOdWFffMbrL4e
FKjfJkmzljnQxYx92XH5swD4vxNXbay5iuG8gbQT8226LtC6N//HTDXyZQITHATl3hbWkcvtYD/V
CLuJNSRIEp5bhv0+bGbx2uLhwfmhwW0PUkryrmTGXkPxYYRPozfHtou7xzzhZ3b+Up2mI6UEZHsZ
JDhM0PwFCEGB0DCLWHh6dXVJxcXTFh1tfoseRNiEn7M/Did4b9uhR4qWB5VLJX0dhRinP11B507P
QyW7Ra/bRp04KW7P3L9APNCCltFLRhOED0kCfbblaYum8fMVxuO6rN9rvwZNgK9Tl9cTj1BspVMi
EmOl6caBj7pheVeZPLdeDHZUfdUEWcZrt5xTEI5J34j6ZEm7gSqMOWBOKAAKlVZS5On7+BqM0Krc
B5uXZOu6c5aRIGIPxdPzZZMAlBCrp3eT6I18rSr/uXvKjlAbvwUa5vIc1YIsROWO3HBOlT4reTRt
HYjD53NJQln46dvKj06kaq1CoOfGOud+0bu9W4HxUV1MM/dTZo1b4pUM56RggfdMgZd5lkHG3wJS
r3LDkQSljX+BnCoCyGRJa3EwZgbIWSnwnPEjBACdFYu9aOzkmkItIF39Ggeqlpjf9OeVWhTXuWTM
/WnzeLuGWFijrv56hZM9CBAsFffjPUdzUD+nHFo+UMeqTkYySenIIMbSXi6xVfoeEpFan9EFYRtA
NI5eTKsRrAZrF4WMqIBC3Dxw4/RK1MmM8x4mBqrXu7JdaPzvt98qKYBHgPIEebFifjkrsId+/Dgb
rtDo8HOGUU9DwgS/nHVC25ID1mvB+TPSinJcxMn7wXeUlwLDFbGHgxcuhXLxMyGjor8vNTv9qy5N
v5ccXWJQeFaVz6sLzNSl38HH++v2QXsvAF/GEwUrGn0kQdmYKGNQqeORD3ShE02yPUvq7PQPke0M
sZa4yghciWf6nhhcltHncoOZjU6L4I2hU8nhhMkrMbYyRZc/PMgnu7yxj26ZjqZhzDKt9U+Ut9y8
pee1m2+Frwj271J5ZePglVJiH9fqmF3gX/L6Ia6sPRyx09Dl8+Vup8W4FOjuv4DYDzQKlwCVju9f
8c+elYqTR9jD/Cw5JV3oOJkP4NErhhlwIwzM+DEXE1ri72DgzT8K5fchd5ItrZs+WQpTqthItwaz
dx6ttcVCTvNOnZPCbzaY+VSjd9x29urxxdx0+OOl06Lt/APPKrLMbLJ/RhSpARaq0ElVDhp0H42V
/mdV6DbijnlBMwVybP2BqILJuwoAYau5ilFZe0uQuhtNb0S/j7gv6IR8X7YS8eBs1ZysoBlmU3yo
kZsAIHp+ngCQZ3jGySwZX8VPFtW5v36ad2+A23Bwqe5hLvnJrwBqtlY+BxwUhp+QMKm4u8+4jUVo
dH5mPCmsRraXVzuZ4vUT/lU/17/Q1dKEHU0W4ASkT6ARHcj8L9TotFHWBNjjuSk8lcrlvUPjchqi
4dfcBnHjuuNgFpQsf12Bc4HbALHoyyiKIZSGRuw6TR/SqSJKhdoECF+F8tND8/w9HJ0J4NSVLvvv
Or/IwxgenIcNbWnpeYxqeB5fuFBiGLk7jGIdORXayepi568tHC9OBxd2Kh4J/iqEsyex+EYyGNop
xSiB0ad/Kw94LUlVbwJMwZAmyd+rvMD4GWN/fz8GdenQyXcyIxxRrrMoLwEqNQmxsICJLpYhAo7+
ZOu1Q0HmcD74ScC6qsKvuXacFgzYRJjz04Mc/H/DNQOdDPZFOVwQLz3DyOPWNb9K5NCZJVQJ+uGA
P89Hu21HRkLXGzIbdY0AZsslcqf+J0rxGLnuhGtIaRR/44m+BnQwXl0rCMnUvp8sFQweJavzH+yu
nI8l/3OJvpWWT/nd0RsZ7ViiIKsr4PLubL6OCvnAKS/ZwuCRi2bbvH/69Nrg7XcTkJxERUWJTxbG
/YjzN262TTkhUNkPW7ka72q/G2zX8x2M94zmzxFKaBJ6HviVlHkEE3h2QEh9zoXhnDOKrRhKCqG2
msOwQ4RjSLSk06YtsXHBdbpEwUMJg4vGpGiJu352eGlwFP62lSJudvZjhtUdNJYGk5HksTRjRytG
nTu+/R5m8swxAU0ZEW2Jod8ddYrfIJDCqO9SBMSz5FXj+RUn/SW1A3g6LJi1AsSIWLuYjMJeF2yx
hjwlr7N/z8qPGJLayJlUaINvijihj8cwVkwRtQSuENsY40EgrA/R8r421VikfnDuoyLh1XgivR1q
KgOYUbTwRTHsEHxskDK1uEqiFbcABbBcIp7q+bLqUidE6ejuXhqFpDa7jSK6vuG4rBUy9AXVvBKb
Ou0YMjNJWA/ExIeQPR34XSnNoeF2T1yNYsRXwVAhOqi3o39YxcIndqbdJe4E1B38j2eQf7UhZ1XR
r8qMxOSNebrivdXOWgpqOldAOanN6e1S2oWnrCA54XYGH4FqfwJGvCZ6yJF4nVPPNsunuJpZ+Wff
ELL6gkJ2bAHAEE+zO5C0Gghl87G05LOw9pXNkZpNCxLQ2z7bOTBmhl6lTh1O35MtTtorWoIDPRAM
+d+4BXRAfRG3zHY6/NYIwWLwGMGXED7kLvTrwZWdi3OHaY0yDVnPvedq/zQzNIirVRUqM5VaWuu6
6ZS0/P4j2r1azM/mjUJwQamDfzBYX0Wlc6oe4PlrZWMsMMltPC9eRgyHwxOLEWE0R74H+tzXbNys
GluthfM+mGSUimqbPAO72NRsUbv6fTMmCG9P5jz+Xm4mfcriiJp1oqvaUmhtyUrl30lXBYilunbX
Hc4fQ6s0V2SMnJ8CdWdjhD918HFjLtKHAyUiI8xLbEXWQaAdxLjrwrhNy4C+/9eNGG/gEcCUQc5H
HbRSXooXR9cTBGsoKMfyMgsj+oL5sqU/Gob9CjTfXgLABFtaSRcHMt10769GtRQ190v5ibmKECP3
d1Ltw2iuSoRGEdOyqsFZqAPcINQJnMNQ65T6NhXSjNWGws7GS0i740d6XbpznKNo5ixTsLB3MBmr
IVhAJz7JJw4g09pjmU4wqHcJ13CJj3Gjy7W5ZvjiXmlVrAw4yLfkfrxGa0HGtkqxIoI7qxbDEZD/
9OZLDWxwfsI+Iyp7RoXc+7HVjHtMzfcGO66uu+ydEIKlRUTY79CpC6Eint+h7x3GynOqr6UQBmty
iyLM8IeqceEyu730tQo9qYsAwfxwgGaW2m8PQ3R1+k0C80Cl1VHP15g2yk1mM38KFxgT1HaS6zKS
yV2C5I7+J2yeqQ7oWcm4W30qQH4lFB1DnTrFL4LkvY723+rKj50bnwieYgFHyEo1K2pPxf2NN4zR
KsuHASp/9QvqjufSmboCwWFMLehgmyB/ucLzzdgPNzlsd558w+AZgUkEqeKkCqeVAZEaAuaG7wpb
8o6Lh2tdsj/wmv4iZAZmFanRorTVSI1aJA1OzJ1ExLMhLChgAR+mVzODe9vLsj4D8kr/LhKiI6zy
DCdaokXdUpYjYT0IJQztVyanAHuwTmJZk43lqoQBqoq46EP6LPFV7KOgJ0IAL5D5UC6UaArLO4E7
gvynE5BVhiwSfS8ihC9/DUKtMdA2GYH26M9k0Jv/EjVWsGuN32mtFCUMskanV62katdLVomtIzfO
JXmi5ro70Iy4pwDbx4uxiL1oz0Eoy3F/xeNERSMmwzRS6ubimQJDhqbMVi7Edpj9UjwwhVNMkgvm
ypmGY4xc/xzitHdzh6wRtW24fvBrZr+4hNh4aAaBilUq+2V8ur1phTxSpejoZ84vW4fbwlKv+BLL
/tn/iImZKoLoDu7SJDmONzbrB6kcQopDptcuxD8V1FtJa6dJoUTeE8AKJOLSGA7jn6kJV2Vx27Xt
n8scPk8G4kz804XO8kH7jrgBhaJEjP2m1+TmUMXnR8puxD8+SdCbGzgAGdg/IFUxElj7uLZ42+5j
vF5SuJTdjGnf6mGKLqN3bIO1or1i/NR9TbjEu61wip1eD2xhFTKv6h4bnFU/7y0IAC+W36zdvwQZ
CfqT0h4/LsLnTkja6QY9Jqzh1kVuFkrMzwqIxXwx60cKLha5d4/sja5XbbS0vglP7gVmy097EQMg
SAPcSqxxxebrJKUhJxKDxzP4197jfL4RozpqkxkVwN6dmM5h5Ts2GOJNYkbI3E42qPv0r6kPWzKN
8dLntPEGPatmA/x/jDOceLylGYfGM4aRLbiKQ1vWHjvwgjERxr6O/dqcb0GuziEjrtiYmMS4ORn7
usI9lva3Buu4SR5G8j3KSwnQ0zOkgwA7Ju/slPSH5WggcOlMxqRo1YThDJaVPBbcrd61DsZRTWiW
ijAdO6ggyO4ZU9D7owNvQZWoDx89i/OF1zBuHt+vQ7FAe/XiPX1PSNzk6JvQ5tNGyyPxJJ1534Kf
VqhHzryu1Cc5ZBkZiZgUwfi53ZdsSJ3qqGvOMVUJIQTK4GnZqiHo/enlr5iJ8kBwDuFLHs0KZ5Uc
0zs2qMEQl295Em6bGEnScR+01ndPJrQyqnb6jk/fV3WUk2HwH9nliiCc2cnGyBLQl1Gbb6nRNpPU
3Ow238aYq6a2+P+Mf3cVAUNWOXl1oboo0wofEvcoQ3PD/pvPq7Vl1Uiw8SENxfij1OBOrfbJH8bF
EyyD/OunmJYrZs7k+y2V3+09YUIZF3qq1u0Fda/rlXcftHhzA36qzx+Joy2uQ1BRYmUzGNFvVJyp
dc8DX2qVFyrxklLasq7h6vWs8GT5wvceMuEplotMk6Lx2S/bFA4wLCiaPk9aQ5ahmaHFs0NUtFgF
Q60031Avp0nSjnaVRyeWsf7r2DlM+ywJt5mPZ8JbUzvXW5UufS2fDk3dnLaMIzEP0r9296SMhtQP
THpxPsImof6tHmx/vN+1ZkD0grVKEXsG+C1qcThp8veTRiMD9lsSDfrmtVNlYA7/ETejgCi4NJcF
LzgSnyDf/LVNxEY1H66SxrndYkSt/FvsFoUq95YmAbbhCuHdeqN/SX1oHYOGIpWnk6RCH9UbK9fi
cjpfjcEviAtczg9/NsjqOB45M5Evwp0954zOtZJq6wN5nvfjf0aMXhj7CIk6DdKpdTbOQHxTmLkt
CndWVnoElVTjKULZR8haHs7//72BgHYgBD+nBbTJgDLhdMC4nNYl2W1LFgQLT2w6LRKY+ycD16Mr
AX+6lEskDlvjlScz/1nZN4CIVglNtgR8CP+QeSoVehRvw/z9EONUKp4+cpfYWCW44YGtDHv4aBrP
O3/Xf4vrHpZ0dPNcU76BEIQSqTCGtAX+8hI+zH2xNBaAxmXAH+LkdcS7UvC3alTCvozj/KMZee6n
Fpq3lbqXuSuLgAnySbRWzIqEwD8mVkwSvgQlHiiz/cJF8NFiH9lA2UUxY8hUKM0dKhJQgUc47vpm
PQuveJbNjK45ghb6A5GxOK+74ZftScX1lMlgS7OCgM2xfoRaz0i8Q16palPuKiVP/pO7FXc7t0ZI
0XqLlxX7JvN6Cn0NV8P8yTZ8TSmRjzl1t4mH1PleUXc6j5VGJ0UMKFcMji4ud5jSf8HoLn5VPLPg
GDIsQPIcO9jqs7jfqeoSj/m83zNoe8UAh1xVW07x60d3hHFlT0DTdntuKn2qpAnxJ7Kn0X+e83Hd
MfQhuA9lBZ0P9+IgniMtl/XuTm9GKSO2k9S2+oHleZhsB8S8r1MYb5QoqJJ5ssHebhKNfouiKRF6
rA8KivHEmWaWl0a4kz4oy42ohdl2UP0gIuVNCgxSknp3htk/M0NsxG2MUMc8QFIkiU2UdjBgirX+
1zi8nWbxrMt9rTAmlpE3HNmoUb6o3QEsADhXbpVLhWrKriRGjbxp/QVZ/DJWdSGqTN2wCAnxGFD6
mIjjwjPLN90TOX07pelHxCRwIuS25Zm4H+1+CZK43tmtE8igkOwzsISGuzzcwmrwId+zstUY/Yp2
GELxIBrpY7BiJTvCip0TTfLgonUGSicSAuJ0j7LglW1vG/RUjAi7v9s6OkGmlBgbearuzEI5PBbw
olZPOA48yxtyutWPxVdXnTwpDU/CJX10npFz8eXGIQ668kU1BKQJgfHE6c07Emv3ABwyGcgqRfNN
P9zUEpdTgC5bYE97r/i9elIs+RK/GMIES5uM3JQ89DQEsuaARBOG019KAtzegpnJbMn/VSbiu7ns
VGSxbnmXfNJcNjK/I7OsQhvaq5lMIlIlohhG2gjkCKydPipy0KbE0DCbOq+UKdmlQwNewuORBd7U
mCseviO34ENR9pC1fNOjucvBTbbx1Xa+piYJrfh16jOurGSR4UJJ9Lz+EbkAz+jxQL38TEnJYIpl
ocZ3KY0X7smVDpqLb1OUg3LhBzLufK6VLE7Y4dQuXpXz29paKjU7DcrUpg71vnvNOKqDa7PoAZx4
Y48y/zf5sV90f75Vl6NxirWaSqYRZzMzn+pr/hyfNAX4pBuLcAKjz27NLcWKRjrPgaCAC9H6NvpT
OjcBqB0xc+A4r2k3IrpYyp1m2T0IxDBnvYbiW0cz4zjKq8ced1MYmn72BSNZU/YMfKNIemcB/lHA
x/Bxhnq3GuA8kkC+nGyMBaR0J+rzCAIwxZROsO633ZXJ64SDpkASGApiEAoaI+HZsGyCBdbGu4qp
SS4HPy9HWBl4a55SGvJTvAqp2u0liPoKtDxMTJwcqZLBd+rtxRk7ItqhpU81o2qqxBJbyOjoSW6r
9JSs8VQoACoHvwLNmwjllOU/WEMgJ59UXiXGR1I3+1EkhCCDnvHbqwsCYa7Pu6wiL1vDsiSg9FIU
tEAm0nt1frqV0Dl4IKxU1yjcb97lR1u2rCeK8dect9I90rqGcmc1DIOT6yAeROYADrGfGCTYtpuf
2DbjUqih9fWRf0R7/uL8uInSnrSS5FVwkwHPAmpiTPqiTCzpNRgPsal4mmR/rYUx28bDlzNIXeTD
w4CC9MsuVQtY3U15jQGiqUo3Zf4Zgu4hcDsMLEp/h4oZTw3CAaYVUfHFKaRxklitJBB0d7u5odCI
k5WbaqVT6HsWyuogQb9/ngarU/9A1aoteU6+MqELleZWUnGq5UQItL9HZbel7Fnyx+fVlDeiD+mF
A80sehnSxxmdMmzsyXL4sSXtHZF5xftKkAFSU7pKzCd8NIjvwSTQJlePusQi0h/qTSfHmUoWOpLr
pOpKWul3m5TM7S93R15ijneGv7zajXpQkvUFa+hFkm3tfyaAcgE7aqCtmf4OETAIcUdMAv5mrVrH
riVLy8+DSqLcGMA3/hpAOG/gmMplyL4av2p+uzd9/iCYfSTr94EDjDgjFgGR+kME15LjraPoRmPK
bGyj8N0cGlBdfnPDxnG/vXkEE8zywD1SdnZ7XkgW8MaXYUjj9q76EOsrAKCASIJf+HCi3wGTPjC/
d9KGhZ12dafElwp9KdhWpTCBh26glKq2WztWYPzkAcUxyc+13C/WA9/2pkHpUaIdChKQYgLmtb5S
XDdcuCCR1WK7dKFivRv0Fnz993f9ml5Zltoi8fmZUS65hbfuSXYXrY7n7kfld3o9htSSHiv3LRgV
YaOqTMHYnCdAQOb6E4kuihPsddj0Xew9OaZhnUN8tO5PsoNiK7BN4l+dsmaQZ1EbZ17DHcX2XCwT
ntJlUsJ4XVqkdhWDBwIVWzSXavNX4GkyPVdspeZQGwnH76hkyDO3BJssLvwUHsyRi8WZL3KisuPi
jsSyjXO4Aw6QHgC/MVHKRlrcTS0RQRh9XHBtJCdxq7YmQas+nZeG/31heHhF2oFldg2G3CRY0Zp+
pzyqWzr96a1qYJu1MW5g1bqoQplsTNKVnQxA+vo2WA+V/SsfSPTiKwYd65xc+PGpjeDaPY9aX1OL
FFvVCwm14JwAxtiwHpzTKJvtzxVObqzPwMQW60Wj5I11YdItt3i7ahu4QJLjL7BpfJ5tpeWV81y8
5iuE3/1/l3OG371t2Wy9p67rdiz/r6Hr1vDEFyWem3TbbAXajrs8LqH9NGq6ilyxmSzRL41GbABi
945SK9EYM8A0wHtvQonItB2JV9gfOwJVtyyBYuDBu4sxfEowK8FLLc14JkAMKXbJef/I81n64h4q
Ef28W0KyP0I1DCskBkS2dSecoEjPxAIvKNR3X9jqtSDLSV9i4qkBJZ1rUP8tfNPbvhUS2jeozDTf
o3KEJndIJSyk25ln9TI/cbpxP/4D1qDb43cWgWu77op9YgIa2rBQdQNqmS35PgpweU762vnW5fP/
GzNYdF8J+G7dX1lQi2G4dlhYNOxHSwl5wcMhVVQxBfdkoi4YpKpte+LQSdGYqB36hj24jVuvreff
+ksbMqt3vXPk/TKr/nDB2g1IWYwhfbDORXWpQD2PI+3SnihcTMk6rLni0qzb8z5hxA+sOaL1zGrY
L2rU3xIs3lJ4wnSgJIGo60TSHxUvxmaHPd1JqAW26/Pf3578lKryU9QBHck+TIa/zyD9JeFSvkon
0B4VcslM03P4zJX4pfkhaNh+cTRTpsYR5XVWRXebHDxsNHTDKcvRF7oFgeP6VivL0cAHqiApvKlu
hX5i3TOwy6CFokR0+OAycMZk1BvNjzYIDQiEc5jXfSKJZsS/TbU5ITzRcTa92XLYrx+JPSbYKa3L
zebmGqPkt8nrVqO/MR0roPsistwrXwB7OfM3CYUPZ8pbu9dW8CbcKlo5qdUlMTtzIHM1lUfTmXOD
E5f/IWAhjM4RZMHfHt71d3wgwyk2oPVjiOz6lJs9ZDJkrPJnRHcRsM/87naW1GdJMO0SwV8v7j5e
Ua7T0DGV6QRPVhjV1HHnBr9h9gXO5Zrg0xQ5QcuWwqtSURmHBk3B8vICIciXtd7ov7jYvXWPqHWe
VJlgIFS50Rf/xNMWJ7cHxh3Xhfp3bxh+vQphH5Vh7doUpnVswjYBbDrbXREcSmiZ8Zpvoi6+JnMq
y7iqMHbFazpkhXSXOYiO9ggRMKtEwdNmJw5XbyQ9GHz47vcwerxwt6fDkSvm49jEXSEAPEcRZ4Yb
ZDMypxAbBYthizxIowEx/EDl2bhvppR4kD3tWM/r14/naOx1DJT9clJAwfoA6PBTlgSeMbiTEjxG
qtOoajE60ck6GCKMrXhZc2XE55o4c87ga8bs9KxLfnssS7KAG6F292tPVLgdeSpSHcKTJzLQGJq7
P+SknT6gvD9g+wzsS+KJpxGgjHfHVyfJpAFJORbHeH0EFIf+b/Mi84PgaKlb1jwCvDIV2dYkdZtj
V1VIB/PJxkblHJkHbl9xuiiYfMmTh5kvL/6S1IJj1rHeWsBxfsijJsPb6LYKRSsTdOGQRYjRzpmI
ha/7IqcFqYtcWIpfFTZioLfRAz3JVpXRt9Vp+x0F8nLqk7QvB++QaWz7gluEOYbBYt3jtvW+ZIrl
jA4EaT9zMwSkYuaPVvNBkPwixVgUyN59lcSC6fsLlKG5sIqIY4hmBQepM1gTN5gtZPqoxPNWicS7
tw7bA35ePLJgpz5hE/F2PzPrOM44n+7ggJ5HsJyYX5q9uq8oJvbWaqW6th610hB0Ga3EY9EgaCV0
Rr4bYh2iXrV2EPduPYciO8Vh7LQ7XFcQi2bQafHj1EqkUPzY+B57YLc9RPj1Xf4EqJMFhtY1WEY7
3Iwdkkz5D8SxLA7ENJuc2sfCNdPz7ID2qNtUQTGsIdl6blsG7FzoFsdxTkCalVDTYMCnZp2rznJP
T3Xb+9FLaGeOmM0LqZTWPIqx8OAiNIZ9UdtlTYooxR1Gl+5RGyibsi8ZLrueurrlSiyGXpCFFXxi
YOLQ2pf3YNAltEscYQZxouwNAnl7T1HZ1boZ8BMWF1/mkPBof+p07EftiGzqKNnnWLA9aRRMzX5n
G+l3HoomaWdOv6FEZML4ky0SvmqLlgHxRYdzTRQAkLhteSVkg3lDHSffRk9Lnv6yw3kQ+sH9jybi
sTrDP5K5E6PO55m+403NPAsqkqfxIJzjV/OLO8XhZkz1uNdAl8fZDxIu2OrhMBcojmtT4U3lZydk
1rRV1uO1n8qEAYfVnDvuYNAuSP/gJpDWL1u0r1aPD1GcFSwnD3oYVsrhav4gVdJ9NnQ9xRLj3QVZ
OxOjnhnxkhYQH3L4yVzAN/BODiGoZZJ/ABhT8ckYZwlgMAHtEIXRM42F/F5fWiTYlAMeEL1EGGO6
Cpr/xMzwY4yEnm0DynE+eq5EbLRIqfvRCOTYrd9v13cJD4tZPaoSndNuHfKbZ6P4D3/Q1k71JGjN
3aGUw2k1XPeL5QOP/um/f3TK8Vj/ynuey2cmKbAmWsQM7hLlLU0ol5McsxEV4lQHSHWv4DbXmN4F
xco5iiKwgKs8tvWnnIVfAdh9XQL6f/IHMNR6Elz3qUrrodsp8e2Wfz4lHEiAIlT5Q3qC8JEKwZ9r
LpQKLDqXEUP8oUDrq9mnwNi0d0YNYm8QdXMuw7y76WjQRt2CVGo/rCfvnRwRb2075icy299FX9Tk
bQ2rSn4jFXygEtySVxQipwv3gGQUA/zHayVBH09Y0JQIT+QVX3s4iq1UgSqnER5kBtiFMrzsm1ne
TPsotn+smBKkecAZvqOfdyKbI5CVHds7zI7aDwrTYDldtrvcc+VfEQeIrgvfU66Gel6+kIpWghaU
MFb6zPRmZ+EwkSQhp5Iee5r2Wr9OyRelO7iVqlLQNk9DRCBvTJwA3UYq1XaFNNxyn7hsOA6+MJ/V
8CYbcGJBKpBf0ne2+5O1bel5+uvOchOQLP/Wus76XpxF5PQLgw10dx4intNeQeGhUV8VcI/FKl+v
ft37X+cldtOX5m2ekUKtN+V62kXC3ctAMlpU9LAjw0Sivpb/nPOjWO76IfHLRW+jy1Dby682Rnau
TpIUJCgZArVc9lBu/haR/Z/oGavPAL2s/57zYJlKkKO4LXG98qnq+LHOec6dI1+mNMoegXJLQxFb
axZcrLFJ8dBE27vQ3PwO5hWs44tiLwRsfgyYfes6P7BD/VA8roC3rNm4t1fSr5LIRK1bQ5tJNEXF
QXTsWq0AlOJ6xEZ32aEV7B1xqrfIrHGZAfdtRMHjvgQGeGuGX93I0neow8Q5TaHtLuFT869k56lS
HG5BBa2W8HHU800NijxpCY+xtGFxt7MJODih/gysJuYeNh9gFwvQBY3jkHaD7D6vckqmUhg+tEyS
G7BkELpEiarD5O8oCwepLb1lwbafSutVc+GgFHh8CZmrDh05n0WMYYfJl8sbyX/uBTq5sh7DLiTM
JofcLN6uq3lc2KKiI3GOEAlE5Ry4Lk9Y2c4lycYrBq4RqJq5Eg3h1z10eS+DE21oahnMUqB2lANc
m9dK++qCXLFUQy2cR3IKeqXtYQQ123F1hArU3zrGrGBIMlH1I4quguVXFjdjqlIVBmyJczb39XoQ
8seA+fw3qVbh4S3/eFBb9CbU2txOKwrDGvuyXCj/FMVgVxSkT7+30R7d3lCFIKidcztKyQJVsXCF
KoYpOAddKatqlslrBo4u0reZ0mJvaz+yjiA4ezThqmkkNgH10Pt5+m9Qk0kASEQ4DeZouD7UC+QQ
ee+Nhy/tSb/mc48yFdDWOCheg8lpuKtRW1GL5OBrqhd+PVkDc1pLv0rVT9OcxRyGm/Oqx7qCyu8I
jV5kQnk3Fc2zz6gVBr0b9AcYrybYWaLJGoWbWxQXNoWHCb0qjlnP6JlAG/ou6MwucX11hqMC+8aP
sPwkpOqgWLtVk0Ul8dxfjjhawsAZvoQi2klUHhiSm56eCmwnlNY7KE1dKdVrcjfCfPKGLnYeBElC
zsi2IhoHApGxALA+3l3K+a5XZjgK+EBpFmBSnglbnrPSW72eBsR7srOZ15nXYZj55QSJRuZ+wGq0
cDDA68pJc3JhwzORah1b+UyA7SAudMCyHtQI2JFW+/uo6Yk90MqC2M8PMGQn8HQ7U9FtQvXlhlet
JZTSVRS076jPIjfyWuTiPZON6t7FlETtdGBHsiq0fI9wGY9JiBbjNK80zwPcQ1ZhBIRAb6sVUe26
XRcAia232wHaTOV+KyBFcx7HHqQC0trGshapqh/xOAWSKaiWcmdIPerfg7wOpCyeOo5CSD/35waT
iMfwecIxLz6fLyrOQzy2fvH+fXvba9SVoPSphn7POafK1BlnBXBOJAqM9/V8ExubAnpG1lfVhOX+
CO9CXboirLtbJ4Q9pfvCg89L95sH9e5gh+4Cct5t2buoo3G/7C8twU+6zFjMIDamy+2NlivFZpIF
mI5ePsXoDH5z+JuFM8V/VCEeL+/Qhm/LWpqB5DDxTRYXDtuLUFEWApNCwCl33dzt6xL8gTfFgp9P
qBoUWKhtbGslWr8QT5R5TRZ2e2oSOa37oTSgxkhnBTRyjVtnQx5cMDj3W7EOWb3Qcw0he9ihlQ4g
ubkRZ/KJbxv11yNdlQLOo1E5GZJZlAFCoFi6tp6HolUwNuDpd3MBGEsv5Gh+p9Ytdw6yvsWcDVTK
lqgUJ6WSkYYfnzP7ide4kpsIa38JneZXscYs/799A2QD2Umma34Ov/t1FGs5jmE8hwo89az0T0Nc
pp1LUFCRL+8Sh08vtMWzCSNokcyaLdpoSw1TJsM6Re1EKaH5/JmcHmdjoNCx3TDqL0iI0Po1cuFn
eByDFL8zS3XZ+WlEP6xBRWNPGcv0ykqeHCJ4acg+bHdtfrAonAuSSQKurWjLQ50dMzLupUKEd6pF
eLYPGd/2fVgn/+C6G5vrP8ju1X/aVe5U6Qb2GS14gOBY0Bh6ltBFrvGWpkFqaJPT5ntBvzNlpHFq
Rb1RG6cimtaWjNkjApSoeyeNx2/YRb8D+GowIKuJX19UCg7tUYhSZXXzxy0O9eAHhFdpSYOf1/Pr
v5kB3KxAyj0g43HpdNu6JPo/THfo679Zw1tr/YLZgQu6TP59yTieAaeKWCJYRWo+tBsQbBC6V9yG
eoWYm0/rFnQkir0rbGYwBK6hsARnjPwuDo+vSexhdc0UY1ewuI8UC4YyvNb54iwiIUgGUfmUekpu
jTsplqXz3ndVmOh//34Wft6nTot20K4ApdqKHoyYGtwMvuwhMXyuCLeDD6X1Ie7yubrRHIoYVL5F
I/Cb6zuOFhcs6dHtpn8et4Fn2EBAYsxHh0gmOIMd2DVQ5qp0cxVcwOZYkWOz5m7FCrmqBO/aS7SB
NTlgB0TPsP++i/Do11yj8+kzVCfaoZdZr+I5jgwU4OfH1uyRr72reU43lKd+Isy65lG9HXXfL3SD
IrmyW/D514FzOI/GMpM0HqogapWwrWl1r515EdPOGk4oXvrD9C5X+UPk6qaEMEZpaOlIDqt1e63k
PdIxizuhn0f04UKR7oGY/O0gaj+qjgNA1CIfOoSCNL1Hcnh0JJ84vbkh/nFGhChEWfRAeYYV/aXj
4urzhjfGoA4EJ6LBYBjtZpdY1HcV0tDcRRyp4GubWuugi1FcVeruqg1qo/A7TSPSWRwTm5/I5FZu
PlWyMrl0h06h7YFHtoQvuiYRAxM+eLD+oOn+HMP/N2/sC67FK69bxY3tkoEX3Pv15+wbSh993LmU
5/WX1vYScqJ8ceje22pCB83zfKNjZoivds/CuItNh8W8m21Gm6FY27QvDTClVGEiFm7rHP5fLpSs
xtOYMJlWbuczqxlUxpb+ZpoJsGK4IZjM1l2EG/x14i2tJIEEu+jzoiDQs7gBJVF03Lav/Q3lb4/N
bvCS0PDODz04i6NcOvNs7QyqYUVeQdrgtu6Fj2lWaibZgPYXRcjtM2v7MraNsrrtkEwhDVGOEorf
QJqpB/7B+hbMROpNcIPfsBND5BeNbCdnVzxV+Ym9llhSvY+aLzZjuotG4MKlklgFCLpa1xpe94xx
HZt5AF8xsdbpZpSI8YiAonvZdszVD+9twZfb+Ty7Emd2iqvlVjxMvo0wGg/OVqpKdp5zD8H7TMvd
PDDDF73VQEfnj0gJU1SOHpLVZ5kKL6JdT+pLvwhl6hd2pd//wEESLLjexRGhZZxGxsj5xlMkB1cO
GGQqsnWXAGBnBTaKp7T7uFNTJnLW7zHHSFRXVA0hkwkXstL5pDRXhR7ZBvd5fkXNTXCdBCSyfZoQ
QuN6sUE/E9+P/p2xR7yilF09ez4sPt9MmnXG9FUZ0hSE0h7Cp87/C9p5MxGoSqCB2XlX0lgly3mD
aXpYoNTg7gh+pMoUwnXKrJLp34UTVqzw1qJgsxst5LcuUh1L3IyrM6VDG/QkaByNoMxxpWZUMLom
a4zlVbilYWfhAuSLlVDKPyq6kBK5VvMDsE76KnNZkKm1ALOJi4D/kRYExSvNboJr8Cbnm/ssnbgq
f5XmUFSY0ts/dUtluKBR+KvdHZR+dJQP7EYOusYutoJUqQhclWbCsvd8JrcFr3vjYTIMoCQgq52v
FcziMmph0FwQ585/EYC9Cjmb9S1x5RVCyWcnsx8WguTNlsudDv8ahKWcwv2x8yASHYM8iwjGDT+I
YSI2EMTJD/Km8iJLvj9TdV/kzMMqhCaPlzgQGdqvKhvHZv7xHWB7yxjkP5UaJFquF2zHz26m2N6U
b0hry5kSurkkKLtfVgv1GJm4s3E1uoGXUrM3rOBxuvtupxerwpiyoWzyQTM8FTW0mbRNPw5YWkTq
kmFCNKRhNNU0oU2lTQU3MHcFkLYfo10xmAlEcJjlN9VPKDmn99IftgCOnGaaCwTqKB6a/iinCcG2
93o20Wlcf3QrVywgqJZRJHnh0DM2V7zyFK7lXRQEwZXo4xGFMYzXSjvBIZGIz8zAR/ope28O7bi3
ZQ9RC26eWcUqhrzo6ktmwBNaF7hPorLCL/BnZSpyOl5UMw4P07jnfH1Qg1vF82+pSIQOydX+PFqA
/7+MGt2pNbgq2ABr+8iKfgzvbRD+2qknpXoD+CJiy/wMVVDGhc2zIPSXWOT3rjSJv0GcXZA0rKYU
Uv1YngGp9XYOlgNcTHMimamCzUZLX1KkTV/LI1m7Q9+fuM2f6P53Sd5/xz2pIrcW/5VxLTf+EZ6X
C50NHg+l8ED+4oleRqU7agouNqJxo5j7NPheTAiHB6w0kV5MG4ysrH4TdyV+y5iEGGzu9cyCQ9Es
gU0RQEK8hiFMSws/RQBTL/O4vZ1KbQV9YWQGgKQIjnpTHL/Khlbyklb90Baq81mCWDP/Xe00g1Pk
CagEzdEM5i/w5QVYgA9wxqdB4D2z675i7hukPEKm32k8j44fPBY0uLxwV1mMC08wJ0sni8rnlAEp
Dsb5/EhM0SiEuc5MyRZEhxs+XgFXI4PSRy6KdtRoq3Fnt2Yz1fO3YnzJrWPyCYE59WI6qC3GSrrB
nJmryRHyxo6NFMmHRIIT1Ks0a9N5PLlnAE4rZmwxn/K9gW5pKEzRDTfSNnQXC+jzrpyR2/52xFtG
cBdQRvtWNZL5SlbAYDEqyFLSni6TBgOeIUkXKIQHhIwcIXUZWwmdVVFsZIZmNpGKGeGwNn1a9M1P
cycv6MZHdx9LGPjaMHrs3jXJ2I7GbzklDXCPd7yszco6/6PLFoCj6wGGDWtu+n0dvSjFCXXoUJrx
GAV+qYsNGwyW0RbHjzyy3g4esr1DEjoQAKurUGJ2YWZH7xeeZUj/SX5YHpGDwJsB0NwugZYrkWCb
iQqZV0FNt73tFHw9/nGPoF+OZXE4qdzMAPHU78N65b2X2DYUZk7liga7PI9qZGPX5DjprF1TSRSR
oNlV7/nlOb7jGUY54srzaaHri13xSvrIm8kZhBR1T4wTsie97t6Pejn7zSQ9qVPC6ypXtHhEHMkd
2Jc6Fx5Bp40hVtarelDQSPcDbK7d+66Ly8UF5V87li3z7Y9oVCjEaueM6xhh8e/W/YkSx6cMZa2l
hDs5361i9NGtXUZEz0ryczkvojpHD/GMjqXpJGZVM7LWsN7N1h3jOtR7FzwVlKmYsYXGmDMQx775
DmFKV0Bsb0oO+lniz4SHB/hzu0awGGmreDp2Fj3k8Y4MBE+LKHgXbVawvWdjL14KkHlGxr87jKyN
UrRzrGiRGFjpRR9VwnNhoOYVfeyxlFcG17ZFKszrzbXKVt6iIM2jZ4fjDAYWmPO885mUxB2CMLFx
iwUlYA90thjb1vw3+Qph3g0TjIZs8zzdVMqPqHppKDzfkXnQzfc2k+86kJDJmaDvZQIBGOluCKnK
1l4xqIYcIYpyz9U2qHMZhFJuK69FeBCH1ddaVkPd+Si7J+jwJp5A1lCzHgDWf9V7/HxSP8YFoR5x
k8X5TTy6SWXdS7dkr0i7KT+oX4Z7/IIOTaa+DpsGjhyYEz/XEp56UCMzHRFbhjyr2lQ3ScJpIH9l
AwtyrBj09UohiTpoXXsEPmxlUdEsS2CnEV6C22FptKL6fhgfeLYpCFuGK7Wq79Bl+B0b14/vDciV
6aosYX//Xum1C6Wg7qxpky/nPF4LObIKUZQYFx0Vr8zFCZp73eA0p/gARH8OjgD3p3x5fBmbXVEj
KunXWPN//Or+l0Zg+1g/qkIkVsG39m6A7L9kxn+AFgDisyxobE0+C+GvBPmhoQb1UdFf+Oj2/8a1
nsdJRxw0UmSxcQPA9qq+OM3zJiPcW1lduZXyuEqR0UhXu8c3J/9e0EFW/ikJkyuLJZsg2IjaQwoV
ByjHhio4qt5iwdrmIXmPFD6OArIDCrefeRax7OBZZ6kPDuweHqwijKlupGa7Fnnn9ypLu3R21V+s
n9O4ux6IMyjIBuBEhlnsfXf69/ZHeVZx4IOh/eXunVFaxPTMHNx+ZtIokt4bJcR3POsvpXsWU4Hs
Yk9k38Mb3bn+NRFG7dzyV7Bs6ABYqH7Q44B8CvEaZ9G6WyRZssV/g82rUti5MgB+Jz5NfksBjFdi
8IyD6+VzXv2PlmZdXUiGWDU58pZjVT+j+OMNtjL862L3PSWvakNwka7Md4WVzZcCweX8Od8ebWEu
obNxqhEjZGbYKV6QfiJWWnK3EBIhyUg8KWifwpVhz9iwPf/JWB5g6u8rZvFE//sD+LjVL9qwcwyd
iulI+EY7h5J0qgFWoW5a0jdO7eXnL9R/t12vIpzrUkHQlzLN1k5Iy+RMhaa2zeC9Iogz8HRsTONm
FOI0Pyq5IvSNVzYXeewd6GaipQFshwJUzjqTcv5HW04lnCfgYRCbPStf1HNfQvzuGRueWRaS9uB9
/HBqvfgkTkxNMqSufM5OSkQC4SJMWiG4tsE/lZI1ptfgnxvqQ6t2qbaALglojM9H7bU/h31sjyWu
ZlhqDtsEEW5oDhz+T+KoMQq5MHuZqxFCZgDC3n3qcHT/n3F6QNvVPT5A9CfLoZx5k/Yyvv+QykMu
FaUz58HajZwu/hzPs36bebADabNdxraiBZvPTwYKizcDobkvsQyxk0BuTZgXr5i6zUjfp6zL3tUj
xpQn1ui2L71AopzMGwZc8EZmQsBO5BYGau9DE/Yn2AMYoZd0IwX9KH5ZfvqeMlXpyjqT/8/ypa6J
91WkCC596ivmRNpINVJk3AFu8Rv/2B/m2mozq9R3Gzi2tiae2Fdy8c0lhXzc0/isEO1Q+23ISIm1
pYQ/ZxqmnugCMmp48DZIV3ZYKXLsTNNEmEWJbY4bQfbGpCPZYtO1pDjfQ81aGTeKj4ogszDQJO63
9dDa0DEu3TE0o47iGyUPkTWlH+KxfP9aag+hdAfxbslPF/VugB9yj+EfttnYNi9+KNTr3vo5P4Rd
PAoVfSxJiK1raRNYhwT4Q7ojLChmrNRbxUGcTvQgEUBhNbaYEhW1tdef8UV1qW0pAALELx+gRbH2
XrXHNIsOtXPvhZ+BjJOUnxUEzFL2YtpPmQ5CLs1wkymhW6DBzJYfWELW0I/94GXaHU95+HzFNOQN
B0SiniNZCZeG0aRPPj0FyKAUn3GSbJGiH7tCRTv+9GY6sF2mhd6cj0Gq/tydc5s9NsHO4Z8+H1Y9
R6GfgpqC9kyUxBgrkS9KuqZmQuZaZig0+jspViXTVrWfudCWsFmxnBP2jr6KqrXzhtRe0nGNdG+9
ZUD02Lbe+n2f6aYrZWCrSh6Flr10HpLPvjoWA4kIS6TAh759pTqUGA8CxLfCfvdrcD5qok9RkIpm
nm7HBhDyXGFTYFONsqvZbsjhljfytH92oSJgTCu0pz4hYU2k3vpmqbZNU1CzfJGgOM5IfAMEDTDy
U5/SRUSYxQ9oiexW5r/Z+tCY6vfuYQvKfPg82NhTQPAtXspGz7jcSud2RcUzEJOL4Pp99TCvLWLx
GujOdzPP9awAPS+raBICjweLUPU3DOtv7Qu+B0yfAZXtADrvI93N7eERM6JZzB2jhwiYDfF7iiCX
82a9BOiA6A5qJA8J29Qrh25zt00di1PDOZ0iv8lrpVeAzPkInaOzKrjYw+gp1i72qRARS68QnITQ
bAbrB1ZJ4/ZgNwyqRd+LDuwp9ujeBWbM+G72HigLJlduF3QN3U4e+34VgNsZXiwuWghvnABZwBwn
0URknfVBt70iu9lPPeLNSc2sc7rg7dyYvFeMnZjZIVAfsxHG8Xbqm3gXXYePajT0VJDB+mBmBMho
/d5WINvYHoJglkXWmeg7Z4ysxb447zq661aZUbh5CnfgXoYhnK6+cXwz5vqj/JBvG1fXS47UDd9s
5rSk4umFvHhsJ2APDTfDo3WE0bl8ewE5WWguoqSWpmGI47EbaIapuPVPA3rhsUmnMebWjapTVNt1
5oLIuXHHLVEzKjw7o4KAtcAPfOXmW0nMy+0JQfoAAIehuJd24oKNM7P4pzBzrM5gGBydkXn9rZ7d
KSjqzn26m0gYLsMue8IwUNuPisDRzoA+ADlJ+Gu4pUXXfEyVX39VLZvZbL+TQ/N8dItn/4Umph5Y
HrTJNkVKO9zaxq4R5jLttVdjwTSbOTiRS3NTTvJ0kSCVUrayaMqF1kkma3ZncpvweasSlgZ5QD8i
mLBJqWfuJTDOQhzbvg94AHO0mxyzWom1EFcMLCTBWcIsARiOG1vMaLHoqcu/I6CtxqaeapYcVskm
PWDzbP0ntCK5oxmo4DXLDSR4rXGt+oTlwAj6e4aPELOuBuEyV3i3i5SbwTZnp45OiU9maYJJPQ47
0Rtp6UCJ2/r56dR99i2q+d16f7NPQ60ZD7qy/UqrH/fr7lodNbaacyBaujjeaSI4v5Krf5cNWZB7
xiGu1xyuRIBLcfqiWIdVPjBaF6O71HSLZ0Qrr4dmBoow2hEQPF0I5Mnk6R/BRSAHuesjGoE90ocT
tuWM4rXHptSKJLowHkKEWUdkjQ/q1ywW09OeJUD7QmtiadGrCjJXRj2Y12gWmDvwVCN969jIMzoA
dQP24UOhp9ORRlZfuxFSts5ai/VslQA79eY9rDM8jQdf2BOebFmw7b0IJ4bhGBKW4s5pGS13ZmOg
iGVTDdjH5nTUFtWLM2n8Bg4bXkRU5puOWDPHqfYrvyfRAxer+3KtLPewssbCRI+/Mb1xkiVtlTmh
WCG7y2re1QylSWpunjsYsMZwwyv38AUCWhk3DQQ5vhnzwrJBy4RAMflPwRkGsnx6rivIGWALscaB
ti6HNhPTLmiDv7wqhEqDNyOs1ufWxssnk08P7S68w3Eats6c2QrJOBFqhZCkWysolX9PdZJA6BE+
XnoIq8+nwTSRUF8YxKXRKKTQop6OxE2pFO6e+wb2q/PZJfrbqIJvKbOp+sk1vVd1qQk6oNEF0bJp
fvppnNSR3j9qSF0r1SAjn6iDTUnp74eQ3dWcqkJTKbGPtqsXsNms8qsvaKOlgUcO7wpXx7itxm2y
vScwf3eCvB361hT0GNf/ltA+SgFgjyRYSLd/Wm15kpWb4hBlAYG/6lz6Rlhnzjj1acEkIVyBGa4Q
MDK0mMFErSwytm0YL+e+K/RJC5eQGD9aCgjseMEUTAssCSOiiC38v1gezOxkdEu5OKPeKsRFtzFy
cH6TY0IueVkgqORpcojephK4eXBOcNUf5oiBHcxcI9RZrRHfkfm2TCUfVuuGH/syh9djjSxDOGWN
hdSZO3DaOpr6rkZa2O1y5A0xoGTUOnWs4QaTSaeSuItQep/pRcI11NlFuMyd41HRwKhP07Y1ULsW
MkLPNsfcCs350vjRx8R+oBwHFrVkMGCEQsQJ2fArRaXdN+ObJ/y3aRiSI8eJVqFsuHn2/eM24q0R
yG9PFUBNJA9hiuv42drZDutx9PRMR6dbTq0MvAuCEo8flTBmVW/um1q3rlpqUYyppztXPXa4vMWL
13Vpy4RLEOFjP6pO6RGe7n+R7dAjC1OOrpul7jDSox3dx12n2Chk+YaZSNglfUnRb53irwlODLbs
RqlgZKIHaE3bRnAVkUqP7CtZxOBJ101K5VRpPfaMJppVHp+ZF0Gq7nGnnubGJ999VegZsfDEN5ho
801xn1g1zj3TzmyUIwruJ3ABD3Q554o3ZMJ6qWhVNlqU/k4GoeQvqihMMPljWLXK7YkANx9IGEcs
BzSXJTtZ0Kj1cTmuqEGv4mh/y9nlUgVjmG35jU2JvFLcrR7YtBqh0t6UQnPfs3YQF9EE1u3fEOrm
WojRF7+M1H6Z1dKmMMFO14GuNos2MvDILh6Mw/t6TFx4L5bmrC42OCP//rjWbuhEKDl0DyXnWtFl
IQh5C05vWr9Q6y8USHdawMN+R51ylS4Tw/n2CeRWjNh0UnOhi7xe0Wgt8GfBrQFsgCNkf2VG51E6
JjRbNtMNCZAoDnFqV41ayUGYlJGUH87ti6Zm5McrhrQffvwM1X6eo1HLZeuFJbAf1gMxldSIC2h1
EIKY2gFdAJ5pOTOxF3Ls6ajJclcKP+Ke/pMAOR060BfhyttQqNiWmf6vP3wemB2ufLScec7pEx2/
KWyYLXFvebCTTv3erVZxILcC5xFFTNjjWAvR5KRRl/7LBjOpX15xBGNsMr9jWufo7qo3sk81NiJJ
iwYEEVYAOAJdgfaZPrB6jLyvEm4qL5MOBIXoMf3lpVCaJGFiO8BXBOe/YaVB9Yuf4ZTwVQPJZ3K+
Zoob/nEGGJ/SBEJAxE4YjEMi8t/SUhLp9mpgmzkV+wDIjSRmV3jCa3fSEh1zsJ88Skym04mT2ULG
DHb8dHl6A/Orxu+BcVeB4AW5YppVoMH8Bb+rCr2fB3jsuWCnAzAjAybAjlrzZm43FqJsSKfkjA3I
hqJIb7pfCpuiOdLNv0vgUBPdf2Ro9YaP5szEF1VoiL1Ciqgqft45LxxjYUG/Mkjg935N65DLkVdi
IRG9Wulgt6IUf3M48synkJQc+aZowY4uDnY9jeeewGOymNS/pbl6q+DSOjSiH5Nd7w3HMyAIwL/b
ENd6W0U2b+zKX42NFJ+czzlAZNk/umSqCcHfPqdmrZQ8kOf/N24zSvI+aYViexhwKNy8esY19826
2SgRt/aib4QkWshTcM3rwn11G2Cp1FB1KKG09wRUkNSfj8c/ech+XLrutzV/tPrRJwTjbmz1OVgP
z1TU4S3w6dfH7kMi+CCgVtQrAqbBF/DyBWrPwcWz+zO+X58qPsJ9f0Def6P6whYp9ZARTQAmEaQ5
N/IJ3mjWGltEVX36gNlLVbpBz4OjMaEy9GIcdHQWd78jbwkis1VR08tY3Qa9d3JxcAOeCJjkhGxR
OVAu0xGVINZ/sSTHBHXjdXZp9NcLVAzrXpqojD1ULT+3TPplUlDC9EhHhWoDcLtEpOKLe57XPi6a
F6Cy3+qXxIkN/j8wO2Z/C17IYfsben4vYCrfOULoj5GH8ps2FEzA+/Iq/cwTjhnLjU103rBIVoGK
s5lNao8oL3e3FFtUoqy6tFlO1HnWdvqpt1BilOW8hB5a7tHn5GmZyY+EPpEPm8UBEbaaHRBCdDyE
GnTZdQhTTKo3Uu7BKui6V+EvTtomdC7M4DU8bvmPVeVlGvJs+6HuXnyi74lfgOGZcZZcRk0fLY9R
tfRaAQRQ86d+6skIce7KhaZDKtl3O2FlS9nSKyXtvxJE49li4RfMegArOaA8om6nifOKeG+OXJGu
qKiqR8mycan41qsDsYM+nKaG8jBC2Z8PYBT8zaiqw6QXsuSI/7RoCSO7IPyakq+/qePDbwSV7k1A
Ff6Qfr0zklDVn52VdPEqiPfzY+UIbstpXA1MlJNuisSJ1aJRalgEiHgUbR5iQiWMCu/xQ50ihXji
qi12nkqyvbAl/xE0GTKO55y8jWPlxmXf5MAA69Vv9FbjVxZOyF7D/tWm77qw1duR/p4prFC55Kk+
4RRvhBgnEJoySDAi1cVIz7qKciDz78/iFp12IpKTSAGNx83vrVlyq6W2qGCp4vewWdA041lg4JH1
6uh53iKFEXqXKCQIp7AZgoJGaCqJYLu3LPnMpCBTvy6gJePDamk4Tywtuxb0bK9C7Xpchdv4xvS1
ZWK9omDgjwSlWiLN5ogAIKQQ+hxXhdnkzFKllxqxOgqIX2eUM+nvxxNvPZnT9Tz4Cze9zAtanifH
XNwd153TVeUehIeIU9NxyRCIAHnlXDmYRRE712NRaZXhhaw6dDW65KVVXn6P4PEE8QpZUcZUzJuE
XVSjLZX/m/FuGaZy6THBz6+HLXp903rgi4HFuO1XRgiXqRC/nYM46fL2FiixzCh96sNSWkFRu8SQ
dVbublV5fbGLwTZ5dBBFPINE8YcooyedLTtNZskN1FvLADnBBMt1ZKf5nnmIB799OeCYQFh/Q49G
8a/Tf4PNZ2Mo5fgLCI+sQVpeJc/uQJPQwbvyTaACXdt1HU+LobLJdr44t7FMBK+wrJN42tqOecB5
vac+ZUmyXHii+M4V4OHUXDHLHnQ2kzuWoXFUR/2l4vFKqQA3WVqGWfcHjN62OFlbp4TnNTNTZL/a
+wYieFayU6KvZ8tvsWGCA8w43ckIk4mlMV+E8foqo7G/Z8joTym1RUvLhyEbOTRUgOJlqqbmInJS
msmXlPkdX0PGq16NdrELkzDo+B3vOOjtWDhBeu4ZT395Ece0TtCf4LuQvYDtTXMJk3imXmYB/tA+
iG1VLnU3+f4bDpyD1W5GjcZ/N2BWMQlxMao5epJ1CnoSWPvh+R8m+3GaRXqR++xhHGP8xIqGa5gq
a/Y5Atx9+WbpXycGIGPV7xRpssKD/s7R5qVFp9N3ZEZnowzUaVrIhMJCnf3qUkygu6vZ2q05BdYN
E8fAXlGg+tM3XpL5yjkCLSP4RGVCdQFATPhZIhTI9eAyMQCGB5tYC4kvuLxTACo3KLxLBMaELQdv
NotuX14zfw6OS1nGjDDvldCCzYVpz1PHidZBGfXdynbCoXNVAUca5la+EobU5nPrd0PRk9MPs1kk
9G5DV0FZMU3L74CqKiJdMLVexYlWo13EE+xCntejbhNNVRTkLdz2FZn/VeS56DT1u90VOJ6OWCK+
3YSHs/0vrWO97JNFjPfqcVpNLrwDj6PAESEorp2NGZxXUOvfoteynRqCp3C1+8gwiByPjk7SPwl7
/hWeWvkdKtiERyUzgNGoAOohxBSOibAP/BgGNVWvvS9/Wco+wA5R+oZjNTIpHCZxiROc0vTELxt6
W5CXqYXmRzkSRQFmbMcpHAQ6tP4539buR1fmFLJG14BB4kes5JDzxZNvLxPmS7ktb10XNVgo61uf
0sWFxTIWSM/s8H3/5Md5uqylAed9ZZWhBKlobbBzcPazWOj0D/Y+qseCq3P3qC/i04RmbMqrLofA
+cfTdgEgt+aP1E93OqGztlIPPAYRiQZZo+JmHAL/jCBLgN6TiZvSWDEH9e8dnE3AX99F8WdunQj1
/4Wa+5izsLGsRBV1N/s93H63K6OLeJ8NNqt+rHnTmLm6UANyY45+A3UQAb87XFpbwqnVALD+BQAD
dB0jpJeo7uP3vvB1ieT1AqR5rjVxYsoKzJ00k2h7auk1LVFnmdqQIKa6ljnwRu2JZiVNspXXmjF/
TuSR49RScNBzg7M++QitDUyJxVNpnZhgiRaaXBR8Mtf2z98zal2GAPsaiTJryfB/Yho+6irQsgVU
YoJf/q70Q3h89XDmAQTNj/5BpWpxJY+HmK36DqB9pvULZ0zOVBNgduzn4gx3nvdhVCvXtWum/w8G
zEJ6oSTHU43wjMv/Fr6LUIXRIsPSnA9yZv62Kf8LcZntMvZ3E77STlUAuRHSca2q1qIezyhuVPKd
A5zcifOxlmH5f6sKqjvVqOn2Q4R7o2M8o5mp8T6m4dTo0YlG6DGYdZdQd096H30O5nzusxCFVjC8
lAY6v5RcTxkcrXYoro5migOSGIYMNfCVg7qMEJebvLH+AS1upG8R8uVO/cg9MJWdF04HnLFGh4Tm
2UAwPf0JIgO9zvOg9h8j3CxxJ0DNPuyedOxFZdEoeguMup+/IjnLBU5aCwOKBinGSnJc1ARe3htU
XSTWpuYPxS60la3BC/sEdcw6wkgFE58yjs2is2WcGEAD6CLBVLM+Fvw12lm695Vk++OZxnj6BdWR
t20YpYkn0f5k3wa81ZED1EMZiXvHz1f9P7SuN64IHiO8ZPNpwnxyAHJDnPQdDrORytwG0E1nhm0F
XdySwAUUTDhu0efTDvv0rISTBiuKVK5dEEvswbKnDR2bMk80tJpHGRhDM7SXzUcZ/1+X6gehbGzr
BVf3aKhwjyI4J4wCWS9FkDWS96QIS8lRVseGieH8fZSjW4KcO1yMeqVuwzA4pCXx+TGcjM3hGCwl
dnlCKhdPolpi9848PfcI+aq2O/Rw0w4fTpxPHfQ05Nh5Jn70bWPswABXtwcc+I4ulOAPR3J0iBdF
wkuqmSywP9K+zoVi/7WtpJMVatMQZzh6xHaGusyNMyoLLZZe3fc0UZsggx9e2ZLv0DxJkkpyg5/U
TF1dW8dtKS4CwPKr01jOG4Yg/ajqfWm4/ZUgvQYevhhXmJmH60jhZJYf+cVowN96QEo/RTi3LvQ1
f/e+/ObCVq67/9GFRt6N9eKDWypEIcFmIGEWoAO5BDNsZk+FCheli94XEDHnoBt9j5lNJzmtF/MK
m6febPXLXq2yAk9YGPQ5tsD2gizbCQvK8LsJfBD8OqJD4kzE6v83EBMzJu4CwMnE3cz71c5dVGHl
WuqHwzBhjJHt2BAz/HKnRVEfFjIrP/Mby8m/Gqsdis9pYjquqdhln+B903ii6e6V7G19cIVY3PIX
4WicXqH4krv6DZf/Bbn5Z37BFhf6zUjWb4Fi2d9mo7bWYpgbjWtl51CU7Iu1ioYjcYfHLJcsVo3m
UY+9JVUnDmz+GHPxQhgntMH5EfJQKCCfbFocvqUzGN8JEaEwZL5Jd/c777OkBCl/5BZ4ZwE+lvCS
y2wmNtD4jqEaY52s+vR+iio+3n2Eein7o0RsxdRkgeqzRBYhs/jmNLjLD4jPIhEA6NP2LtDaYA69
cVGldhWDZzu9IeFmh2J60u692Uc6dr5mui9urSsalgBHGuNIrgzx5TtzQelAPqOa9Dg6DWhxyvnD
IbBccjBZZIq1t+Jv3cYd8KcFNHJnEoRSxJmqJiz3wxf6C7v2+ydbDMdZlGXQxTsAN5oX+LSwX1NY
KDm9vq7aL1CISPGECKokl3dNQz5N/09uaEZFaDxWmFCUuJBXH6vwkCwyGWv9Msc64tmbdd6ju8L9
lWvgUxpkb04MgzM20wmZQ/5Ws53yFo/tS8rXLRIQUC8rgB+uXXb3XXsPiTM+62Ke5THBWvuNMvjC
+MnE+cl+sbgd6j9SFFhgshQCNTNN4ffu9k2aPSY7nJVeV7vkXIuFiZopRF1dJWYOFkLXP3h1eCeg
tqNyAsAkkWozXMmYIzenkcPD8RjLDEcVniGCt/TDvRqZvMdMDl4Tw0A6kaR7qedDOHAGFR6muJ1W
cJs0apQzpQ1TAaHAHYPmu9UAhB+k2Np/Ec7aJ7l6X2/5I9sDcYFf7ESK0pjGATfzE29WONbRJqG4
iYKpPJZD9eiZaN8keks4O7GJ5G/j/S8Vmn8CGy8yKu1zxO2d8GxNrpFf3LQaCGX9CJPdVeDOA4Na
Ur6RQmxDH7ysndqve6QJglU/cah2Y7r0T8I/7wYNac3oHWPJDBlxninFVlQb5AR+EWYPRZ/81fw2
qhqJMbPtYQx73A3T2we3pQCHFLMkxvhCithIqh0F7eqHrewABZA2cPGQkQ2PzNsAjMrVNA4q3LeE
POz5b6Zu3BVHr9L0UvyjZV/1zUOXTNineGZM7NV5QKU45C4LYXAWPaHq15k7iWI45k6aqaWcDg06
LJ/dv2N4bui0t1XGw9emLnJcgGyH/qBRW0Pk/YMQPN75IhwWPDQx3gauwgx0Q/g9VFcjT8SHO0kI
KDAopjDOIanyi6KF++2lYCMpq5lX9oVMarVqsbqvWsNd/tWNDwdplEbCGXdH1XBb1teW5iahhFmh
v2swxQklEdQ79+hSkHukGDfmuGvQKh1edfQL7YWcrh8YJeEUSad77p/DpVBnH/TyxX1kknin37vH
3bNhrlUluj/6DpluW++crmYW5JYEp3DvciAGjhGS7mA4BPjhLR9NwN9OSDGvqHqTRGH6QCjFt3rX
y1Zum5kOQ1+7QMRyMjs00iCfhyG3WHb7DQ0WpSsm5rP4yI0tbIkaKhtSKvaIxFrkHkz3YIWoauZo
6tf6Lr5DyxjnqDW6/LnycRYo8Ebos3Fk5Uf/Kx2EokOQsNiNuUyqTxeE6Z0x9ScQ4PPVxDPlr7LJ
SrbfnssglDYPktUPK2sovNLBcdrGoWG31mc4FzOWUtyVG9A9jqYt96dhUSIKgudc1KGi5zMpYct2
5+6YoxKIFG8yZYeHfvutHW2kk1uFkMWuOlhZH0HnQ6hTjE3feBJFJo0nW3mSf14lmZMCN5IyTvh1
8kvCCDiU0GDUfB81QMmaR9YRM682zHm09ZBFpfDI6QIEFmw18Dcs523aBQlK9nmxfqFrDxf90J58
LcCzLbac1PFJzOzBJgZfKnqRnSv+xuMNNBtFWyi2h/GeSplZoIinhR4tWsJJqanEvt13b81eAANx
rSwHX6kqbfgwmeGEA3Qd26fnWDrp6hcJ81wCxL1Mb3hFogmzWZ2VkpxQxO7w952wwk3g7TyetEaO
OXDyMjcpt2uzEydwW41B90ScvonvJLeZVE/pJk+dq6j7KQ22E1bIjRWABNxN+kl2SB6MspBPmjwx
u9BSAnlGPeH3Yse7LpaMronPG1PX+z2W9GFjKLOjvvPmOPlA6Wda1LgVr4sxLWb0C5sFA1D9uRgB
8A4a9XiSnILksvI0MsMQ3axtysd6d/RqSKYSekSNhz7d2Vmld9bcoGntcWhelSQdodtlmdPzLdfD
P+WB8/ARcwLgfaX5Wi+6pdwcDpyYy9q0UqhW3m/eIWCktvU4KtpPkjnkyLIg4BUpM+JyvivrXY39
0CGn2xHSIYhW17RJ3VgTNbkMR5ASSHBOEwnKKK2Q48sXkKmpSKv9fv50P4XerKj7s7d4XxYvqvWV
m7eBocKDkHrOZ7XM3SlTwEotJHgAl33rjgBk2Pq3eUbisiTXOsP+gbdDoepW27aQTiCysQMLhrwZ
Fhfq0zluXqG6wvoMQ46TIwys1nTQvlkQvKVYW7zu5BiB0XN8n/CeBTMtSUv4DG2c/d2s7KQHiZv+
20XBGtxTbYhNPbz0roY2ss4aaoxgveVhalmksutBeLzicBombRU7dToMvv70dLE3/6JvZvewSO6/
pE8mx/MxYDLErawTWI70gXYDisHkY9J1j7EoQkxHTa7FvoByDQnvGq+24Kq6vEx8MRTHbDMRep9J
VGIDnGbhij99U1bo1UHOe+vJliE+EJ2lNFhX0dXeebFeXsaFZ3yej1nnW+olDoi5tvC6LZbEWp+u
vpdPkMy2qu5n4YWh4Xk7yRxQUSkzcwsaxfMAU9Aam5IpDUzB9TTGWqCeUFdklU0nYI/3K8K1e25S
Wz9zyRk6cSLW4+0CyC5VUYnY3VFgekIFsACXQWqD1u5BNNArxVWUClULXbUNF/6hhpRYcDgaDwrd
DbLL1XEqi1LzSlbeIrT/quWe3fYwG4Zkfyoh2tkmJe3mTHgTlhr5+x//x6ENNDdky7Kh6QCL7G+J
NGsV6pIshDKIb59FnX1zlUrnOKQKVe5cbjxXEPsOL0IFF4TIkxOr6o+I+DVsnU7hZoTkWlkO+2tY
S+bKadBUrbad9/W7ZsYODZ65W2dkA0kpotxqtoeYKNwjpguvFCnaeboJG5wHzLCiSGDX5DD6syOr
P/q1hOU1fxgEEWWoIRYfDxtO7zvf1CWvcQbGVX1NAjHDt94/tza0SoZdcSWEjnPYubUFPlkgV2HK
pXsdIxpvg7FzS2HaAlVfAxcLWjFTo3Y9i62zWzMSG8RVNHyxxqSq1+tUyqciBuW1r9LzPqPysT5K
a+qjy0RT4Z5NSIm4JW/fNbZnGLKvu1bU6nSO5HB2jf3wW9SX7beutK8NcGhwVg9FvPyOS7PgYhKD
z0tdt4AMCsSt6zkcU+ynqBJSdPR3tFPtlGww3V61TjhXWNWDQI/FFxfMFfwC52X/yHX9gcCZ5VWi
trm/32CabhDqH8MSmpIoEC821/M/a/h1t/kFz5H7nGbVvy9OIia7jNTu3kaDPz1CGxecCcXrBif4
RoE06pUV8QXK81hjQWXxMOGnU5zlesDhbiJpjeI8nIGxCsytNACh8zYvqnw159aU+erre9jAqyHE
E4Va9vf443qRF8Pw+Z6xt4XCBRqMeyZ1nm+/xoY+ELE942U0z4QDfJcIo6ZOloCF8zWwY7SsbETY
t1VygHukikaC/WyaN84PFELsaceQBXsffvX7kCtZhlsEmVnINIBlKyhfhnMCG/hmC0wWFw1dVFE3
SDQBi03L3WXcAJDmQSKHyoQF7byvJdlhDOOA/SBF7UtQMkBK6f+HPeorWZo3qK7wucU94KJNriM3
4nCKh6K4Rh3AMwpBTvCJdDrrswG8AyWo9eOEOBrxpXTEXqCi91zkeRiGA6VdVPDkq3VjVEctROk/
f8qlK3FIKvILj7Zj7t6czebALtTcMTy5d7k8qDmS+LH+9kgSaXZckNlNCj9R7vraCPojIvv/tsg3
6NseZ57cKpqhNIsQppF2Zra4vOCoZufw0fW31y1lnvnUXBS3w3BpULo8Vr2dVVUPYUEaeRzRvfnF
B/FOMZ7dZOb0x4oqYblVYy/jY/8GewXklXmrNpVo92i+it2iwJQsnQKxL+vmrzkLev+qLrTFkuO8
hBepV2s1y2pSlgzT092HrbpNWqVGYUBFjreIIFOqbmuzRyBzbCt2rc41NkL7QhUuUmhjpKWB2Dvz
tkPGVoe7eM5XYR33iFjvPURrVhYgf5mfvBl+citWiOumEOXu+HV1u+VHJUCGQ8mpVRzrt6bR/7Gv
U/zjXW0mki6nml6oo79yjTESRExT8Unju7Vst7o/VrPtzAUJbwL9S1eZBErgIZDbaFw1aBSfY5XA
NeAUKZNeelwpYu8E0GdFkwqbdRYzzJOXb41nJh8XT06SxcUim3IANAtODAtsWaJUt8pTiWlEfTi+
EUV08TtXh2zirVvMVDrWwSYzEf8Sdh+R9YlTeb8BbCfPBCtixQ4InJDUh95tbOtBMoOqbU2ipMLj
ge8EPWXyMpdnV64lV9GXa4couxLnt2Si2JEms/mQvjon53HRQsQNaBxMlUbL+yNS1N8rFwvDwIRZ
8zR13QCIpX5kS0Y5b2ivuNBGgKjn2ViuJ0zdtmWs4B7TIgybuBd+2IF6Mp3KYzOSwCJxhJTE52IL
FT7mJc+ykXeLtjtKHNd9aZf5bZ7fcMmrYOqryUxddYswP8Sk6UN3cIi0VyTBolrSUsGxeXDe8yuz
aCHvI23DkB0o++vnBPlUj/quMpzj8xqKIkKIinPsVfCwr1wQlfcl4AeGKQgawD6iC2jwFAiZvxvW
fjqPrkryIeG533EAJGfJSmBO/j/7Gqe/RwQs2M/0MaianUgmmM6oZjnklYAwoJ3yo48Ev1CwyR5h
n98d1plz7HL4F+N9dZEFMnGMdGeXBT/QftnfQcmEj6FPM2oVXRCtCBox8b++aZyT9meYo5Gucy/V
KIor6TzTXPoq+XNuEsTdFr2uQWzxZNqx6J5+viN3TX4MRjEmnkk/PWHdTp7LnGJiEUoPtnviInsx
33+AieCWFmpNV7p3VYpSV8Oqu1dUW/IWENAyE2MpXyn0D8WbdDex6jgwYCnwvQ8nS87GRvsYPf7u
QIuimig6AkS8xX87vOBQgsiC/CwLQVfGJ665bj27682Hjx69uoseXqak6PsNUgw8oXs2jq1/TkzM
2YMbfSz/xOVnhkgKaR3kQuBIMx9Udz9ZEqzpOQI2VHJz2287gIhmORktIB46ruZ2HUbOCNmpxXJG
9yYZQob3eEc6bsg4GNCeTb4Wdw63j3DBjPFumM3LEmf6q1mJlcAl77dJFzJbFT9jDY43N4n3Xk68
CjF41qZQmz08MBThPZL0Fg/NObhCdd1PgAgVEqI1DoVUX8kOGOznmtmoWgUj8dsNyvBrwS/qYIB9
R4M+ORHSJiStXAr1hz5h3OyxjV/uyVCIsbovQJuVfSjMykI3IZxLpU/Z482+ImsqBF2Ur2YbqAu/
f4msS93JpQUjxRJGJwNl6V8Y5C+OwM+ittjeULXaDoG2Y1RLPkXz1KHt1WluMSbA3XCaaLYy3a/D
owptr4E/VCAWSmg1VBz3R7BGM0TswGNquPwU3ISZ4F+wjKkPfKpg69CLU/BNGhkZ1+C0mC8oYTJB
0J89NwfJA69/vQU6DqGVZApWKbG18+2d2zz78QuYXBHSLNjOlheiv0rGDx+LuuO+nnsQrOqmqyIV
4Sc94xlaRrcyMUJ7rBXz35KHFbB3ndMDXqg3JbO2Qnb2N5McmlIgD97Tf9uMl0LdD0osCmmgvROz
ZNCE23iQMvW2cJgLPKXIhGuqlM3TAN2OpqsVfNHCCGkDRVhdoZYCaHR9sbOxXPa9pmxZE8uHF2Gi
QsucrzhjF4GxPj9e0neLjNRjVHdzX+lttUamDF/7wmy3S4OpTJruo9mPUmMlmsNDgRqMveq0UMU9
K+hi00IrL6XCs8IE0+n1ZyZ915mdf0HDnO9RUY/FeejZ47dhH4oRp2hLy7Wdw7paYAJDrTJZOeQa
x0M1opraUs71rxZYGTytVL2GowTIi9stW+hbPY4P1wfAkNngBm5Iia0FsMN+TT9FqPyg/gQ+M3nw
B5KXlgfnCFd44mLpsHbCnt9Sl5wF0tfy2VRRSqiLBUIWX5c3OVUNkoDtgyMYdSqaTjRezqy2jrV9
b7A6xQM9PYHXPnzopqLEpM+k+hw7moSuNlYweoEiZz/v13bmxfs5NBRpFp38TPl97ew1sJ+ZoCNd
rgy5mxxNdNlM9GXjERLwoEVxaXY9SNKmnVAs2iYE9CJHDCYZ3+P/P5PpsXeJlF7JoGGF61gh3fYd
KJ8A7q0egIWxg9b0AI7ZKY9bUhF7Hjdr+GMhRI094zYwEZrmC7BS2kADSYQXf4lpTUt59mNZ2CFO
jdWulMKSqnL2n/IMihxBJVpDMeLmUC4Nb5RoyBmNOwEjA2sBi1NDGmVjyP6lZ3Oj40IkEpDdXR+M
fhsPF2ZwagHpnxn8YX2THV+u8Y3QMNbA2qGnh/DDMetFQLDiAy0Wg3Apq4sgks9M303s3W78C+CK
kBxRpsgjZWjl38oQkH9TUu1fpiz1kR8ku6CDeufWP5VJMiC62wVQHUeStxRiylI4bw0c8ycYvGrr
eVU/Q2ztHKZOhC+/ye36eophW4KN6yCc7m0JTyxO2V1GqZv6xUStE6wT/DBR9NhtU87jbNImX89K
N9QMzAxFGhZOeR7hu93lMGqsQ+99XlmaztkxsgnoVIGHrxD8RZ9y3wT/XQWoJlazpbH5HpFY1+8v
x79D3EeBjYrNmdMTJ6YH/h1ccHcUktFcjxb0jcOO+eCxuLj/j6R8pkmwe5HK/BVb4dsh0jZJtseM
4JBRRWMu/oAxxcanCWCUkGvmQBvzSPzWBqwGRlg4gu7Pkw5wXhyh9gMtFefvDLiGUWbQQryeXqPV
m2AWf3nD8A/k/tjx6B54KSgX+NUhPak36YZl7qdlnbwIHyNPEQSLcv6XprKCw+8QytjH2lSsGY35
VjK12EUE3O10S/EY8NId/Ia7VgvsETBtWbzc4ujJAi2aY/Ikyp+FcXjfscOvH9Gnh2s7SL3+YhCW
kKR/Kb432eVOYt41/9zpUlmIbzsLpPD9wnyfmclimSswXj84dZvGB+MjgKSthEjGDq8mSopXQrnf
6+iHChAf3gbQuUCNWDUW5NQpAMAjKA+l3Xm7oDKz4sZ2uLslzdtX7lFlSk/Agfk4NxOVww9SYcs6
OBB84SA8iXIALnC3pK+qF69twGnjYlD++FiSHTteInsNIJ2OZD92irmFDgAUenAKWYlthwbNVAz6
HmcFkPCPUg6LBfA7pON7rg/hmIRm1aOoPFAx9hHKKb5Mw3AKVsdEkLhbKpLOOrXUUzArTr+nuN/f
fT88GG+N5g436gGQMZF9Re38jk3OrMZyk2Z9CqQqfClWN4/hJV2G3fDvIIuORs3PJVfsXLpv3ukh
RJqPoJZ25Ht6ozRKfOjNM1VWSEmsoS0MU/Hn/HCedhsaMtqOLj6hNoyNWD1xIcnoniQiQMBj0Na3
uvZgFFVlSQgJpSlXdgGrn8ToySOHa0+rBLy1z3OTmm2ARo7G+V6v03Av91hx2KI8TOpw+YqrJpBq
EE7y2dkohayF4w+VchUHgGqpzbPvS2blFDZhCmgKf3azpdd8J7rEmhsZ9ugOXcG5A8/Lm5rGlRpL
WkZxC7XFQVZRqvLtzeS7bdsqpjHKzh3LzScOQUInhvORZ4jhAXOWVtQq/4GVkjJuVKOJGf4xt9cn
Cau0N5Fv7U82D8jJpCXwgG0Ka9fOJmrQrEml06pQ7AwI0Pp+GMFPq1wvtC4+8gXB4FPnZPHQubR0
Ct8E6HyTtKDWe+6NPNdIDU+GSKh/8l3lwJ83pX20AR0pcR0Cs456ErtWTtmUv7nRXqyZ6iwO41ks
+YfDWmO33qLU19dv8P+zogpZ8dPP/woMqUb7bQMyhCkJnbaZk8yVTJavHkNSlcJ8I+56QuPstkas
bpuDVEpuj8Fv23XLExjnFvRxqENT0+r2zbjoplLDNEf8SaH4DHE8ifd7NO+rIPGPeJvLLI8OAmbF
723heqMLMT+GT3OqwYTLaG53M72h1oB97uPFb3jhF7Ji/uShn2J+k7itFbsxPKnZL+0wQ3ROVeku
T++CeRf5j+pujcM/jIOOZq/hhQ9ue3I7AdHVXoQBiKK7VJvryz/XdZ1hI4V+lhFz/6nF8Vg3RSP5
v74dU32aNsnnW//vK1a5nU4bo8WPFwJrm+gNXuVoj79mP8CGtPBLJb68Vnjw/gLex1JkjSckls+d
vqHNCc/3u75wJysYINXmVnz+GBcSScxqr/SFNtQEyAvhJy8BUPdwd8Smwat5BWYpF3p4CL5dVksT
XOjWCEXu80EyS0rPX55RGIfCancd/eZ5ujgZjlFox+AixccphOIiyqW1oCWqTxAfqyAVyJCJunWY
sAAYylbD29i4BBJ2i4SZ0+avgaialWD/y244jBYZLAL2D0kjKp5QAqtzBtnCR4RxlpNXeDlXsWYv
WXteZe1RLraiFJJsN9QkanEBOp8EgfhvaU8MPP0x8qmbpL5okh1e5/OdKQmBB7kn6/uPHYYSlAH6
CzbTs08psj8Hjg3kxROY5qB9Fahs2jWWeLZ/W1ezcMVql9NaZwDoOBRbaLdTh0okR9GQdMlfbc0E
97oanCBVD0cP6nRYDNSmazAzssaRIXb3PaTIP/kA6NesuYIosnvMoZi5ZOVF4lF1bilKMkvQay3G
SXzoUpk0u4n45KwoquLvhYmetMyKilK0MhSpI63D95IDoNBpueHdxne99VpwBW3CKbj8qcYo9Blc
640GEOxpHaQMm7Fbrrb/u2cAt2b71ato31fMr7N0ND4o+D736WyFUfd9wo1g3jBX3n7vS2wdAP5E
feWr6vmiWAyR0spApPq8275bMC6W/VvDHVEzdcukV8rSBfkwYUcMV7oiFhQYPviNNl+RCRmSilza
bggD6ef7JkI1FvmiQAllQxRtlLCeHTeW/B4UPgoXykkBMplpykK0AJcYEP+SPuIuEFtsnfKcGEnR
cq+F1FOKvw7HGoAXeG0LMajaHJusxkRdTMw6y/Vd0XcqtYPm4M0Yby7cATUkEG1DGfIOs4yzMG7h
4KlBpG1oCqHtKuZtWIYsCOkDrDcHm18E4MmEt9Z8/1rud5QLFStNX/jSZhrU3b7qk8ySSoErDQMF
7LfKTnMGxf0lRHl0vSK5AojXb3Q3ShczxFNH3N52baWRgBxPn+IMLX4pl2Wxdl0QJ4aTNmjBJNyO
+GImA+zh+E57/b+ArsZ+BSD/FN+QY8ALnHUjQHXsyI8ApXZcpqKNHgMC5pinv/GkY8niR2giT4Q/
UEwnk+qo33XNmEpxjWj/X/PIV7lu8tAyS1XAz4qoBg9uc7nvmdwG0ij+Sg914cyqp0tEWxU/BNQl
nfBgrBKL+HW2iT5Mm8bogvCaZTZGoBu2RKqdNWTvNiNyPntjoqx952cyIb8Gq/h/P+20/frmxTli
Q21FYqWJmzQdtmc8VpkwuxPj0eZxe03tfGSjlYvRMGE7O12xT3JtTG+eBVFBCk8kin1cT+Vl4/f1
8JLzLTdSUuigYg5zL8C8kJ6C4Fsfeap+vfALHvoxp+JGxTLBerOFBzEt/pwJRBPPFUeICrDvrgre
WoP+bQhZQ1IXAS0cEKmtWOin6m3cMG4amGX+9vJrLANN0y7HS3/o3o4nl3QqjVT5l/71V2NzLeZK
mIe3Af4VlUrIIZjfBjY2PreqHWFBQVaWrcLv9xtyOWxN6XYHYBmuS+4o0++Kc3nTlLFJJpEBcdcz
P18VDk186IKg/rXzqW+40AtWC3GCZz+YJ29aj36jZCn6eqn/KBZWb2HojyEsIhaywHPXV1huu4ua
+UBZgDEwtLDZsts4kDpBiSxqk7NnBPNAa97cbRP9ZDIIE7HGIvjUFxf2D2MRM0Ag1wRkBZGiLeg7
srPGlfPvC2yqH2IJvHp9FHtLo5dlyoVaWjzWxGeTDI6TuoaTDj9UlmDztfIxgnhvT7+dRO+9a4I8
9Ke4+PmNtsett4Z9i4g0UgK+iSqUHVSd/PSr4DivgFMdqrSOUIcA0fCPPK1SctfLloY/JD8U7cEa
3vcMSXn4klJ/tJjzuazsD2dRiBKh8w6UGSNlNPcFaNVborvXlsvDXMWkr/6JqdkHG/ScvvX7BOfB
ziWajQ8Kgv4QW77F5nyyNrVgh3OcaSo8EO/DpAo3t1uj6KLS3nLIV1TJxJpeYp/QL5Q9M06LekTc
29zK55VONUMuvR5Xph5gJ/BWIbrA7XlDQadC4I+MGwiFHXkaLRDiNsGvlLnOfuxlLYyM2z6Di1mj
CgaWyLHkKdhv+QMqY3bfqKjLXsFSK35vJJcwbdVcChdhYa7oUj4wpXLAWqSUV+Yv1Cly0Ikq7ql+
wPROsqWEZ0yZ1ZMo44Zamf7ItMib4Ez3kfg+zpTH+jrUauoPSSFawzT2K4+ltsQ+uhF9sE7DjlLE
S0jvy9JokShxpR6DGBvGxFkEN6gpCeT6fVuTcEEmQWtrE6i+lBIkvuhgT9Bu3AQOAP+ba9kmocmP
JZu72MyF6oO+PPPlOrj8M1Z6Qmk6zGZkSn2iJrHp5oNM7wUNvuRx/w9dvnXlNBdbNvDVGe+IJwBB
zsSQjSPNSqhBGh0k3l0dvwXghTotDIoLfaRBWcFdswYqrTUyAut6lHgwkmDEsYoPBej8sXO+xxGY
nR4eCVkEmaxVNRFwmBDdWtVl3ovKmnEDId8F6Ic6FndZfMKz7PjFRCbUmdGCZ4TtYjvB1sB7+DUF
9i30xlbFNTdVmhSjWg7k6X1HjXAjnsNU7pgd7BhOu8lTd47mV38TLkDRTrXK+KIOdKJyK7YupJWp
NG/0zmMEg7CmFEfnHchpbrSaHN6R/MTwB5D7zcVzn7YLF6AciEQ2vv3/F07T0uClivcT3gZjie4S
Pf9GzorqHXGNFpmHDXVDOg7Hm8CER0vMgtBf3SInmWs+w3U2qm4AAprW31GiEp+k786KnPT+eb2d
tG5xmbP2bgpb6U2IZ3gt30ZF7zmcqQOPT1doCF41sFpv5tI4BnfN0SmG2Wwmrsz1Rm2if4V2/zzc
4G2jVkCVjjzX2k/HcsQ7dlxawk+EbiQd6Sc5+utwc833dpLsUSh0lx6kPv3rtYpoLwiv2mYPHJz1
5+bPBebhUeX/Zo3eI61ZwuG0Zcaiq4fGxCZoiRXeQxnYHvmvgLS60rNQ9Ofr1uVcdmm3DQvCAb3f
x0iN8vjS1BQ4DByGfD9dk/jGY6Gxw+/vm90QvnFvvIzn+dJtMKCKOAsM7zLmpzOTwBQsrDeWPvEE
IgMaVCRlT6ssBJq/ed6s7aEQvsUMuBDYPQjJOk4F2Q+ySJYBjqNchzvaeNYaIi31/qJbjiUPlotx
wYkBd0Z7SQiQr2Mv4z06AguRg4Ha/gam4bIZR02tVd2d77v3QVhc66V9ExdrInVY/hIzepKcb2Mn
GcZIr1A6kpJl9NYYgHU7xNn0qYI0IpR5SDjymGsAnT4uZhWjEveA6TlhLAdU5GmYjOQ+i1eE3+e5
qqQpx9GlJE13b9TKwmeHUzq/tbxJF3WgyxGcuuM3QE2seIB71EyqDFrf2yEd+J2iv7W1CTDU7U82
TNSDyTS2Ps7wd/4dS7MdtM594Tqe9qhkSkFyIV0KpMJMxGQXItRK3pXAx1Q228RQGzkaoVGaOS3o
F19+oKb8+83nNQIT0/rNOkeOAKmS9nNi493ob5Em4sNrpqMZ9flCMXnQydOoLNjs1F4yq8xGTF1o
ym/MpECSWVTEK+rmcGKZsx78lDEyhIeepV5K2/r1AonAFzH+yVFdNV1BTJ5hcL+HpIhpbk1W92sH
V7RllTr5KSD9diT8gSdaDQqHp7p1tDeMWwmjrkLZjmLuJDMniWOYKGuPEtpYbbaZb6JfTULtNYju
g7obAuW4fY9mYoT7a3THmTuckIFVGkmhmyVzrVznQNaG+QilhQpkRJFtjyQ+n4ZFvkLxQkCJvnEw
rc7tI9QdfaJ85m0wGQc+qgmaeqzMdsUqNCzqyX7KkjONGn0z5hoe6l7uDNZZW46PcVJE30m4thFH
Q5r4gkaujqfQSrhN/j3vNldL70hPNY+sWhmXEgGfE0rZEffFqpGA8ICLX46R6AjCdIZmjLDRnAOd
fs67s82PAVZ7J5Y5Ze4WsIN4/bRpmn20Ku4aGv84iVX5EGxAT67twyf5I9LzfBfWD3qfc6V65zYg
89q01wseC7kNLilWnjeiyBvxw+X1ZO6kGnjcetLR1k2KXZCFNKuFAh93tp/79pbRbieNbPZ+4f5+
l7+u+nB7xL6t+8X86ZLNovV7xhLmn7/E5BIGub0IOYamLFOkkEIE/yEN35uAm1RmUQMUE3PQtj9v
yU+2Oi57Y7EuNJehDoO3y9gdd66N5ybzcUjsAa43WAtuVgGGqbGF6a4C9X19OqvV8o1NQ0dRx9Dt
ttJKuXDSTEB/O0jk6oJC4xDyHUYt7vkKjypDV+vH7l55cvkp8wCEn03TojfADchdUVeY21LB/oTx
/ZyS96BxFfjZ+6JdUfn2EDxXG23dRtQ3g/cVbeHCdCB0OrFSfgTceGhhSB2bQc/iNaUHRCMS5xlG
ECtlLJei2X/4eZI7YBXBZe18DsdDxi9I+A/of+VZ0Q81qhRmiqAF+3u9foFqVSaC5fJlj1WxiaMP
Vp/flCqBMQxbiO245bu4RkiAgK3R/kNia1gdRBUo5KY9MCO7JTXKs8y57ixbvATAtvvt6sfZv/KJ
i9qVvQT/vkE+bVRw0bKrF2fYuB22kTPi490Fri61n4/f2dCkjHqYGbflSRvf59+gIpKXrlELdgDW
fC5Ysfi5LUqaJBlNEYBqOqlBVqyVUj2WRNMMlIS6b/ndZBOBL8mgeaV9yH7QeNGwp0HAxROuaRBm
DmUXjLDXntgASIyAdpQprn3PxeMkz3JvTkhacWSgClL5LL0VHpJoUTaauhJPGIQWiwvq++pVRmxD
qXC3bSg4IH7ZAfs1iOBBwzOoy8c9HgP68YdoBJ54Wb7ScQYdSFptSIqkltuJaKxNx8qS3R51Oyhe
HpHrGlpYzLEnO2lfa0ArEKxkBtNRCs/DcetzjtJrjGW5gTtc6GJQVg+8jj8+GDDjcEzR1qLUfrmU
IwH753xHtBkLznIcvwcvogWppfG+bLlyEoLPSMCwv3hXautzDXbbHaZLhyiOL58+MGBG9DvBQvY3
+epKERWj/rsdnPC9baAKeEew6iNMEqk0UddO0LjGiNRdM+4a5/SnCC2mGjuV40sbZUVpHmHW7Bs7
mHh0PCRmOlHMb2IOb+fb1BO3XAnU7IB+lv7XUAv2xly9yBCJOoGWpw9R0USou44jKuqKiZVp4gT/
xE+7IqgaALaQUWbY4/PH5LpEkrb1xA4DKme45XSU8zxyEpkQAAZ4nX7JJapMjeDs50WlLg5iNdvz
rf2INKJiSLRNtSWZWoFtYxcvMH5VM0L/Z4Y6RfN9bLq9t1TCoAlC+xyou0Vr5+TYupN2on50EaBi
dp0SFnhxa+5HSQj1sgUd1qJ9zaI4PgrRt9bzana/VSlMugLh6oW31fX8k/w34qGANa10HnQ6hdEy
kNG2cEzx/zW5YkYxLg04K5SsZvBCJY3T9pp3OcSa2iNbZMNTWTRZTXuqwN1ciFb3U050PWqCpWWJ
22VGN4cmBP+5yMpcFvOGgn4dKZxvqko7BU2YFvo7tZtL4ez40jx+tNxYEFr/Z8XG9JlD1ptEOIbN
dbka4v2db80SpYkfttslwF9E+kd/RC/y4jw8Qg2hNvf24XiFLCqG/ohbzv/Gcmno6vISgZ0eo04g
oSGUa8ko5Ja6t3kgVDJm9Y+RZPuMoVYqdw6JzyDpgaWAUmlt+AUev+/ZV5NG9k0lkAMqaggMgBOf
nt0dn0wpbJQvVhaMPuWhbdJ4uLDdlA3gVnF+ZCVB4tOm1wK4OCa3M/jujbd+eXPAX08yVhlZ97I6
yyga8aWFTCNy4bVFfZJqRYNe6CNXxFg5WLzs3M/kOHHwiRajFZWpazFpfSiEO5RufaLI3KHV0Vmu
rkI+JmqvJbh5yo+dKEkCPBysZ2vW25HURC7rGOBCdxAqzlBJbcCU1Gfm1XT0aVbz2SeCcOuvX0aW
Ls4uIG4iKKd/DsVx6w3mCyiEfbrhdKZt6L/SJ7GmEgoq0Pop7mNKxv4Zy4VBhIlT0pkLusL8ava9
MkeW1NpISbbuUjSh5XQfDsoJYqmkdcVuCRTXaiVwx5LDvszX5lBq3KutmxUDpFypwrGGExkBy1xB
fgcG19FePKiKs4fM4uVZvPUTQf5fXwtL3gpmnoNUYZIBc7X/7vPiK8i0DP6jgj6rpmV17ESuS4a2
jQFdIioXmW890d+AjWFMSE76JonIpRQgKsys/sCmSvB1lmnPFvvqrTgrN03vyz/idPBJBXQyfG9p
pAOrFujKWe8+v8Ypdpc8pPPe2eN9OubG6aL1MqCUTyGcBIQmnZoHW19kj/gjGvxXZPn4EcjM9dg7
MrGcKm9o5yZGqm21vz7s/ljUuzeLF+wwQujY0JYIlmjQv9jxlGGrLyNRGhctFw1WA76o17BEzaSR
4x94QhYwoFD4kqygOifb3FmmIskQCiqurbRMufczCCjjP5GouZSaDdL7XQsl/Zcv9KEND7nAFobj
ra4e+Df5Q1DNeGo3iBPnhOhOwY7BP5QRKt1gQxbrOSY8yhc/+FOA8Vvd1Ah1OLWPFxy7d52F0iS/
YunPGfbhbChLLVnrOyiSjDtjl/T44EIPukTaMyBiz0d3vyvZ6btzV6mKe2LkryoLguHJhj5rn4rX
i+o53+wlRv/8sYvNnEPg/OTvFoJrpAitLHPvTFFKozan6IdB8qojmyH9i15c7pIy9iVJYnmCuMzP
ZE+PWNNbcJEVPHdVHXGXAvYUwuoiZz6jHuFhM519/iFGrP4Qq3SRyVG6wXrSYcbtN8UR3mbdctbs
uyS2UobPyhCGnXHQcebM/zYztt5q5aoBkbhVOv8NCu9034xAoeDCv0eyehUrEmbD0B93WQjhBFYQ
8XRJHbZxdTZVuzFT2OhpLN5dj8ah/VjQ184X+0LvzhaUE1DvD8FieAbrqjy2dbkonlgzOSJ/NDG6
eSJzztg5JeOPglknsTB+nnBoNG54P5TPu0dZMF1rbM7SORbj5/rhtzFydL/bcrjFkGq0mZDA32QT
h0evsBNvGa3FqPe9b9LnkYjeO6z2eDi1Tt9nV1O5ViBDyb8ndusUIAIGN9m9CovVNQe5cPofQRr2
VnxPyLAfpBsSj1zIjdKtxKXA64+541/xbvqO4RRzuM5SG5qfoytVV669nN7JaNl1DSFJAHbe5Zce
6J3c0oTc+rs8zCAV1If7NNVX0GOG01fFTBo5tpJ/PCBsTnLzN7uCoXkEbYQI7avYSu6y7DUgk6eh
dsC4IbvwB922z09OF9fpe7TMSp0CGhsQ2aZ3DI5icZW+3nK8EJCcojXGhQLK7gnMyEOYo/X6hjV2
oBp2k9/VXOqanCAn/o1aBp5HTU/ijBvf27u5yEMTmQbcpyFGUNHbY7IeWHTzRBBsDlTJVv4DpbBK
ML975CXE+eZiu5XkEe86H8zYFzbx42qjddsIUcHzWNXrQqPZCec1BzkZgiDKE3lidUk9ufI0czHu
e8LoRY7qAJQfp2ePsmtKggwOAbh1m/73coMN5M5fctPh7Jf/hpEfaA6jaRRZOGywc3lOSS0NoLfE
3Fj1y3RtoMk+rliE7hg/f6oDGPxoMXhJg6imTdkfcZx7X/neOgRpFihD0tS+dHHfWd3VoogQ8tgd
RMFJaFZxUkQDHBqTQtfjehRUX/ilZ5ZjDG2Vk7swwFalWgBFZ8s/CxGynAB5PxpQ25UgOsfhWYES
5uPFjyfgPbPJBvS/FEn/78NmLkIS/YRE9p+opSoREJCq9Xq1o5bXMBjiXx34lsYV4e+YLwOTCdZx
BLdhnSUf7CFDgTZz+KjoDpMtXTyJ+G23Z/XhG9lau8aVAYw9wNjoPQuPx1VO26W/I/i7MCG8uabb
4kR7MqzfqgBWpv6w6K47QfTq4TDWuUkoYWFTGjLip1vMMD5eFFpzWeByIu0FkwUUT++6YQH3pn6g
4lIkJZy+EuP+dbnWocb2CKUpEq04QufobQLOA1qZyardbVDkpC8uws2hKm30dsJrkRPbqdWjOo5l
nt6xHEIkxrBiqtJrGRBD+plbOT9okncALEWtcKQVsPgtn0gLCH8DxbDJj2ZMeyBkNs7WI5qs872X
2agal+mY6XrJv49o13nqU+L0oHIQl+kF6TRX9TOkeg08lpRJlfxeNFHXV272zDM/8PMYKkcs6yz/
BteiwO6jKXS+DnnUtLYPTbKVTwIAIrKFYa/B6YrUAz4EnWlooIDIrb+IVM/i2dRpECwlZK/TKLA1
nYgTvcBtNtUIgREaOLiSfs17xNH4tLhyiuMqAHgQZ853TD1mMDqdmYppd7VF0LD8OGo0T6L6mTjM
u9LZKQeJSC9rs5R64FyAt6dNKR5OYwSmUYAaPTAhKpX9wgxTFra9ALk9WI5kju45iTUwZ/uk9zZ8
lwWr8wXLqsZ45oLiVPLyb6fJdS6H7FOati6vbZGF1p7JLhxf9d21xFdZ4DeSLr/+fQeUt+VKZ+kA
sSgyZ7ZHxhCyhXVxV4raqpDHfS970eWV6hZyXoxuU7SDGrIBtiHrmiYLsr4h0Nuwqys2zuBrEPW2
vwV7cx2xtdpe3+7dD7c0LutO0nBbYp7Rb6F1QrpP9BJFMv+4Z52H6iDls6gWpj7RMGnYi0qBTMYO
i4OcaP5Uts2gqcbylEhnrcl93X4Q9t1IO/HFxI4wUTEX8XonR4EVSrzQic3SIPqvmCsi70rtpp5i
Xo1+q2HaQOE4IcdlwzO/RscUrx5Tpp+x3+8uO4MtTyswohEdCW0cajjpjixUL39UBzBvyzYQbnzj
ffy/unOgIb9sOCeF5JmbW2MOZxfe3NLwi9E9T0MocJYxQsVmtOTMUafGATF3wAbOIu2bQ1d428q2
04bd6pI0XCB82l2rFWsNGCKQZbZWWYoolVBr80y15NpQ9kSJIkhaLxDG6GE3IqpjJIJyYu/uOG6W
LUpeDwwWwdogJnbS7jLQVTjlqmpXz3OqymaxUoTtgnSLEhcT9aiuVOw+GEoLVlVRFx+BUVNPtv1q
hE25D9QuGGJmQy26NVMgqpjqZ46M9XhhXSowKFOab9Heaj6qJmO8uvGWEXr4YjvUFnCpqhDh9Rxj
yQJwwbrMEGV1okgHq/M9Hwc/B8Jp2SBDqFvFeOYRyUJE59JZWqQZ1bQDIS6kVl071uWL1BsYztVP
3e3DisHTDtkcDNRH3YorruKl6+Bp1UFlLVAybyvqP3aLIk8UU06KmfzlXpo0WSyaV1/4vSgHrDa+
mLuiZbpZyBRA/uLyDyqvk3AgsrDmX6ILqGJQH21PZI9fFxYKsIoV0RB1ljKhNxxOrgIfzHC6RNwc
jDDGSpEo88yRpispxEM0Fn1vRcbWfN9CPb4MMti0Eh4N2l/I7WpYh3ZS04qel51d6mqnsI7arstn
7gywzkQqKVOQgeTTtIVojRRaVzVSugXT5DURcjbPOfcbdhhRkbEytjI5iAF2H32GMPTqZHAKgwVg
lFEazkRYkyLM7NMnmokct6kFBf0l+CpKNqk80foPBRVZwxyO+RTVTg1OMFE+9Vv1KtOnuSh4//Eb
SaY9epf1KxZT+pUM7evS/U/XogNp5N2dKfVY9VYoP3KmQ+I5dfCSa04t+WsbTp9TbqcyVlBS5TAe
1sN+LXk2YPzFT1dUAWXTHGOG5oFjDEdPvadDawDsZUDuRaw8trMndzV+YXBIyDYl2in0BxJ7Xvet
rDMeUDqj9uHXpNe+DNIT6vNdew08RW94AETIvVbG1kdymYpF8SkWFPLo6nh59doeSQxlu6WnyrZK
niQGnvE/+eUVY4XdUMkLb+9bsj2FWOw4UIYWQpp5nXxkR3a9KECN2bglaAPSeYmKLASF4yRn0SKD
7zGNJXHcsPRoJjt1MQG0sZW2XCyYRBUoI+pJOeqnuSuNp8zE+7BgIF+hmF7h++5+nhAp9rjDjCBR
4BE9XrBLSsY8e9Cv6mB2JEinI6N2H/+letT4ZPno63QD1ckHENEuENOs4fhQ2d0r2jqfFChClSNq
9ANe3UxswIj4vQfTWlua1MqrrV9zi5pfzjlVeMPint+eqfj2a9KxZ9Kl4NmeO2qG5NNKV34kw7SN
OCqkLe4uyYZ+CZh49313QvzjMgmwCKxJI2CN8j72e6nN//nG6a30mdQ4FnXQo4Mlj2REHMljLAg3
i5kX6xUKDC1DorAM2GgZ1dDY0hEcyphSGy2Qu7whcT8hlpSsbhMbLfuzA7fBjNP3IQ5INdNvQBon
541quowwLi6Dv1j8lT66kA8c1EU/ilYTYb0kWqYalQwSCNYjTiH9oWcNZWrmT4ga7+F8M/bQnguT
IWQXsBwBqLJuHilqB02DPIndroWUUK1ephvMwK7VlOasag7RMw22BRnR/JUpyQfl7XUSTm/KdaEC
KwyAI0z08w4Njlpz1MJJ3+4Vk6fYRs4CX1uRzIDe+FyTwRcYC/vjApUsmODcMFZgq0hI32fwMmKl
gNAkJX6ZU1ckRY0VlgktagDOG4mRT/7YQ+xC+5/DDmuQxz4e8SGlPV+Epn5K9PwNvGJ//PTme6Gb
2qY0gZDzbW6kPkYtYvQe/xQ//DJMYPCBJ7ieWSnn+2SZ4HcPAg+p/eqhCwD64NfAC9WaNSbqP49X
GlV9AsLFMw0IKYJ27WXBzJ/UVUj/oW4QfuSop0uAS//EUpPE3qzRbypIX+HsHaPe/UEv+/GJrA/H
llelX0T9CzRdB0S+vyRfj/Dtqs5l6VXEEqR39JKAXfMglXqbSC42xwX8rBF91EJkLTyK1IUTplPb
XQR+frdMYC9wIaBfn1Mkkj9Kz4S0GLU7PTGsz5/PoEe1eKXhX/aklA71V0fQww7BBcIF1NPUtU8E
2xcDoFjp8Cl2jzU1x8EtBUKOlctmTjfI69z0rLc0+G6fmVwr6Otvni+kwO61HCfkX/whCvWnkwXd
oWSDJw6kg0OoGoHcHYgVW2igTvYnWrDxM31H/TJydmT01S+6xyeq4nFuSYZULLoTOHfm4Lx9+Asg
I6Cn42oMVd+C4ohEAqAMSAHMy53xdt4BTUSaGkOY/4ePw0IgQ8O6Kcl9E/phSrkno+OpWcnHfC+Q
FG+hjNfbAfsz20aK3leyv94e2NilTLqOFpPakA6Acy3Czyn5IS3Bo7fhXyR2oHwFqu2TGj8HX65I
k2UlIc1DuiucKZQOF2n63PS2fDtKLybIqKa0nY+YJO20alAY4ZINeqBqxjv4ZuVuZQYlrJqR5zYq
JCPSRy0s4DAbhVAwVsArRpN97tqP92pdtL2iNVzMGtvL4YgmulO7tKy8/6VWkOXzbokKF5mqpiK3
X6ug0fjv+wOGAgtHXGYN5gomGvmeQPu4r+ozPB5+FgMUvU4yy2aVoksZbfiAcNkg/Mwv4VxbfnNT
K5FbfoH2a5KMTTuQz0zP8Gynhn42nV9NB1120LqaA/yMtooJAocogbzDKmFSY+Hw8wamTDTbE0JX
2NVMb3x3rRjsDjOclpE+/qiw6CiNIGlspZ6HiPpsgDI3MGx73tZR/yw678Q6oW2s11p6zNRkmQRB
z5pMVxuzs6QNVQLaLaZ4gEdak5un51uKkjrk86KarQyTxhYfRNY/tvoCfK2o1E/JuJfezX2On57E
Bh8hbY1ckexZ2E0GkjFh4Vms5vCJlgk0kzKoiKigvomTWXKX9tOsQPh9yR8rRqZL8mDJstViecWE
ZC2p7hk58fRvuOBSQzG/YOvjnUIUzNbju/hrLAW1TfbZbCOgK5/OVIJunzzrrOugbBcvPs2b6pqV
LqQRLzDO3lodaCwMl/hz1e3qmhU/YgoMmBoLUpN54R6+JWSSUDBfBfjLScce+svQ80K2ZKKECtC9
2vOjItJ6VyT0TMdG7T0Xi70Yp+EFCe4UFAlHu7vgWTUuDQ6j8kgVQI0erHqsyUqchVNCsBlr1196
OjCLEI7JeBK0pZcDhB0ylnriWO3hpokNOr+a6tpQ/r6f54D7ow40MIyyrfPxR1nss2+yCKNijG7J
3/yhnFELOGWSu2d5sKHC3btbFEjtiStxws5kBUl5JiGqFV42zOSDCLOa2SjnNMyzC0IAuS1saeag
gn1seB6FXeqF2o1/P2+pipkXzuLZfkhXoZ7ClfV+POfIK8tprDDXI8duYFW6CTubmfRX+mo1bkAf
XFG5hWFh7OdYY2xNSXY5CiaIyXl/fSR/Rrfiuo+Qs3RHqfbv0Ihi8mQnXvUHOZ3ZDRVwx2QLMjV1
m9NNMEtvcD3AiuHqcSCpP0u4U2e+mtwB62HQDEgPkLFbM72oOYpU+DiWJhQNDAvdP7CfeDDE5SNg
OzcFZsP+ofW8uCAjV/9GW2ljwX5WSZH+MvoN7R+TEiMcraSl3p/0u5lzgNFH1I73m1GcIGwF0oqX
YMdWcJoRHAkh3HalLX7N3oEp9TkkK0p/HHFqWrrnh2K3nYBkjqx6H/k0LgQsfDUQldL4l5HmYfZi
IedM/pUYoZ44EcnZtOUBKrj8btbgIL6mmvSoh2lDV3hHhXS5fZ135DoMtnKEDXFuScU0BeKtR0d7
R20M38Ex3ZeEVfNyAEL0TZUHDBlLDunPzbB0ckjHpz3o61zrWcLdC+jQNT2isNckJjz5tzCb71G3
TAxOx5PiNEtNOpTm8IFTGoZm9qXWsvGBHuJTQ7kDwfOav/7Js7l2q/gNUmBabY6P9k699x2uAfKE
Dbj9dS+NoQEgkkIBwhVW/MOay5BDiAaeTjS5jAm3C5xFnRiKRbSu4W3+iF/hqfzPZ1XrK70cQ1Ze
vinny2APIbftcOqA+UEbcoX77DOJSX+np5u4ICUNMUc0CmR3PVjb2BFd5tPCyMnVqf7qs1QWcNhV
+IP8poMtStqRp15SuZwYek/IsWjJXL+sokhT7oh9kqJCidGihEJ0WUbZ1eRIHD4ANfaCihqjakr/
5SfNyCuY2aafmkwhji+TVjdW7O2xIccSYMw79JGEqqp0FmnZB1vqbcxTiYKNqR7Y/tPcv3SQdMhm
T43QTbxNtWs8wcwq7B9H2r9ckxwYCdjW20MvIDAxRulsoZnEYcZAyQbqBIl/yWAoVDHPc3srNdYU
eyoL6qaouL/92p0uvKbi7yPHCvPCxzkdcXRGnGxBZ6hD9hEVkc0LgbybgXRuVjPq2n7ku/LKGkqx
KUwBeLgcMmmUTaLSE6hblsxbXOU9ntHv+qLdtI0WKNOyOMGlZIDxP5LnLBDmC6+U6UvbusqsRuD1
hB1R4GvwgcGM7fRKMIvZl/n+kFTZ6JNRmlzr+8G3s/R7VDWtrHqrjDoEXG+MNS1UtqLntLF40wOy
PEhogBUSG1esGKvX2eq5efQbHcI0UtWZCn+TdSwO2r6q63ukchn1yj5Dkd9r9VSaV5jhQvWLpof7
/T/qzUz51U162Tcj0UrXMUOlmnLHjoV/j11WtN5KCehQkC/DU696pAZp8blqLQAidZWTk8ZlkLcu
6ViHNpTWUX7xg8bbJBWpjv6GJr2vmxGCYif95xGMv4xe24be4orJhHkuS+RvxjbgKK+dBuFMhujs
0MZjQCbKBPwTQhe1JDSreUz76g+VRIzQcDDPys3rXm0cYUzGL8ceBeZRpwIQcvdgKQdI+O1jFk5q
o8vbLFO8mnL7vGrchzc0rpk//Oh6RI/BV93rDXuhkWewesDOOyBFhRkVhKuQqTP7S/9zXi5avDR6
IoYwmsQz2rAi2kfS9KuPVKZB/CVOx4IxfUmFTUZa223hSSnYUgkYCIb2PpQLon8Y3nxktHoXRF4U
Bg3KcssBA77IZ2H0/3RETOqFHwneMHDwI/8xpLGOKUY6eOs1wl+OjBMzF02RaohMPJMzYv2uvlMA
ixzZ2DHyzOgURUMD0EhdqJDwv3T9vP5Mul45cyvmn6DDDNtkjBs5oum7t04xjG9yKfNHutK1xskX
q369DZa4Lu4Z1EDtdHZGoL/Ljz2QNDabFRGVpYbqeBgrmMgXf2bFP1aiojvlU6d8ypMK8O6LvnjN
VhW4YzBbw1jE0sJkP+PvACqoj0evlRiAjQutDiWJafgAt3LG5JGL36cZJ8AJpyZW4hPqvlH6dWEk
EIHAwa9qrz77s7U4Car9epJg6I+brh7t6Zp3iUsF0K5kQS7dcEAVUfcwRJcdvJOfnifUFADCAJwk
5NLzYZtTwXlO8mPbzXFgcnFCV+1rHMpaAmm/SPnZD0LHDmxqClRmDiXJ9vvRyGFK7SCW+/H5vdBa
OwHZVURGADTIJ0Z6jpmX5YzA1L2U++c2AYBMQ3H3HLnCU31IEaEz5+jjBJb4rO7KS/hErhhX4qyE
Cg9Nk2yCV4yOlIOWVH9iy/RkOQrjZyur1X0D3pwaWthDAo5hxWW8Yfqjj5ljvLlVtKkc3tTVVDe1
vubMBSHYMO1zVGNmFILwediNPQc1IsFaYw19M1yzCVHEmgEBZHBNKM9rpYZvGxy55LaeDeBOGRg+
N/28UsHT7nS0uu+dnx5Mc0cjl8evnt5WBQjvlDLVSmRCQKIckxVrgxOmP31VVtJVzKhGoDlnauQp
O2/sWHFWmaCxa8jgFOvBtRV+y6vDdUSaW6BIW7sXJFc9YhGjt0pdHgZVb+6ARLI68JLHUX6r0jNE
hhmveRlX89qXjPEuoeKX50lxLB9EYDsm9oYSZQeHPvFwqhyIqkR/i3Q+9Lt8wZMBr6v6esV3lJN8
67G0x1BHV6b3+tC+yqfM3WFsk8NZPZj9aG/wrGJxHm1XKak5HqQ4iHGzVJkuF2LZuhtEI2VxrtTn
/uxb4YelvNzfvZ3OkqSNQLmJntOi7MwA2AYgdEckq5RpLLOinn5jcY+8PgAyXRcJMIJQmu5rRjeC
Hvkdo5ht0TZ72j2qLJweXdcInEzSc6ku5qft8RvuD6lXYAiuK1LPQmPgVlPqjvOyRhJ1a6ts5Ol9
CYAJD5VmXlokuw9MSQKEuPRnE6Jm/hGPIUslxyJCvuwsIbrec3fDuT+Kq9N8QwV9JF++R+3jMIQt
bonEjDPZ6Rigzf0YDH/925esCPDubluPK/2/JIBUiEEe0PamxDdBfHWTxgSXoFyl5owUxLFsNnxF
VYpSORWB92tqoiieWo+l4peIoLelB46AukmnrfYXqU6yzBfkeG+BXSaRXXcSu+SgurD6G2YFrSuD
2q/3GrMWtk9wC3+QfxcdJdHiQWje30pKnfCpAprhruIVeqqycPTAE8+9II1K2yONsn6ZA19EaOhY
u/6oSmuqsZ21yknNoxjebx1HELg4RttwDnDUJdKJT8uFA1SEi99RMuj8+YCj+IkJhcXoa/z6iQNf
NIVrOfOQnz9Bb2S/HiaVOpkHIBVCxsqG4aMdE06zetWDZ4PPikMI0ckF5yDa28IQC/TXq8SXCSLD
hYJLYtbc5aPLN0cF1m8I702QM1SOqEzqFFUOeGAW0mPXNBeMDJW3zQvs3OOKE/2Ud1rFIJPb0Scu
QsiyPlGLeHVaUrXrTIX1D6Yq0lf1fsY2KFhYf0JJnkaIugp2bzHUTyWFVxn9/T5D560NL0zE3eXa
vugLX6LX8k+3x9xcuzOqCH0DuWfLqHUd97OtLwArKDt1/FOmnQ0rA/JHHZ8QnvKjCduHkz1qJpmX
ZTcGNXgBWVorKOOh/XlndjpXNznHeWzabPN0HEvK3e8FymIX8GuvfrmSI90mU9vEqEW6m34W6ibj
Bx0aWi2DfE8t9XCxr/d3ocpwweRNPqqgL8a9g8NiJn3GVfCgGCeGxdcf5L6f/+0oP626Vz+7lWHu
EYJeufj/bBAlTSfvS4Fm7jJw35mv1vtVpkwhThMDmg/hJnlOLbDxnaAXPr4uOelTdLvAS9RAj58W
OJVUKimtmXLimq+Sm/Ee3qVNSjLtiBZX+D5c81UDcB2ysF2kclVadjjmBDvso6pgpHQQCS/QlNsN
61Y1jq/48MpjRpppYqvdCBdNnbldOoGnx3ZOq9KJkN4HQXfbfgXPMY4G9zlSUfnSpMqGWejmaHvj
K3mCdJxigngCEc5hUWemml88lFTTFjVzHp8x3osK6Y886jeDe+hHmm+qYqRSIGLnG4MpaFcRE5zt
Y4oZh1i3EhAeOl/b/B4pt/kcIq2CdRAdVuz58c5EvtRyqXggCcg5BNPnRtffSguc7UvrpaGP9Mlz
b+TJ6Hgr7fF4JrzDPx0n8ivfpLdfZlYtzVhPGth5du/rV8rC8LiHcLBph5nieBOFQSmilRryNU/O
Ut+Rq6j5zCPDH/3EYb0BUixwwRfgmq6WrMOzIrsrxVJvKKY1TZdoFHbpKbWgtUTNBRi9cSzfoYWF
LvTT+BYkpuhCyHUUgGo8a/43Mh9QNEOuqJ0V/kQjZWW6OT6lpQKzY7PLmdfpy2/1pdrS1Id8KPD3
gUYdlt1/bQJ3VEx1+NTTB/xW0LSIg/lccxPXbcNk3XHCgkl6jIFcwhhZa5dwhA+l11/4+mPmJGW1
DDEs69CNXnWrYD3ifR+YCed8MDwt4k/hRu1WnZ7K84F4k61ArkHG3FSU8/FqCWR+lSCX4YX298n2
vjicRUUQJ1ml6VvYZhA/gnyDJ7t3wKDXdqfCCJgD5RD/DBKtBpyYylwM+GYCfuWh8Vj2pA5g9ga2
LKibxkF+Xx9Zgl/frGJW5gyb/pKJ7eX8pf9BrvJqyGwGVlcwuyTdtvGIVUN9K8E/InON1HBOE+ur
C2bKgT7/aKAjuX6kJdk5XMgsihuTqDHc1I9wkS4P2EVQ3f/nxAWOqi7NiSriL+s80Epf+wyLZzU1
CXznPT2Sa6unt66qwnkOu9gn+H7mkyeKQAf1/MSvOY8qn+bxZ2dhPkctbrnJwYcJeFLXRx70iH5l
+Y2qx0/tIbTw9tJEcbLhkko4CN58TpZjRTlzA8qeTcXphkZHYcn/1HMYRgW4SSYS452GmlUfcZEg
L/wuJ5n1KA+IWfUHtiV539snWZjwPgg4N7ViMCgPR2O5ZWuVTdL1MqHNEI1BwPiiDIqCr0Cu4mYN
x1Hq5zwx0/KDiqy6f0170vwg5mBn2VBUGgPMTSkwNpNZiag5ATOjQPnTV1sjBBX5m/VEvVWr1ffb
N2x3T1kMON4flJSdbp6RzRdGi0m9ETO+F+KCXeqBHcOTsPRrA8txb0Zg1zDTaxyMehCXEyGx58i6
qwgfvsv8w4e7kPAX/AhRmUQvZJeJVswjk45SK0kY7zVCS2gLB8z+29WeLprsSEuPv/mUsCEp2sAT
IhPkQDZw0N8fQu2poq6jtq0Rmtol4E6KxolqYAkEZ7zjaox0Ge0Lgy8lF2bB2dq5x5GVeThnyYy+
/tz/qjkpDttYXKWAjyESHEx3D1EwJMfCVSeF+zNtQ4QcLZkpSaAYC3c8MqR/pmnkpZzxutrSKohk
OMh1Pa7+868UgkR8AzfuyzBJdZQ1dIMeKTsRutTnFYZ6q/kOeMcq+h0NyklC2dkm19wYKTQrt30Q
8MFZooDJ2Wtk68vt8gtpNbUDOEnZQkxV+GEZWMcPl4wlrUszlz1KWwIMxnTUSM0KUTaQqwmzTqR1
ug4GRLbuj3DzhlzBabixFb+Xc8tytxRMz5YIMPcU7ZiYIjFIFkuaKwyP4ZqkQdhw1Ok3XAHZrjUF
usF4zCTtH6wsLa7lpgK1CP5uBVD0DalrwHwjRhI1SW4mutogKiVj+rF5AwqmCWaBiz6Sdg7zA4xs
h1cyjbE9QZ/R5NTrZV3Cl7Zf76MNm/z/xapVNEOfg5eokBNUifXK6qlkSrfJLfF6W6QJUJiWdSv2
EcuGf4efx3DqZvSkn87UZt8eBl8fUlRRN6w7fR6fKIBaad0cZuxMNwg1qE+mslkAeCxQUKUmZ3fN
Lhmg7CKTYpAraMkUmQfUI1BNXCMQCpDI7Z1kUMT+IKuGcpvnZPVTNnRct9YFQpf8YkXDaY1NMRui
Ch77rWZC4cZiQ2UwMUSDMa5g4baM1XBeUJcfjgCgFHU9CAz3CYshqtkps2x+zrbV1F2u6ey0zeBr
05wS2YJ5xEhB6lzlpm7uOFmGFQZBeQuFXPYGoTsbP5XdmO24gs/KTqbQEEe1051yg8Z0rEYwaEXD
xUhWbLxmawwdw1w3cBUke3oWuuYSCTXJSKP+CKPHzhW5YuarKFwiSjuKHJ4XCIrBujLZkgMXYcke
HRZlI4C8t7d3zYtpHA+K/Rst5V8eMGfXKXD46rQ8lkOespx2vVlXWOfKUwd3XOgR9pQ5tC/1/ndr
IJ++ICc8LHz5FG0XW3noPv4DymiEsHYy7+pw5/TtssfbXmmablvfrAk+Na7AA/wOTfKq3Z654mHo
s+Kvqky23gvIL+7D11AQ1CLZjLSduXMISVVUWg5t0egS4QV2D2Syp3ddNkBQ6fAwbhZcG+Tg9FZO
3OTW0D9TsQCZpOYb9lzIh0HXuqHyMyGGJ2BAFfhElaygdHLlc3RmZsiMPORinGACyJ3cQwAZr40s
eXFkpHBV+xNeUtskCpV+6xI9PjkXPkX4VncEcz8NzogmfDsz0/Epzy9EzG8M0R+bgLG3Dlb8Ve9+
PynVwOsRky5kMYreXdwpfCLwVr+tw5JZvbwW5axfUjIlVJI4R6rtikx7K5Po+a8QCX0tuuWTND/K
0EhzWwdzA9Yf2G7yNlAVbM4QmU86J2r60W6wUsvHKlKNaig+pFcAEHpWyHSUXmGNWj09i0uIjdZQ
JFZ9xPbeMJ4CAsSsLTCj+CjSz8XXjejvnBSo4MeME3GSrmIrjEXL6vXScIxksdRPFL2e41veC3kW
1zi2cv0Z1Ryl1LbNcI53Ud4qXrAOGWU56ens/jX2BId09SfAUM5Y8EcYWtvyo6ND0iwA9pkrwlOh
ktXDPwk3HVyhQu1UgqasomSOTVcKo/1jqGF6BmD1PzE62wulyV+a+7zVF+wFvlxPI5mOM23UfAR6
+w8sJNp5uhgcuB4Kgl027SjJsHIXL8pM73lCxPYxHdTe4n21qhT8Cyg4ekwvxUMafPwblFrUTzNJ
5y/Z/d0ODXaThXN8EnqNO2+mapykCQ68F5D6QOmwklFGArDKxj4hh+6HqxqMwNi99l8MTpZzYpt7
MyliXEuPKEe6Fg4Y/CjgjnuruyqotQrVIgYgr9hVB2JctRwx1vgupcUfwWlGPvITaYeEDI7lxzZy
n37nPCtf+U0sDKohjHKqzbh38FyEVFSt1LDu7PUzsYxwfue24qyyVXgfv7XXOS6HfZ+qvRryz7hi
M3rGvqgLwmL9eaavDmFNlvm0ZI0aIkNR0tpPBDtOctVb2b0aLbYhRvY2NcU5qItZy52H+yy7Y34R
3sbZgGmH0mzsO+Sf2Sd58opuSa1XJlI7vMQsbYRsxy4Q/lgCyu9aFR7Ib9IdCJPnRvwnD+jVHrJz
DMq0Br9XeVzlPLtnlVezrLSM2/o0Qb/SM5/5VjmE2G5waOWPYgwmjQ/+EQ3R4sSBjnSD3CURvokp
Hm+mGbFj8zrRw5qp/q/kYC6xz/+3fzDZis4PhviR6atTP9CaVdbv0BkDNPJzgmwwjuyjuhU+IvQ7
E9Q0eOTcqVzMCiOHxDW6bvvKcuTKux3iGtQt1v+2Evb4adY1ZUBvpam2VAFNaaGk5LBf5sTuXGyE
/N7ZSl7A6/bvr/EmE4WgECMSbk2N/qiq7uNOIeVLhKwvqz/3x/+dNWBUB5wtRKpqHU/ptQ8Mza4D
N2/Y3jb9WXFB67wS0MBRugYvbLUoR7j6UDEG3dZuvT9cjzgAuIUV+BwwoKdeL6HbSTRY8PnPg7SR
IhDe7fPtvvH2IV86s9tkfbVsGmLb0hbLkdZH+//59K4nW2Lr930Gfm3F9Whs9Qt3PGaiLOQNvBYk
oWKbIQxHK8m5IHBC1dsYqeLj6bXyTj51wrmieDqtwAYW5Q9/KJWHvESh3Cmobj16TMNWF94pqCzg
QAP9evoFzCzFTHyL1ILBc7m3TyLvo8HZviJNNJNauV+MiNM1OKp5yj4/9X/qyr8fUlS3f5P23HaH
MHIZCAv4WNugLHEGGxG7Tgc+s5/sBKJcwBcvk2nvsLTyhHG6LjW//FI9G3MQ4i4RBGTlOc5yvqYH
HR2+a/GVe6MHcC2ZaXu1Hh5MrHQ6cNI+eXuzJBnjypmHEuRQnrM2zvFcvnlJKKQyIRhcF8oMhSFK
1xjJRxas+XOA7JhMuQNLO+sxAEuLsha5bbcv/+0XvE/kviF91Rlkz7LqB1R5yZ6aUUJFiFNSTRRj
y75LYWhxLMGk+x5mezB2Qk9Qq1cNs9R4OyRXMiWufVt7/a4u6Pw9qbbeNbi2s2RVsOSqmOW0Q6rL
0M683w6wv/ut7YnXczRGUjWK0uX9B6A7hg/a1nLvIiG0qkgMS6hOBBjxpjxNd+BRxwz/i53qd1D/
Fb4xC12I4LjiPoTVEnIhXesI1vtwQMwD6J4hNtEB3ZDU4XTtKL22zQVTomlI0fQjsOxKLw2Emwaa
OAOIZAuRzZdLifQcQ1LR+U0lEgX6sZuned8klApWljyMmTJD9tx3z71QeynbzaEllAtT9+7FdF4K
0LsHpLDc0fLIUipxUjxu/EPq9Q6/IN9+jUmxeMNK3UQyDlrordawSy1eLg0QRqOndm0X1anD/CFn
DQ48aSPKiueM0LYteKYMRODI/KeBjcxxJ9BimujnF3/p9MG1HPlwooW5hMkPhtg7oja0l1+WL+SG
XMqnYAzsxIncb3Ea/mez7+TyqrGJYz0Jb46ZduIDtySNkBojw7cwG0POpWoLDYc0hobL6OGgzSzh
f3Kj4dAhvALh8KOCEjx60AVVapTGF2WCArcxuiagYVVILFRcjZCMLiWGvTi42PEj7S3R1j5rwpZR
Oyd190hhwB6Mk2HQb5ahHLzYLGVxwUVGPqTrnHWRqh8ADidqtP3chLUsPTdheLoBajf5HX7UgbZN
EVBwR0oQkEh2VgIceX4pmzC7/KEx9WTFcK0F590gNXpZTErUSLTkJNdS5rjE+wZyyTriRhclsZG9
COBgPrkJ7nTuJm0f5Mx7tW7nqD9fwKFd+FaokJqeM+6eKrEQtq19+l/dXbuv5Nd7+e/RgMF75gCl
ZWxCAjIAUNcoTl4V92g8WeQ6aqG0eycG4MFFwh1JCg3JPbGQAVNR4ahzBDnKYMeEtgAw8L3xnZwB
CtjASym+O/04seThZKOFjW+nMtpsC1s/HD/OjoPGQbCEEQAGT7XdXo5M6F0kxWwSHPlkjvCfhEnp
vA+Ng4fyJY2OKHWnPndYR6S60x6GCVCkwTaSakSCbG4XCGYBvY+uH1iEzSAFXUYMXneERzHw8814
dqniK2E2ijvYWzuQoe/HH+yFtKqD7h1TU/l84iaX8DmmYgW/sUcLlFXH71GlbKO9UKab4Ln3DNYx
jYwcSswECvmCJuaNCLTT0VV5V9Sl/u/q2o2XPVcyB0AZ81I8+IMJQyk1df87OgYx13JkNR4LJqLR
gA+cfd+x/1aUTtD4bAO3FPI+hGfunsloSIHisU6t80Iaq3y4bGbzry+XsiVJkpCscSf4GLmA3Zpv
QhUnlMXwiKaJL5zoQMflCDP+cnc8p5f+DDr1ff2ykzB9meq6S4ehYL1F1WUiu0j/yTLP4xYkKY3k
Le/aJMDWIQnxLu0l6SJ0xsfeCXYRylUwslyamK5IfUvtJuqA2yWSr4EUY8mqaPhTFSZB90rJq8rU
hdRVxOKxR5XqM/P22pErhI0uHD9Qw+EtFLpYyZL34ks1UU9OSOe9B/2o1c9bWKXFNNFNfdpgWM7Y
vXum6o5U/mTJY9wN+8ZIiGx3MQyBKuCHJ0NtAe1W6xMq1U+qB5sWXYXDvCuxHkzcNqILpoaSvcB6
It0BKXbUoiwZjCuVVNfxBaW9HjTy+Ya60v2YCdwYnrNG6FybUceXErJM62PqvatCNIxVBf62sv4G
CuXzuepBm7pi/TB1DvtUukkjRImxDs7DYLwox7Ugnf+T+zvb/YavEMYzAtTZc97QXHLVXfJMi6+e
IcNqGbEmtxPaNjHO5VqLrWSDwKM5gZjBBpJmDZP6xCHwCLq5Ud6ZysEE35myudIDSKDZnvFJ1N6D
NUQxEsT2c/TDO++fR2LDNawN5qp9vmKiYVLOzMcCHW/0rpuhDZtuw6xRTMytBAYbfLlEeFVj2I/z
nXeTp9cAwkDveucM9wqXewlhVLn41UVUj+b6GbzFU8qlVlJnDFMpm0+FcnS9EdKjgBQXupCnP3Xe
ZCreROKRrCeSYEL0kISg5rYDIetZM4o3ShN4t7rplH9rliVqLdaboaQrvO8ZNFYx7AsCPLaYVpzU
LwCC2eQPVwIHBnngR99waI+by3060HmGvOpphiGTMtHiYgjBylB0EghVl9kenlm5Wjy3q86kum53
5eShVmhmn4bgKT5f5JnJ1ckC3I+br6MJWoVc4Jn+1PFz7RRpopqyXkRbH/iFBM2NQSpPnOcscwtc
xWKKNSBO1tGTkYwvGsz/iduq7oiEBwYXR1oRYJ206fn/+jV1FVJ5dgu9iALe2QFTv6kjbj2Nr++y
w22Ph6577g6HgpVrXfQSDNvex5ylcITvc+eUB60w2swhmrvIwwNpLb167oVCRMgoxDpvLgHz1/Bc
aoDmx3BtJonKUZUu3ZQprUIAbZGYKPjMMPMkAR32CLZr/33RlEyzBIzP3yFyGrA8wwL8f0YgEnPX
ZF78mQEH8unSrUZVOy6jRaavg4GX0bExXz5cDi3wVKSMJz01dVqy2CYKu7pdVa134hiqoxkK8CN2
ocLA9monoRh8vCqe/mlAupottNQUhSxkq5zaZ+2Lv14hLA0CUYuIwXLTW2ookUcSwTFk46SuCWwJ
yiICO3AptT1d9OuF0pU7D/NiJ+4l165QTZOZvmG89BlS8eCWanAuaBrxnNDqQ92N7Oeu3Xs7Puyt
/zUcgOxD+uYljOpT35wsrB0N9wzaOICYlsoQcVVNnj3TqgPDAZNAzqiVLsCDf8yLoECcXw70Uvyw
HhLiUkV0l1uOuAsJPoZw+L1zFrB4Jpz6BiyJjB/3v+/yW+75OvkW+af2ndmNAWaI9TqTZEVuH/G8
TcjVjFvzJEcvICk0tCPjO5ZFfwRbNYo8/LrboB47l+zmubzSHJfSy2K9IjmpTOSBtQyxd/fFuaBt
w9Wv7DBuKRDK/TRZFPgaFwzXiUP3Pok4fjYBzkTRd/zOzZNaEs/Is50rhspersk2kds3lmn6MzwE
Ekn7EdoRjVhaZrQDzfr8tifU1DfNGdw2BzXMeVQXEH7Tj1Ghyu+UuFh929bTbfoe14SVISE3iIfc
3OHvcfjArtzxlc6od4c2t4TrsHq7enuxJe07Sz/rG8g7LWS6JKeGWY7RoL5d/BjcbH4KwG94lgqD
SIirv4smQ+iCW+mWKFRd2CTnuEc6Jgnf/u5IBcj3Mh4AWStPY+Llk4pdXASTtHDy0j1EX/Vi5an3
nMG84wdQIYyMm1ApjjwgsAv3DH+HXFfA13orRnDlawLRfNDLEos4MHVur3qbAMqMuW6jcbevpHSq
FzMANH4RpXTQusM8oMCucEa9p305YOfEGlGAkG/auT7htm/jWpLjfHxMvXsWNcGBAL8qKQhlzIcb
50mMVpHysfO+hmRA5Rlc91tUbPhG5wHtx6OQLC02XgoaonS5BQNww3KUxogklF5S9XOo+2VRKupG
2/NbJSshTt5J/cg4hmxYeDVt4ht7nh7/qnU//scTNp/lG6L5J915nahHAg7ZpF+gNcH10V+KpIoJ
H3IuGEESncorQAqFkbn+TKibfdsg8uifFlN3xUtf96KwAoaWM3vr464PzEZoqdHLL7ELXmYztayu
aPBMdzPakmijYdR7nqVjviJOkyfhWjdxJgnizGgYuWzlRp2t1OTUp7aUgXg3JWlqyQF+Uxok1C+0
rzIfKJrUm2UFxn1/d4fEhWRynAQAvmeww7aRZOjnCGcvL7eu5aZU2p+xClFoGNu7ryN1GIGJ4dZo
IUgYRYAcAuoqslCcasnYrCjA2NQbEu7kZ0pfWQwH+fHrjma5bKXoakzjuTnJRXXoBCC2AzvUZIVs
5qefnluWPhn4wyb70DOwvjFQ1A7ZaB9xbXuK3lilfYLLVMHtyg4kpqL9Gw8Wkr68aG0Rr2Z5wVzy
a3hX1R/3QlmyKRHRsZnnqs3dgJuLyRb4a5CeEoIrWQUf8zRT9WWisN1U8lRLFJjzfXvHDmNHABK5
2jySVp+MnwAyTFMRaA6txI2tEx1ekyWPI1M6C1epaYye5mhsdTbjA0UasLDI99L9janCIxxaII/3
QfISs6L9+iwWs/SywYsAhUyje/xopPYP0tgILxqae01r0IP+FxhautxYvoi9KkmIR7IaLTD7+J8N
8zgVUny3r8lBDIxvCmXaCq9eofpu02p8OLxy7oK+qkiTiyGe1cZzKatcGLdpNzD2axQGBCtlvg+C
tc37F/KwdpYkV20mmjdKfVkHe/EC83b3pn1ngoiOWYAbIY/yjmGo842eb3MfYuLQ9wsqXRFfFEQQ
bKgpzp1S8IlwRQnODplUmNq+151VYrxWQe2v//5kvK9C2GvwaNGsmLxzQMaBCwA6D8HRJ8orbi1+
f1mZtKtAnza+PAKTXrhqDvpckEFZbfraOmYkmp6y+WjilfOTMdZOCWleVsaobRSxHqoNVclx+GqQ
quFHJxunod46JG8Ahz54hYodLl5RKWU3JfGqMEdURN178KU3c4xHfmca5ZJB/BhKf7pVl4gekBpi
LM5dbjMAwOVyj0z1lGZcAvkm2cf3lTs4hdfGJV8tccxMuaJrBWdIotevypkG7VTB2qFKWSOoeh+Q
XJZ7a9WlqW6n8OfKtaskFKgBVPCl44HZ6KAE5rsdY4rAVkneNqb/VkNTS+FdZxLdgzglWFm1W5sB
aAJHTzjDzgzP1LKnedDFOpoHK+rUVQ4kB2z1FikPRql2FTu53yjoU+Ye54+dXiBLgsbJif5I1kbI
9jSpDZLy89HAP8otSmMhrJ0Vlx+UGeopd2BXH7PpKU9hdwT7rY2sYBb/QQB6ZfLvEVQFWNRfz6w3
k2lXr5DRzRC7nVFt1khLTC5iaAsuJedDB+EBGtcy/YuzWN3/lJHBEYpdi1u/OAQ3Cb9ZAS9r0tnh
qPLFVukPiuBCTv39mR6HR8it7fNJzaWS8rptDCkegSIfx/POoCGkdi5MrZ9eGm4mvsy9HAkdSgEE
vEDlD/5F/2mNQfH4r3EDeakVLK71NdsN6MrQUxA9F8elWhsoEFUQwV+3/S0Qoa8C5xRf5y2SzI1Q
WwFBg/a0F3OrohZ9GRnauHAxV+wqA9A/lrs4aaSwNIhwjKQImBB+ca8m6JQlW138RWZ+4Gx6yDKA
ry8YL3B0CwQvqJTzqpTlhQ1TTd23m/TexFtmI2+Bx/LJTmgopkjGWjImgRcneQXNzsTKMxb6BSVh
YOlP2icOnHGCsECFEGff5RWei1QEeXuUUzbuzm/cDugdBXrwg3tRWEottFhGs2QE3pOP4ADa8vPG
rJgubaD/68/k2m77gU2eCg0O5PkngXBPILKaYFu3e/sqMUzys7ayVEmNL1VR2gDXJNjcMrVfchuP
oa5ll8nlJmaj37V73FxbvcSvhAuGoWmxfLBx1R1hKClS72hlL547oa/uXL3tyTKqGrT0UZA996Lc
uxUtZwhVuo2DEbuYpIWzwXFPCJCuz/gCCguhURoPty17s2WKOmJ/kp6XeAv6osgSFiMIIv9Oq5lX
nJLNpGekuLuTfcQATF+vEnXsKEsivPId5UWtCw/gaWpBkhox8+pKqkHcT4/o/NlMRAGv3NsGPkOF
RuwTp5p/x6xFBY123nuiejjHeCNksyKFvTzpotGQRyEdSCziCUkaURXMgTcGzsxCCFw1Q/A/c1vI
2YeR57wlU4oUko1DxZd6N3XOKCYjWPH73nOFVhULvRdPC9ROuERDhHXUB4BzrKuRAfZyIZUbyf9M
exrRY0XTMIT96ZQdmleV/ahswQSP0PhHRu7ZFKF67/XVx/BH3taodzmh6Mw9CNWYffviDcIrHTXU
yut9RZ4/UYmd++RC2ZD99IeI4lqP/MV7UGTpHQbvipm4RgBlCwW2PRNFG4Bp/p4PAoX8hyBJ3v7y
fmi3yCDCwjYr9PmGPBuEzKHxKBnbZw+mQ2GD3eWhMDVrMBwpA2q9+6iWAGDrYu14yUZKWxX1/IL5
ir/HLMH7fzV5EmStXf1yOlXPxkuMTPFLHdc/cJamRGXbZitSCk4ky2WNWFbVGGZIy5jCKn9LIvKS
2dSc0yylmQFh7HrPBasZEXF7YgQs9FpsBXv0v+mTQVPqLNyCkbeWOCcZNLruwe5BurSvYsMabDmn
YudYVsWa8SWnOziMKj9nue6yWFCMr8uztQzG2CcVzpk+9QeJERbHbNzKiVDlxrzKX9HWdG7iDBZn
XkV93GBAdgwiGI5TTmlXTOxrdJc0waeFkckKNzGJGIRy4hI3013lsf7svDOrhqXGof69w15zAdNZ
3DbYhVva9yVSC5tW4ZxOrJGr5DZq5R/n68K6FpvfghboSWZZEdG5n4wYtfbZl5BGI6dRRh8pDYYr
k5wcaJ/qkcIjOH2BP1h+J05gdqX9rMJDlYLKbrw2XfY8ZPhdK6dphJNIycuL+ofef83oBsIQs6lg
YTYxzTUOS+mLCbt5rgqprm6AB5LyLdgqcbvm853koDBC3VgWxz+Rpy0ywev7kRmFAdh0/9ubjgt2
rt0rjZm2NFSFlnnsMSIC6IO0SZW32OIDzo/vbLzwJWsvQ+rQ40CnusCwnSW/YkfaUrB9a0vR4eqP
blCOGgviQoq4OOZkQ/4qvUAvdPJ/Rcy5E7HFq/h7siHXRyVo3l6GXDXiAEgUn5/xcnYubMWsX0RK
b997BNh3kQTriqWhuNm7YuaW2wTIU6QBt0hh/DXTDKXf7/eOeoS57XA+DN1rKkYrWiY9xFPEpe6J
o9BqKetyM/Gbyxo2prIEqrYhZz/eLMGfkjNgKge5KyAH5iMPXw9I4LTXUUQppiuM5IL1Ltwv3kf1
DXr5KrU0FKPK6QiITHBySWMKMj8FGuGk40CpYS749qodATAju4NCmtZL6nzOtawbhGbd1P0V0sZA
JLav2hCUBhQMJ6vo67XARTkSWHOecO0WIm0lEYlJiokH4j8o3Tj9qnuUxhGx83Zt855CHwmMIWri
pqCQos7csBd+CRmtSkZWTP7btaLrPz0Y5CHbyu3VJHVbX24byEChVhUHst8UOylGvTINsOGYA+Pf
2hBlAE2MG3WfStu1t8RNHL5C94mCEHO8WBPQFJMuiaLZuSa/vZ/8QZeY0Y7GulPBNi37Wgx1uX94
jFAUCUfcAWYCREsp+HWsZPmBg9LPuydqoll07+nFZn/TNQaaKcga5DZS+nh1IyoyDFJWsaJ576pu
YwVUg706yukAvpLH2K1srANCTU0Cl0/vZp2/ycUeC1nwqjazp7+x9aHPboiyF2Cn31U3unNhXofG
5Mm9ctfJrmvUAP2PUIPsES0HNs//DMdat0KzoQ4s2KhddX5zPtVNhv/ZrOQCPrNcllgb/tuntml9
YtSmGYj5kv7ip3iFvxmXlkm8I5AtEcnI27VFK6Dx18bBLGqZmMlt4naCesTSreESDNhGT1XUYIWe
IluKpG1flqsngFMp4BmHxoRiYYorrH37r6trEdiX4Uicgg09PkihGkdXltjV/aMiK4ASWtIK5q4e
anMLn6Rms0xl/9gJfCyONXGH/qKwFPkjwIdu1IKTXkjqpoDAXIRJjM9zrhSgxF/Ky3AQ4VzoC14S
+SloHySY9B+T+nqnRzuu8NGp4F5RZA3q6Mh4txviGxjWcyhGxnKu/pGcFr0kg14whEouV//onyon
W8FBgDLJ/7JPedVTKjzlmTVHrIT5+DLRObF7GnFXBh7a9NGT0Y6JsqbtPRh2yfO0CYDg0KM3z7A2
REnDZWc3O0wSHcpPD4AG66FV5k8/kHgm71g68g+TqDCcLS4L1A2Sq385ISo7H5fLR/YhUR+EcEPo
acO4gMhKZepmMSUg3ffWBqR3NjWQUqpGIM84ki/mnsdrmrau2NpDGEeO3ycmCAVXaRSCop8XFx23
3gWX9V6bGNLUvrCZ7OVfDqh+QrkqKsbuSSAJjnuCp6FLh/BEpJvqMa6E300cpr7leDIrNCTaUFC1
UiAj66sKY6dICSAHeY/vRvYxcbiPtQcOJKoVEobvNflAAJlYP+IbLwimXvAhoNo+02UJS91TzXX8
GxxUa+0x6FseD1SxXqiudk6n2YDDrwnlQyTR4jCrjqKOaOWRF54kvcX1eIAgiOPexrQH7sHiQXQr
J8Ipk3YxdDGSnN5c+JyqRx3ioz9qthshd2oBohRkT6sbwUw3NPkuwUFMCUCdR2mroCP/aR5KZKJs
7mAz+p36EfG0/eF5az04sFWUgBV1tmLdi3TVGADSuJb+8kgBtYJE7KFYhHtXgZVpY5qSkPIlBWxy
+cH4fJEl9wyqzv2hT1WR4cHCsTBCc4YgetAwO1T1ouO9sZujRQZdwPTEmR8dUEvg7ESStI7G4JeL
Q+DLkxe7M/1tv2fw5t7pgWxi7+dU5bYbdUWa4h34DAnXHahHGLoXzqZHbeIHtkFC+oP7bGl4Lz0D
a6S/2T/zNP/zEwC9JxR8VArRv76qclpZmEg7lwHO0HGjphwoRqpf6Uvdt8rnncLdok/RLzbZfVDd
nT481o7oQ+lIvc7vYiKNbizAhaL3mdHwQawrylYyHR0Bjg43bwosyEPq44dRlnLCKADhdnAZX+A9
lohQysl7AKAk0/n2OWJzo1V+QdgHd63ymtlrg3cXFH7yuuCqiAZpfFanN7mP5l31sH1XBZb64nWt
k06927oRSmeg7pxnlCiFSuvIsPMlKiuceP/nYOqXLZHxZWpZS5OlEG7kZgg2HlyBMsCeO6brQCBh
AZ1LoluYuYWdHetxbfjmZqNn13SDJ+9VHSN1PunLSYX2eeeGYfUmQZ4Dn2jyP6fE2shdzZHaVQEz
xUYQvegrUE6cwHPKCZRiEZ92QVOnSe4S850sEnHvZC11OUdBD5FWq9HJEwZTO6PsbsdRqoVg7fCW
/Lc4YWJJ1gVSG2zxv4GJfPe/apGfMhxfh/hwKEBc341I/fIodGC+LnSvxYb7rXVJPKGwHi1mFTDJ
+PjCh+RUmlu44VlfrC8nHMYkNUOefsGLb7KhPfblHSmbuiglyhhzOo2D7ezWxj7OAjIRK7ZeARpr
rmcMPkKrW/sDcD2vCePsURiZCMBMQKGiEyLVCMuLo0Zem7R5yCc5yHvzUGqUOQAQ0G2JILXoS4yJ
BH7z7afQVdUOm2POb1TIvGHBgLi/w7VqylmX3FtRk2vrX3NdpLHzKTkb63DfMevAMwazeYO8R5qm
8bHVA+p3IZN8X3019Ru6DH78HHgTAz722GLcDNY0BtvR2/OxLD8syReaN0ph71Ry+cWIpqE2P3iO
yWNKn5vFngkJdQVSE5rFCSGjw/Me9tB3+iGy5cqMXDelo3qyABPGNDN42kDaTCFOWHafDy9rc4so
FU0u8VPNpzNFebZuomNt/X1AYpgAC7ZK7SefW7pgudZsZZjPEVhdAjI4qd9y7Wa2Ibn+t+oS1nBn
OAD1ZssuJdTXBoTy539WqnvkXiry1V56xiTYyeI6SXX8IY/A1lZoX6gy+VYFTAnIP3+ICmgUNZmf
dtX0vEipIxqvtQt5hAKuL62pyjArlB1IPRMR8QkkSGxvO9bu09VgKkdKBuYQiQllo73TUh3vtl9h
21nv62nXKTo2uY/fDjrjTufL9R3om8rkTYsaqkPZQaWEpdUSswvX/RyETMXxPIhxjfg4zL+TDfBd
97BpQKRlJmH9s2mb8uSGBwpM3Pr637XLnw8O+mmfbpNPbuCqQKYvhx58w4aWjMvJ3jQd4pIx6zTw
mcoN4BrSdNFNlalUwbbqdNgA+ukk1pGYteJTPb3VAUelIp5tlPqLlaqOGpD8BIcNGdOwvTPRZxOS
sTKBuJ77J3YOvTC9hUDTSfZEc/RJ/vpKm5zIjD3Jlh86BMxauAzxptkZ3lPmB+I0oOf7Y23rZ+C+
P9w7PRPu3iK7/gerjUqV4uFM/j1vyYIz3MPMeNZKm1L7pn5hHp7qaGAz7FDLOtheIAmMsGzsKg0Z
PVt8vjRzAjisNB2y+KJxODencfMzniu2Tj880i//jIQS8bo669izuxz6aGfpdsXpB1oUb8KmePTJ
4osm1YwutzSS6P+qXI8fqB88QymFgsec8cMN/WnX11kV7xIk2tTiov1Gc+RoXWZfi391pvmNKgyg
in0BR3iiUAtcO6O801htg7NFyLCzrEeRulwgtGxMGNMfDb5MZGLlEPu1CVgEKlkGa7icoeqAlLaA
6twsvmP4W5AlyO+DFgJ2f+8R9VTZ39W4LewFFy4gkOiiT51Mxzn664r6dvub070nFgtz/K1ASPwB
NE3caBV7LKHSm0hugDci3qzH491yJAyz5cvN6hUzyJBwF8ZBr6KRIVv7DAoFM5X0uTb/MkWHug0K
diQVjuQNGj88ohOBfmcx714x/A/UAzEjLGQ+WeYiubs1mlUcNCNQ62M1PKhlad0/lKXIzNNglrbp
mRchr6nbr1B/7AvuR5izjbojoSP91NQzeBSQCDwZtfybUi/7EcZ07+9D1zz2AmgQvTBDcLIqcDFL
lCkr03KEm7enLt+h+8oq/+rluiMwV88RFz4LD9qYHnqXXP3sPq6fm2gsMO0+ssQcZ+dqAw3HACqa
U70HbNWYqEBYTJoIAgeRDoZGJS568N5FONImhRGN3QzXiU5MB3hF3AxQosRPa3Z8K2DA3+chhK/s
SX+2jCyB6GaLWcQarJo0xVlp3kxECg4r2vqK8bJYbMB74/HB6LGYvLp80v9Ms/anOhkPL095YOOO
XBCLN3mj6THnn6BUIXBVnkFJM7NejWUHtqINk6e2S1iBDMZXbcNh+qx1bztZ+0NU48sUvE6unWBD
d3xFgNKGxpL02JizNF4HuLp62eqym81ZweSNcGKHUmkiAlb4u0aYsSk9okm9gFYOy8gFmHqIleka
RO4b9Igs/ucgM5k6WUfZbDOJbQIc1T0KyLLwbB7gIOgJWu7DUPKY4Uecbrb3gkqFEnA+zil8WuJK
6prGTsA0gDa0reoN1ZitZlGISyTyW/QRoVXY39/+N59jErAUKF9OofCzevRj/C+hEFXgvMyByonW
eYB/7M1m7iJSo8hhbY3NRYy9EWHWDTUqv9WhpYlqUKMftAwrriCvXkna1NdGl6V2aDBqVT51iace
/FNqP1TTAYyAm5jL2V4C523uuLkVn7GRQdF1R9TviWyPZUpbDT1yCOkZUt0oBoSvBBYlq63Ne6Hr
QVgvRy5J0GQmV/3Lhqmeohlp6EVkIN4iRvh0lXiIoitCF5tA7UaEoPTsQJjkHv3aaHlDQhN7Fi42
CSpG1wQcuKmF3nu9BtSxM4yb5CAEAjYkxQBnogEFZ+Q/H+sQ57lPguOVyIS7uw4wFo+NtgQsNNmz
+4rljYccka1SmefeyRFT708Q1vVM5B8BChKYy5aT6P7YbIUz4+R3zdHWrSl95UZpv9pxgt5uLrKY
wTVwqA/L9MSjKiA75h5gBdsBqictYks3GbpG/6Xb7iOwU+5N9n3QydCyedyYMcU7fNnXJH6OJ3F+
/5HokZ7DXZ0z3Pzue4CvfN9JE8M5ygkPKngqNQmGiQi1ytd/D4VDUInaFib/gdI9U54Hmj10jr7b
stZNGBCDgLAM3dLhHnlJYJqZOuqIl4nZ6ypwrXfE0qSIER+dteQx5BZWPiBnCPCTthgQ3CHaRADv
QHDjlUZg6okfrXfaeDXOzA/3JvG6BNbpeHNlkqZR1opNrR6OVp97fjSHhZRKW4L/hZtubXpRtlbm
hSmylg6WvmvDw1LIkJLUeYGTSVjpNwdeIyV8xVxeNHAKI/jz84iifhdt9g/GGugkJvt2hePf5ydl
U8G/KWUA2VPIwkWhKZ7RRjEs9aUi0qDEbCgj+OFdWZYgXEtjFSzRC6QueHCZ1foM2KA6ZIN+P+Y+
+zNnQMwGAKRvfm3DrZ8fqeIhC0KiXeHwg/9dbRlJ1xG/iz8FaU0huXmiqUMQu4F8b3BsOutA3CWp
9Y2KwtCnfirQmqTeTYaMVtp17/KdHjDyr5Kcf8ZxyXnm3WKZ28qFluMXPXlJdmCG1aAI/teJLn3c
tx0fkPqCJROWDpWH/bX6SgTPuq2jhm52vyNh+IJRWUQ6GLwE1Z7gZaoWy8PFXNLPFh2Cj3YBN0GM
lG8maovNtY5V1Epg8XR5ptxGXZUltyyPv8g3935PheEegLq/ASdQPcx2+D8OmrlL5SgKLSHP69VN
9VULr127APqrVPbZMfhvOKEt1nK6e9UvHASyeHVSF0EtmtSBmPrQSNLxFJphfoE8cXLR6iLZdHD6
qADT19Vub3bb+s94QvZiksmkBCzqvTkczpHEO+yMeSS21O+TWdKzolsd1z3TG/A0YQ8a9TMqXOt7
ndKkm8kNTlz8g6qBTknFGT3S3ql6+Dpd4sTde4Wmse9/ccrZ+z+z7Z4UFyDyKMSynqeuMjJsYDXH
8PAggJLT+RTiWRxlApK9mwzSpQPrGULdFNvQ8g5QWGVoJtKmlVjxMkdZQLOAUwBaKnL7Pbky1lzW
EyxyWhgs3NUGDcQDhpBBN8GuOQuNFMCoZImsSkO54JVUCzZTdMfPumsuClp5w4w9TAMKSUT+jMpx
tE08AwJRTviquLeQXoBxPKoBuZFbqs1QiPFYp3e5Ac1ffYMgTbFOFnMXRlCIIVfb4LwYbpNrn/M9
nzdlEq6A0fBrtmDwHS1O/Tzp1RvQ1u/N/SMagHI5+ZGWIBaGEnE6KeP4fSE5SWfyhRVKM9u5au6r
xFGRb8P1+hjBlgtMXRW4mhaqrklz8h16fY94FhyJCEeAp2Gps61c/ZoBGMjg+2BIWDDwR3LumhVw
hcO8siRFhABMKsH2/Nw3Va2QiZvFa/6HhPAyq/kx10izK7slG+3XPbPnAl0WgPR5Y1+uCyw31Jpn
+0j4BtnXJyOX3X3t5c+iqNjhpVjmTHYl3ek4ptDYKbc1DA3NQsTajvbIkX5+NnS9mNpDE5Drlyus
cFGAHo+8QRiY8lbctDhbOYJiMEWJNp63+UsThe5xl7Yginhm4kzPRmWV3p0O5HW86sEMLyYzOQP8
JMp5Rqp9bUHgG5jtrmyxMGN8QvUSDgvruHN+BsnGQOY1+MaY9n2cgXsQhazdIBkfFocaAj49ly6d
L2UFLkJVT/yIJgbaGjePCPO+p91+8xdh2SbKumLu40W/ySG4XTmqiWXZ1r43ewVy+IEL68zwt5FJ
2iARRZSiP2NHnNSnFtHwjc1apfmF8JhEx+aGgYDYL/LfS+Ty6vTNoe4xw4EmPzdOC0YnTD26xLRt
L3p4dpLtbF1Hp6VjyjigYZRD9us5WMmBAEKiXnTxiECOOsqgK2VqV62oiAlZVcS+4C6asWImWzSG
hxGxPPmwTFqY4tRKZNh09g56Q7au0UrFeBUJVIkvjgwVASWg2VsxwwBvp/37qf+OyqzyR6jidU0A
mqU9VoGHv0fE1YMtJ+tvwvI1ND9I/1kisOR3JxjdZm+2LKZQWP36jg0YcUz3neHqQoGp/KBV46LJ
E8pjBQkr0Hfs61iIJ9DQyEGBf8uakEpA9nb7v/SkX1D1jlz7UjpEc0vTkJCpzzjQB07gTTRcIof0
AWNltzgnXdFa4m0aO8L/ejjcb+p100ZzMIZ/yYYkMDHZz6w6az0d62PLBdAw5DX3KbbI41bkjYgM
ZSfi7owAzWvAJ+Vm91iFJ4iAf501Ulh2kQI/STwJjubeg9POOjtxt4DZl8s+rzY+pCiO0C3i8b7g
CZQy9dVj6V+Ngxri2G/5tMEdP+K0W+1pWM4o3eTCQqt/MwW3vDbMpFg0AfgWP0Uxe9bbu42XbMIB
dzveXJ6k3LydskUmskcUmcEe46MrdFF5nwy2eD0nEy1Te0E0Sko6MGM5CYSYCfSlVezyYhljX0cP
WAGWG2TeHqPzypElXJEtjLcXZqMTn4KCDP1irKX/U5yEd5AfAVDYDx1LkNsKNZ/HNr+Pv2XafEDt
AaAmmbx1xDCrK0tq9ISGGZT8Nmemcsjx8MdN3f+++jocKiD4S/2b5YPOBC/Avhu6Pw6rqwLdUMlA
MLWqnvKWyBKvB+xBGVpP+QyejZrGgtHLLLw1wdiSGITUhit0gdNYaeUN3otUcAyIRY+SZxauSFsU
nb7/A3UF/owBrrgBmpQo5sRmn0DJW1/Tfs52ZGTHapz+XfbDrxA/kFt9ciMBIIMvDci57rCrr9Ma
vG/kCR9IPMTBvpdexy8qLpnaoLzdxgiGsH1gO/+v8fTad6v3TOYNOVw2UOF5pCFk3cQtG0BfTUVR
reZ1yi0KoX5DQFLIADheMRuhKduF02oWB11cnHCc4Q38Urr/eP5e/bN3YYGPkkHWcZ8RsCOghfk6
m35PSdL9yc7MWLbTUha6hSEUJ5Rigby+3XYuOUePUilVvurjHygpK5IBe58Uanx96g9bodXfnQP4
nzgKFZf7aPLjRKW/Lg3pY/coKBRQYBuhEVTvQcLL+DLbMBh30EZA3YsWjB3Ra/yLPF7O+c4+x/oG
3eCm+lJEUsimnfwDXhc71pdoJWE0NFe2TpLOL9d7iydqN6d+3KSFEHA36uiB/oKC80GAwhn+Uyi+
08bP1syOunxDlVHFNh5zQX+/umQQKUq3gzea92fv7RFG9PuQyqPgAtT1BIVVOtQA/sOtPCdDmEKq
YwR5jQBaLP7KCo46p9KbESRS76XMFT0hS1uGytRixIeb0JwED/SksDPQEPckmA6oFjo9ULD7/1dH
jFS/tf0pJwJbYMhQ9RuQG5r/hGDhfImkowhB4coOnGuQbbmWgXNgnk8ms1dTydIzW94RI1lZxieJ
scHG2q116P+wIRZG5jjxXs0AHPfh8KAc82q/4kfZp5AOcCN9Uic9gcvXIj/+0lyfcdYXwiS3ml0y
1Sk2e6uLZ+37TKVcYuuabiOt/XT7oRlcDTzlTMLF+tDB0/zFNg9Cm3hqkD4lCh+LTw7jPF07XjDm
QdglECr8x0Wyq49q5ttCV/wUFYrWNluxVSTU7SpTy0hknXbZiQHTDzvVHYWVWgQOMR3CjnEotFMQ
k4jlLwWMsGC7+ct9AtzbnL/j0F7X535WwZUyuxX+2NDqSu1+LL3okATojDIhldSe33BM83vHbWBM
ZsTad8j+oRag2jUeYcxMQUUaig/OXTtbgpkGzDyeoyC9ZNYXXmgRg7blIGPtfo8HMYIKxHWfYaHy
4mmA5IkBEFUmuZgvXuNfa8mMLw/ZwkrElG8lw3cbgoazhW/SgRfrt7O1OJrzFTdKwEA1B25HSN8D
wLioQsv6XGgVgVPc7c4JXtvJ4yN/M0OGUvRzL4avuQ0I9TgiQHV7A8uzXhC7ACxlsWzCIQB+MpOi
YlwaHK99QzKPZg93VG0kXNiQ0Dy6kSsuyd31OJsE4LSZMw+AwUJaCoEFk6KXRCgpYi1AKer27qA/
wPy1aHf3+/oY4N6AKk8hyKJ+YIRJBiVp2ijX9VvtQXaeFP4TbOcjwB3DKTKD0HrZgn2QopWv3Ymm
t3KKeCc0ziihc9n5tTWiC85z3BpIL/jjNsr4uii/tzERPxdXiN5hVqOy1+nW+iUxhAE9hwgqHTXJ
ZZOmkM9roPXTmZcnpCp5bt+Pl08Th7sCO4jHs+coxQ/2iRXuUyorY2jOX2dM8MMiwy7gZd00SS7w
ULpNqtN4HFHiYCaqxQJY0BYEPlb+qEUr2UUZZvRVijhjvYZnC+eEHzSeCuR9lXlYCKVSz8jJuvh3
vwdcuGx/cwqSRQu03y4yI5B0qFeqv4YgUOHHfW4zvsX7cX2ngHwmkR1xUaotrD+gFpUg7NgQzH+U
9ZinljoUbV7Cz61LhvK+xVzJGElcP3Laxk9BqIw5kD3r1dsAZ0gKLBqCCczsLS59dSY2pt2XQBs4
pbPcBVvApi4BLRAU/hYKDYzBSKZ1It43k+k2wvqUnwlo+xzMys7GGRXbpGAf3yEbesekSuen9NaR
rlAsbAt2QY0z4gzq0wZsdwMZn/kPeRScpBHEH2FHHUv17ANknMubqHK/hPjdI1gQUq+EFsKqawhN
l8mz95+GigI8T9rO4b7aeLLmkEvfz1a6vICoBm20vutjTqTJKy4O2LS2dzsv8eT+s9XSEQVjvWsi
gnoEtZMlH17jAzwsXDwFNjSg0JU0Yw0ZibzLPdPgo3NlTzxqre0bwiHCCSLcwuUMgGQqxc9jkfPS
HHl4XJKH8RGCwXr4loEpu5Pr/hKa3LM+JBNg0yxHN4tBzh0e/5mo41dErBRlG55tMO1guOl56zW9
NXiW8kp9QSPb4zeyj77+2wHBWA8EhnUd+pTe9OhUDueSkcHTZR2jRMCb7XKJtZ1su6x77KLYjl2b
TZ3i1A+eudRwNcAD/luIyIMR0ylpGxRtb4cuZxHAP9EBfyqIHjsvegzNGufzjXIwE252Lynwh6pm
krBEyqDdscLdousrN4/dLjDVMCPBdc+Q/o7OQ5iQ8JAYkMQSOWKSmO27s6TxLBboCVs/vdCFhppg
LdBYOgehTI/8GIMVeRx5kVMVDze31ZaGZaRXYeNphNzHtYcg4JuFAC7DdyvG2PdNCWVx4u9zf0Ry
xuZ1XJWrK0Z0P91x+GgFMhRuGRJ5Z3lkOOga/AQv1ZXxa5syNzmU916k5vK8eHlSZmExqgb6Pxxl
xOenkUNPAOryXW16521+Qj3JEG3boDWgILgdMpD9TaIBpVJcNBY9CoXnqpri1PkbuqAmwTqSM5aP
g3gNYnx1SUd9SU/cgKxf6yOSuNM94uk3eRy1s5EHTO4/NEgTgBi1sKiZbSMOstxQX0ckyMvAsh7i
TUKDrMI7pZqCv9SJnKIp3KDnyUPAuCUgLVCOm8atfK0bAOBZLL36DHhlbHEXK0NwSEjnl8YPMSPh
Y+S4hZQq9MhjGWjL3igC3QNSwQfIXrx4SR1CPTGNNe+pAwdLpBa2HbuCplbrVv/oB64EyLmojYJh
DXWjP7OiPAkJaAy+EBPBuaZ0YVvXx9990EMCEm99/qJdCFTsOEB9TbmQ8f0JQHVD1dDvEnCCczhc
XdK8bXp2gU791sBe6gDLDtyGxFjTY5hrnW6Zy6In2Poyntu9zIfXEH8tbp97PR4m/9SLxpR8p3cj
FuUBeVAtYY+lFX8JCvbGRtwr+AzYKQKlRmTVOnBR7ZN8M3y4ZkB2KeW07KORXQWuMKcJcgTUoDtP
kRy+xJJ3AXUQtP+g5V7HuVKd4d29MG70tnejfRRxlMzWtd8OnslbJh4bdOCuQfzgSwmwPyeaaPLC
u3a2ygAjogyIHafOaZETHd2L4Q8b6tWYXOLo94lshYqaugmjw2kDIM2+UaruWkmnASoTpVmX65g9
yFHdlb9Ut85nauFpwbPBolw0SqOqSmILATNH1TennhFZsRjR1YT5EROQIUKLxpHpPKRY06OhQTuZ
F1HI4Y31/N1PvUOoAA08aFPott8YYu5PAY+Ve2Hj3bl8mqBU+MEOkI3eedVgDOHt7ZprT0IXYO7G
LmKRMNsFFw5GNZPD+O9hSparxOOmcnaVEFFjOFRweY/NY/eB9Vg8rQ3mxpq4pvWRXFOqhgjp4klN
x5mjx7RvZ/7a5cgsXjAV+9wot+UV4obX/PendcT07mje4KsEwi8fH9u8Zc5jgdK5B/wigoq5NFya
8af83lbprXOaFnuAUelhWbBvXXwK8//G64ckQE3JyMpeZg8VTfEHMsrYxyV6km5UmhXJznuGHkib
rVHuOCLEAZ1ReHu5UkTR5pZB1lIP3sNlzsmh0siIRgyP9MazZiRZzDAZB0jhoGuZASbarCjv37lE
b1RuAJlyvq0bHcTgr1JJPb3tXuH7OLxYI5N2zPZsd0+eODJzDolFiSjlj/lBYTGFI1WNse8/jzm7
9r/+CR2b2oupu3+lZEEiTgV8oVngOipXSJfHTHsN5rERIQuCiy7mTQy8X3TbfnFBdl7i5QnKQrs2
qCQMs/4sMq4moAzrpzE2nTo5dbHVJYAXfmTXx1Tw5zVsmn1h5CHUEhiH4RPhq4K705M6+mcs3v9I
zhsKockdRg6JoX8XckD0dI6YjLKRRe3z54O/7ahvAvGLnhhs4B1W/0LWuOLIX1HQ5EB9awJohfNL
XTHub9jZ2RmKqaiAMzSOH2c3FqUfYOPyC4Cvmp9/A3J+TzVWb4afKJAGIsVUOSvFVDG9WnVOZQxg
B6WZyImKM2GcEIwtBapM48aXS9FeTVPUy7Z896AjmDWNe01xRA1d/JWuYWhCzO5kOg6LeuCpn++4
PUH1YMqHiX1Aa672dS5tmowAdjBWPHdRu/DnTRZCci8zsX8OiqVnWYaekWXnH5V6peyocYtURbux
P0DbvymNgVSZT/n0zdWhBuqFxhr8w+dX0i47LvVAjDO4cNim7O3LvAo4hmLSsYerIpSWQ715yL34
lbogfqV98Gq2L1reXkeNSDnYeXG48MEf5EKBWhx6y0sdxw7URrxBA+pMc1xErMWKzz0Pxw7WtKPF
If33H0h4SQDsf50+iolxfMGiviLdn4pOdcTEk/h7Cg7rDEXVUgdyh/dTwKWIGzrrYFJ9dm8fPIJ+
9FjA406jMIZaFw8yjsPuNLGU/zopTayT7qsEmVQFbhCu1RzojRI2T73AfVLUG5gDU/3wpSba7ijf
j8tC6gnLpObdqIWio3YTsGufuVtnqnEMZzeERhl2GkYswlCe/Lei6FmVvCA1epV2syQgeSG2bmSQ
Cdr8n7db3jWNpuLzRZxpR0v61Aem0ew/SYopwF/aZp7QmLhOl6atN6dYHhmZ8NDw314ZtJQcOE9/
OJb3Vtx+0WYVhnaCqiEaFre1B2HET4t/BDBi7kG3peEGLGo3puRztQjmEkro0QMDh/s0iBTlzLGn
2Ym+OX1VZ7Fcs07qI3waRkM+5njAer1gMXa/7xpK48112IxnHyajz7m0YJMTKcg55MNZxoPsB6Gb
EN37cfKCW4rKbOTiIJt7m+UdBnklowwOw9oIgFpI1u3l21qR4bnmA/XsM73B/jJTLmeghja4S56Q
qjZDsUP+/F42T9bE9vv2w8vuDI0mScctdlz0NzsTx3XxjJP7scD7ov6MbvePUjEqyB+UG6LZzJ/2
V1WioAyWzOgOKSUba9bZPE6ZwFqMbtC5N87uV6n3ikyuE3thdm7yL+DEOYfW2+f85+SGfoqZEmDP
Gfx7d3CELkGiN2AapeQdmmYi7/GVPX1q7nyj9sNcH554YhJ2QgXzjf7qwd43YH1WeKHs3rU8czme
qqh1P4uFb8j9BU9fY5MDKv+VbQWkC5+8jl+53tNRzvdZ+3vEJkiEtFJgu+o5mhLLXRebOdSy7ZI3
gENI4hDuygiGX6S1I8GtnvjPN5gmotdUesJPNdRDdCrYoljzPQGsU78X4NhNcMFeYA6mSFYSKRCT
QE7HokB03ryqzGYnB0OEeBnwjTXmYdnrUODy7quwx+elNLMlNXgTTK2yhsi3qISlFcfvxDbab7p6
xlJKPQylQ3LRyj2Z1Rg7NxpCtHxZuRsd6QZEetuhtU3Nvsm/JkNGuhowdc0F19DGIDh0B+/cbGI7
oFL1Bh96IhHaZ2I9vG3NDFGrOsQBkjPKgWPLhY8bd3Z0Ucz8kr1O+RnkXfgoUILkiZLJIZqQx2MH
EJxPitx/JarKhOdGt6hkbJ/JWaNbAfygdUeF1+37nEXIYTvlYkA6h2JbkoDx6nAGGu4x7K6bY4Rn
k0FdOdHGo8gRIdj/WnvqN259xdZOJTolXmlOGKCdhN5ZHYS/s4lpUouFFseQWMqwkKT6rJoAhk3k
J8cpyZ9IImhKVQg2SMYZLlY0RG/Vxj4GxS4VUz4izCOAxc7PIVSpJv5FqE9a+w9tqdp3/E2z6jzY
C7FQg2jsSNzirwutqDoLZSH5fEKKhv9SiPtHUfj0P6WJCV0S4ai0kQz0hM5AsIuiEzbv/eYa79D6
b31GGSVBbLxfdJKeGQAeSS4Ot2ImmPiPpOb7mD/xjOy5MgcPK/LHaohTTaLmayhDWaaK/EN6lA3h
4spq9v9x8FPMmtoGHvm7NSWQAPooT34cpVz77eHXGyATyLmZISkuih/cq2/ZQUCH0qtkWcn0JO+4
QQXtIS564HU19kRhr4btmp7dpZ6GgscEygbV2hyja6Ld4639A4bDQ6ARPSSddCILLdznUGJf4Rvi
YqjiSARHXurhg4qrcuN03z5kXyskKTu2hYtojFQn0QBkSZzClAtKaCSMmI8XANAhnGngN2HeBP1x
BotMHRoNC5OaZCqoYALy9TYnuOPNh8wZlIu5UqkmYAUAo/xeS8L9X0tkKeS1QXkSaU9GoqZjjDm/
ZMJYswPVnz7PKXjjsGEelMxIUHIRgYfGvhLyqNkdA093PeX1qYiDDHZNz5+C+ui/86I9sXaOd12f
6zeGyZxoazylxGilFzfkFUJX9wGvfesde47J6tmwRGMvbVRM+WDMU8N3nwDAUwHOXm36M3EC2k/g
Jf1+bnyElxS9DWCall7JcUZmJAK2VERAXl/QOAs3SSM9gISt8RVigCrdTLMBPvrqBgVWXK+ogj91
VzYhEGqLBVgYn/Pvfeat2YVpSEOYdiiFbdMmY3/Gqq6Wc5o8z6+BHo9xCbMQcyd2wt8qmB7l29//
oCdHvoJrrzWE8cjjs188UVbKVcMPWACP9udfPeGxFSpa7FIsv21GWHNITv0PbT7HHtLTBqctzFhg
CGL2P1zabJz+/wm9Eklj//RHGTAwpJEZmToEUI5YUQyZVOtGKyLQelP7NlwLjoAf7yCwoaAxBvxV
ejijr90aTuRirc89Usq0tnYt09wCIXqf4adUf+iA/Rl1UB72NuOFYKezymJkwxJr7i91G5pOrU9S
LbChY3FjSVFcJEi0ckTGIY736zsWtqoCQPVGXTJn/hfo/HBwlrrX2JHtrRDLE/6Q/DP7fgjHmqBw
lPrmSyZhYM85IucJUE2ag9D9nqxs+9rmTFdYy7IJX5EXU9R1boQzsx29OCGGUnnAg3IkJJJCFVEH
6oF8y5q1BD2sTixHWGWj8Rq5ITn3VA1316CDqYpvZpq3Bw5nupSlNWJHisoSYjC/C+jQL/hoO02v
J6v96UMs8szZ5W0kcCTAAQGl74LOxX2ouQRRqN9hPn3KD098IhZtHPhVo3xYQ2DvAJTVteez2OUP
tvloul7e7YfzIWuYTS3xRccjwniwNvkX6zwL/r02HUNSkZcxOnPVJhmg6zpueILOpnlHvOzZtUlK
c6AsUl+FouRRcg74S6gxaTDoHPxujzHI6yj6GaUDng2pwaLYkf01/hwhwaRm5p7BShyBd2FlB36a
ulMScMrOjvgr26qU09dvXvXh/R1gwb/zRBmm4euYPc7lMXvTVKEPOTFymPr1xKAKrMPS0EME+t0o
TVMPmaiV0Ly+d+AaZt7bGKZ1321IjBVNVoWkVCDjnhZxpPIxoIGL/CcOLOp6KTkH7WfMR2kMz2si
6kfqLQW4WbLOWMlvLngs/QF+qvC6UCzKLZfRJeytsNf+zU5nKave+vTiWoEe6YlyOVW2ElPxlSGq
BE8AbnS+TR5/AqLO8oMkYFv7yG18fPn73IRQ2yYeUM+Jeb2msg9fzbSbYU+ZyLE6ZwFQAagBGoND
VjQlarTCh2oqRTvGGwbjCJtP8sGX/VAFmSgLso104TK5CP4IbV6vBJKb8qNaUDghveO2zNw5WA2E
V93GMC4KYEtOzJUO+JBGT7/j82P4FTIbnlifLlunMZqfVuZOHU1tfCDnbHWgYNAEUOS59MWOPPYO
QDdoNk9v0sqvLCpc3GbLenR7Idu7mwlN+K/Y/AWXya6wQC+muw1f6rcpY7g+GaJAmUIvyzEkb9l8
C7cU6qNVUhQArz8hHGaKLyOLRs6BeBVPXhy903JZxNQWIdOJmMb12cqBvkksL+RjJWKBpEGCdwGZ
bMfoc2GYO6Y5x5/lPtYPEb1LWFn/U5bF2gHDCPCo5sxnBmlnZy1dN+WiAfycc3zh/gfMt6mIW0W8
3LkSUk73M3IcKugKBHlQXdiyHJdOuKbFDEFEnEoRUeqJbCxaL/4oz2Y+4Gh4s7YPNcjzQqtFAsZw
noAmMq8yS9jG9UPm/faQYho3erxrT/LeiZs7dchTwYRiD8BJPJIoem0px8VPrYseatID5h/8vrUA
wtfLFbv/1bpJIbUIsR2kusqIFhnNJbSw3DU+n/4DdXCrW+H4Tp9Ho4LS/SxDsx1SR6KuCL8UmZUu
H8sVQ6u0l5nulNswZ3yCEd8EWqWEUUDA/1zGWbCs8X7V8KK/baxA4d3rQSpxBkgr/iuDJgLSFdpB
F1Qcx1YCTPuSJvsujixrVFTLLvV5y9qFMS1R3YE9kBbhinbTszR2oYzJugZvabjyRJO5kUU9NCiU
odOHePxzgA2E5bBQyOTA7Z+SWd+V7LhrOq38VKaLFg9EETo67OaDfCtsnocWs2USco7JG3Njl7qO
vzYtH6vDVptoAI9KatjTsWyu494Yzl+YdFVuPC8HQ/89DX/2H5FWsPG6BZIexiwjUEsWuw6rgw6c
GR5tqgFUdLhCiciLddVe+Q1LGQA5RTMQ6seVU3t80VGFY2FqjUA7mWQouZIQf9Q9X2GlvCezGmOP
uyzXRDQCLULYRLkAG4tK0WLPvKQ4Gc2e8QGxbBzKHjQjLly/gktdHeO+WjCr8VVxgX7PpuPDUeuK
R4o61XjwYNwTX6umqBEMzHDeEt8CAXQefBVg4aLS38u3bCILUBuMa9JM4RgjZJimCqxunRANMEpk
SOa1kjgvNRVL9fAvTlkZbPY1IIaGIZjpPt2Md1/tOM7METSe8zmpwGZfgP5ncILYOA4pKUat71Uc
XETwFHdCqeXb1dvujox1Uxz++0bGyB82jWQfhVAU2ahXTSlE/Q4CFk1m17kzT5bMkL/u6ZNxJGH6
rMM5zz1SmhuI1/XrPeUkXtLGP4XWqqwX4LPjLtAZheevgqM/HbvaVVu6Z7c430gzzJxpFAm3BzJX
hlvO/LbGSIfFHaJZeqdH+2/QcI8rGnIufRsIOa862nporwpyVmvsWCJei/VGa7U2XjdiMeNr0Czj
cYdvb9GTEYofuoT8x3/XsgcN8mdOR4g8KYu9SlCX7JlsDcbTD0oahah6xXeLOoeuv0kptKh2vood
c1SlcqwU3xndz+aH/VtQ6jZMrBWrNgAGvclMbbCCFaiuaPaO33Z8HspKrZKKhYMCTKqqFgGhx+48
VoM9wCaINSierNCzYODuj4nNs12gNsYnAU5j/vuliueFWaVYseLJAzy/G/ZmS7SZ+F6N3IMkrEzu
tqlPVKy2+f69kVRU3dsl4paaeAYYVGeCrfSCslREfPeA7EbcnoOz5kiuy1kzwQv2stqQwhF/mW4l
bjj426k7qfD0MZgr7D9G9c29077DtnK83t2mDB2fgg4tVPrLfV9u6roaB3Ez8CAtN2gDzwcA3UYP
XvmrrIL7lA7/CcBsUUEA0AURJ87rPQ28cHEDqxvmIo76jKCZDExvo4ReK9wgBgobqbus+wdWUdIv
CsF7O9kuI19iP7Z7wx4/QGbJVLZcwgV3cECbLT6HBKm2ecW5PXpweyypKy6p6l2GFA1ZQMybGTt+
jpLUb4fqh43m00JLY/e04xoNrLZxOIRbTB6TYQ3VATZH4W4JyAOCEqocljG8vFvKhi8I/R/BcMuO
wuacj1obuXl4Ador4pv2HB+gP14NYNlHsQfRvOGSGhcv+Q54jW1C5BYkr67mlitEpVV0xMC5DwFm
1R/NUMeqJ2QjVS+Z6ZifJk/IHZSplcNP3TbyrV/zP3wia+8tlxR0f1jwOYX71/UYHCAtIw9fpYxI
TiJshdIQrvhsNIpqwjJmdg5BXX12P1l1NFZ6hN8uaw05jY/VYC5hEyjk5uMiXoeZw2LnTAhV6MF3
+9X3Hz9jgbueejELb1M/YIRWwk3AcdVXryXCSSbtgRNoow6X+4lc2xm7H9pTy0JCcdRBiwzlOPoa
RG5XBKIya8IVEO5Ock3VNQkZ5ppZFeAVDNifnSM3Vzbnh0UfrMNHGRP4fcDRhDs9QWc+4q2VBwvx
HoGfIn/NQupbX7BFSmaEsB6TgsxaUxL7GJa9A0IkIX9JCW2EYtY+P9A+H9GL8HWNPOI7GJswPXdE
FVM8Jatgxbi1IMB15PiPx+tvQqsgcb6hbbBBLKOJCy1iv2y20tHk5qKnw7Tdv3rKbI9JXn2XAdgt
KHiQ+IvgXnpgmJLDyqgtzV3FZbrVM8Mib72bW+2foZe1MDIi5nEB+xWhMemdW1pwQgG8BqvvVOCD
QVHvDN4pagxlOe4qM/jNGPGEx8tpqFWTzoNBp5H94cg5usvQWddW9xAhGM2nro4M0YoV91hcq8RU
07HZ4ZxTim6ZDr319NdcDIe7nmDfO4v/nDFzzuyfVXS50xhX+avHlEEdGmoUIeTJpFaDBFiaYrAb
/dMm4z8bb9Iukzwi68JF095xqex+ocbdW+XTbs2+ENKFF8JYhnEQV4/KuQcVpuVpOR7zTxyUmL7T
llh0LR6VvkjyZvJ2BWqCupdEI7swqoKaXKd2KpkQeO66vAaD4jWMmyzrKyMPTgF1honux47AkMVX
09x5vO0/izbWKk3Z6okTH4Qnqppca3R/t8YKoc7krfIgW1WmDJfdQ/LjEGyi7bsjBQw4KIW5cKtZ
bE2J2X7aPaIBCR5nr8AMHupWRG8cpbn0unaDZlaYl2v6yxFP8LNXhzI29bQpmzUscfbV2yKWHdnN
eXyvZH2n0q2H1xXlg/jMDXjV4VB2dUiv5ucRQmysJkgIyShmPtyeDTifBrEh/1ZhCoqtEPvt795z
hOUdw/dFGOHOb05ktibDTc3cYrcw4HyefiRQf+q5MxOwtykMR8B0uLARN9nhULKDQfxBKKAIV2LZ
GSmdeb9tqfXztiC3FvGAIkAS0Xos6irrxYbUhDCRq5Lt/KkrYvyTlXWMuGcXEw1eqkKTF58FxUBD
bxtw21CoBZAfKb91gYN2X0LVhk5YUR/U0DYXa5Wqo8eJTOJI1d+6oRXxWsWjqXcG3udCGajQgqj8
da2xTSDDtGbsBZR28BfDMaKLjCEItn1Ltj+Td7NCyxQ+7GbywPYdvMPvePYAMLsbNYDzrE0iZARN
vWyOk8MhAgavTM+TLzSeIHcC/AQ8YsYo+OPtihude47QhCLs2jQWW5LzCq8jhn70TExPB0UidbhE
oGAlZsUNe0ro/zsesJ96efHtCzTekI8Hf+vlDrCWSPvmn0hj52SLC++2VDrg3/Axjb12a7n+pi/4
LxLO4bzhUAZUNTIpOqjMW4BzCGELGcVI1CTo+ghyY2TwqzAGId3RadW8rLKVQpDNUygiomP7Konv
U6rinAjdcih7CAcpeS/tFbyWLuMalrNPzSa6gS+nt1lXzuZIlKHK8ZFe9Kh0WQFzcJ4ypJsF5+d7
qaSSTd33p7duiTs36tmQY+ul8HFy7dyS9MuM5lDrigfTGentIhzAnoJLnIiO015dB6gFkcot1lmQ
G2iVUpM+XbzFO7To1jxfs2ReJve5vdoDNLZlaphZn/LqbTthTVLv9ycDh8zEuX9isDLY5qk+wBLT
TrMHiUlbQ5txL5HY1jUjb6OYKg8Vul+GuI2GNcuKABgvbUm9F9avMuawPe1vbuHPaqW8w8t9gG71
PZNtdPlG8Lx17oz3denqCsVXhMwa9YovgaY7IMs3sQUOeivBvXyp4fF0Kbk96F+Ruu5cYy9jXUbm
5qpDijOkX3yjky8Tj6zUxHSNPGC0GsSCqhmimp6K7nwZkNy6EzXJbUdqtG1L/KPOxQiFBevac24Q
1SquZwu/jOcBSSrj2IP6fv680U+FOtbR7uFzJNPYlQ7U6R7/OuRncj9svt7twBQ8zGEy1sBmT6e7
xlpDfkIq4SEOPaMxOX6tmNuWbhEPxG4+F4L6hDd2IYiPKfoi04+v/KJ6BehApBQv8TzFifuzmg1a
ddYpqstGcRS7tNbMrsybGIE9433fTGlvMjofMREXLKwzQubdZ5kqj3jnWGh5Qfgau0+J8SqIqExZ
akqHYbtayMtQMtSLLVA+DzXQCx9DEoDpgOPzmpg8XvPpn65tR11YefAkf14SL59k2sHxBo73MtXg
3ZvsvUIJb90m8Yf69ZF30dugE5QwW9mAgpAftQ01OwTnQE6878RRhlBUmjWYUt30yyRetsaNrOTq
Fk/BeED/dxXM3QXC+6twXSD/usiQw+xNVd/7p9PThWTuxj3/5RwyBT7mFbScdtMreph4kEfqOxjc
ikjel9pWOPUsLTN9CMa0k4ADsM7Gtsy6hyD+YVnGaYp9xKV5zetL0NH6H8Cu+peNY7y6ap0WkVpY
8ty4arAUowOxvdxUKRYKGBXZzX73gYoOfifjuJHvQYQdmdMIdb5MiunwFbryBYItvbl3oU1DcHgo
LmhBBKrf2NTN7A7jbOkxqoCT0S8Klk1TrKz/+/txHkQGeJgimhepd8VX+4phNsZSjBVsR1WG+ztW
mKtN8Jq+FiJjQn5czbl6DYORUPt34LNIZ7LMlyjwZwOCFOr3uKDpHte0sqryBZ/bCnEQ8iODypUG
GWoZR9hNFIjCZ7J2S45yXCh7OJW2gozDlsq7UsIrDu0umfNTlQxEDpgHqcMnZBMURzvapAfjKJg7
sMYNYVYYNgsPxa5NP+84gvTuLfdT47WysVn/8O8PrIqtzLdqisHQRlUF5QPaAlHnRTSUUJ/2d7EJ
s1IimuXQK/SyKSgDytZefMCF7HdJjceDPvneXq4EpHcKp4xo6p+JV2YzJdtV3IMARew7hhpx9B5j
pwQO1NT1f+HGtKyMKZwEVfJilCA+R870bRNa4qR/jlkmSwdr8F6Rzoy3GY2zOY3rS1mXJ1t/bHIb
YKDZfysUDBYGxjypbGWL5FN2H4VMnD5t9nLenEKkobgCJwlG6QtZ7MMbW5KwUc7lbh3+YgCWNA7Y
TPasqXmbR/f70EjVGqWyIsDRiQLOD3SAymjw3dhqM03nr2/seST205ibk/CISJhb50Vexbk3uPPU
aUhLsBtEIl7zXK7oQxOng2f3EtAv/3paPO0e0zi7HuNn/SOmvg7XHZV7Ebe3G+0nnckX8BUlObox
pgIlZAxjtd3mrygO5HbRHX4TnICghNkGzhKBfRZIY+DBAHV3Ao7iJAhYA6wTiFcFsJcaxYOjKsZX
QbRv7c1+JQSrIMF4OV8HjBbzPoOljGmUGdGdDO2Z1+z1V/c8d3TTAmsQI8cN0C8Ae8kzQhNcoHjb
TFPR/DzqAhUgJLJ0udkEMxyUcaBL62aVvGQ39/ULgfLvbDn5uYeycGfWK6uvrOWtWMlau7L9MpFq
Ysu86hiM1f3/NNyppw22CiL/G1YGFhw+p4EZnVG88TQ8Kmeg6bzMrK8BLFoDDMShkepTOaLnIGit
bo9f2HeWo29H9xOU0yxDJ6/7oSK7qJlLpvuQWLpyA0cthRXDK4BS2aofD92Tnpzix1N48KMLZuKi
RHYrSvgQEGBO6NIPLAnRgIkDh1lsWg2jOXD5gqEiUPZ/p1WPdViE6X7+oogWYcJQC4S4yRtUNTPO
hgV5pjr9b9m8ad/odsNWvXyt4hBOyjEh6oxi7aoOq4O4tlvVMb2X8JBOVitTI6lvve065k5Sv4G5
4e2l773B+EXqJdZwitn52aYe8vqN2IOJQOUY0j1dW7HcophYeLKqT7OsBXlDdgNR0ycyKAANR4p3
xT3PwnJUa3BNaO/PKX/uOnEd6ntDBTkIZ5/AFdaHsuWagXoOxNeUsPqoN6PUnjv9lQSsLr9QwYOm
KtgX4WXevyoZ8TMufbGT9rKF1NOJUCOgUW1wZC7UxQ0KYEWnD/L0Ns5baqx05stEW0lH5o/xXWD5
7a2qwQR7Mm66QBKQSSHSwFbg6FWRUC2K9Ahytsbz50t1qcK408xn+E6sSJ91nnmpcB7XcLyqNVSt
qAlym2hkqB4XzRIL1OVqly1x+4+ckZNu2Oa5m13zax7Wwz4VjE21fFGy7Vin5vBsRxVvxSGA9D/W
UUs57xFZlbRbwA3vHcEovnTMjFEFQGAAisVNzexmZEU4qH/iWsLoupnJFlt22MUX0ouz2YsKGy57
Zb1Jl2bO3lv8IaToWXoKLNxHUUy8Uaf6nOU3D5Fz9MDtPq588NIWuJlT06W1xj7dciGX6J/T6bx5
uc05piQvHY08kFDbyHCamRP6wM4T5eP1G8dvYDMTkSm7IAyEXIF0Lu6KziDpcWq0fdbiX7TDCLxA
p+2P3JvH2DGTxE5Az0VCPa9pkt0vxpYvurn8oKgotyuAOSqIfvilfB6sz7B4hcodhz2mYd9IrWRE
yPH35z4YpRN4FtVF5RUwJZFJu7qy7+UjyU3fo6ZRcnJ2ozRYVl1aWoJLvV+LWH5o2z5M9DAUwBSB
ifljV97akZ+xIDx4O9n6LqK8OGexH5I8tOIbiDDl2WGWY7xA3z+yIQgIPGdovScvpg9OZsj/9HAY
nwgJPbcRQMize+jLtnjqX0ThfESOyvK93nzzXU3BcoJBVgNtzhbyR4gsOfNVU/hOe0lQFZ/4U38m
tOmcFcSfwi9nRpnV8o7TnfHqO1w7AbrSeKKnQGeZWn5Kj+QU1PWHAv8gYunMN7xW53b91416OaEV
NGPF7wIgj/e4kKKblvS3qR7I/s9LauIJi1rtgAzfDgZVndGYpTdfIhKHUYTDhr46lg5kdguEzigK
Nq1HnpY/pUSfTP+TqrzSgTiH7DdXhnAuF5DCqBE0O3LUMz8dIYHZKB71iPBr+B1mVFf+jMDC0Grp
I+PHn3FuXmkL57oNLjnlnCRhZPCxbA6D8gLuTxYLTUpjm/zNzvUQa7kxjQ/zWjoyR2Pqca/cJCm1
JkCNQ83jZwyd/JuniQdpwbT1JMgjREKUoTkDbrjzYzT1mYYGQr1nNBbVgUaS+3y1UzooOJzWY+9U
yudFV5bU1eDhueM+qirtsJz8TEEsYR8V3Gmxlmnv5XfV/4wgqVsldhrL4AJQfxJmu298VP4tdyT/
rzM8rGeCK7bKQTOwlV4sArIHmYwSQZ7Gq+oqOKoSeYScImbhwQjfEnAXhMNCRBLpxrqz28WMUMRc
Odyui7tmTBCF6UsTc2jOjyok/jEDUKy39kpKT7mvgQHpecArQoQ5au5S/MgOJ20Po9pZUKmn0448
NKJCrq/cASHeBitKwoZISwJfQyIKFgNf7aQN+KHzffMIHAPaCMksKJxa9ddB/BM0sH3J5kym+CK/
wl2g0wud+0p0gLMt5oEDUbNFAc4FRfQL17X8pliIWauvo4RfjmiTUS+glB6GEwEkbuxG5KAAIf5J
X8ly6ykBu7lMeb4aArd5Da/cT7mmjAru4vdNa+k3GW0zDHWWKJLGmg0YNYtFhOAVkWooI/kqleHM
k2ybmmJoD5MFK2cfLZ7zctvJvgr7SxeaDcE383YfpXDEyq49sS1WQb0J2aMk5wz7mpe9rAlwOZv6
MCDahsTJw4DgJ7dAFvdVJz5wWXvQZ/KW4xu7zKtsLaldhKOmG+YXrwc3uc+834R5QPLiHVcS7Yzr
tDXb0tQtRVacOty5Oi+zWccUB4aQcYt/xYIhLMJnmaIFFCECEDZPyQcvGz5tS+zJIfq3wUL3bsic
Zz9KeGd951RhD8brKfawK6IcVnCHMGraFpgWvQs2B/N66W0hLMSA43+qT13pXOiPwVj3NxkrHbNE
n9jNDf8jqp+V2SnTj+dahuhJsLvAWqTKPLElzgLlkdmYiAp21/uI8DUEWXWVDmQ1noS06ttTUy2W
uPNZHDG2RxCP8REwrWX51GUuQs61ZDmQK/4O7pBt89M67IvfYcqqDfd8iOdC/FaF5FAVWwgHnJ7A
P/wp/5dpVomFIEjwMvbUTO/ch6wYQuyKotEEpKOo0nPmhr7XJhr5rTKUy5plgMjLOZCZRbI9GbDF
uPPMLTz2yStW9cpurJCBXFQMZUT9MP8tnkhr7jZ5bfUOs2MuqNCSXrmhE5wBn2XlL9aoXU4pBWjk
fYZJz9LTnwdr7k6pyL0oMIkiluYkn43jGHePDdE6GeirnqkV03fc61HBBZnBcOOtM5vd1Qm1GzWv
oYzBWfr8KXSEO0vXj4v03rI3pg6uNhAM36rSZF5BBmN3cwg/W4gzFZe6PFQfRuH/qDZiZUIwYpNJ
wA0tLUYTcNqLkjQGNFNRPLmpmEnQ6Ug3qkQaTxuVoVOIymJUfOzIa5zY0vNQ1OkI8xrDYwcKeFAZ
d8/9sJeC5r7gW/urnkIL5awC9HuVoLgwcx6Hm3GYWnlzJMXdETwIXetaOi+AupQHeezqrQpDT+YL
nde5mpbD5HFxvDrxUyvJNzlMh2T88/iXzGBY/5P+c6boMfVSwAu1jMqzfT2vvfCiJCSA9Fn2Ph15
nUsxOAAc8MWOVt9w8JVRbUIct6MHXBIGOqZQwJSkbd+ys4pQWZvxc07/HhKVvDqTbqsUceIJrHQc
mueE9vYR/ZAiCcFSGqtl+c7JTuXVd76+Rx76kPEI7QHPke/NLxIJEpyVtYLpXjeH6KzSOYsoWYwR
XVZfV1nNhwFCQ4b2FxMYKIDq5+b9LrPdCT/Wz9eMB4tC01FJ0eyJabJoGQlJtnOLk1I9VRy0BmRx
gUElPqgb18+cqnTSwjNtG17lDL/PHgxa/G0sS/eYJh2q2/CYuRBoe+lNnkL+/yfCRmaHi4NTEnUq
SuzvX0vsQMmI1HPOnOlOMJUOsRIxfpjYzJCriAfRTfgEu+k2Ez/vSXCsVK9iqp7Z93MZ1rDwGBhE
Pz5E8Q9xwXu2H9CTFGl2on3zz94jgoecXCNOVVrr9NcO8Jpt32sHgYpLK1cmDTfTikv1oV79LhCp
f6lYYr2P8RZ+MwoV+WZELBHBmggH3dpM1diohf/BIDwFhh4F+RKVCBj8Eo2LIF4HRwCtYQ/yOgf7
zfjSDcYW69Y87xNExKWD2lCgfMNdaRzYZXQ8aA86Z2TxYOUiDtZLEXyLrSBaqf0OQyl5bBySjyDs
g9gQM2+Gx3ALpGLN5gf2RTUJ9tXeq8rws7/mSrh4zyfRU6dpC3DLz8fNhwerZlLtKTppw3JJbKxF
e7hiFsM5K8JxsVsKZD29TbShU9RhjyncgkOUkYS824vXxYA4loHVedgeBLrp79PLScpqgtxSKN35
fvTfswQp0AT5TaN4fQmU9vBls8z2TnKBzPV+yQHuXXB2UFYhz36oefLYGhGHMKwRTD7hu7wKeW4x
UNf5mk5I4xn8O2tYP1IV0UlzKNKFO/my0QdFw/h7QNUhwSJaQFbXUpE7pLIOx9SP/ctCrROFmyFk
U5x1nVGjmJXqQCagNWResO+uwk7PoQR7X1IuW7BnEM1muYU1aYi7+uozZ04MxIkKqjCFZIetAArv
xHo66AuYaKztxpT9jQ6Ebxkyi1yuYPsWhKJb23ELQVhzZqvOYIJQfl4FTvitIBlaGYjL0o07pR20
Xyfn/RIqv8KFt2DoiYq8WnDNt85Ozd8v/9QbOPnAGfRZcri59EN31G+OSJryjpO3HkZjoGBSgCwD
1Mc+b/xmllRrrglee8nx4ljTGYa2XKpucOi2zkkd5Wj1JlHepalBJSKZ16SRydDK1bAmu+kSPjP3
k+lrqKcpzwxs2qIpF7hMvxHT9t3vbIu64oHkv7avtjuuxPggrbWbaYb5YHED2iJ2EpRsfK+ytM/u
k2ANr6dVVvUhEHMdiXfMFiEKx041xcf/5Ik6A83LheR21QjAJQERauhTqy6xtfMKdlgAcl2sDJip
M6FHU2W+nlZ2RK3QfbfTZTr0kXGm6x+Gk5SIQf4HjYpgMbtucIiVeVY3jfHpigt+EClxL87ul4nA
Bzs5NCT6aIMqzWLj6uSkoXyK5E+DLi8ayUT9pnMB/Pu8NpyfZ2adc1KsreTUuD9OWjBnvU6HARfL
KTfhp5D5O+ml58TvirvxRFanY6minIILfy620N3DwgWgz6Gu4wRiRjHQUcFZIqnBl2+FySr/13MT
yj+w9+BVax/9CdCHB7LqxV6n6V7KgAwh2U+vOZbjlnUAhLRs/neJ6Dmq9z/uZp37hlVdQW6SIYme
nyDRnuGJUQGuT8IKUJFfNrL/l6yGKAujDKucn3QIYtefh8i3ftC6BH3YT3ZgntRc2BvOWRgWRrfL
1HuPwOneK4cvt7+Sm0lqLKO/D28/ib0bXY8jWRHT/3Rrwphh7vbt7bFBAdqWRZt1bzYaGquobAzD
AEEZlr17lOxVtCiURaWNDO7dFmHao629ifkbIH73N+s9JxfXzsMTw7xiHWsZIR+qMDeJ1yUAFNrS
mBmbK6jWvTA4Gxe0KVVtPr61UK5Zgf5B6oNegSxVYzjruF7YJRBqVBhTKVWL4YPYVnIOSfqkBFYa
oTUKn9Gom5L42ytxSrlCvAKMOOx+hupBz26MPliyftXk+bXWG8dg7NpH5SdyIRDrgmq9i4lF9KhJ
LPBelU/VOk4IJBBHae/X+Sqf7ZCVeK8//u5/+RJroRGjuMbCBKqSbjRbCn6pW3SF5jtnG/EJo1QB
BnbVmDMnp/UKqnxTrHQPUDgnmV5IfZUM7U8aYLfbqN8V6gjIIyzOpT2HaOyb8v9qNEqChXdu+ZR6
J3x25AKHPcEDwK0j9RU3M+SAA9Z/HNJsuqODAfFrZKlmH7MDyQrwquc0oN4+KWFtzzzIzHMiScHY
77rhzJ+TnEL0sZ/yqleGRdlafiijifDLnZp34Dq/iMQ2RfGXjS75SOOF0SA5zfLRtxL68d32bJ+D
KE2XpYNg9+85uRFRpgzg2VvbqA0LY7e/I4BL74KWYTTp+cuKmP0auR28N5BDaYmsW7RUjw+e8o8C
ZHTUU4i6MMHJRttP+AzZdN/Gat02cmEHVbMwJwC2YqZJYKK5H0lbAAFY0RzNYqq4yk5IpYikiHrt
3vLJ3//5UOpevXvJGw5EmASL+zAyyc3RTVBwkQi+ZcgNJX7paAdFRJRfupO1lkHdSGCexArnUKkb
kcip7y7U8nRMUt2CIutcu7yGLlOuKpkLHGwd9W10Ef6jAqjihGHTCi70JAbum9uWgwv7wrYdn1Sf
B+vLD+QsCmeOagdQN+s8xTU62DDLhz0NPjei7gj1PQZQeYDff2ZCnQOWPisqmqFNZBmoJz5qOPht
l9885igtllvrLnn8H/32R3NdEQHb8wZtOcMZO+PNPPZ9fyVEdD11gT4Pqr9LByliBsGLJAB+BNFM
1Ncj3VbutrTfciV8KlIelb7vodGAwFlu/s6lmZWM3sItzJK/HgJWR5qjQm+/uFwmd0uyg5lsACAY
u0baYCG8+Z87o66HaItOPydMiUw3ndaOGXaaMus1CsB1INrKyNGTHLWb7b7d5Gv6O/kPZKDMelrO
e8Re5cr906c1qW2HKv35dif8+aFA4eZrv1lTYXCe21WchQtyZ6tec8dcBi34WcX3RWsY7ilXJcfW
Izs9f+Y4l1VlhOEMf0ls4lKX3bW3iIK1coCZnhS6WS5pQsrUVUrAi9UGG1zVyZrzT6+euPBteK+Q
yBVLiA/PQrrIP0a5pKTbLkWInr2rcZIR9XX508DtsDWmXWCP/M98bOPscWSHLnp66eMQpdr+hiJh
EmYNuC25j9XEg5JW3+eyiz4qMbd64aO14xLfk+dcPPjaCSFIaONx6+B8t54JNlodFzslO3mUPGEC
VgtEcewQPim/3dP/QmxxWcbHlVv2j68KprmGspcauHl0zYvFwLwS6J8FpbbFzPkmZy3/8+xE+LBZ
tDRV0fT8mc5HTaAdMlqZWTBBSVRuisR7oRbh5kkgIUkfZTO59FPhuyjQw1PLXG8zLxaslmlHVsfc
Ls58PAH5OfKiYW7Ndwy03roQzpFXBGtBtMkCANTTqYVM+neEZZVUT+x6bAb21h+izaWQeLL0rKel
NRi/WRImehICNMyDjTmx6TRxQ2YqtGM5q5JZQAj+4uQjp4yK7VUZ8xYUOnhdvH0L1eEVggDNy2jO
7NLg8R+h18dW1F3VGbCIImSpW79P1J6QXf8BM1E5Qw2pMEJXGaEQzlXs+HSDiHGpgfawr8iwNFv/
c/slh6evx7reFe71ahgiiTmil9xa/Q+MyZG2m+nbdvDy15BclL+zLvBRh8kMAwU9K7a73XO1Z+WG
ZvOuVl8BJlIMUX+y9yEsA9akvKLUomy1k15eNI++cvJkg3BqUpxIRGm9c42+tDbznwFRaf+367S/
/UajRii2W/YJYUAtbxtMnMhZabEXTgVTGAVaC6yY0uU/WLN8fXtZRLKXnynmgTm31lFVJpcxpoS/
2u8Q/wLAqXGKRW9ylI5+O/9OnQfzviuu0hrcRFC9uHVyTw6m/qvXjD+qIm8HEDNmsiCYxtzMOvmJ
P+KbHtzx/yxyboJ1ch3mD9BUNxAmFAtGbO0n47c11jBBXOgWqRF7+P3kc1rwyQ8lZEazMziaezSd
a38pUGE9SqcLWz6YGu7ks4Etvb/OJs9Mi66A89r0HLfUmH8+uEgtXM2KQIisJ1bPnUi2loeB8bwD
4tTvXrtXzIjrFsLxjea7RR5/7tpwAkCeFW9CIZc/8n7l1kC/MWAANFi2w4kibwL4u0DViN6zSV8U
sesczpy/YsLRosTavqTA1FIx57LNOSiBRXqr6MF7zDANfJTXYUEvb/58DwL5C63n/W4tyJAgdbdS
sX/8KZhRIld/eBm69Y/jZDAQ55hqb7ueEVJyLpyg8Gv8OmPqoJGTMJP5hBoFWdFrTjFkbGQQrLg/
O2mI31igZLLszht3kGNumuBFhq8V3fvyFrg3ggLEtzRHC2BsPPwbEI0LxMxWRd6zB7c6Y7LiiB4w
aSyW6DY38lDrr+DsNK6PZgdt1iDGiC2C5XvpXvJPSWYMAsY6PxCecsZ+rftCLb584Eijkf1Erpxf
OIKWkphIuKvzSWam/NuqeyBvGlGW1xy4i568N8xGAeqZgnzB1DDhcnkajGxi4l0dGhO8IOcsfccX
sZIyykryRrvM2MwagB6qWlSvPbX0O4/XrV8HQOG0RE0kvgiWitmpXI13hDyVSe8PR+FG+vws2Rbh
UZI+WQiLsc70PgDnrzs1ZQqLSgRZcfH0+wtwYCpTfObY/MGbihhlMGRQfGoYUrZ3Sv+LIuJ4j2Pj
L1UsfsFM/z9eJN/FiiUaLx5S9Zi6VKObTX3NK4uD7AaPs+fPopcbywHYb6BLclUXa+4LGqgG1GPf
wW91/+4UqM0PcNWneYsIP0S0/wM8SWvhRuFPySxpHnZafxOSBzoUx6PLVKLRzz0PTg0C0gFcUCpl
mVCArFd9iTLodVhF7KlerwbA7sT0q+V/dQsNgWab1geeTQuw+HMG6LFMiiif8g2fIz33riAsmbT3
5gx+FNy9ui1JR/eS6MfB4P/tBZXn7h2BiECHnAJN1tr1SRcfsIChXQ466NCkW4on3XUGsTvUHpuu
7SGq/p77J9cpBlqQE+FHdSyGG1l7RJJ+45SWkOEYQRfqkwzy8wDzdrPklKCLBX0+EJs1mMZdP/WF
h4bbL4eFRrE2cvvEUi+hEzPEV1vv2QZMhGk1ScNXx6dm9p165l3AapA+Bhr/0E5HhVR9wiAEEYEs
zNha35VwbSzia9IOFMZtQcdQKevNlnRGom53PY06ucR7mCvcCvU1e1Ao5k2qb/ulIvEiaTE9M+cu
VHcKuX65BjY8Xriz6KOkapAp4d3EkJJUcVuWfKrXbNTkpP/8WyRVybBtgQe8mvvCf0tcxPKT6/79
LKEKeW5BoQPtkWTsplr6a60k8hUJUkKPKPX3MEt8RB0q6o4PAlqHVL1Asofc8gXmwOVSXHLZoVDK
WLdm8p+gUcfEg/Y+tj4jqeeJA0ibkl91nFeReq8dQNZIZTmB/7FX9pHPcyQPALhF2e1iGWf25iBq
SQ9LrDGTd6GBI8RP7S96svRFN4w0cELFbDAmfIAlntaO1BD8l4GX5d0f+UeY+KYCsNnvXKSTndIH
yakBvx/PHlCiSocZCmaUSn9F5ChPj3H5gErJoLPuKtdL3BS22D+0Q8Six8N15YFlCW0Ak0JH7rNZ
NETtgTZ4g1ThHtJCN5zy2pDzVsDlR00oCr7Jl2jUaHz8SBh7gcxIlUQu5bfXd3blsM9QTLDZRmep
WjRqSETUpl2xN2+S8oqjcthQWTf5tD6yYcmVQGzg6NDI1jq2KAtB56lAkqaNPUKDMV+DjNvNeyA9
vg+ihZNK4badR37h3kr2Uku1S1t9vtH7q8Nh4fo8gm7g57LQHBua+sf82/dLMQKwsp26wWCNsT+A
PtNY41+53jR8KZq7NSMAmVlX80QLxm9AoML2GVPFS5F1G7qhlXriScVAAdNXaCpwBqdyFymCYY5R
6exTopVgwOpCBszvWt3V9N1zp8ZfjrZquvtS8mYpbUFNNwJ3oLXe2qUUxTNhK6zjNud6nRL6345G
VquhN8gSppnx1hwAgC1CfWydhA/tgJvPKlvPIpmvR2EdUCO4GgTCyfalIuuztfM8SFx94YeoUikY
RiEj8S2DxjPXoU551SQ6b4nRKHYjuisDN9CqX8uPT/6Esw5cHlUDilwHRAEpsJ53c/Zpy07uVWfi
SHUM9V3cnC2AUESSLf0trV0p6HKzAHeDoKUgnPwtLcoLe4mRXcYY09ffXMZ1lzPn4W2jbAlKAvts
Vueee3vJWBqQVskylqLey8WIQCQObMmh5DWwypVO9Rzy9I0aocHp1KnULmXR4EZ+YRAz79VPK9Iz
D/7/xrz6guVEbMkmcuXuXbF2a3zL2HcqNfJaFSYbpl8lqlK3pSFWGA0MQ8/3ptrirx8dtFNO5ViP
cvCqPzyJzXq5/khGT9tZ1mJ38Sglo4/b0dv9cS1RzNfw6FR773N0UM/SEB1l/UUaEVduxF7L6l0Q
vPKTz5+jTtC/ihbHpGz3aXHXSAsVImp4tYvVRU3omrh9Gt595jkor4HRXa8uz0mIXvlF/PRJJR+A
hfUexmN+WiDWe1j7Xjuv0VsZlG8NH9CPgtcQCdd2f6w1sCaCP0SLhriDAoCXasUiLV2i1gVuHai6
xKvTi+y+b8RHwqQgRDvEMLAK/KOQJQLOEB2TljDmjxkcPtEtMgsXDCvksMRByjOFIvnuIzSAnbW9
EJ7YfKRTakFHlAGB9vsOJAI50vgPIA+KPphU6EM+lj5IbCXqz7NRz3J1Km9gWAGnHDJlpuQKJ0eG
+jfJan8BY34MtNNTRIWUvnRTSfTnQ9u6NIerMRyfAgx1GuwTTnpbarG+VS3GQ4PyrAI4ipEeDXSX
O+tRVlrMT3gFejqkAByfETQ3CrsiR/IO5m8Xa2+0D4zxBnDbwnE+NSUA5EFX80zi3B3t074rtv4h
X9xzGlpVWin4msxrYByTUh+pH8x6w6WQEBYxcxa4acgnA3PqTeANdahKnQiwp6g3zxxA+gj2flhr
txDH3eM6Kfh1Z3Izv8z4onc4Lv5DJ+xM0xfAGvn1awdDqGhhuDoGkZIvzM4/7Wr3wQmJIb4xhda2
YM5zbgWdHAJ5YB8XctJvaeiTKa2BznieyLVmZTUSbN0oKjcTQj7oyGxLeyU9wmhZfqmDoHfvdFaF
emLGTZECGFH1HCJlUL8jQQHMgHNsMkyx+ySlSGsP4D74Ebw7FEPyxWGfX1dqoMb20Nx+hDvcnjcQ
qFkySWOhFny0fHOR1T0CJPH+swfGlSjBD0U3R8f7nbbAmuRy+2rxlz4PKn0vSpJ7uv1k48vGCbcu
DLcX7He6JKJajry0+doLv86QUs56cm/q3/JfgJF/a/AJZF9/wjx1yXYwiSjMonT3Z/JBF/KVDOb6
/R7hziFhKX9Y/1bD/eo/9yZgqz5HejYMDuQtVX2AUyk43tGfF+aM04hRekz5Uedb61ol4M0PFNp+
9nkC51IRkUXc5Qt+mKz2cJZ6DBXxFHYvLyNnf2JAAShkWWCnx98nUQUUk8Q7qXUfXTqWVHDStokw
WfvtVZ2ccoPwT1+cd87iuYKZZ2m93PKRrn4pVnyJcMCCecFQiuh0JN552uTnWkGDIwtO5+EIN1mq
hC9xUA+oF/0zawyK4x7oto4WDTJqJwIvlmD69oL66vz3DjNAJCFBcB9nb4TAN3srbteMi3ygNPtI
1rfVnuIXcq5aw5ru/UvNyLjUjkD25Hf2j1SPT+UOKD+bAU41vRaRjFrpduUzLDdAH4MMq/xY0tOR
1mH3NFZ9IuH1TsJIq1OvzNn14CODxxnUApcFE04opApvZo7CNSobQgZm/IEcvhVP/lpvZWXg/jLo
NW8WVMtB5N+Kli29gZxE8mFomNumgqmQA2tbgZOOdR+PGbRV0KLAD84//V2zpoTgGCfCx+sgOC+/
clhc0leVHVyJ0NKpD6tNGBWt7+pBFZagS6T/4YmAoUMNQjXO0QLUVMVxCWy2hsQ/uk3ZCDkzOqAm
DzWuZa+TOQhhGDK8lLKug/19RtxPzjDYEZ++GQRCDkiv8nqSQCZTAHvP6KS01SauGfpwAQFDHkkq
/ni5IQ7I/jBOE1tY953x/m9SKlmaRtP97Ts8YCgnlZhMACMt2do3DV7tq5ozV2/3A10EuDXk38xR
2RNi8j36yO2JXO8CrVeQNV05/LqGHBu1ssLA98ZLc0mZMRJMhsle5CwxC4Gatp9XPAWszJvVYN/f
fmaZNF9Qks2YCqWEEp2OcMj88Utew5ygG2wNGlM6QHpaILdAMuQ4TjLLs4vPiHKgn4qn1jc7w6HJ
cUhccexcvwvmgerWVvrQqaQY3S3XH7v7VB/xGWhJKsNXXeX3R8RZtr+eMFVZivtlptAXz01iDysN
fRQliJgUvnRgI9fYonhhCct+EzZf7OgbrygiQMD8OPjVpuT/6D6rYRktY1o0ZkvPc9jTjJFTy0l/
NiWEhlhdMCMDxRRgWHzDq+B5QS5QDAzuhICyoaNZTiyR6hPzRm28yN3b6tp6tv8QJY1e3y3KI3aQ
pVnb0UOCPlv+QtoshzchQrx/aPbwdAyG8+lOWD9LJZBrfOGzwn8r9PGumMu1LCm9ESXrqqC//iCm
cofeZIL+AujUQsLuccAHuW6NLj2H1/cB9woeGR1jI5o4TaK9ffZUSQE60tSf+J9BCLyNcHJvi/pS
jqqsN8oaUv/xc0IB3xxVNipBX+D7PcnoYNON3yIV56k+tBu1jG2CPc656zppyQk9u4YiClZq5pOl
3V4rgl3uoRv2EG9FOaUbw/JJH4Ej+4VMdhu5mOnoiGBcEWqVbDIDayKOoYPlqm6j5RwXcgFG5nY5
7RkEVMDoo2mKcOoVFvj511gJJ3OkdtBZlJPWsbW4l8eQck9+prJd6EoleJ45R7SBYoEJDNNIVqhX
rVOYbBugPyECJd/LiCkXjJSlv4/MlYJPuNYoQYgxpC8ZW2Iz3xopwpPhfV/ZmTT8Kh7sAPPiOPzB
XliLc2DO/0NOEyM+4MHzkVh4Uj3WwYzUDSN2TTvo8YgnV/SaA99kQOpkyKvTOUSjUk/55L3OqpCx
J61/pw40GTyomLj7rO19h8dQIa8DV/gr7wA/+dVk1Fq8SsPr89JU4z67OqGAXqxzyffJrSYGxjIw
5ovbRs44Gms0SGbheqyGmV+JmDu8KpFxIRiqlgz5a6hUp4W5WWBkvj4F1adSHhI/PtEIsyM9eZFM
Zf4S3/Yc+36ueJP/wempjft9S2zuLH/wSDZzciw0W5nNFlN4waHGOwTBh0ET273EXjP5FuZgmIrh
04DuPndulCnEOWPz0fh6j2oNKpJ+/FHB25rAEsp3KwDXR0SAWaxe7I4PX7WCUuS5s97XtwVgPPkb
wGumYwaob2kV7I91QQ1fwW7D1AE11cXRvyUIvDNyGhWqw0++pi/v43COqRPTg6M4ID7FL3JCGuTc
HGp/h8lcbUrzHWDDj8JcWq6A0e98DMSI32pB9XybHzCEPWiuKQFK2LdAkOAwk0eW9GAaUVgGKQyS
E0l/XJRRMLSSKZTAG3Vjzb1ZQzuJAgfgqYJo9J8vzzSvdcIAMeb7lJParWWqe7JaII4/B9wT+JV4
6QfHl8MRWPOMt8iva96ik/NJc9Mj/MN9/qEEym6V9QafILcimxoRBAsl6QM7rSvjXq53fUuz6KDv
EtA3yNQGIVQEr5fezLFxuP8ezrKxwvBpxIjfIjtFSXZ5N/HwBfTjy+cVXyRQz51ZEFY94AZOjazf
y4Yi4Ob9FSQMxY0vf6YvFL79hOa4BNSFuh3ic7x7HWSPU04cGVgLsNn9GqF4/c6n2MI163lNs+/G
c8ySzmZkNlr/O0FQLmgHPGpyCm1+FRTCyB6cVW/GaJb+Cb83L8cL076OZ7DOLoZhg8GnR+9YJN0C
AHtjSqsVJmj2GLmBrA0wFnlS6L8+ye7a+v5+Fh39A9ZtDitezAjl7accbBccwW4rn0wLErv3PJoh
ASU2pAEJgSljce+jPVhFEKQ3tBzo9qGUeAHy2FkveDRiSk24QttL1/ZfhaBABLNXZMqre6DHaDlG
RLG/CwF3pEsIcKwLzVdkV6xYlUFosVDNb96xl67qkriuVz26EmXDH3rvfSi8VIgXDqnPFO83UcnN
i1jukrYJJkKKy2VImx+PsZ8khPcbBxUaDG59D7rDtI/ZcEZTgBMD3lH3JjXJimLN4RKEbyjF1G4a
SRZoxCZkdiYMG2ctln3Y1bSZgtIFBfyWvCsil+/UtcDTBKTQfEx430qDrbiMYpOS6aAnfS84mCtl
iL8OEU0h0kN/gvtczzwAi7c96sAQSpBWghMTeL6B51dnaz/Los6Jk9UZSaDxy/B/T7NUN8uRth1N
sDdJmrkX1l6uuOLcrNy7SLlf9O4eJFa3167zn8WtXl06gzyBkmkq7nHXdFbtQ58xBKLAs5DkZAqu
yPAI0vIJxkXTXr1J8gW/R6XWFnKUwebLd61+KvTLj70O06IKXPpvxLQyGGJTUq7ljO4ykW7RsY3+
jediPn+f3RNF/ZM+R3FVEhlCDKj8dZm9OZYsiNFGoC90CYweT9FwZw9ZK0Btdy/+CHQFlWDJwRxd
oulY8ewtIgvCxL+p1Cqb0mOoN5c6rG8Jxjek8XjCdsPpKd//8zD6sbe8X5kuacVTk7phe84Arotk
F+H7ivav2sHronfa0l4jGjr8ej8XMC69GwUpXoxABP+cHzl6T2pcZuyGNQQd2IGxldmAlciyvXPB
MLnuP+9zzeeAvWC+SpYiH6ExSnrbSDUX8bv5C9vEHnonHwpzW7xYlWL6bxm6ZkPGhb5BIQ5zBgUN
sWNFrEnRDnJuTeKKAN1v9vuwh7FW/9d8bE4Ywq9bkODXn3NysRLhfI3ewq66IHrLUWqslHm8B1zQ
0v2TFDGMeNmHGxLyFgFpEsmfLbyscBPZmxopi3hiEPS5LgbP1CpdknVAQmlnqhJp2JRYZgL4ht3y
6k0S40odlKvtQZ6KFsqU3NC4+KgX0UHjyJ+C2q8zzB3+NTVFdbn2ciVga1Ik26HqWcttDXkt9qrY
CABS863cY/qCghMoREKTyiKmp5PGXHMn5eZvOyAf3Pi/EKARSai0rfjkDXk8fWKCXfjD4Ows7mjs
0zUJyJeb2jx9rD5s9S493E5ll/nJr6X0+t3WL6OfcqVa6yBMnn+OFsUbSBL0HYgkhD3/SxFuNYXv
QezvZQyeEPsICn81PztndW1LNZfDlRhJisXncyKz9I8MWKHfF02oPJYcPTsuDMkAxZ29OJTVrtXw
mnIeb6cyj41u+EQpOc63E4iVzfqnGJOS7jqhQ5tCP3FKNejZ5cOYjJ0qivXCbtdRyjya7FHXFbaB
1szoHHSXwkZYEB/Ft2msmPu+EGxKssBjrUaYX3xTH6hBqFZMr8k2LKgtZxpxqKThC9/F6QioTR+0
L7vk9XHzRYCxjPbt8E64FM61cYRiGyNKRrE3Zgkj8pgxgnXT6SRK9HXqQVWrZ3sijbfgHy+rzvel
HfejnMg2xzSWnsS+vM3bD37Fvzp6QmnN8PbL+dmF94Y0MQ31CLl2jWRgQswo1BLxmCYubHCsKa6I
V4gZhMcFBGxxJoe0jMYQAaQqNmk1Z5wy3ejDGu1EDcyz/AavoVFHGPDar9JzUXLXrNUGIb0zZ3vy
3wFYyyDmyec30k0nN3eY0BAh/3Fm5Of6Qo5f5AiY2Ay5zrGOSFsZKuiNz4z0X/YSFx2FsZh16QDm
VU3igc+ZDWS2VmI+StvmzZe93g3PZU4+5M8uPZfeDnXsmY9ofQHaDx4j4unoWA7n45qAFOKes/xk
NHVLAGiaNGWaArkKAu6AcEUu18jyHM/0TGixqWi77T6ZwsnmmVa+ycHHh+LceZK4lzhV6mDofhMt
mRfrJ9x8vtpiCzOEh3T555mwhgefGZwSEfZIQ3NK79fiVRaPb78d8HuHgPMpbweVvbAvWAEMKlmO
3HB4kmIryrmy/XJsbpsQ+y1AdBRScESxaXQLIV2ZkZlYHc1fk4CPoBQDHWM1V0uKg3Cnvg+E9MKY
2oUlgFjqPIRjipakNaOt00wjniRzzi1oFtLbaBRa2478ZJzwylgaVGr5KC0zdPsCjMf9as7IoJ7j
Wr2H0ZyfAWHULf5Lv1TuVMIvKnaejcagR4SxsiLTnkARNtTmjU3BRlqTBYF38FUPKz8YaEKpOVqW
5xF0sloJLDbCFmTmH/VPY7KN5b62dRbnTQwVte1/y+livHqa1TSioMSamsw+hT5kvXLHcZH4W3WD
yYRRcHuhmiwPDe0GS42x+BfTMh+3qnh8goh+dkGDXfo32LQwkxq1W1e36k8T2fFD2WNSVBA98HQB
OLe5UWSWdLrP6bDvQPWHdnXcf8Z8unCtGUURKiwZILPKn8CtZZ1n3Gc0z8+UP9v3VQ91hJ4Q2ZBL
tugpIOUHPZczgFswBtxWU0LPIf3bAWqNXBpsioxf8J/CU3OK4JX9zfkjyHk+V+FEvHuXy0ld18q8
axQWCY4KKZryfbc9g+Ccl7nRlWE6CYghWlRSNd9cu1VLJ+icFjnk8O6eZ2zO/SMVbsSmcwBJKnKc
GrGWQtek3xDKyj0d8QnEtRf9EnJiZ2swxDXEK90ON2zRPocHawN7VSw/4uOzEpuHjvNhw8qiUs0g
qGP1jGxmCLf/I5kjiUDi6gC5EedlXtNACHV5X8Vra3QkdoA6KVBftmSOyfruZpAfbYBI5GoWlq/q
2HKlGgvET/EgofnJj49FJeiR0B+T4JXcH9oThldG8/6+JUr8FmwvR9BHy042uPaBPw3Cy6TX47Pw
C+SLbzI6Mv4mWmEPsNugwf783FBOlkxYoW/MjMaC9hbDVYnJ73OyDxGIwLKJDhkcsm+MyEl/KdWq
H34MhUBvjAKVzGvUUVlzV7PIE+CPMSJVbDn8Urnn6xRKSTdnaRP8GdI0pCajHxjTg2MgHCojK4ab
IgU5t1oSqfMJE0O+UsCkbwcNqqVAMuWZTll+OtamlieGoT2ICI812nzyoaqnV4o8vlqzFGeA0ViZ
QVJyLDm14MWUGEaZpUq6IcUIJRaDWNCgvK5E/j82wnsJD2HYQLvPahZ0dG1FT3htUePPqsVz2Cnk
RYJfwbEImeKRH/RRlaSeiCY8msbORbwubmrsX0bJG2hGByym1QsINWU83vHZ+ohriQCFhAV+shwj
OCD/K5dPXXrJuL25H8f2AEWmAFNsJO2FUa1IUCCTEWAfWqf61wqX6Xw5oykzCGvoNVcoOSxAIX5I
yP6eOnCmNSirEtV6l/gAPlziO6G7jlS99yPTy23RWnDMzGUj7jUWKMaNbfVq9rJolOmLZY3NU2BT
S9drqBMPtNzT71ySMhlHH+UJ8r4r42NT/bDRZelIC+2bmyfbsLZdQTyJ0TMDljBcmYYS71yGrjnV
gL0UaP/vvIKakA8pYfEXMCE2NexwcSO05jSrQipjZOmn2u92uQSNEIT/yDQjFW/q4GkTPNPgajdD
swlevLDcBbz5k9Ax+eH+PcCUxU2XZSFiEenJKXdNaLlrNGbpl7QaqV4KvNmtRL6rqsC+dHh0vxol
QHdsnDWvm+9nieaH2i233ow6/+STzj2fyaYazdf74RlYvVKA4jOlYZwLXTZvKcpEZ6nu6AKLoX4Y
mXSn2rFSiB0RK5fdAKDIB2aCmd1/ta8q0ScbtF9JkT5S+Hy27UA/l6wZ+fW6HAuY+M7afXEMFDPi
RF5rL5e/GEMuLnDl1hBEudmyny+4nigoQteZNUFJUsSSUFN1jpyzy6q306JmLUfWhbZyb3U2/203
uhzTv4rXPDKfQVWu3Q6SJgBv3aarCbkYL0Ilnm5cwAXOEf03xT5+VgTW8oAhcpOadwA+mKov7Iyj
MENufNGSsi1ybWC23Nv4CKd6jzscndGueEtq6JYqsSnTyqj2Fx6T40XuQmy5d/r29S7m3iUlJgWr
SJ1W9iEJTd9sK63c6IpFvRcAJkwGDT4alDTxaspMhOmIxZP+YV839Z+lvb7ZxkLjUFT+/E4BsFFg
fdX365aWZolzSn9LMvdO/i50v83+f3jpKuvLeQXDumlOqMxy7ub6NRuVh/Jk7p3YiquONLQ68HBw
CMGDJlx2kmY0+ezYXj8A+z9x7jvAS7uDSIrflzCcE7QAB2mUJqf3UrEjXxeH3YMXZe5MPFvOQtvp
g1Dg1r0D2gatS29BkMPJ3PYVBlJErMP5kjVswMiqBy/yXbZWinIxkZb/z5IylAJj5wdDJ1Y9KfLF
2/lkca6ZoXOOAHGfiede9IFWN4tv0OqM+yJAp49vweWXl6diiKTAIbdUGZBHM6bTEx6Yi01kM1Un
T3hnHKaEhC57Ym8NhOMcRZ533uY+irdkiYjAA7na3+fnXVVfX/C1WWhGuLtZZsOazH8WfslWPjGr
3z+6wcyswMOiWMzrrScNMMpVrWXkNnpNO+UfPhnp2B0aBY1g5ELl1l4jm3mHZSLuuzVAj5zvN4Ym
p3Mz34WmnUIKGEYUvLwnt3fGQDnCaEbsydW4aWeBHA5P+SpZa9fCuXbdrapkVPxu9x1rArqXK82i
Zfqt08uObKtUAyKl+T9sgOTGpIdVZI6PiRyUK6502W1Dj0rahJ/amHxWbn/9tqOQJHPj+S0aqExz
bEwNku0GSzRgsJ0lGbUVcdjACCeo7Fm5cFc9lfQgg7BUV3/HOkb/EYLIn49eXyfJb+Mmb56k5W7u
+kyQiWWMAJxmxEnaAxJjo1QWwoSP19X+hsDzPYjsURVSYa4ZizbS9/drO5o1w/e8tccHPgy30RLc
OhVaJQFNePxckHr2ditpPLrCzqkqr1AqCHaTqBIUfE3V0V44nptMfHElSZ9IdMLmqAPwixKuxInI
RIkb/IZBwxZkC7sdFBC7oCQibverW5kKXF7Z6qtqcxEy1pmbdxt/ote3t4qQJweQbTCprDO3h637
EokkbTWML5BhDVyPgQrMgtrllrsEEIadzOmelqiQo0hNZ588BwoJsXfzEzII5xw5SSpVkX8fupiR
AAJP/DBxTPr63MbFZ2QzFcLzCXbtw7DQ5GHPqkNrGu9T7EX1RPwY8f/gLMQj2YPIIUWZn8Oh5H8f
K0vasZsZz/ELoeD7RLP3mvA1bV3+/3VVLCfT9ZAhYmc097TdJbEPKig7IAD67f633074H4naA9IS
fyEaL55cMTkNfMI0zaHbpON69bG7HwAtB3UiWpVCViIonY6r3PxBBHIwwDjkjD8gzWhTNfqSQs3M
0NEk9kpm9TtYgw9XqXNaLw+pojIdbSXzmNry5ia6l5iMnBW78q9GB0YMpfH8610Pyp0OArrOUDm8
Wax80/dYqUDGGGu6VxI0SnZiqKqb7CCd0Pa/WXUv9lSnt+FdhM2rxtEprTpepFS5B38lzHvjYW8h
oLjkQRXQDstK3hdR+T5b6QJtK3Rblt+YqAPAKB3UvPhU3ciPf0+ZvWQ817y0FVM1ozkjdGHUvUwv
yktbVIHKgYVyQRPMIySwP3uGJct9QX74mJJrK2Dvo2LY/XU2bQo6PADRUWT3GxqpNcG51BrPW3Bh
lQT8rGjQs3ljxnPbqlbiY1pgSWAhyI7m9YzJQziyYU3uzlKgyQnk2bsD7K24GyAkP1BHzBN/e2rJ
umTQqJ22AJDJN7zY8PHPJTu+qe0VZvYyJ5xrH/n0X8J7u0EG6r8ao7V7CSURPRo+/JQYrgcxK8E7
2w2kVO49FA+i4dqrPezjdFmJ8j85FCpFOkjOzGebcH/nwNX5FXofUl5JH0N9AYrRV3SLUV0dzd2A
UBthbAWX0men6wF7c8jM7f1Gvn1gpnLZQdbaG3iwxq0veB7viEauJn68hTiQ93NN59xETg7o5DsE
0Q5BcT7NaEMX43c2pp30tNxLC1CJEOHOw9uv/PCMU8BxxfPUmV5G1vNTjLrl0Rz+cyPu/YDuHa86
XVbnOOx0bBj+TiceTm5PhXnv98AgHi5GWZYpBu5lEgIi9TmDVFcMcQQzBLEtH1/iWxl2Bd92M35d
NLJ0yHXMbEM9RbbLtYiowlIWeA8n/wU5YuHn/IVPDqEhyodUoQRC/x8SEEDDlwEZu9pgdq+XiPfg
p27mt5KC8u+3aHq2EusGsY+g4/lkOOP5x936BNIiHXWm4sjQllo2g5BuDpreFb6GZX777RidVpKm
/HxXKpM29wtZlJdv4hwnIVuYruhfHL/dqSd8dUoT3wWsHdLPXzoag6kHQ3OuyEzUIKN1cA+1GP1Z
If+OuYL9gpMWlF6b/Lcgdmk6yuB1INBNhPtL26aQIyHuTGHSKq+zK9xAliEgNuvvCzpq3xRpEvUU
hYi8GhDy1AxoenSuQGWVSYpfUwy7UcU6QLwqhKj6Luf3d/6cxLFNDTciW6DkyQRxI8pjYoSrXrsr
5fN6rcJSCohftndEuxBVFggOLfeGlESUQR2iY+ddvZdE8qn2oejtqLaMsknLBrEpAmGiTYXR9FPF
fASwiuT7xkorXVp5/2jNDafLa/qe8Au4MwLPXYr9OGg2hIjXxtZ3rq8cF8kv/R3dVtGjOnRuSnd7
bkXHyRJdCyV/Hlqc79Om2qx2V9AMw9vz/xO5kN8WZeg3s9TSyPN+et5RWt48ztkWlWwFYT+9/gtp
wbHZSByCC/c/t4LVnVFSpYNshmfWfebeTLSkbkpTmxf8+TshBfeUgTdsQdVFsL+yO0DYEzZx7Pg7
t2WlNx+iwtIakJLg+QeEKELZdARgX+qmR3D0tVwqSI8Yg6ng+MPf0FytMLxfeeNh1unT1rpAnS+7
yoM1C3U2p6PyoHSJIJNrHAWxWAe5u5SKHCrKDZ4Q+Nd4Q9tnBqG02gaKGsgPESgpIdH4kJO3Adqj
Tu52mn3U2/phPLuIXtRbwBAqVlNQPP5zOv+YNWnQHHGJ3ypP18zBsOprF22ewum01d/P1Xqg690v
odP/JQLsmAGw3E9biRPg7XaQ3pgib5IxVmEcWcNd3yLG/KLbrkxq1ZcODtD8HP9ZUWTIblT3+wup
INaVWSFVXtum1DFnFFR1UWF64Nh2ZkiibATPL6iRldxyMBoyRM6FZXkfym7sh5qYyQpLsEurf5L0
4i7OTBI2niQJdhCcrYQtMLDH2st1ncoGF9lyyKCBGeiKYRVqTNnxxqpt/tyLJPgiScsOwyNTH31q
dpAYQq34E8CXA4m7Jvle358uumgAh43Q8YGyHe4Rgcd2YHLS8154b5RST/SjODL6lxGyEjW89hf5
JJFeO6s8hBaa7qFcbUsdlI5sgR5l9ShiNrkyfDZccAPDtLnrl/p22R+I65WSjRoAv8/MeJrQOlXd
ROTck7g979MyHwvsNNzTPFxr1p5g69NIHCJhKdBWkP959h/kOTGn5UhPNUT2IvqeIHjrnepXJECe
tPZvm2lKOUhe7UANkGGKyArCwrXoQ1Xc1vDTadA6sp3ibcfsENopgU8YbaZNQTSdMflPD+XS9CY4
CisoMjqhSiw5I8kqXdlbs5DbD/vzVIpwNWRR5cNDs69Q0ndSItyI1DZC7k5OEQLHm1bkfm4UgII8
a/w6VoWYBm+yVHCCsiQuY9ZWk8dt7w0Y+dBVzvqC7nPci0TEpCWqdghRQEbQYyQS2lUykhW2UKz/
k6tj4bexk7QzWuFaan6YuRz5MqZLaoUqbVzzm49wMHEAL0fQkF+dpbofmKWlw448sN1oKIqUs07q
zamvUPnxfWEDw+lfL7azhjaLp6rLWAytwpG/obPBXmlsAalIKhN8nFa2JWQlSaf9hdrE3Dol1FaT
XL7D84cs10XOT+zRjs6NfR3AUo/LK8ZE068FWVj6Bd+CFDk3Fcrpo3arS4Pzz3WSRDgVG8o68bGX
cCJ2domuCmANqdRWcjRmGG/OlUfGJVKI9OhsGYzh0DF5nupKpVniUwDbOBvITyJLDyz45eGYREIM
eVdv09Qjz+/zFZrx9K19HEFRpb74Y3Jq21bNQQkOu0wcTuINRNMIi2o1kGSQJZyRmeCBZlx5EuXM
dvO3YiaXtuIdYVAFNhit7HfBzh2mj6N6OcfXFpeV0XpjCaeAgzLTIKzclMR79bT+GXPFoDxC+3VN
lxVDfreTsU+X9yBaQp3xxqyuVwp+bsjbQkQXR2Z+U1ytR10W+zJ9084jvsgK4Mi2N/WtgWLtoA58
w5rDM5P8bmftuIROqRbkhlIi/1Lo87GU4w09Ob4iBI4BctNe1NUPGUinvz/dBorE9OT5mYG+qhpd
SvgYXMcNdqTr2qry8VzADpNJzIl7m+gbXymZC4sR/JhQS2vKmtPLAtDInUWZ2cOJEl70CxNzb9gd
BaBN3uArH0oqVkldwH/2+ltbQVh1yf0v+hoYOroqG52PEr1ahJXGn0CLPmT5BA4pY1GRpbx/auZL
TJYN4J9ot5OEUJRA34WDse9AAWRjwFSw34cI5EpoN59NLSw+YNZp9E4mqSvRGu6E8/BpSsK1pnlq
Y97cZ1Lp4NoIDWx5bzwXu4r/inqAOfFTP+3CZKZfzSih2vkAv4Xw3+DxD76HHwC65v0MGkFQVbLw
nzzWtT8BwBTgVKykv7lSkpnRXMwZv6OrGpvyg+I5C8rdrj/uJLErwRB6D8N6x00CU44ybyVJLGQR
JXUj3/Tt8YdwqeWWavLtjegdKcMSybjrhDfCBFXYNyIQq/u03hcDzpGiXwMJkaqoshmhOJE62dGQ
N+idmVB+EXxMHgdO6Iz0fQ8VDpbb6vwfHGvwoAy9Rciiq8fo8qxp/zuD5EeCe7dPWB9pzWvhhswr
LcgNJgJIkk/9uKJTGeqnSJOgdnplwoX6Oi6fEXj/fwjCBq79RD3DnoHc+v+Y1n6ZF/3yKnPv/2Po
bSmuKtkQYhkSYLD5fBKk2VEQHf+uCGuLwJ9Y/qBDMaM4+D2RNxDkUMBGkfD5BXbLMfny07C0lm1p
cEhevxeoEpHWrWaup2WbZ8KQIf9ozKr6Pk8LGC+w7M50y15X3BOKzI4it0eiMfpJPVfT/qxo6k0d
UXPsr0QbzCd+LWsmKNOdBMP4woBzqWnvmg4KaaHIpSVx5Ry5c95PB+nILl6Rlmcv4pULagR9Oj9Y
OgadpwX1DfSMFZYk2tg1TMfVipBkTWYUi5oomSvPANu9HXUXm8veFuNWHvXq6iBZiIqmkCox0Kn5
41O8C3LRotKnxqi9ZAwbSizjdhAfwYq87plxokWNgHx86KAmcpxftnrIGPfe4auzqTX7cOOGiarI
pA1l0Dei3wd/6UFwp8Kl3ArvmyiAzBkeN25IeO84EuEKzjar+w3eL7SL0xrIuS28GdZLSxZjV5iK
lAEbeY+fj0EO1KKQjrBKjjyuhZCNk18iJQv94bKkbs5vSiAMZ1a+Ht4O1tWleqqV0VNOucPUR43g
P1jAmlFjKI9O6kXugLMZDC1oN2KyT2wi0qshr17r/7YYWy7RHveVA9VoMyaeAEvwaITBAy/OFpnf
Kp9ci/7bSudLnJHsVODtS5/KtEq8YePCxgOV3iqu0MKkq6RfunE59QVEYoPcWKorSI0MhukrwYea
p4qlL/gCmxwnpvNZQ1nG1lPv+aUXPmZZZfNADAYM+OTYVDPkufQYY4rNJhNXz9Xf/716+Av/YLsX
SKqGtaCWVyHdmuRicHK57vnGBF4x8O+B13wKQ3jyAOX4LYyTdRC2mAVJT08CjAfmXcosSxT8R3yt
+ucej9AHHJ/nlHh2I5lCvTJ//Ec3JHtsdBNbweCSuZ2Q2RPmZIxbqgqyEtBBMopWG6XZIpCfzQv6
WbQT9mhcr0Lo2xyQwkwAXqo6G6DL0dAuRA8Lw7KXqyM0cZUSZj86No03yTXBUnGTZdHj8/ybh5eL
LeHiQLrJoat0q+u93+WdwVbC3ZqtKWJB6IaBMUy+DXkudgOehZThX65jn+Q/34C5DqxEn0dPob4H
g89XkaAgRtg6u2JVaDj2OR25GgHvcobxLLuMWwL8cXU8fPhFtWNQTsA6JMDLBx8FV5dcSOtbdlEW
1zI9LvMeb6i+Rst1X++S2kNQXPdKrR9QN7Y8gDxWvL5W1sk9fD1Ou7MUtIWy5ez9VgapQyQ7n/Vz
UCzt9fRcY1E2SLLMAvVtG4E07PM+kMTcU3fourTcYtK1cOESm/rdPpfNuAvb/Gs4EJEATGVcAveb
YiBspwOfODf8UtHUpXs/WYDY5Ug9lb870eB83nKeQLoS6FnvaTrwmoqwqno6N5fnfzTKdkXQuo2H
G65FSEYSCy0/uxYwQ5mjfq8UmNG/SgbfLijTpJzPTgWPymSfQwKEDDQjnqzyOUEVJWrsgx/eb+DV
wIhAeDWc5BvXPvgcjtBfWx6HbbWKl+O75Z0ghzwWK3u4tPiIlM2vZ9N/LJR9if+4a7gNOtCFOSHK
gospN8ulFMg9SDVXVOsm/nF1CGTbJ6jicGg2D/87D1RbPBJ4ggKLDWd6n+i5NQinphEdrvZKMf9e
5/CdtlgDlgYuUNEDa/BLzrJJDPo7PKVlaLWddmNN12uJLmQXFeFad/XobpkZS1LQ12vMV9We+b4Q
opDepzKQGNttd3hes2iFTT4942YwiIg1P3adXrymoDJR8A4H+FOgiahTll0clC6F6iilrXVgfhz6
o+WHHAgxPICVzmFj5zjPjbXxMHehHwGx34HJGkmEwEFUukxo7rLBj/CU27GQpI4tEm/uW6TjOsTi
2D7OBA0U04FHC4duZQ0xw0jVd5C2KuG+qkOV7KxK/hdUZ9g2KeJfc5n0+61P3kJYzbzqmadMbbf5
JXiz3Ls62cnzTBWpOPkZHpMdnbhwjfarfDPWkprVxB63kn6wU+1mjos4MROgcxh/2o440175lP7V
VqfaYh6WGFeeaM7g9M4mgis4zCaXjAQ28VMI7FiRk1rgvIzqeauFRAknzaKn6R27RkeKZtFUCWOQ
/g13THn7T8ucak8aXGmaNz8Sc+128gQO2sF+QEzgqTkTCYD5qProZh0wIeXnwjip3RNEXOtKyshS
AUvUczgHbplzUhp0J4+2fuHDyjQ9Mjt72QIxwIc0L1vnbMnq0MR+RxbcKaPbQVGu5PoOSjIvm/wQ
60cydCFezyyJSnSJyhKIvMT7c2lT6N2ptubflZGk7O5XnJuhlWaVC703lwULsDjXr+rVRoIP4Cnz
4mhKp8SM3U6UBEZU0e88iCparpTOH+hx+vDe4K8+YePzGRWB+HBlXpKn8cKSPWkDpZ8iK7XIPZr+
fJHO8jy3JSB7+0p2A/ZArfez6QqItCdFG39eWCtrDMdWLZjiidOtXV4nu0WE/xbywd2x18NwHEGY
LoFBeUW/VgLJcM1TAfKYysmoILAVvFa7Oox2LR2QdCtIg8OdPuv/adlXpON6RL8eJmLeddeuyU5g
MwLYxm76jKd2ahEpbdx9k4CXSPaPji+wLs0z2ogIg3qgRWbKshl0jd7ns7CoZTiuxihS3gmc0bqi
aIgf1i8G8SaG/8L4kaqIBpd92udlpXZwzVcdFVOfVrF9lUcJKq5iNQhSZCmIS4gbnHhHN7/rgkt6
+lNz3vXP8soKOK1mqJCgQj3ud5O5xwEqZ0Jh/sjytVHYiXIWji5g4k5tME4JPmHs+fDxCeMuUdOW
/DR/0I+1ulAQcbkyoNRFVswmjDQ0CJY60Hx5AvBTdgD5WMi2XUde8uU7ZuCenUAExZi1Qo0hya53
03hSZQMQ67bfo3/YThi7WdLGGfbn1BcesFcTUvEzltRLE4jpkbr4k5DbSl1PHJQ37SjBERk5XHJv
KU210s8Zji2JKfdBv1GwZb2EJX213Fv14ip2klmVLgvhRYd8iUYNVYEJOu0phIViOVXCs3bY8Fhv
ErDUO7ehByH9rTK+yy/YpS9mgUlXhe/YlqAy6C7TZSu0+rOykLbODbx2K5ORVNg8lX+w86g5hPjv
cP+2CTAA0OnyNvILhEPNiotBR5eTHlxgaJ2ng/4r5xpsLCzrkXq2Qj4CmOggomfZ+OW+mQYTOKrr
pIqb6oKwfBbUcFW30j6s15+Mrr4yW39xmeqDuadJiNhMm1JO6HYZn7Y2Ks6ZAzGd7nPNQ9iZKeM8
sVtqkvS7Ki6cXuK5LrWjqjMdB0xbYF0BLGu90lByHn73bF390hLmHYaFZn+qCcr1g2Qu/YyWxnGv
VBtHa3iqpbk1jxrT1hZJRxGq+m/U1LR1EVs3+yS4xR5ixfcz0R2kYeJKaykYzttuRfI+uoyRFz5G
bc1L0eojSPTomV/1/Jf9VHIJALqp4Ii6sCymOPPHf1WGUXKz13Bfq8RaXi81FSVfX2C3Y452XW4n
OD/26k9DYSZeye17bIsNA/DyoOSvrg3GLd3d/gcVFX/OPoyr0hQT7t9J7J5s0BtANlVdvzsD1w/l
boI829wRXLbzBh/4dstGmUpN3haVDXrG4dd17ssIU7rE+QDWkKkIF0NnVauHzQbKv+/n1iq9FjE4
Fu2EnHEoqvb83LCABgAp4jw8zh4ZUMghqxuT9Vrls4mFtO4eLP0gj+X7fhN0fPHGqe79WPoxI3hL
PbP+rK6eWC68u1rPoYyNZnCjycj4KiMC5B0BaCof7fCN6OZl0Bu8p6cVD0Df+cVkXFsYXB5V5qhB
Ou+0QESOsS6hajs5qIH9BISeHNJAXPt6yuku1PdqZsJCBDUbAy7QjNXbdgV5d4X4eeFlMR8TTZsD
NIZ8s2NzyE/yzt5cyHxXN1h8dUrOK3d/Ip628A1v3gDiRUEIsvpYvfPRf+wJ8cnzhZBhhaT1xXEW
b2Hd+tWhAyw1L63FrcWPslptFSghrBuD/ggLChWTcbqu0IyfHN2hzsviFu5+5XWQg0L/yKCbh+1M
sozcDI9orZ9GVmuOgzgVMm7Jv5w6OgYnlolxTvizIINRcdSdUS7GkK/V/ZXLR9LswwACDxmffHr9
PVCsu3aEjp0vVomMnCreF4tDDRqeieLXzKG6+UmT3DKtXkRsu6UXscoEOGwnDhvCIwXPtCQWl7H1
HQnDLT+lcQdngDngifSHUyMfjPKIrClIk789FoHqqvr84Dk7m3LvYrdkbBhHfPy+ij4NVEq+nXTK
IQPx2/adUv4pCNMAc8wObYoFtuwZuXr5Y+T2NA1/mCKniLx5viS6Z1mLvMLnB2YdVJPJOjTLEuxd
p80XcNIEui+nwrBCBiBDXPkCz/CyrE2klrB9qU5jGAdHl88RTOoYMjw/zG9FGUgpEtaM4r8Wo+Ac
RUzy3wIqSrAGD7QpWyHKvfO8yW7/xWKCe2eeYPKz8gMYqD9Ovs1CVeoJYdy+zs0iFwWuq6CbZv4R
yhtjpPpbE7DU2txEkgsuQX26Fr2agx75FRy4F+cj2vybcndVsLljdJdbblDgK9+3Wtz+kYjoduCd
+b5QxGw0tuCl+fQmVj+A6e9CCKEKa32qj3RZLKz+J5FL1n1pGeOkndyjWQh51hosJAuOTBm11pSJ
O+n8qINp7gtzH+Taa27ne/BPkzVhDkl7N832OcRAnCSy/iVh2+hUfuZ9KbUT31LhSmh/zUU9OSIl
62oiG+5ZtgrxMq9n9tYWHystQnOZz5w0Nw2Kh230zXeKQSPNuTajRo1IBr1PGazXNe4pmjIv7KuS
kwtBsnVs41olLXtZn2mYZwpIYXRyX92hLLtl7LCSdH6Fh78JcRypbX5AJ6rhyWMzwJ/mH3wgM5Uu
CfM8gbDF5TCTVRo1byaNbvndki2+mpbIP+TPQtXYiFGzJT5jBuVN/nU4xU5l1s/kBfY8GNp87Zwz
hzLudQ+7bS9s9KMqt2UWUH9pWvmMp3PlKyu1UtFpZuyTI0oZKVNnrwHovU7nSrgs1qHZmNOkmand
+tyuCZbEhKmd61z3I9KMaOkzyEjmpFystTN5avCvHgz49xcoCgw7OIjMfJBv/o7Z8Oy9ux6Hfe3Y
PXltMo8b1HawRmD8bV/meYiz92a1xvDPkXd1/GmrvrkD0c/pC5sFXPt8CzlQzS1LcNgM96noSDqj
vR0leKcS2PEg0n9JDrxyrtkTLJs0JvSPnmphsxOjHt6hwvpgHInnN9vSmJgwzscht3dnR4r1JkIA
/zuGispRm1OFkdH41mvsEjhwHC5eS3gOeeJl41ip658Ld68D6ykAIJGNgwnDwqzO/w0VCK1E1O/q
ng6y75ZNRfZ/BfmMY58OW3+Z2c+gAnWcwMXnkGayCRVZ8ULare08Udwl9IcpmUAh/OOT4OfWuEJ9
E2LytWbjdcalVxM33yQ5F6HCoKvE8Gz1gadNm1IUytwm0ZzUbNONgQLVZilz6CZ8wXKUVyiL85Fj
w3th0JB6zb/MvXAgJcfmHFf5WFxS/4PWn3xSteIRnOrM3B4+1KMEqOGBKzah3bsMKw0Xrc7HOEoE
P+HEie1Jw3614w9PF/0TJb/unl/zBIuQXj3rJL2iWEsxEv49lasWEmwC1DZZodL8eQaP9ZK+P+On
xoZI3uufbN/ieIOiLUAonwh8GB7PYrTlz6piBcVz7nzbT7taHlrac/sM4RKzomembZhMBWzMJr1k
wtKxwtS0kN2O+5ScwnAI+1ECqO5k4EvD4f1AnFOHyNeOdzNRD9iAzol9W9nC/yUONINGdMbMI01l
H9I0D0wIjO9sOcb/3Q0UN+8eUM0UtvFLhUqBVRlsOlYLLiV8i/GQs52+r/i9NY2cwqsi4AH7rSUK
U9gZz3VDIqe93oAR6od54oOrU+CnrK8ayIDMBqw/w0071rMjF5JboRtCZnetzxqa3XYu88EU7RGe
ajasVU2wMF1zUyPMIkot9IGTf0XKqnIJINejIE8umX2HaxWnY7thtmvcvxbFN0LaQBg3dwgMnuaj
iQ14o//SdLJqsvzEZZp//2ilC+Q+VdHNW1VylvrW5S7GMIe6S0E0NeYCZx7QgyEypgEyHzHn01DC
rCsBNPT9xV3I2GKhiCvHKQzZNwsaTLlh0BXbgZ8ROF70L8gUV385D9u48yCTRx4hvahaJF5AQN2Q
KIZPa/5fhvhHpN4+Yviv3MMC3oAn+tAiVADxm1FNFiNzcJ5e0B3KSXluUQZzdC/ucAwQMam0WWH+
qWuoAusxvDtpPMZyFKKuuVSoR81bhlVVKIeHRPn+w3w/r9bVg6kdAVjzLBqGW2uGp8ayc6H05Xv5
eokd5MLREuLdkLJtuqkCLIXs8n0MK2Y5sr8nD/mH8d20BSHg0LowZ7xQVC4aketSuMZc8TbCkrFk
QB/QEqPT8IR66traIsy3rBzXqpt4CvQOyd+Py9zJA/N25PYnpRxEWAgXj3Mp9be34kpuw55vgx2L
ISslvIi76Mpygo2H1qBHlRzJadrccUe+fZVwFwO6HZ5ziIuH2ngciH0Xm0ryAs/D48gOg5sKCFWg
1mEbk08crmySbGTu6xgwZM+U3qhkJ0tT1yZtk/vF8Qpv0YBAopJAz8EBeeysZ+tHP4t8NFvQM0/Q
HpGmQRutod+n5G2pPqZ76SkK3Fd7Ovqv2Ko5inJaCuepftaMcMx0xkUAJ9bMThV+6UhzRzjTv56g
7vvVdLMpNYfRT11k/uW7D5nyyHZ5EZpbpw3nNAz1eG72AqA/bQDJ/Q88URv5nEluaSAtcrVpH15J
vbwxPUXgczv3ApgdlefmsR4+fsYOubx7ibBrlXVIFtAXl2S/4wvOccwOLhZNzkkiYc1v6pqmDZxq
9VvVXyavYeXgs5PUO4t+twFYIFAWGjOVkeaAXyjdg3++xCSlrcfRbWeAzNOhWDkyGLzc/iVCTgdU
m1945Thw/zbed78+uEWsS0MR7f5wzLzy5RtD7X7FacfaTlGt4k8R0eAGRMTzK1ldZJwO9fBabJ4u
ljP2ezz/wdFUqOefpmexOyudNoeFg3U+sdBgzBxaEICE7/krLpjU1IxovmK2rkt+nnAB4CDu4HqY
+q4M+dpsZvABZHRLmEWBEteuc0codh4r6ouUsQBJK9QIZ8LCqAsyw42uFXCMK7OhTQBiXPlo8KC8
6bPu4JcfWqmiIwlLXZhlXkAmXs1R3fRWg0iXQTD3QB2mw018AR4ObLLlnMxyZivfDZ8ouBl4XLlT
LNAp8o9mgnftqOB59zRvjO4LR0EH4ISgbXLtXhCErDF35t0Mnz06OYKkcXCahlDcm0WPRo/ArfnO
NqbE40GpfbDsdsKxFNm1tQif6nSIWajVminJ6oXZUAWjhpFWEY6uDDQYW+tpm8EzWrDIscACcr7z
UucxdeFpYZOUYlP85J5AxI3DwfJM9NnpXQk03DHg0T+QoHyydwvKjcMvg3BXCY9FWObWEI3+7A7p
a0q2vBSN3Jpvwo10SpOnmIlEytIHtEMfvEIcVdUIYO3HsB6CW4LsKcqKyS9ZzVuxmN7Zv+6z4++H
LLt4QtasPTXntHjnvEngV3HwHlQrDaut7nMoF6BXzEPcHRrS4S7KZdeybAvn/T+eXD3AFYfZL2cE
W82QjpGpWIjclLXYLabVQKxo4j4QexgGFeyxyt3xzi/uIySNMPmCkI+1mkphHyHnQNUHSbxluh05
qQumj+MCEFMj9eMfUNp3R7KUbdyBTxqp+oI1K/5zE35eyU2ox8bMLtHekT32z+TLoRbbG7eZJlK1
08E7PH9YUZjrDNKFWOnBi1aFw95czS5mtey4gzY46KkHeJN8GtzJmOPLgNt1Swl0I8hD7wgCKfVv
Ay45MeVBKByi4FxS2sLexOBH90h66FG3uSk6Yt1cy2VLneSNhurUawprIJLg2J1kgUH9nIimE2kU
MGPTwc70Fox+uDnO1jBXPM05Zmyomahko1GklOImKwfbc/0IXUff9fgpH/9iqD8/XvV9krYVbZx+
HRTCvAj9JFqzI7Dh39zCU1+tTVsY/XZ81GBA6QO4MEOaLfJyIp6JblNC+QO736Hw/XN5OtTXPL2W
fiC2FsybxIWewz2D3WeTR9Ih54px3kK1pLgl342Abouwcz1nVAMMV/QIzV211zK+BtvEEBb+OaTr
gPF+6tZ5tNtaAWjlQ//6oremE+Vk3lyChiEDUqebigD7AmEANrkVliz8iFYn19a4mATgnWmBKt/B
l+Gk+cC+4cuuZ1oQVncprw/xKI+PYHegF4GbOSeKLiPjrFIKK7T0vLTKqtpSTvrMHOj9UEDmGtxD
Upyyrt9pnoh+gMWKT3qPTquzFFQBvrZ1xoDVtzQo2/OxX0mF0Rzn8SPO8cnrBQnfBnUkd9e99qE4
v20yppkRVSDEWx8FJPYVAeuHE0QhSsacnnP3V+xqk9NgaLu8KhFFrNy74rO2zOT08HY9P4cePuDF
iPWOjPrhlUhampdluzT247tJET7aAuCj0PDEkWIAaAk5Ob/BdbP/K2u5WVqdt+2mLTGf4/CD0zEA
sjgXAT43lgsat2mspcmuDp8BrIea6g5dZgmqR33ghnN6ZIbW+O3ius3/iEvBxSH5baP/W0qrlrsE
eZSZaSGrp5mfvAO1REnVDW/zxVt5eptdJZPbt0hLKAv0/nAkZB6SsbK9vHIHt9tU3gclGBMHTTUd
rFW3PBFTwKqZzg7npBHBr5LbEi6SWBdH934hnKw+UyCWHipo2/vtUI84qntf1+Ix+QBwD32zFkoH
apIP+fPlyB9nzOL2QaicBvnVfnAoxprI/YXO01YX9DW1pj3Ali8nnExOXSh7Utwzt2aOCSsaeVDJ
8dGBnnSS9v0JHCOXyoajP0w70JH8maj/OnQ+7BMCODYk/ZFZykVI1byv0fE5HV4U+zJzQ51BUAmL
9VWVieruXZ5clcAyFN8aQe0xufkJAojQXLFgFZIIhCwYnDRFig9anA7nmQxk6c4Mnrn8OofJA90t
zInP3Zp0jwNCTKMRj/Ng2yIrTsJqP7vKXwkbvncxYoG0Cf4ui4xww1B2gx2bihd5UXcgpC/AyWrB
K5zYF1Rs7miDundoTL1Ve4qFn5KUdKBgUv3Og3jbP0FzMY26cNbvT1u9+KiFG5CnVYlPPTpTw5lL
CDnQ/3LKja4sMw8oKp4RUo5kobrcP7YT6GWehdcHD1R56meVlmskQnQpPD+5BBIAyHtC5P0DKCDb
w563CZuCzOY4y+UBxc/YJKS+CXgcEG7MIeUGh/+mr4XLCtyfgM9ytE6Fw6FpPLCguzh3bk6vjnL7
/ImGHjBMVGTMir2eXIlU3O/FvawIRAdeI4onO9vKop7QloN289h+YrBgMepAsPntTy/ar2mFwduY
D1GIketVcyLWPk7iRAS2yGGfNCH3Dj9mUXjPLDoSPyIuXKZg9KA2JyTZt5tqNnq9zn7qLcggawNv
vUI6p+DVGUu0Z2e21+1vRKX+pp22b93d2TU8BAA4sZCAOCyCVPWPWtqM1GLDfFMbWgxrYxsdoa8O
iIYvdU6whMU9btr0zDgDZk7FtXRrHBMBCfUeriifE02SSD9EUxJnrHpXV6JqSODmWALFXbOIBC04
fHzIbIauCakDRVkCGy8AcGPjVfPe843Xk7KtbFt0oklfnZuwjRVbRAGiQyZUTgPu7sDdYq+USwyP
ABjX1aHcPcIawUcmTb8P6eZIQw5tRx82dXRJ88r4oLCAtHvF95YWzpAho/hZAgUB345OXbGBTzC3
HvGKecRwI1rWdZ4V+65ksaObp7fiyB3y4aWil/e957DzWpMumLu2h9EffEkCBBb0FfwI1S258HAk
Xh691aWDtV9GSLFlmiwncgL1Jw1YILmpkDKXJLDvQ2csBEKgY+Dw0n7uQZ3E7HIcM0kG/2DTz0Kx
y8AeX8DZbgUBnT7NNGDliCglh2j8ejiKcjyjXN/Ac8BxF/49t9cuqfZe8sLP2ybczeJhFd57CdAF
ALaA8Nd2xglLT5+VO4lzIqEJofleIT6kakum6ipMmW83NXu6ZcdGIU8TKaN5wpjGWYCQ4AtdMsMp
uAuqidf0xFBASuxHwwObM4zutNqJ14b/HKNAxSwPItyWZpGWb3UD65GZwMpdv28Ac7v2QUrUm/Ff
5r5dbYrnLl1zy6Yn5qRU19hPY2mHS+QPB6/mBYXZTI/+Yb2AN+35J62IrrsYqJtP/3XLmDVAwkDK
QP99KQgVK+2LfszFOA9vcox7vx/HTvYpjRhkJqJjN/jwAJdlfyOG+o6KQa2HY3h/SXAddXGC0H8b
AdSgtc6t0L7/USg9z4pKqycxHN77/jKwR17RsBd5+mFf4rXaS97jXgbQv7Qw6Ry4rDaQt/+0Ocny
qhaKvoo9uxKW8tibUgsL9UGVyt5W2VvVUXDIsGiyqGzPzfK5DEQQbbRdgF+XwoJ4jm7zUP/1QiDc
WP+1Ar/BSNDozHXUv87GtcDdxemu+xSiCsGgcy5eTrBjPauZ/2DSLPeGFW65GelgSOQuGrPHS4CB
opCbMs5T5l8kjieFfxGYb3VJJqf267iCvGwHzKALg1I1ILFxLFXVtrisDNUxrFE6EmQR2h6mBzcj
g4OxtZp+L1croyVAKnNK+eI/4MyCoZx2uzIBuA2XS85HSY3rJl77BmOuHfHDo1e53KWZAneR0h3C
rGcUpRjPU6iXwZgBrWEUb56TuEY+moP7XveqO8J++fOtq142TlyNGb4w0tBISJnW2VGQbSM3jF8c
AEQhIgtolgadUwSWJs2jj8u7R8cEzjsXqhkwkVpvEmL7CjtzKWVpzzRjtksoz5IKeCetlJEAPU31
JnzyLMunN1CnJt13WAz5SZgrnMkkKRaeNhQAoBK7nBV3N0d6nobHHSymniZmzV9XN5QhoIoPTSmP
rr3xJpjdbbjzLYszTZrmq/nbmHMsYSMie2bkxJ5bk/6tKeRnUsr7qRVUGrCx1n638P8u3Mnc5ZjC
CW+ZzH2+vOaEbXF4Czoc3wrcxCaH8S9EbSWl+GWyuULQ2ELXzmGELVY79Z1XO7BmmTKzEfERbyX7
C1zHVn/qxba9BcQYeview9tFPzVDAWPE+pU7ONYoVqMr22vtNX7sF75fNs5KUVDf/YnuAe80WJOq
7T2FdHuI3x5popDY8Y2Zfe7i82oM4n0PHQ4BFQ6e3ykxkW8slmhO8L2C7tcuIKlWbpNklFRqLh4K
IHIwcTQw5JXUuyJdhFmXmIPjQFtCdSjJFDjbP9eIclc/fhH4YRu2LLQBeiPeG8JprQDyWGLVR5Er
d8LP0VbIFfb+KJbKTRcQNyR/XttLaatvC5MN8Pj4EsXGbQdVsKyDAesv20bF1oB4e6SNu8R2Jsuu
xAN43lDVE6pEnX206EkFh1PSc9IlG0v60k1kKGzCsKkfS66mMBLfXC+6iopJeEvOks/6obzg73G0
k7MXLGARk8AVlsxAtR2KzjC8Y14fOkFCgSlgkmxnmO3Y6JKgA24USihP2/wuIOA/wmYYs0lF4kih
LVUnkLzq0gZeRkUq8V6F9y6jC3re2tLGLXmpZ+tciL82roc76vFCW/dTWfHXMHy7RGh1hxgiaKlp
2AiW9jJMG9x4sNsL+anZSuKU/uSQ0TCStiMyZV6SsamoXR/rcuDeMGQLJlx5ZWcEbX+ekO56fSVa
g0Ozrgu6GtKKQ6kVO3RYhbrRpuZHDb1ogVE4VEtNdJrzxra8b8E/CjfxIeDbiDpHSqSqfcYQBmsK
fEuShPgQE3nYna2Oi3O6qgHCKd4R7gtr9NuHvMmFboh0lL6UiqUZ85MpL65NDC8eT0y6oNptZIIT
GhXOPI3aq4ugr/31msmyPy+kh3m4HdPRD6zHmo1x49qBFZQWjeBM+AXqPct6NXwE5AMDdpBknD+H
vWFaIatJ9CwrzeRu+yUHSS6IizxfOzl7d9g8oDNE+gEAGey9za5HamqaE8EYkBwreBoSr/JaCeqZ
mWG+YRj9Y6yjCYEVe891THWlT9z9+Sp1GMK77aWwVwd2vpRW2Rc+ZU9ubVdvD76AdJ2FwYfV2OZg
fsBBhVQepe3troW0w1GtEvkYOvBj5CDN0lgLJd7zBomj6iq/Jpb82BXVRaIhiv1kp4wlGh63rNk6
3T8KZ/cdXrbgYlj4X/mbEvaUTnzLBtGN3h4vkCn+O3J706rZEEOBoe40gNgd1IYEUBH0DhwQ4EBb
tpX7f1+qnEW8ITSWHJglgKG0LKNOwEIaKzZzVSUEpeHoSHdZN6lpXG9LFX2EQ23U1b6YzciUpVni
HAHSO7QyrA52dPdZJ1PJycYy15D9HvU+E7yg07GQCCEdPgFMiexmE5kZ/gyug1x55PtvErSnfOhW
9QWwxsyhQ3JXhAhHyCUcfmfEdonz43vD0TZmEbjTys73phcHrBtHaXMA/HyXU20Xvc3CAmnZAPtt
hm+H5FutkcOFSOya3mqGuTiUiTk+0A3I7dGulywdzBLEpG4w6OB26Vp0YVQ29OS8Ai0OX+su0OOo
XO3okCEKVeyzsEovCLdGmsu9dAiwf6oXdDrowco+jgYQ56WxLtZk5mMoiGzZjoy67EryoTzwTDBY
9PSgxgBFar5AgihNsmRiwsztR+aUeoOwR5AYIuiKNwZCrvryxOYBRCGQ0KAkf1auI+ydIJq59aCT
MEi6SYFtlVShzqnr1LcLnafhFOmUai/0qaOUFIM0kzYab1s6BX0n/llNqEIpGhtUnbOd+q3kO9uJ
fwzkmkofXO1doH1b1mduLjgRmmdFSGEjC4ugtvvTN1HuODE3udD8E9zVHBTLIGUDT+OEp8Jf0uwK
4yVM26HNRdQzsuAUsZ7AdHwQs5gz/fwQ4MX6BkSb7ZtX8H24ka2+z7kF5c1NBNGcTE0l1BCZXeMh
BbBkpGU3TRzmRjewdiV6Lm/oZm/9CC6hiPWLrBsNGhl1VwxkyYnQ3B6/PznHRXSbRmMnNzOxYE9n
dA7pOdVcIb5T6rFSPZhgcWnf3NEVDGHUsd2AmlDcRj+KUKyEEEMW9vEC0eAXWijH+wTp08ypIIhV
dAvH8re7NIyb4avWI247gU8zLI8KlSyk/l54FPDlRUDuS41VrxS3ht/mXfxFPBUCkzJKbrnlWTaV
G3z1VpyiozqE+A5MDLqQJJpLqjYZ3WDCcWWmQ8ZdAmktPrfQaqc6DKyPLAUeqVKt2T96goW99CIV
sT+lZZ27LtjkfAoW363XVggzQF4jpLJd5woycUrDF73E5PBhPVTNcT/0sCZYQbzfpMeQa8VveDPS
xN6Il8/mj70yiLXf/aYQN4zVJoej4Bjy2wGCb1bQvTPWnS+xhPmpXJcRnlThiMmF7A45tjzqCme4
vcjZNJNlhwMVSx7kPakG4DOwRMVc6RPtM1lmvL2iQ91RtgTveAYxLfJ2MJYsmtnZ+L6GF6SWNOzM
udsIppY8rhLsovNeNJUAyQwiHimV8Jtdk1jA1UXjP/oHhyNRKvB1KzeoZfFHxjF3F0PbM//r0nuX
CqL5j4bMkmZpZJeaqGYE6ZGH5TyD0lVHL/MtGh0eK40k4mOUB3bD2o1LIk2Xb1Tz2VIzZKU4H6ZZ
JgRYprPzOfOLCQ8Nqj44Xp3Og6wp12P718QM8HCk8QtpesG5J1m1JiQP2V1bSeNH3Gctd8pdoWCy
zAahZTdkMs/Z8c++NDHAb0Jh/rPSj2V6r5tUZLMvEV+Z9ohSpmfDi21LajBafXz6A0VuS4PFUoA0
xcCo+H4rrpafteKoiTV57DeOBqnz9IWAJG/y3SMpxXa8f/xOCDzw6QRSWFKDyqbg0/ycZRsQig3C
0l7RyyLgp+Wpx5luwy9UKiFO/AaWPRSpErZEqaVe3vGaqpfRmqM2ZLwo99ZDY1Cejqm6yMBOJ+R4
TOub0SR8GR6EYwXkgyfrl6HBsiKBdL7ZsH/Kp36duusldHLWkfWT8xHs3UYMjbazXjJaeoh3vRsw
O37kec+ZetBlCVd8MSIBDJ6tFxP2qaulcqBomLtwrl6z7EyqFqmNUWz/xtWg9JcWNBusVGkrCMQu
zF+7CHyHS91qhfBZSnEGzncYL0WX0qXvxWZphddOP1sBBWv64Kpukyx3tYEi/1k52B9srFvJo+ML
4l6n6UCCKuF94DYEXFvow1WC203nnYeSRtLLGB3HAg1MO/7G1oFJAvc5Q3piE3yX2+dEbqQGs9ks
CBFI6wyLSnWlN1352kWnZMCELeK4nc7/DqaCCO8RIvWTZUfyr//QEJUO97gNvCXrFZNAoxfpFqKO
+7dDWYwbTqkI+H/0sCBwgP4rQ8rHBGjeaVOfiotpL72PtoJtgHvKQBV/BaCaZy7TUcGmqCM0tWd8
B3n6V1xbtxZ1KeoOdKmGN79BvJfWrVZQiJqhACi0Dbzl4QbzOIEcsaT+jl5J6Agl7N4Ry4plWyOC
uthcQa/HFn8cKyOUOjU6BPViJfhdprMGpepTd5skthMTU2G07WJdDflXs6LjP2FldejElPk+4l28
IAsY95Zboolaw963UbfJ/2t7LBdwFBblteBRzTms+0gUjRoaHycdMo6M8a8nPrMtkebFa8Gfxf0I
9ODhC0jgEmoaSzMFvMoTBhNBik1tux4ZZZbyxEHLm5/MleQe4+bv+JHeJx1S77Q+nBI/BnxnEGnc
ixHAoXiZW4F6x2BjqkYr1DiA00WeARTBaw8AHO8wEKNOwYntzYb9jCUHcurhxAEJc2wSzfXEzBl3
jrwO9TJmWVoNwWwpjcWm3hWFhZ2NQFBt0RwZ3yLi3VcTNZogrAXDfgwvXeBC2RxJ0+yZLcR7q4SQ
z410XqWW9eUMDGTf1eWNm3rlrwi90DqUjhB/GPWoaJPLXoMsgxpdbwhEsgIV1AA80IraCeoNAW8t
fDzatPZAgr5Lqc4q0VfSr3jEQeNX6Vt84dqdE++AYLjkbDiDEhQHzpM2Eyrb50XMRoY5N03a8PGQ
bxT4F/Nxax1J4fxaQg+q4jK47ZTwumyDdi71/RyFgYv0RBNUf2mKw+TI7+jiGSmKiKrzjNItpRNT
aLv1xB5hYf+9xFSVG8E8Ilf+Am2SVlPNcdWsiSTj1jWq66ZBCfGFJLSM3GUjbGPUwi31sSQ1D1tZ
O7K+y3v8WAdJtE3qs3/RL4/3L5Nd+RnTdrwC4B5NDRX5eNYst40C3mUAFS2z8TEr7Sbh1kmC99bD
Dz0t+ALyj4MmUwt8ttnAj/g5m9bgrmu+A+bSe5I3ZePkseAvR9dUhU268UKeVMcjvEnlLAGd0h/W
jWeUOH3MzgaAGXVdHwGG+0dLSrJiWeXk9jja2xK3JlqBYHATKGAQh1FKiUmL6y3F6wmXbH9SWB1v
jjd52iPJBObPTmzi4GXalL84BM2yXiAP4YkRmrLI/ow1wf9RzmagypHGNbjLD0Sjhprg97qhHXdo
N2GNOTdSnM7wRVKuwwlINslWxUaJJHOji9rOlOhQrlVyG2DOqyk/o0O6P1f4TNoRmCwO8N8BLUdi
wTQss6NcscHSLp1dgnKfbzSluaHdfsN1KNMud5RZaD1qREcXNEAIwF90JbJNScw3PizhiMfyPYQx
70Q01kjAkZCaM0JbEQ7RWwYZbIxlCYyAB8JilWwOExHk/w2jWFo7i+v8Bjh+gYcWHz3+e7O4wCq8
7Smj9xxRkzU8MKg2/D3fcOAjlkbgJ5j15HlHd8AiVZe7Mg2wCKJNOp07IriSBWc5O7S8CpRzzrFc
mA2vKv0d0u3yB6nSdRKYJOZyA6cd4wEhW3vLrCvOjGLKb6cHm44YmyQ6ceiPqBvC+s2PuwwSnIIV
1PRM+qBBCy0v1tNXuziDWwCeWXiQrc5nWWunanjVm1EEdV5HEjTFBJf8Z9Cy7qGtDoaNQSY9SvVE
7z0KSLpNzz2BeGGGskgty7A/FIf2HzCqiJ47e9GzzmYWBD9cCievVMaG370tuHUaHCWrEemJZ8Cm
N9szXS/LpBaSW5dyHqps6a/lOOccKV2QWa5kYdG9F1ltQBRex8OlBhl+9UGiJ/goSWi4Vq8mlwg4
8QupfnAaZRH3S187Zj6UXLN5XAFDjmXbwLKjftKgdm+qmgZkHrirR6ERHiJRIDDQj8ASwnjb+p+M
tj+BvVncklHt5BaBAGVXtuMXJQPdcQwBIGrlp+BBSCuHutg3Rt/QyHvIsgPNsPY/2fsKtCFxhszb
VZwJaPig4bNYXs4oKcviGtFdncqk38310ZDHlj0zhLHUkvtpvFwiiRz9eto6GOvCqxgl/UMH7TXC
Gi3ylwxkAffyCRxAOnjMkxL10ShR9kHtp+e514FRA3LM9Ow7HXYcvTEYL38aErnmwjKu/CbaMhZz
Zj5UFpzRc3eBCX5B9oClkKv7b52JcOgRB+gqmUQOegINcfYoY5zOXbK8+YQTmy8dhHuGfpbdlEfG
8sUEeCtLI/0IxdZiBG2Xg7i2RbMX5ujS96FOwK/h6AIRDNaYRw3/NRhlCSh4NwLaFlivd5BanKok
EykIhCKvmqolQeg/jX6hFzyOz0fo6T9H46tA6p9WkYuZMianDMkdBYn3Fl+ArF/wOw+9vY6oYc+2
214NjupObFSie76xzbOzK/ZKeyiFja2np1EKLc5uUW3IgNvNKiuaJla5FaX9uN8NeplHGcCaFjzw
/Do1rd+PEeorFJ2rbokR+sO8OTnzXZvHzW+GZEiqW6WemigqL9lV3ql54JB1jWmzxfoZ6qfML+5m
9YP4X+RCUMIgtNqS3ZQtMk7AUQwVP/gNigFRVXgy8hrRlfOWl2EcgfxUlMxkWdYKm7tUepxcIFiW
+5/mVFIW01ntyT5VNtRI+uhijPA6QLOt+Akpq8kBCVUQcJ6EAvNd9FnyfyhbQPLX4Tyo+vP5My5Q
q0Pz74ucQ7eLr4P9AZeER121Kv4f5WHB0PHYeWEUUSSnJE68vND4jLQfFSwIL4stqWSA89eCTKGW
adNGmoTig4GLDyCDRK61UPGxSwHlBsEAYItU+hkyH6/XzwiFCNJGAjcY/lCXSCqrUxyLDSh4dp2x
+NIMTGaNHEioaDYg5EKtP4rO3Xgj+vdGcfJvZgU/7q3mD3nFSy0NprTjxuSeeOLWCcQfpwcMhIuD
Z2td1RALdGFg5tLpKJfv7hKn857oSnGNWRc8FBAW57FRShYiyqi2gAmllHN/wLKAvnfWbzZJakYm
8DAN2C8nfumOrRwYUoZlNohTDLIxbCjVqQmhsz9TKIL6tbLxBd7ifnPteaL7uYaEz1Retv9z2Q/M
XwhuiK/zSGm3H9N1dKwD1yzsG/yWkyY9N/hXfh8S/vste6vq0m6w3cargXqFIWalt6jDMUr1R3lh
oaQsCmeV7PML6vu9yDo3jqKmcB2nHYz0jYahjLOsU+AD2r3xsIRebyyzFw+7pAlhhMpCJGbdD0Jj
V08b5JkCdzuBcSW/r2aaPpCGQkJu+aNNcTpeQ9/tSBUI16aWDgu25crW6NcCkfDzKo6tze688CDH
Hg4G2XWA7IQX7715oKiGbiOhfOljnYn18dmc5ZQqvIMAwAR3tMMcq9Uhb7/CJD7wa7DheXTahepD
QgW3w5E5f3ynkYSDypyO2yV+yWdsg0x77g42LEu69mSOTHDUCYTim8V7pUeyuvqHzThGz7UUzDhs
SfXVVhw3Zj85sdB2bUAfoX5a+0Cn3b8OoB7n821ZV01rv72QX8Gl11ESdTP/cXeBsSk68H9busDp
6YRATctu3gAc+SIEfOyAsf5T3sQXmcShZfYEqks+klbJ1O+kxmYRAIT5gRVDkaqw3HNbRwvUHAu3
Qz5GdubjXFg4zrl6Q4ZsQBge30chIXORrFTuImVFm/dAdvj79MLNN5AoR9vbJEwmOh30txHz3c2M
5xJE/r3jg3lVxmQG7etigMVPUdnj+DO5D+JwMP1+AuAm5tgq5UnhGf6E/6b42zLcLRIH0qMQJqag
Es51sJyY7tkzVSFDIMHlzyO+O8KUjkjEztrP5OYdVZshb3DCkvcMvqCxcvRMvMXG+jKr58KsdgZZ
w1fPt6xHAFXi23WzAy+jNfZrtlyDV0iEsGJlOAZDrI2b8G5NwZKEsiZeNWjDDIwimXaUrS7ToqCa
MjDeiguOlXYuVs/qb6Q1NZETERVKuYKlRbM76fG3SThQYQJUv0G7G8Ht4yOGXvlj4b0XwYe+indY
6bVSt77QW/fUpRPAHsAsUGQNV9T0OPVonJTypJZfdT6j6WWAVB9ii/EUFelAeMYqtFZJe1Gtt/Kr
XTY62VPsa6FLuw/4MfAr40joAymOgfGXaKZlLFBMplKULMLV++PDgjTCCOkOmL6disYPrzYY34EZ
900U+AowGYoFKRwZAptPOCXF01UqOd4co6edtjEEg9AqtGn2bfKf7vFajql7V6SABy+ALv0ofT0V
2MLSxyN5dYLSOemfM09hHvUAA+YwBCWePJ6I5UvSjZr/oZaJby4DHIFfBEQcEaXOzNsW2CIVnmpW
7bLd5KunRVGSArmsy8y7dLV8jvt922Lr49/z2oA3C9Wh441gTOhKtsusBNNcxyWfMSqv8TOne5Ab
EFpLpFdsqOxWT0HU2MZHkP+YTROaJVvQDpeb5KN2nDBkBKMfVQJLOy/ZyAap1GKcVUnk7vQP8Q0r
Hcx5QpXN8hnI9b4g9wrVfLC/PGJnFco/Rl4s8lSMxYN9SvmWMXnT5KJrP0mteytpYpG32d2pq6dE
2t0LCv1uw8s7Xrk8OR0TT/6UbIiIajozW9fISzdkjeHj0cIZNzi3D3dkTt0bNZlTB0F7/c4QGc5H
u69+b5jdezMyAMULraYwVyMAIQchYhe4Kfzvph4sF0ujGKyY80ZaM1jTqPS4JMNCLVvU9w54VKJ3
0jAeFNOGWyH5XanVYehjLUqRfk+zJwDS4YabChMqNie6ft+VUnry2jBD8lnY3HV3xRQGlIWanb6E
Ecbl2U4+amRSmsT5Yn7Xd2HkyUsij270Qrqkc9WaNXR1IVwiigyYeuUQR+Qd+Qicx5DrW8/WArYu
aSji7M9zKNeGREUJKMtCKYus/PxzHS5nd4301H+JAR9aYW6N4+QL2WKkht9u7uMGC6xPWvLfE4et
19VlmCSO4sFqdu9RO+QxCuGev9az2J8prLHebPv8P7zB/AOJwa38BvY7RW+Yi54xHeLKjYrPVfWl
YZuVskJFwrIZRtxEHoWMvE+SKjVX0NZdkvS0t9AkIx6EM+eRjX3tRD2TcmIVrgWx6aEOu5jsWqWu
GC48WP+4ZiDah+7MRJBwBZhOCPuP+7F2N8SilhD3X0KIz3IKBO1myc9dCMXfr9Q8NO+R48+lCCIZ
gfi8Vh1dsuxjqgFtW5xPDQt998UXQ4F/Frgb8T9laq3z+SH2eLw1KjErMv+bw1GySDtzt02dsHAD
5F+8ZtWs1PXvQqb9kFwxL36p5uiv/fmAczXu6cTIKx+bB8oY84BWraNK823uNGZWx99o7PYXTA9a
N0HIp7ev9TZg7hj1ktIsI/96dlHjA+WyLmPKjtQpQQJHgP6uugEgr3aWaqfa8K91hER11sXpnTKV
GMpehUgir+qKjU3MfR2zPXlyTx9845YJd/p2jbKPo3vxN1KAyojEzVApH3aHMHmPNBjgzaZcL2IT
RipJCtDTzRM8hdyg1voQcR5zCTMHF/7LxiFGzqgqWsInlyP77wBLFRJNo+0z45bECHwmhDP55sOF
9dmGDtR1nT/9x6DPS8JLraE+8XVgA5zNRuOq+FnyvOt5fCWv4ofTGrmCK5/aKZCUVzJDK+kmYPrk
807CUBqRoz1PxkBTrBOasdobYV+KdLzroDmyMyBtAz/LsD/IuWQjyCPibw0AlwrdZbb5zi5Mgywp
DZBIttJBWSukrTUeDs2Q7ypEUnB0B8G4hdEbwoNwmS8EltQ8pYKf5elrwLbaV6856ifwHInzQQYW
hVGRa2TFgnXqWY8HPSc59q9nJuuvefgQ3AHvEOrQY+XPzPHpWi/DFjlXRSZlyrDoFwh/w/AHsX2d
UtAVMMIKRLFprFNBaNOac7GdzUcb+Hn0aMgbo61V7jh7bPPeGJm8nEHyss23J1dGkSQ9bG1KWFz4
cCTPYn8Qx6l1BHNHjy5rjzzGrzWUXwrAFwE4TJGv0P85Dj/tMygsEQnr0fkZDNx9fZYjOwTUnXOi
1rWCvqnSHcjaErsMHEppg/cQWZrkgFk08UFEqIznC4OBcuS00mjAARO9uo5dCXW1pQ+mEnM/UJCD
Q3Ir95cG70Xf0DDXn72FSIflsO2uuv6R9KLE100bMTJ8ar1Jg1af4oB4Grb35X/en2JKiVMgabZS
UieTjIE97tr9CCXFBOFgIHlB8+BtqKAs7qvW6g7byOi/FXoFIEmbn4TRqbZXX7b0IPpbo6IOI4Ua
bVpWnSjuDfDKgeD/lVHvKEpgmFRQcMX0lP/xjSmLBpmK3dn0zSMWLe62rCWd+dxC9S6+Xp4rk/tC
qRMLzLb+EUgM7/BjYcwcC8qwvAtwDJkRruXA9jTMxav8OEDTSJmNIXtFeXM7gZcbvHu6zn6uVx0W
Wq3fphyVBc2L/z0fw/SmiroiJo70FBGWl2wPD1Ouc8zPfJosTMbqG8jiNUx3yqO85SWsxsXM21+e
nmWWDhEqUqHhlU+bTf3Qbi4qdjoMMaTOx12rDsh9sB1CD8iLKTREFzOYvfVEppiMW7be4cKZEJfp
zHv1pb/4GrJ3BGQB/KNlSmvcCaByXm4qZFTjPNtCS5kI829vjq1Mg8Vt/KDspJt8xzCRWKkuJpnQ
9dMrO8M7eiiRYz4ALil+6OtGZyMUHuOkmKI80+pfzUO65Pxg5P164IyVxlvzNey1gPnNsQTDH0h0
48NJzyPjmdO0rGiSHIO9NxI7OGILiXptv13F/0sLTtXx/5LPm7Z6Sf985D8jASfkH+WwdqKfEvn/
7Keolx1ISfO/u7A6NoxTPolICcLepHZBwlRL/9avgOoPAXfQqjlHtGN4LV2C25d4zzK9P+CBBCzE
wAxf+nVuL4dvc9+ghdOoPdPRMnoRPJZFAK2+iNbD7QnaczSeKRViiLpdaQH7Q9oHJ2DQ1BB4aCdI
55ooM5qHISldREW2YdMbuSG7Wap2iPAa6FGgOqfOyon7Je7awWJGxw4Xn0o3s7ggP0vbny9GdmbK
6v/207gClmbfKMwtnYBUjzDEoUEfCvQQFFcSt43Fbzhanby6nXHiIj2SguY3QQXPQi3bA8QUW1zg
QXHxQK/hRV5G7TOtKY0awWckghMM5md3gioX/XjuMySplPlGpLJ6XCOk73sKNgcV8JAHo4me+Opn
vwAywN4+vaILdH/drnJhA3vLQ3vWykOf/L54tM5CL4cdBLGbXXWw7SeczIF7jigpcm9YpZgykswV
fmGKAZgFTa8ro17Bsy+3+qlXV2/wkR9cJ9PbdJuZqH5lQD581JNf+B33YRo8eAMt1L48KHElyM/Z
b/8kcq8/YnNOJYYzBLLrqIoIZt5Iwe6TjfzZo0olwlJrQkdVDrauumIPq5wOvo1jyiLaSY4Kx21M
Fmw17pdRLn/wZHFLIyIFR9oMguFZGpCqYxCTKbrdEuya7+oZbMoWqwYsu8n6XclvxUbJx2MoVCOx
UND3KfnyW0TtnYzUZayXmCybQU79/esXePAHs8J5CnS3IeBHXWmXTdqCO/K+IjjZXFgA3JSWM/mh
ljM9ttfkiKkmHwRU+mwHA6oKsFsc8JnchdQ6uBZu3A3hXH5flJJy+maKTH4C1qWu6x0G1vCL4fND
TVaCAxsqJTuxATYeDtltMw0RzcaxTZPnIxyIkXIEk6qcJcXLjLs8ovxfevXKwriX6CMz9PL64dHQ
sLpKyiDVDEzoK9FZqyl27llulXZcTw5TAUm9mNlRNaEl5onTWR8sx3rZk5xJd6at9byHg69JkTGN
8D4V+9V0QYw5Kr4FlpVYpl8cZX0KTo/ggweyVRe/BN4Srel99a/J+iiPreUDJBOSFOrcdraHXcah
8ssctBnFsjR9uHocMH7XL7c0aw1Eghe9ibiuRHWqdZ25rQ80IDjteZK5TJbYv6iZUlLtPZLRR7Xs
yaCbdnQxCEtRif5wta1YLtw8iFBsIZN1XxFKsb4DTAEGiyr5GH+VZ3SW1b7YgKfYuKotfhqnMGGf
kTokVh07iSEZz/H/GMALcYhJWbYYCuzrCvSU/lDwVAtXnKH5cDs6+Atn7fPHWIsGqKyCHEdgnMWI
gHOA1P74TnleGKSIiEOKOXam/usbkSlWktRLi8fEVHLuiQA6iAQ4y166AO4Yqji5Bo2gGm2a6sQe
O+1Tw2OIY7luamh4BTpjfTyE/iBXkvHFqJkKjx4slEGfZQFMYlvwRpUAAhmYC/g3dANiKadTgH6i
uOmVzro8gMaeH8pQ8RyjDpvCQf1Vw5Cpbo5tA9a1+cO+PqoJnWcAmOkVhK3QDTy06eTx1bzvARCI
UE6GMvgUOZ47BPEy8TpSlnblOlfWacTZaY+jKR/jOo35gD678ZE40PbfQhbGI3UWlGs3H/Erzy9K
c7j6ymtyXqS07mTda7aFkvVeFHuZmwSPs1LshumXliwfy7U79qmYpgDaw6Prg5TiCdHgtkroRYeq
j3FRy2XErtSO50cWTO1Z/dRH+16NSECrRo1ynMviRaWphuhq+CcqbOT3iohqd1cwmxY0FcB+sKYQ
FMPBdU0m1sSD1Wm2uyAVjkdnMQq+f95G2VGKNVJjsDAo9jEH3PnvTjabz+37vIIEN7TXRrOeyTVZ
PGqdRJBiwvWrrSrnY3LduilB5wOKZv0bHbd16Pkdt1QzNEUgjR/AwaJxjYFG8G/ICz3kfbM64LHC
i3WeNaS+5KyTYlIENJByjW3gF6XjaahVI5m/urTegllDGvzKDpOI5lJtypFcjj2hXNSkgO3igwZM
m2E0ioBCi2i4UHx71hgUSZBcyks7JN9O8UcbOvEfW2xDK04l9wZlpbF2zP5kdJB1dk8Mjc/18Ch3
oAGVMaHhxBZ1huiMXyFDpWOQPDC2BiYwfHofFAKeCHmKaNxfvlcLIr4Brk5puTVd13f7S5BLaTAp
4shFsyaAdFi76/Y5Z3lg/EsnlJCYusN34XD1u5qBTmXCpg/kgSAPfK1fpwxVeEhpAE3wQOvw/lkA
h81M8ECOFtzwoveye6JEyAihcyvE+DU9w7hlwXI8t8DMSg9T71UCvAf80zrfiDz10GtYxs80bQaI
sfm3P32fpg756XXDz5tg8aXBw5/VCO+nyiYtgaHD+f1Is3VG7tgGiYPoXSv41dqqh8h+uKFz/2gP
/Nojlrg1O/kj5dTLEyWsTeJJ63ijioej+LFYa5jMO5nWWApe8b/+Rt+IqSIXD41Z4o0zIXVburU4
tV9r0J0PqLhkI21P5spMX79J6a4QvuMHwxfattjTxbGc/nk1IAxCvJ5fz7RyNUbnheuf9yZeDV4g
4bJnh7nJ8GHiwMfvQM6iYEtGjIGaGz/bGxWx7DamOw/x8N+JA34CqgFDnHe+VXc5wTYw1T7WaoJq
5iHrDVzom2zgn75oG3wVQBHkgMdzBlpVXpEfFk/jThgw5ovKZjngb/mt/DsibBG2SiiCW64bd78S
Xbso6HRkeu1dXqSgTYOMXd3/mWH/f8aWTqdZ5g3w8OZRXeNlbwmao5e3oCm3oPcUB0w0sSFwNP+j
PkjaAQ/oxY44HcxdcFpEj4mVWy1Bclq45hOQYRGsSbldNVMyJLaU1h3A/1ckZ+rrzCEre7Rgco8C
HAaSMrE7RatXWa9B/Y1/hp+QS8J+DOn4iwMUPhv4dNRENSNl6VizZJF/Ylf4mv5+5WIqdASidT68
LD2NpoI+7IzVSsgJ/D/d+lEB5+trpOG78K0QJDdrlNA+nh+PU+3V+IxySvjkW/39eACyUQ9aOi3j
s/rx3cnZlIxUd4Ky2IobeNZisi/48+CkC2/3Merrjjb1H6xbAT9bkGA68tcXtI/tZkMeRNZKvJPT
fcTvzngks0uGJk9+MBEKF3CtAJSsZkQDoYbwZIQiVC9NvFDJRpugCK5U9HJ7l2sHaXRoweYy2DVg
1+CDt5BEp0J6FdjaztI2IAq7wT1E+SI7T9djqSYtsdA6g7zKigJgcXHky62cXquGysa71Lu8G3o1
h8avVdspkagBg23LbXv2RuyifE7GhkIkR6kQW4VX3rcdh4dnbUs7cckVZv4Xx7kJd39P4IV+R8Kc
l19KzHo30IB8zgkkRmNKpsMzIy0jkre6L8Dwaraxf/ruQ/2GAqoL5hxAejwA5LknJmrcJvjIE7AV
9pNl6N5oDvg60zpEY6oxZ2tbDnpW1OIPChkZkkYaqKrPbRPQq7WPcn45O8pD4a/sXBqrvOGQhyLl
PyjLc9laulXZZL7g6bMMAHLjk/31LLnVkhEEb4dCaRLrkJoyPSSzFbisA6fQIdWQHBp2GkcM0EHi
q7wanocHfW37Y+E/RXSujuMBwvWGfu+0aFkArTfqPDg3W5J6hkKaJptLHEjbC0ZzWF/3Qp5ZUSXK
ku9Xw31MzmqE8Z7CFcHhBJTWQwNYXvG7LNqo6Or5BkLLtcg9BamyIt68DZ27DVi6W0jnykJECoto
heg1APdEbMbXQ2Vrb9Huti8OkO5/IxfOyZ9gaRqTR0v43ktSKeU+WdMCSU+M6w7Fe7fBRq8e9242
br4zGQCicRSaafLGFqI2qJMjk0PwLAG4oWuCKdZxh7K2uUvY27geeyDPNFMIJiAWdC6cEniMeLis
mYUerSGmp/qQlk0+gMlM1zU7L5CHLOpW5dU3MB54ixIbymYnNLPRNo6PCKjSMTGA3Gtv1ZbmhC0S
z1lItVlajEnOfoCOIoVNHH8y2r/NASAhhefwYjsIAWrNhbCEOEyTiuiSjb/MXJ0FzXNcoPzCp7pO
hcOx7WS2mcdy39YR9JLXYU5iIdiQO5QTDuIyXZ0qAFMSc9pESXRtOetlYGDdWf9D8LYQODrjCqS6
umf9djsXKADTK6ly/KckVA9+95RMokoqIxCeHDK5ww3ujEppeUqrCXaH1ZqUNHcojkkzceWxycJL
zVcOZVMd+S5SF/+BesOXdI9SFoQ3YdzErRXviqKYIfLZXotc/BWnpM6HPQfmbyeOcdDG8ahXFdTB
ACbDdbp+2vvZSxnVw7GtasRhsKpn2m1oyrMflVehvQNS11JTP877XLEOzpH8eA4kkkcE+KXPZI5m
j12q3glKkU+7OgxVGASXFMZeHqBITLVmH7RFfr+gXnznXtop4ZBGCoqhhnXvE8fxym8hPVWL/7G8
8dpmun00sZRCmrlz0MuSby8nyOUNcK8wgOsgUMsr+u6Ks9/pL5eyCJW/E8+lgNi1m7wQb7R92Dj1
aY3GGOZDfeH2JzzLU/JVLVC2DmcbbDO0V7TrcFSwBW67l6ny8D6Dg4+QhtAT7rqGQ51TbGuoQpGg
8T3FMh4fqs34BnDxbPhOWKG83ig18Uk3hExn5VHvDqSL0x3I/pvjT6sN90X3cfmVgJWS3IAuuoD8
aD6YxeIHfQ8zwEtX655uyYHHDenwQoDrEH41Hq1oKY8EcXXzMXaOyu7AmWaqm66cam/pprF5zci/
AOEIhRd7LDd2h8l3wOekN6BSNJKBQE6Hf4MJQ+a8q4gij1sqKzoA3dEzynDpTk8MUylqJ0iXcBg0
/MbIudpkgjemYvE8ZJhJ6CZZIg7SQ/CrlUKsuHNtlOz59fpiBPl+ceEzqgTn+EtN9rYFRXk3D8X3
MLd1KHZNErOL5G+hureMGrwZVkO7Fs9FH+ipnPoC2Aj5jzSapGqKWQnQlPi56GvmzlG1XTbTjIe/
WD2WvfIEXWrr/qXYnsezLPokLoaDMVp7rURHikRb3mN58x9PYOdQuqEwQ1jmt2QkJmDkb0+rHVgE
aZq56f8sXVpGpuSDXzCayemswsXvwJ3JzHEGZBETmUgTEF1792ZjBvEZWWBNdtL25+SYXU5gPwH8
2n9QIE3d/8ixjJccNqdnwaG0M3ADCwrta2z1o1iLb7lhs40OPMVy0NbkZV5QrqDxfg/o8d7eYUqS
3G51eK6LBFoOGXgWHjg0q7cNqSbMfKfgUpUo3k7pg+I6OVviphpugVXlqUjcibdy9YgKw5C/Sz0W
7gkUUIVVhjtr7t4IdGe+VfmIPXg3jZVzj3OVZCq/HoTtAGtc035gKVl3yFIVLLi3OiA7exg8pURB
KUuLe4pv3DEpRo9w/pbLc3IkgIbeCPqjYW3ulNSVC+ZshbAEJui2GcyA7Ha7I1POitGRV03yVPTQ
ugE0CBnZT4d+5R5NdUTlOr07RcXwNuvYdTu2BDVGQ0cydlrvE6EmlkIXde86ZTX3luGVGXJqJXIY
5IA5+sLxjAYCsOREaOXzbMnMdyGXho5mTjKll24qrG9WysAzZDDrKje0RG5SBM+dCONkMJF+lfGO
XFBu/pfq4MDprFgdxfWgb981XXfYxVe6y24DiHJsDpeNEHzUVfA1fDWyLCohA2gf1wRv8nxHD4/G
V0lQMMQTJ1LBmlDeTW3Asxk0UyqESEXjcQ5vu6Yj1EJ1/q2bu8ptnN1OdqFLgDOqUV2QgyvEk9Ar
mhcHn0lpRh+8GyKfGZhC5CWsmObENISp0t5Owar8FH4ST5B+qy3ncZihTd00aoweKecuND0rkJlw
G6Na3CgpTe43aUUv9qHsI2OGCTmGdJjfClg24Fz1Uptk4ZaYk3vYGGFieA5txaqwShJ9LwDLScwQ
aywNPlOc6k+9r5ljTeLqHJmpbJxYK32xn3dJANUrvNdCirtEEuAo7/HjDT134NHOfPy8GRWibXVn
P6Fm5o+DCoNlhDAefWxBr8ZCnd/P1CdwMHsJqnlxteWZG1Oi1m5olhXJS8NhVWG6b5Ef+oGTJ/JK
ki72ef0oN4cDpRFwRzzUBGbv5JbD/BMLoRzS/eiIEsczzrVmncRAGXNZ9/CXnUcAn/0pBMRfpSOk
dE2RkfoMyigglGyJIwjHjVmeZomtd6eX5LYkA2opYbrSGe8C+e8Ix4azlhNbbLXsCbAWttQCVbLl
0zAvXMfDdm2kgb3fM28v8ryiN+O5KU92ym6hqdcImcekabFZ3HTpxJdGpnnrxRSiz3JUbt5o6QDa
oa7hmnn8LYjkvLpLqGO6hyRHOC+zWS+P7u5vDpfaiCuKg2m3oNw27mixxreiXwVkJBX6YZWxVkfB
Jc1H43H/rz70wUKX5GJyltHMq6hKVtU4IkHlY/c/96aOOs69yUNUboX2s4YS5JzxH5eErBNXYTXN
2ydF0u2KjtQEtxAIiVVCWt+rsv0oFQjlQ3XKIdOBR6SPsXfe5FM9ncgA3IDc0sNoWBzpHI5pffmg
xqUPylf2aIKDL6zogoI24/8mJ8jODOq/oZ7bYqgOnjOpox9w4VT28ZoDBBiDJ1xvGHJS6cVgKXRk
UzCXVIZuthyyJSXWpxQccyrq8LGEe0YH4GVdq8V3OhrShbirPA/VoCNG5ly0Ku6hn3o3pgwWYaTk
P51vMi6BFM90XTt37WnzEBjEWIxV+hbl7ICzpLHy0HdIO9mofZelYraUc8weQvX/zcw2sxmMP4bF
LTMlov74cxFOWbd1bXIDdQlssLwzWJK5bbL0Yo4rCEG/Hw3QjBuIvoMnYys7HzdhtMTj6rzjigHA
/lJHH6wGNOnmutd4iREetxXK5R+oJXQtriZtQZGwcS9ZVqQ/swURjY5aAtgxchG2zBtnHGpjekGn
m/6jyPz/UpBeV528QFBOv9rDJreST/yErXNh+Lx7IRFWS4zeZp/Xcj4PlJ9FP850U9hu3f1fO1Bo
zR9bMhBV+Dt4qREgXEeKayFU9tRLxk6SCWdiXqiIe5iVLX/p8ZxyiyOMtyV8r44jWYxvHLeqZSlq
D4YoV20m8hhJMEh7wOlUh2MkMdjzR/6prQswPIttfuDNwkiY2IYUFw5hvi8DS6Vpk4qWFqpDUMrZ
zY+RxcC9uU9XwqROSrwfWsmRniZHSQDysZMN46TB1dwtBRpsJ9p55GX/W9i1Kd8puGQmJMssP2sF
C2a/+KjfZIlTVAHM0eI7mH6VHrOsnF60sld+L3a3Mcooe/xbXVROMqxDKXCB4FOt0Q/XSdHqmEkO
wqj+S6DPvARQPv89bkF/mo/cX5JJsY2ZItNGJR/gWEHvTRTfJTVmMpmfQXOyyTAiHBNzHVUiEKJi
0F3vj41ZlJoLMYvnDh1Ya3e1g3aH0XoiYkribXgZxXImjPjSfcFDwc39WKSmd0qDyo9/SV4wLA0g
Cn04lsv/zGpmKaNwhg8NgifpQV0l4GwABjdksVyfhS0sw/ckj0vqUkRR3pvLr1+e84eLhqjTPkLD
OVY4fsahfYRX7DMgTGON6GnAUaGNHlhG0A+P6e+kUa3N5PD5GMjkGIaAWrhpkvka1BxBoQHKamGg
dyB6GCftDsuHuaABtJZ/BdCUCuj5YleupdpE3FvVWdF+g1APmNOBXXRJRKr5PK9Uj4MKccM57wEl
1hSpJt7518Pg1+RL5Em+hHm043SuOxESgRnbOo/lsbn8PVllKVGQh8ibtlkB6wNtK8DclerkHd4G
V2+NccTUWwsbPJgUF6JHG7qLqIYuS/aZ0xwJA9XwDdYlcCck+yPWnN1r0qi0q2zrKu4QppLLyn2K
/+fIA2qfq77R+mYhqEhWFbZx/NvJVsb5CTI+rSyrGzm0eE54a7B9w4ISuUi51KcpBc3YvQquySV+
CjJgG7uIuFrKjTi/xTMY7sT1DnWgOBHNLN6/d3/s2fF4p7BGH5dVavMbUWDM3xJ4Kq1AbU55iLKL
Pewbqmym/y+aAufBIub2TqypVw9G8yRGS+mhd2ABhZ0a2wHVkLSeU0j+gTzI1DiEXhorUzpWv+Cu
oS8SmUtb96w5XNz0KPD7kPD+v5TZeq7jrgindqtyVe8gcupogAsxW7KFDv0ibQpkZcV5x5/iHQu6
ksk/xbkJFVpEFNOketdKKqaZT9HBDrD5tiH5Rm7Sg09Y/LZOV3lfQb9oyh8xeo8jPFeql+HiqpfM
G/UJ1MEPt+I8whEq3rxDvaySU53xUVR7gxh0ilQ+NKAWHIfY6zVO6DZsRtIAGsHmSvIi5/tzT5uI
NynfbG1VFGUTCkjGSrjqw9lI81IPq0D4TJic8r7LM3e7LsEfiz46pjBuNFiM5HPr0yGl6l7kRSub
y6n2j8kXpBSpAWGZW7fBu3Isz6iSEp9ed7g6Tv4+O+jaHdsD5yiW7GR/44mNvj660eZHhBLLA4hv
fsB+bcq8FnBNLyLVePoelQQ7oXQoHZ8c/vNen1WLyskdCBBHJINDnmKgJFTf5Fg5gEBZvvWyl51x
lU//Pz7aMb4vJXOcFki60zFSHPdB25hWhqRe9LOIcPjiDFLwg0N94PbA4T2m4nBbYJ3+GUjAlHsb
MxQqHZB4Tnprni8IAaYedPa7YHOGc0T1v+/DmQcWRSL1LzFLMjGZkNz8m4gvVbDac1nFYCpf5jXj
4655MOShCA+oXPhwkgRhF9mW/JcBnmEm3R/lVWnjap/07uK4/E/JOCUKd8roQVchcoa8X+JmGGuI
OYwirU+RE8nqfECMu5BEEFyLDV+B7T2LzVDLBGj4acBXY+QSpcyjoGFBqKLShLRBI+1kB9yHP+lg
WPJdZckW+u04QOKeOx8ubJav/C0XYczd8NA3HQpRUdmJO6DMSUzV/nH3+j/PNTUNvuUb9vV/qTKZ
wgT1wWXjYx+4728+w4MU+FVhCL8/SQq2b6cTf5pvbFek9No0aPec9kl1f0mfGT2pITQuEFEP0fD4
1cHuaHlIqRqR3CVf6M0C3woYMrAbCPkfRcJXt6yMFafMezsVit/UMQNdRRzjQxJm+jQqWtowIlGC
OApgH1XuIj5NOCXKK247M+ngtyokmuFfcGBaPFasGCpgNT5ApqrPF7V9ZARWUERgzmS5mkAlbEys
IJpvu7OnQzCqxIhzraypDoSqYsPgRn6gyAzobBaGVnlEGexR6hTvQwjFiGg/UmEvbZ7K330Nj20T
d7i2HHikIqrk+f26XhXW6DBTrvFYRg3krrCqIP2StO3D5R76BaZb6X+HBKr02I4MatBZH/C+vS1t
zqHZhCnnOgFhHq8PCQzUu0UQ+bpGRs3zhwPdMMuJnP0Yl1eZrVd/BvYm0s3VrGW5G12piORlNABe
8g0j2V+u7TCclBJIgYm2VesgM7oOi+4piiaq3N6mHWdoEnkB62eQptDlxijmlSCJHGm2xqKz8aev
jYLpe27Ndu9dedoQtHoNzsLIAUWE8u4OrXyOLnvfH9EfQS4T2TmSS6NQSLKHImc7zjedbEpNRnER
xdahu0BBROJ8PwmgIwD8zDB6BiD3L6N7NrMTgz/aLi5frlVt+jv6q9E3MCsr8hSdIgoOTbg0ww/b
5VV50Zj7aVdB24p/D1kI0VSPaCPedmjJSeN/1MaYeHCIUtMhBIMPWm5JTyOg5hDn15SCemTcHL2f
sDKXe+5QpOgtcT+zSx78E1gjTsCH6qKYT5q02yeEWDC01OD1pP9FhE0MQ2UbSA1Xod0CKGwfyYs/
BFjwECAX5Y1f1oFQvtVnKulpV4hjsAGsNWTladocV5fuEMdB24BfvhQJnoZsf8IVHZGRmvHXFxLI
OSa1Bh8FoZ+ib/uHCkEL5kyh/G8sI9nFOOiHdAF3mzu70PNBC/E9CiA8QJwdnSOPW+/U+BXhntfC
Wwoys2KYLJJKwLm74e8onZ5ZflVa+VCdGWMs2yMv0n2wkIoD2eyyx/VV53uReHMwXbvGRqL4hHDM
VmNweu30G3/juAr1YSB73pKzc+NSUpOVmfPpSQQqSmevM13+EYG6/zUsbaVEGDioVyAzytkzaofb
703Q/koC5lDkaYON2FXfHkgJX+4HLBmBf7Th7wCiE3zay9QGiDNMjljrG49+tFgSpkUogt2FhMWF
09hZ6BTzORERqRpOxDhQn4UiNF/H7RgTz4vRam83vQebt+NP8wzyucZeHSXQaQ4oa6plwtcIfGw2
CxIJGcaUqcrx1uIkoxpcnDFpmCjfJruZI/lgpC+fzKLfVzhcCPe7YEgW4yRvC36zsJs28bmNodqc
XfiZwVP7O/sn9K0HimX4X80YlOUaFWbuy+cNgT58IprwKQ7SiDawDygbjUCyYGL0xwca9AjAKyv1
h6ZOh8k85DpgVUlhSOWMUSfFu8qKFwhLhQnZ4fZTnL4W+Zv2UHxvm4DN+qpGKchGODlzJW7uaYS8
jbQwaiA6ffrze/XD+zhbfito1ZkEniG4XfaO4iM3NPxJP06bHlWMVMe3Gb9zBnDgXq8JQJt/uDVA
xlRS569rXfFxpl/0uQ7A9fQs4AITsWEMmiAp6yX6chcer+gM9YpT6BJqTBSiD8TuXte7igw4SvCn
EXHAFWg0z1BbmAd6/jP268vVEbIRTn+y2AXcOGlR4UZ2xmjRhk7VHmSxDCKxZxzL8SuGRhNzofds
f1Ipp2NK+0OuQrPXqUScxSoI15qYl0tcN+55ttTZ3vR9l1haitFTZhm8YSnad+OW4NcttF3VW00m
XiJG9pj0eI2QHFNHu2DLlHgR1FTp/NEeuaXJLSpH8jEGb5JpnwYv6jXSYRCaU59krAhUkhhidh8V
J/lHP+pYQSirW4KhNxi8p+MuQLrth4+v4fs17rLluQS+N1gGmUhCgoaUujoR3cXbuZ7s+zUCqGyl
xgdKWNFXHAQzjkHOXMNQnLQ1AkcjunFmnQO567J0jsir8vhe3/AODkQ+ipCNItdpruOeqXLBgnPm
tDVGZFdDjzOsWcIsvoEvs3ue+/6kUAFmE/N7ml5Ix6tF+F8Z2weEf12lCgd/oXq/3tf2jmoEkMuq
7UkNhpmeunGFDdvZCYFolB0lEsLjqpnwVFc4T3ouAMNErGLzWeEKo/4VM95ovYkvl8w5rg4Y6TXd
Ih5rcIC8M2Gktb4TJRaiX6uTN17GeOnS/0zsIyVajUN1W4lQCF7kDnUoiN5YoZAH2ceb6yXdIq4Y
ZL62oJbD9dM8T7igxpZVmOFjftKtpEqj01wCH1fT2UIpgo3aMdE93IArMOnl+gPawXbAjHyHX8KZ
VVPAJN9e33+VjK4bGTwdipTTGLrXTOoPLsmvIWcoh77iBjgkB84sMqFOR87f9trSPJgpv/rX/rR0
4M0I1cPzaUQ6eOocN9pv1kxDqVfKnTtguwbLjQx62lFtEykBt4+OMNgqfnxtLFSSEKGAOH43Rupp
czx5/ZCqNAj2x4VY6tEAw9HOm2+CQpEwv2YxsKcLUWBb44rnxEL6QKpFr0Qllc4r8WDSJRziWoFp
s1tV7k1MKpN2D8hhBDDYq/BTd4v3mK3BOei1g6uVVYFXIG7xy1gOCWDsTcqqQLlcxcLqP99IXcRy
WYJ082+uIU2jgQwRRt9qiTV741qTuz64rJQbw3Q0CmZWuVhqJ/rH1Ic7NXL0o0Tq1jXyKHMXsmpS
6E+ILziStPLdj4bYECn3T2TE8Uck+BVL3iqwGoONUoOGRPahCohROvXAug3MV3JVIdflYoyoPivH
sn1F2TpANaIyn5iuTuRYzPhliyDzE160kq6R6v3bIepw7JpVJdZ2yTghfY/z8VkK5TaiGtDKxWF4
JGa50q8Q0meYf1MWBsuAjAPqrskFA+iKBjysKn5J8yLl7k+aPwqA4xUJskiVHs5jbHhY9NvgFu/f
69FaAQ2RPLq3pB9eD6pYPWJ3Vfg1/BC3thK8062LpjYPRm6J/nqqC0B/DVbE5cq00oMCC92Lze1B
WQJaat3/JU3OLa2WRTLp9uMF73WMz1+DZGEVFcuxBU4Lf88shgfpBnWXti+Vk2HGKtq80YfUOonN
StOfymCpVE2cN6kKZECCQ9E0CwabnOZyLqH3SMRUw7U+yu4JQS0DUkzRyv1wMN58YeDPWavV9JgT
h6AKqSwKgK71XiPX4b0jAi29Zs0cKdXUjiBRHCHQnLKhJq4xxjeHfSbhB6A61u5Rf8OyjDfpyde3
8AlK+lw/Kxkn5+3AdpNmvJSjQPBTkJXWXykwEqUcIzrtfupb+HlouWECNGCAdtL94s08+gvqn5Dd
L+c/jwSvvdJongcAATGMp25oV2KlxpduV/wiZRvVKs+baomuiy2QMNQLlEO1UeKdzUpCUka+isb5
4aEFVN8kxCTik91+d2d2kYGh0zE9ByQ+1FGCkpA/Iba/0qm8F9qIYIHARJg4yjI+YBvtSVj2lGKO
nokYAFGMjABDF60MvYOFqNUAxbRdA9ug9nhaKlzkOlIdrI4yRsiI9Tpd62iwVCWyf9jO7vwhhu+U
aundy54aJlExt6WvYF8ULOlKiuPITBeFCi7x3fHvYSAMNE434g+xraIOdPwe7dmWpU4JEAZOq7pK
E7Rsz3BAao/Hx4wcltPnWn/cvvjcAmZNSy8QBZQr9SWQ/bj2+uz3cz1LK1l+EQq9zsibjc55Gw8z
TVOVciALwZtUeiHValn0TPW/OHVuHluE2/f9E9ahi8fSO2yl4r6jNpo8fuWjYKd6ESqlwj0896tM
E/NYJzuwu66hcEIDfIDs2NTnZuTwYqE6w/Ml28ZNOKbVal7bGedGAkeU40Z/EgkDojqCd/kr2nu3
5UpghTDCuWofByodo5ynMw1FF2lBurhwxwKofY1RONk7iN05sZFAqj2Xm6sjiKQ+HXwL3wu0fzHw
nnubF/unadFxaOFvOwsMVY3KWUnNsqMwh6nXyrbjbDyh7Vh6xFTFKAVroLF3iBsLzvs+RsQY2mfc
+RJ+wqy8PAwW/HNGhIBrOSvSUbNS8KWmXvMsyiL0OMVvsve/MzwA6Nrq4bIqiitaHzTJxtrlTGdx
T7S99IMuT+I/XtF4qtKN7hkxTAdcZZrzBgi5hnjNhVlhyvgMBZZ69JDfA04BZ7r6Vnd9OdFGBLjA
mWarHXsMhOR+H0eOrJBn9M9LTkvixa/ROr3BniLgiThExGbFI7Bk7WElCptnrEn9MJt8PtOzuivS
FbMZEXAZyDdMh/V6H1bbsQra40IVDWItNI1GbI/U8RMfxv5hCcrty1OOjJ4ZGdLFiwZISXXO2XaN
TGtT+/vXdocGjGT4jwQ2/r0dYxYWPZumCH8qqtwWO8UpDoFRpEZ4JHwHksDaaF8i5ObApeZfJZ6Q
tHfqteW2qIXQIdjn2ofEl88Qix+xIxylyYH8k8GRWb++y7n79/YkeFGQReFXtpP92M/vGHbuMvQF
o05VIAOpd0b6gKFcyuNtu2KZ5OP6r1gSr7DgR7pAZEmRUEiIDMQH7M7GFjlyOpnGwvPchOAcguzc
AAZPiHBhDgFs+cMeJiqIafuL4hGMtARZFa5ltr6ZDkKlohPf4gTN+jgfQ1DtZRUlyHkYEjUA7Uqz
WUVbO5RPbvS+K92m4yV3IOoH5UCRIb8kqF1PgCg64QcPes+n5W4Px0soseWJS3gIT5+AMYRxGxlT
PnoHG9rOF5r6a34WNp4EcpsB1bN/9viwBSRWWvZ3EEHKSJXO9JajTF6X12OiLPtyAlbBQj8iV0ir
75n9h506Zd1INznYot8KxocBFiwrqO6FCrJd/t+F+IxhU7P6C9+8yzBdGXi46R72beVBpDSoqzFg
St8E08hqx8HogEvvhbza60g8biQY+I5QxeoJ2RzRLkutBVOLB6sOvroZiPS9jFFbwDnPwnaT1Bnz
GYDRH5skltLetv8lt5Sw/Hvo+zg/goPpjyTTsJXrbIFQlRlnz7HSpDrUYxMpWNpzML0kdO8kb4IV
eSJ4dJGL7qJtgA9IathEVKNTRrbwNhmIeIroOYR7ck0CCM1Owi6T8iHbTM7fW1vd+GaDGLBFSS2c
uMOUeDtgeCMAN1wA+sdMf6OmnY4ewwjE4ctvNp/PKkAvKHm6L+RR8LJ9J0IO1O79QTgnD/X2zLvo
T5IUhcHdmGg2AZZiXNmSOIavXrA+2EBNgq6i6VQl33SDZNwf7hLyLrYBrFn0eIVyCGFI1tcAWbbL
IYWTh9WfeWoS34nXfoHZpgAlR9gdrdL6Y+Qw8PcDPEmFd7rsO1rPf35EBOgglLGF51Lj2TgEGLC+
djQt5OBLjtZc7S2MEx8xM9x0ZcAMfolokKTLAb3tyncU+OiSwlFByP1/OplJ2lpOrqGjYQlARHcQ
GjCVxAfQD1Na0vhRb4MTVEMkXEE/ijK/VIiciKaKSAEv7n+IaYYPfypZ59d0gsIPMj29nFYMsz2k
IjtfgdDgvNQGuthx7zYqz+/rTUrlRpTCZDgjwZWyCGycV6N9Qm8wdn3D2pI8Fjox/U9U44rDwY37
Buwo0i8Me7ZGnkq2Df2TIeIgTrPcKr4sfcSA6/sILy7nLDKc+86Ry5Cd9bxnXFsyL0dGknp9UqdL
erkxfr7RF1uJEd2Q5OQEoTgo63uCcB4EJulcVXVfz0j//XRQYHwNIMucOtEjiqgvw5alyecoiVH7
t7D//BX15CTwpIYHM8bChfkHRhKrBQpIL6D+BTpwjrP8Jt2uv4InpaDruNq3YyOjoi5uVWkXpFGJ
IKQxFxC4gP7ORQKJygXLQ01D5Oiq1jZiBQw5odhq02mRHjZgNawRYhErQXRJGrRrdZr7uumsO6sP
ewaN7F03mfR4N7h9LQd2HecmXE7vQ9s5z5DZzeEb0bVG9ah+uvbWayT3iixHeAA1ppyrrmCf35qq
+WiuX+246X7bS+94h8KBCXTM9aFxycn59RRK6Cdda67fZ10w1Bgqw2DdU/gTiuHpcmVtimvVu87C
48deBWHQn4H82tRRu1H9xDwvvROSJqz2qpaIxsuGO5W/sCVYbAkhrnYFBvDZw5DtCoMunD6NI174
ZFXwpYalO2wUZbRyki4TFgxU+RZSnvLHffu+OvB5YRj+5xnhWPqBNVILr8WDUKkui3xFOiQBvCn+
B7JWvnBot+ea4nZplWQkap3i/s+1gPrQob5B6qQUKUhg0pYqOpI38uuJmi+4KPaOVl5DcycnJ2kF
RHt70YPmrH9MkdDDtp2CREOKxrv+uqcqWV5JV5T8wE7ilYwhcoH8RKeVQmr2gH+Va1S1ntmqye4i
hRagevTcPntzWsRoO06wIJEFrjp47nODFhlFoFfgMplO3TPRTj3XufqfA/Ezqcuk7ply3bMT0gZk
kxcixV0SatL9weaQq0uuT/OtGqWOeaj2+2AbNAm7jeQ6aw9onLN2/kpxMpKI98vMQC5iRwA8MjaB
zCu4CTbMbHkEBVvy2ri0UAaO87GaQ7VRBToCfQHjoOKpnBdDJ0WkXtQgzJ2VKZKhcre8l4dy/MTS
hEy2MFg2QjgxMYXNvyckHMOyuyjGaRMyJSU0SvEeuBD/Nj6/GcQS9RE3pQJtLbD0NZLHQb0ZZInS
AFUHImv+TbfVJYLdmqnSb5ZtXGpgZRbabsTldzdYtHHooo/gvu78m//RhRaro8q2brSYFhuPC9bv
zicWW9qWURf9flBkD70IwfWb9xejDrCnBjcJEoowO6Pbr4ykGXM820d9YFrYgtMPdCrxnmf8j8Fp
I9iHhZlc2dW2HnPkEBGqwfQ8gFikM4I2Vz4MBwFuR0t1wpuIOhoqplsh985vUQ+veCRKIAK3Q8jL
23OAkU9tDaLgVgEXoqqhkSyrpNHi+i4dgUJPbpmu2FQss7sQq9Ypbf0HqjGmPX9PFHdI/rmRoJx4
4YdTcwcBjV+6bHBv4tHwPsL7rXxQmn8v67RiDvFhFKRFD0gbndheEAg6clLxqdjBOIPqF60vuXTB
DMmUZvl1jMNtwlvE6uDtDm1oIuQ2+gEp3hT91yhwxbvhzgkmqphOX+GaWOZcw3zWVMROup1fWdO4
tlhFOvi5fngpIqwQoXu8iCKv+GHuRK1jMTAk+aIJeaQ9mGiLXLsOzFZxv+9eiYKh/DJw3J/U13KO
ql0qd3DVqCltY9QrsoM3X+f/9CtIiciXUO+arKpnJW648Dtg4EbpDCAzpb6ykB4J0DNNGuyUnizj
FOdsM0vdjzr91m2zGWCcBAMpiRwnNM0SXEb2nddMuqv15MKoGxcW2ayO6ooa1r3HcXNQwwJ1pJjE
gpwVocNc8Muq0cAFWVICnrQUK3uE9eYThAu0c6rvgot1/hiRzmiyPp7iGxJjWMz2B47+VoxqbZTv
nYCtZu1xSmOSLezZYKXqyqQaIBxpj80Oz2O/Qmb8UGVDJXARQVZ5l6VYHu9ZNkRJjf/AI+ortdHb
f9Lke0/KIjo9nosgRo8gAAumJwBB6GRfOaTmF1u+rBK1+02wrq4C4s75SAx6Qli0GTrgWWPvFDu1
WyzYghaBTThA0XFRMHWrlCu/oKYeseGDUCHgaWRC73unBj3xHCW/CSMasMtTdAZ2q7UahLXDtiz7
bZzmzFOAEMoZCZbsa44JL0pPkQmWdXpzX73z45JxtaFFCZocLScecJGb6dq3UB6Lq6j++g9t8jWG
PaEs3RjoRMtA6T9/HPmntDeZQqEoBx4tyJNYfWvzms2SnC1D3EcrrRG7EXBUTsj0F6Gz1gmD3FRn
mqVqLqUeyFAJsudYM1dlyn3qq9vWt/DynMYF1jhhfUxemrybA1XVWh8Eunil4NwQqjk6OUD0HCiE
L4DPLBBr9ILPl3b5WeZmQ9FsKD92qT4s05O0Fiz+sBEtExIHAGXWo7adIDwG4c9XKOAsjTNJKC1c
8nfE+jTzThX1P6j0CTrC1u4+6aI8qvtDzt5nIXv0x1Ud1W9u81dMl+AYdPCUZ2lyu+D0l4gTsaAL
OoYrYcVQ7W1EtY1PJ7JHZUHWUODAoBcaowuwtQBaNNCTI04WG5cWmcbKItQ0htlxU6qJrArn62Kc
0amoiWQ5VuNZ10K/tefegJh6weEhrI9R0gfxmXwbiyaUyRdCzrJRhgACB4+/95pQVKc05e+LQ26y
T+IYVLbAVzDhDvxwoQXCjM743Q79lGBc0c/HpRjz2NKDgMiA/46R0ZI9xR6mB1QA6eFukhyQ7p5/
YY0kgivQlqkQRI3DvxP70GfMfz/LfSd72uyZuAFv4RsZVU0oygL5gWLYrYFIY2aKaBxMIq2rT9za
RWUJQLIceQvA/N6eY0HHIUAQGh7FJGtcjXOItrpYX/guF1dtkYcbfiRfLYjkkgov4Q6261VkiXB6
+afp/bijSSXOxL3ZKZNkGo9szhoEcAQ/G2S1Xv4tNp095XZD2/7HObrrNgzRy7u3UYJms8KETnY9
/VA4I3cxscd2b78+P68P1ZGYCpNlylKzw+fJ46e/Ink84B0qqAoBPsCGGXJBLzCK2iSOn4UPvya2
mAc7UmkDP23pmTUQmbE1jyDLFw0BocLSYyjr0/HKW08xAg98kK2AoItoXs9PCAXRY6dt56h/9UE9
kGbn80T3tQWFW5Gty9bv/D7xBGCQDe/cGj9BWp2H5saz1c2tSqm5nKKkFW0RL6D9TMzKLK9CqAh2
GLOt76TQM92IzfjTUKJ6OgcR0UKT/laWNqxyCbe5tl2aQHZOrU0S9Qiq4BPaPuZSc5ZvavPyrjUI
YdXDX8z8NbgzjZZmVVwX8H50pL4yZ3dNuwEI8BLIPK1HHZkeom2ZyxRHStGnXKjhL//A7qO/3Ers
/r/Cseh7EqOyvICbt0WHY2BxnviIu2xQxS49W8xRbIfxkShj+ee/qUULIMevCJcSbcvY4r95vmpb
UE10lK3z3GBmlFpHLUQd/FldNX0W40J6oXcZmclA1LpPw81YukmH8btv2vPdM7zV3BY3ceV752OP
MZ2w4YF6Vd4/oW8VaegA4R1jqseg8iSzSA4h4jvR+pTm3fxdrTqQ8BhglPfc6DnIb2SVkwE/5Sr9
4PiqSBJY9gi3mNgI0AHLAbTcEGSz6WQbAlQZu4FQMLT7DuJIPOeSxYXG89hn0kj4ZJj77lMS17fp
YkqkdG1TBdiLeipj9aWsRlVveE+sctgCCSMLu2T/ERVTU1U72wVsCFIvIk8FZVzkw8Ceii/eBu3v
VGML58bgZgymM3eUdxsu0t8hrODpHv1x2jmxY870c3/Unbk9+iKqYznJgIzpW2i1B7X7rjl7vr9N
1a7msqdHoWICn8RN/DznkkmIUSvhiY8y25B2D+pzuyM7AswdMJaA3By89NP1YPHJr9erFrrk/4Zb
52vY3mxRQGuj3TjGZgfxe/hUFvQVxIEr3lzg9HIpZV1GPMECvmdCaQkKUzFIawXg9PSvPKA8zCTH
qyiX8KH5icdeDofjYItZlZ4BKhtzyvPxA7xbF3GbZ4E8nzdsP1UUESUs8mgwrP4z08mGXT9TC7tk
eRB0kXyBX8dfJ/WuxgIThFOsV77NnYvY6lSYaygJ8jh3spfgIUI9LQwq82Wyx3UyktFJberg1A1C
LhNE4Y4N4OWjbTRNtBy8eYrMHKEV76oc6qXBvUt57OJiHgAfDJsnBaCK/n0WMnZVLrYjkQ/9fIRx
lBLmaSVQzIgehh3EMYzMt8U2Q4aig82pSgMAZHz6jcQpTZyMyGTSOXsNpJ2LXPPS9by1iDf9FCiI
o72aWS2a9nivzdoBGIpQzNp4je76bMsSLlO7C7cXcUZXWPUWpRJHuL6AYLyQlWuKh/UGdqDXmGgk
CXDkMiVTgyOEE+6JzQkpDT8XCoZZQDNDXYJqjp1UWJL+SMDJ447xsp4ML5P02JwjLhhU0r98GfRt
9fevlQ2RxSIwhUxugBwsZFdRoArVUwyYKPiJsBhlGpuRitz4rUX0FJ193g+vWH3pUoaBV0qMMgdn
NPXSAbFzvGl2C1zYFFAl6VTF5JpnauI8uqYEn87qwrQD5n8CiLCsNZNaZMHCvbRLRN1sptT5qiKT
vMHZjfDPMYELRFhX+HOEbO2FaYbppD2sRvqPswi9lC2uv8sY1OiP32MsIYUhOnAU089ulcf1wnYx
1KgyzymrhCRTf6omv3RTNGPBOCt5bPRRnRUsMKoJJkwwA0gWojqWdRB4RjCU4LpxVvfKJDkSkbLr
Kgix2c78Xlxl/6QMFdxhv2nFHpSkFAmrTmiK1P1vC6I3rTUXXKVxW3S9EsM9iUeV3rVa4gLciVF7
354F+IackOa6Fhl6jQ/+TK5lyGKsC/7fll2mBymKo/axjNg7gE+Tj3pZVb2q97Jp2y3ilbgQZPvy
PIEqJs6IWrd8gyRvIfpuPnD78O16yEi30F6AzBBtU3yuoBsOlFMdqqACIBcp6oXWh+VX43s7JOzy
AaLzk8SIWcIo7dG9QaTFX4lRRBiZhY33bFqrxcw2kFB5hlJKSFuXAeUV7YGWLQ9sMGBpr02NStuf
mrT9oN8i4BGyvDZB/FA48B9pns0qgHlMpxaDQo/CsK2itSed5E5fltojKYjldLBwZC3qnT+RUES1
NsnvTern8aOx7DwhwBC7AK2RepR/987cHk47uppEgvUsDc/gXuX0M1zFapM8peRh4Fq2ySlfxn+5
CWbpikPCRYSRqtdvGltaRoz4mOWXst6qi/jcskSLeQ5UbFkxafDTiIeJJu0265+smLoeYiQ1wmwD
+31C1dla/SD0Bznl1zAOesLM9+ylMSouyNje6FqP9TL/+8N/mqiTO/lOKjA+zyO/Nkn6GLEKzkh6
FHAGZ5X6x/00XYbnHOniUZ7gdraY7/fDuzooIPJRgjIdjzM66jWrcvc/s7FYjp62/5NFh/iWkTI8
BAQtrVo9bdapU4usDxcuhWSLSVd9ppy/SBJ9jOFI7eOPAAUD6gjXjFA7j1zz13MBkTmT6ksk4V+V
geGGvKNv4zhedrrYUcfQPrnUnwVPd2FEvwhSALkzjj+BJKdVfMeVz+lOk2xARhNvka8a015tI9SQ
vJHq+Ve0OAIt97xnMbIRX07ahbPxHbsk8r9gd1blGkQdEhpYjSbDIeig1CUKi/5AvfNWK7WdeM9c
236MbKcWLztEUwkaJpqbacJRsyPChqB0dkS7e9xUR3rhuB9MtfTeS7QoOTdlLUFMsIVtaTYGhmP4
0MitkiAFsr0rFsqEA6eOS3FHBV02JwIySUafxgAgqlp5gvHaVtzOePevMGObGXDq7V1mrfn5HSCo
mcLqR0rWSroSNEZgUKWdWcLh9fflykCt6WQYE/3hJtMqG8NzN5egmskspLrFmN2UovIH7RZDg2bE
LXLlm5IvY/DdZgzFxsbtvXXUg/QLHMVueVizaMzu8qorXvwsRnTL29wh1jNIdTH28B5Dotu2d+ct
7PNbgOMzaBPkWuUNBbt/uw9uJ7nZT5L6i1RO1lie1QUE9qL9ix6pYKwIhN3AzxpqUR/DDOzljoW1
+fNLOXU1AhSvfQRTtVZ/gOfyJ2LrYnm7bk6Ypct0dqn+R6LbF/h20YseGJfatDB2Dw2LPl1z0jQU
0G5oGa4Lfx50yA88HqNNfW+LxmxsWafUlaMEdmX0Bwlrwvc+JEUE1Sv57S+2U2Oga8We6PwRJwM7
B/OtJfEzCnwB0pvh1RCMnD0k+3PQuiFMS04B6FHd+AkKEp+pgGiaZeKb4ph5MOl7i2Xoun5Qdd9c
BPKD/YcynDOOU1RW7bgLRadffrx3TYz6g/GmOd2dezeLuMda4WyEtHAvARvBB3d0FBwF43d8fdh9
cqLrjFunjL1pD2hfokvvsZIs7e7c9fu5l27IR9mjo/U3l1Vkm5XtKvwunXnGRqgD1eglgfrvXYRI
lMis2Sy0WZ66OJ4lgIhy9a4lMixnIzCSjXleGId3rJSVqct8pmtrHND3D8kJPu64YLSiZmQR9/rp
4KVMWJAcLdhEzdtmzJvyk2mlwK8+oyFjfzttdN+X294v22VCI/vlLXTb+36hgskzGPc6SLIa8tWo
QjmE/d0dppxgsiV8rQDh1GwgbOVbAeq4+vO9sRe243m4ptLka7t6jA3se+GB2jmRSVw848XcQ9WD
Qa67P/qzxQg6UdU6SUtWBiOjJI8/6a6U0TTwR8pMdGmY8Mnt5B49TMp44QpCUFABl0xfRTGlTiyS
lQyUDVPJnEZtplNpYqHktKj1REZuxW9aUzV1x5n6S0qn2nr09vlJeidDGfRDjSnooebZS+buOT86
5Lm8ekPHaHemz6FkHiynSYxBlhaiz2dMgvmqtfdkAYY1Gk8VQlrz1SvOo2NPfMpHnrxmoPn82Fpm
jDi6Suie6bfLTUhLo3mZyfLTjO4JsN2V8QjT+YlJNcocIlzobj7bdJJQRK7SSL+sX/+pZM2bO24O
0Pn6uwAW50B3sOogYNITOHSkouIXo9C23Z9iXjov5HOnLu+apL0D6X6N3BDcNg4CeF/Ccdohcc5/
FCWHQQWua+2Y8J988CY8ehjH80zAiF+LQjQ7ha+aCgQo2ujGMOAuSxfbZn1bejw1viVGTmcqm0lk
vwMOD72Yw2/JL9MzouLY8R8M9kB53WMG+EZqfsjLThUvuTWLfvMBrah+rCgCu9P8gNJhKIKdwkwD
k7xHVv6JhnWY7QLEJTPyaqERJEs//eydXJzrHi2Me5quEhMWW9Re+PrDTBOOnv+F5cKgaagrd+6J
fVTI2vTB7UcQZiESczX1Qg6lAk0tBQwn8QBcO/CUBjPqz1BiwiblBh2CU6HsxnTOH15nZ1ADeG7z
fESb4USS8f3aN5XKlpmUtJZlSndh+jLp295REkcOI8a9Jgq+798UIGNIFknDU0kJp831xgO1pzOe
gDaB+4IhnIJgPT/BnKTfbHzi3xb1dLM7Ghh2xLwsnVX8CQpOnMuTbE5lmRnkxw7Xj5vhA7ELjKu0
P1IhjF3cmhB4UKJKyivPFM8OwpiqgCsBsRPGJKhVJyaqqTHWnLlI2Tq8wIOjomVAwSpXGSmNUTta
jw6pI7QM0M4mlrDxSBfCxtZZJg5KRFJgS5T0vj6qqKcc2npbf9XYMdrrxGNfF7u0vhPqxnvYd7hd
LoKIHBImf9/iLv/+e1oXAqaV7O36B3krqBYYhe7hFNXJz+npt8eE9S2XBgC31n3MKbRzV3Wl5YlY
unWTtmoz8GfTt6Nv829kKgueB/tkviPJvCuRycdxfdoJpJV1+TNQcvt9HETPBrLBFMRzM2AaEe9H
lMkJqZZjo82ltg+PumywILmXBSwhtP6QL6PY+oT9rn/1v8HNJiTk9CJe/rbpCQkMDb1924ZrQggx
49BLWGEBu8WxLQt+pG3IunOWwKVrf4Up9p3EkK7QK/Ag4zTANMMFOtujMAPkGa4WNL1+h/kdpP3N
z1ZUAZiEuIa59oszvmkZe0G5ywwDOlYhITKbWfHjnKxZh3EbXEf2vxvLppfiUFxkQ986hKr2eV5z
sFtMiOBEvbMu3QykPzq/8lvHin3RfQqP59M063IWjol2zW6lqx8Wk5ux6AqJ29qgAHKESm+YPuvw
KkitMjn6P++b65MIYOVp6AySRs5HQWsTqwiHGy5bY0FUKnOqli80cwwqGKC1FpEHl2rt81zHMtAi
45PKg4c2Ge15D+l+KdpYGR02YFi4D5A9jeFeN8e8Z56POMkXnrGwaPEqj6xKzQnyWxakhGMZhES2
YLPcCl3rYODv+rvwTv/2JOPdenkwBYegDU1Rarv/NotB/TAbOwD/zJ3Hrc3BbIadvPExJ3lEzeU4
zmoREjit9HtIyb0LEB/YdosfyI3QkLBvmQYlhrWqYa6ZlAXkeditOxQcln3vTCIa+cdzhUVQnlYz
P/LfwDd4Z50QI9POhDA5TDsC9Qxnk7Wb9TsU3SsVd9T7PgapCKZ6WXgfRiLwQ04aGuNGiFK/oBEs
rRt4v+Xa7/Wmy28VNDXfURa+zCeCDAa3+WVzpqJiWhYZm4bmRXMjhCeLFxHLrrhyg5oZv7WYSyQY
yHO2D2TaJ0bmSre/ei1EHGnYSi3muv7YMXRAHbkDgX2pS4xc8c3VEU3tkDNOy/YdoBXaFBdvo0A7
yJ95QvXhRQF41m/gcu18aZ0SCI+nx4hYiDWzjDozIlojyweZcbrEyL02YZ/zX05ONZdZomazDp3v
JNcftHYoO/vagkE89FL5jLoSV+5fYQ/qS2Ai0TgrZIwGjQaz+XRaqmG2Sadfzw8yphl/Ke8aQM4B
n/JgTRdOsHWtzpWozjbfLhmP+d/y9UM0rMTeODl0rB34NpoaKYtVQ5zJjn3in+ICd3x7USNjTYxn
zIPdGmkfcLeGSM5Upm+hhLXOmA7PtvOFTMxL+dYxZoYjAgaIq053MATPchlXwf4zLtTkYkHbLen4
LRDXMXhq7A8pn3pSSAl4v67I4+0eUmgf/G/BK5x13LBanc3SK7TRtyQ/sBiQ5+I72Je+im/SXXbA
tyzpPLBXmX1zMp5HiW3LEaT/yMr1Jxu/8fNmbnGC/61u2Qt0xsOevuegf+eeqFfPKMdHN4Xt8D1Q
UHMVxLy9b3WvbFayQ64M0IT+ajrssyZ5XLmBD7KS1Piq5d73/zMm49OJjjGbt4WriuU7YN131O3H
mwKe/nZptABo+Y9M/Sl1SQ8zgqLOAwi4obzHGjDB103CyvXsun+iogUSg2EJqc0ffMhhpOOnSvY4
syQko641ArxRuMbX/Fi2kIiVpbG7pIfJ1wuTZQCd99RmKX/InKgFm+50iv6P/Ha/uWlwDtMT8A4A
ngNeE3YJZcUSx/hATKfd31M5bT+zhN334uh0GXf+/UUW9X//yqScf+OObuS30pbiVlAHqsf9cvq9
CMDr5iZDhWxtyHoripIO6dSi6ufYFBCiW1j36uSf9NM6L+69+whnmCVzAhXEd9T1lX8pXONdn6VX
U7CL6FEnCSEONGNjvXq/xWkJmm+fn2k4hlC/7Z/x6copAiWsGlMWP+rMkFPFq5bDZ1VZqU9rchHt
MfqClZpCXn7NqyhOCZpnMh9H+0lAPOP+FU1F2y9dJ27mbIATWcq2SKOiQXlHX5O9LcUwXrWJlocR
tOwtM9Ux7ok6WegxlWbPluRi3X01yr+RP53HFe7Fw94CireqxjyjZD382J7NX/C4vqAXWc+yBOgP
00Tt9JE4VFs8DkG1WWImgUnurxCKkv9Nt8OCNl4Rx4+y5p0WlBKeGiidJWoO0VseD3eKRrHQkzc1
vDpptfXyvGjD/Lem8dpw+6SRWIj7X0Mew1DaeC6XvgWn83H0dYknW3X1Zz8pPCiYr7HtSHN0+hbL
HTsfIMoA5/pGrFGiDbNkT1Yd45xoA12t1eFKz8r0rUK4LLDVwI71oQ00YSR+8zUufwngp7VzA8hf
Mc59eRD+GMpTV9JsNfz4x2lTPNyRxCSPL0SlmeI7u5UkLPMcPrBdZknmyxtK7vz/q2ck3KUpH6tG
1R6rshkUVUmbqY497D1Hi/rgIMGQrSorJ89mWq4I2Om4gNYDKDFkyX4xX0s3hizzScx6B8DlVWKw
dXDzpbvGtBRqYB/jS/RNOWJs/SQkig6yE3Rn4nSt7EDotJ9PYnIGDu8wDY86CmMo3W1t/67TGY0r
JMiWXK3OVWDDMLDIg5KXps3bS0qHpl/ut2gp4hNLzf0lGBsIg97Kj97xKRlbkj3N/dFHMnI/M+6f
+abCMDONHh4ykoRTk0tBlvqAtn0A8xGhnZRx4ygEjE7HyA1ceWCA5+utS9AEz7e0gKH2OWjhZE3+
3vgWWZBsUETLMfWA/Am3xlb4RcIbumEyqm0Tas6MEVcUIeP0AaBaLAFYccu1Ss0vjpaB0uFqxMSp
DG/sDzV7duL+BkTLzeVcTNbaLmps9i1UgCN5JtzCOYTOjFOW1TTsLYbzFq44s50RHwH9blKmtJal
sZRHbf/Ceze449dxVwG6WCvHe7H41uZNQUiyoboUfWsNF1t9WwT3mxW30XU6TIrFgFigB+2ZtGyr
QPKvjarHfQuQ/fBKnYnwian31tG0fuRdhs1KXjkLNHomxyqokBNNq2+bm/TjsK7LhGZSDZrnsXWX
55HZejn+Qf6oKoEz4R+wNExjmF07VZlViUU7jk7MYEMUtYw9ydc1zK/AWNZETr+uIFkl9GNFsePj
opfJ0OoQrp85+BAWtrUkn+UGHx8XhEr+0sJ+Yr3u46cLWzLmrNQ9XEhWg9FajOzgRUMm3vbPg4m4
qyTz3Ph03i/FKULrRP3lcFYVckN8itr9TaFD4kD38NxXMxdYnkZEdecNOqmSNVHXKRPs9MdU+Ipp
Cuwdja2k/Er70xQpz9cuCU1f3Q/HTvzHkjReMzq1J1djv4TljqU0UJJ9m8rMdOjayJstUr08m/Q5
6pu+AjLba/TL15dGTo8Oxy9PK7RuMoO7P0Mp0KQn5DzkUvfePZcg1irKGD4GXAkjPG6vNDyjuGCp
T/g2T5BUWNHhx3eNovvVJFosrQawYqd4+jHfbcFH4FWO5My9csDBhYZqAQ2YD10s2BfJYaDjIirW
Cy9jRc8h9v/r1ES1yPVZPD06TCziMYYo49Mx9dGlKSWA6xed/QhL5qLKEfrMnC/SpAzwrZYXfaGP
zTpWP9M966YAx64SQoCZLg2bD93dnSR7W/2kHu5rv8bIgODLiznPwA5BgPsV0DBYyrdLG3DaqSvu
19lkXnQcTXtgoZ1WpAutm6coivzOmCXF5HT1EJpd84xdjGwZbA6kqapmvsUq50i1BUwRTHEG5rOE
jq/s5sRIpwgDeqVYh8ldvoAaPaFzIJ2fMxjnATSBg+aDhP9m9zihgXEzep7o5JM813N3PcGMCs+X
pc+7Dk2PAGCFp7I5+Rchw6wMIbgaqL0IWA3RBfC13EEYhGCxDQJv+aoZHnu0IUrusb8WGNDk5sFV
FkIVpoG0MQbVRF1VHzJq4OIMRQJupptOr7LWk51LD9lTqdgm89a9lEDHdeLXCCS71ye/GgNzmSP2
aqmpYrtFMjpyW/4aR8neHlpOFNjPUq4AfVQuIZ52JS4I9dD09xCKLO9wC+Qez3dw3/uDigOcdB4v
QciaGrKbWvS19MnGsoDkO+SQRceWyPi/b/tB75RpIG5ebLjPS3bxmOj0t8MCAge8d+L+dN58a00v
1YRMFHbgVfFkrpFuQsDXBJN1F/7THdkISgXY9FJitDkUNF/CxNGl78epOAO+C0JZ2MPrWjm4IQNI
WLYKTBtwYUlO9TF7LgEZqST9l4p2xDaukE3C7bHSM6Yc1nhSfw7Syvj+PKyS8CndcE4+CySPbmB4
izcrrORuvLm0usw/s4kjfYX7UjcBhgirbeaZQk8XYioGXhoR0Sv1QUbqC9upEQslRapZCWlhR07X
+Pz85vdB/7D+W6j1aKhk5NYoHdqUgcYMbqm6RB32zzAZACseHTaeqn5i3961ibxSnHweoLnQJQ73
yyXD+wOHGG3Rj+1lxzYOLojKK7MX8xPH6JKG2G81TuOCowbRoJKFzSAq8lViKe+NwdMdBg+jPEFN
VyQYSXPDWPVXKvv78ne8uRKq6GuRdy6bULWvZV6Wt1/YpGwIbv+gZmT0ErwodHmrSILGxx55Tgic
z14tfuIwZHvb/tW77H9pybamrEBouMWNlGjc7V8utngBhw0wLH9UerLgWskHuR7HP3MPyO96mvbu
iFlSwceOn6RCylY8S/uNbKZnU1vN6yP5OuXELcpZOQ2WEHhF1bcGEX0r3u9Qquo4fToB8kNbT3kU
z07WqQ3OWCJDvK6DYR5j5n4heLW8PgkV/yjEOcXFrjrHfmoI9x6R/6Zf9kLd6WjiGPG9v25uQ/P9
bNcw4LKNMw2998mB0ng1wShovU+/SBvIhCxdbmhNJ0ic1Y1B3xS9cEzJR/a46b/NqOKVFjYM83mj
gpKJPADjmnUcu95nhy443Hv++/JCrnPq5QFN8xU8HrjUCbBGfF7iCVrzavqmVXDv65sxwYQY8+iP
0jKnbWs8I8TXWy61FIZkg5n1f+9zZuq0x4Z5AAzrG6JNxX37Ukys+f+wRzU7iozgcGaZrwRt//ne
o2gAonaH9ejl8ScVhkd0S16YvyW9vossMpOWEMWMfqEH0mmyKGKScKFojCf5pn4Qv3mY2PUtYmBB
x5mCQT3WLciXnIhlLtCJW7RvUK7YFEXvulnQufu3GkFDcVYNJshlnnsqtuWrxNLGn+jIFsPCYL9C
pgbz1Cx8TyI1Tzgg6UpbMKb1nbdeYLxCOlmiq/U51pIAKttxsREIC8DoFK/qR3P0EDaVO/Ph8vMk
WQ9V3LIgYo4Wnlmd24AWe2wdWNAQH33MD+F30k+uka1xJzwaC7F6yo7+f6f/4c4NbGx9V8YLXk7Z
EzfMgUKYCpP6ZB+y0t+i5s5HX4cXXXP+kngvO8DKZJeNsHkZ+FzAbbIKtmwOMLGpPhUpTyyIqRoX
Q/+NDUCr8Pl2z0xNmi3NDngfyANbCl4gCGIjX05zsYCOmda8gdWUFG3XcQzOTdxzt5hAHGJ1oKfH
bQahdev5Zs8MqghyY9xcvK2fLs4S1IxBlSzCgqnkFv1A1zWGfqpDE9YLvpgvfbeKrt1sANJ2hZqt
2l42ll5IWOE5bGYWVKc/1WJUXIfLvQ1Eo76WEXqP7Lgz9xN7zcwjxylO7y4xKSx+jgdWxVYhcvL3
ZPUTUBvqA3lHGsvUEfLuaUeodKCM15FHCQ1qkcgmlyETzchxOgeBo4zznijYDfkS6znj2/AYY2yx
uiqRZStaoBsJNe5pBgfrCJB9zo+MuBgNFrhVsyNCrAoENOGmGqt6yxbeLN8qwg7gCWfIOgNHtscC
5X1JR+tZWhM6LN+pT7iYiVy+MerCA+8wzujYm9d0C7tUOmuGrS7hXe5sgdJQzJFQB/Y7FLT4ZRiJ
79zsDykmqRv12iGAOriF7VeRYjvvhpve2TrMlxR1kRsh0+MzPRfrQnx+IAk6K/ji6C5yfgjoZBfN
AiRqjK/TvzBtjHqI2pfj6v4LfT8RQXVnK3bPGw+LUUbJSHrRzpazdbB75W4bEjfgOpkrRSWlsVe+
v8t1TJJC4fieTxwfZ9TbvEgieJiT0WOa5bRujntl96nihI1v6hWl5TlA/eebNDsTbieIp+zFvR23
x3+fv/MjHExsICqHR6+99SjgivVgknDVXuIotA7zEuFYhB2Mu3wyIm20pW6ftuZUUBMzTNw+4v2I
agVnGxJEg6ldejqO4wXDW67oH45OgQG0tN/Ed9VcyWeWa1uXCyTqVdj5y6eKkh5ND7FM13NhrfqY
VNosHs4ZRSROvSfihKcG+rX82kp95FwaCyrt9OJ1q3Ci4tZcBAHPq/pt7J7GUjzH8RmXXbiTFtJ7
0ZzZTCNMbkYUSOH6ps58fmLfKa0XCNWMcAf2iNZAB5VQF9jWdOSa7g6XMQ82dBFAtAJXt1Rn66fJ
muWBIa3i9TVHTYB72KrcrsPCpmyKlKQhR4sEG16rWASsqmy2gPa1bFfsvddCRWIbWXzU6jo72v0i
5u0llDGiIxl9iBftuMF6FoOWkt8FPBB3qkTYvXV2l4b+dZtgrUA2pZ9Ql1Zl6nAb1m3ho4PIws3S
/854dC5cIGKNcJzI611qJtMGxnagKeE4C79Tx8KFHztX3/YJQTmmf6/mYu01ALs94mF/LBeGdDbK
7GuUapmVDZgzxwQIAJwRicIfL4TVcTKi3rTKcJ/hFCUEC7AVF37GijWsGDLvEkz6ktw/ujntPrw3
LIw86S+cjJZlB05PIxOPdlWEStV3C+huLyvvgQ+mOAeP/3/b8NlrqgBaEJXgdFydHLh8ve3azlf5
eyTc8MIJkODjKCNP0HK3trdMuQVTMbIRju86VF30k8CmCuP/mg0Vj5TzbcwP6bjcicxEYCEeX2SY
XdBzZpUN5n/9JhmmKoxpK7EIX1aAbZojcb9Bon7PRZ9Gfa207gpwLLsRnDPWtMhB04ka5KVwshvp
e/vkh1IlBZXydpYaLpVI0+R0ierydRdXVkf/evvftdWLlIR9wed1cPckwoZF7BN3HpBCS9+8fBX1
IDo5DIC5L0Ychp8uREqGdpKLuh1N78Qm+EDec9jOeo07qps0oWLuoogFtN3rBN5HfD4Fe1cvoSF+
SQWFhYMdwkZD68KzVfUmtPenNfy9ww6Cmilu1h4UeFGVgTCACspNt9iR1bGe++6yAk7xAIfYHZSu
zBoP6yNXcyI7Diy2m7cT85+9PlK84cymvsFFtwUapiWrHRLPwhqICzec7JyCpE6Go3iKZ+osq5iV
a579m/3BtYloSgdSzvP5px9HU8YWkKtf4Fr8KXMxkiOTnLr5zdCkOqDFkBvVO/HgK7tMrTBNrqha
872wlIDT6j/9o7NZT3KzR5fNsdBrJ++vcE68an3M6jlctISyCW0Q+MrckDfGc5Q4OXlob27Zk9nr
zAVkgm0tAbwWmOk6RAuZIUZnDyAws9X6B6f435nTM0bbvKAmMHajgYcxilKjG9u5rE7gGZSx0fLk
LYc+n2z505brBdh/VgKd25LAw0InIOntknMB6ff73P4/ruRi6OYfMq7ypoISg1W8UNfCCvnuck2p
qHLSbPT2N8cQZ48ws31dilDoE9MRldVEvI9Vx83M/g4wzuBkSSKXhCOj/TcAbFdD3Rl9xgss1Y5z
cPTmGdq1UOH/E0cHgUkzQaEBDot3jQYGcQ0N2MQ53M/W+C4fxTIznaElgYd+akvuJdNKEyIaWhi3
3s3mkFefSQ6pwMSNeU28NhzmTOi3tNqLcrvw1PGN8OmcpK5pmFrw5Dejsf0GOBIuZ3xCO5gCd0xl
TT3z07ppkzY7KWK/8+xjDsV663WA3GrFVpWJWqvEG4NFtymQpts9ydIbvfC1CVjSVrrR1pqHsfpV
JlUv/Tmzdb2NkKURWBSM+Qe7CvhkaAqxiMn+n1T/lz2D+pdDJGkjHj6UamtDLCoiO52Mey5JQPQP
LapU3t32UHXlKbUxhcbf/9cV4sG+NlZnnejn6iP99DTIYrvP1sLwBTseE0JZz6UEH1xw9E5/NZni
SAahenM0Gd9WHZ9Z9/fB7em1MkZvaLE7yONGeM8F+urWZ7sjZ/8qURY+wi1Wof0cHqbdOwLpdbRD
r8T0+wY+7+6MMgqNYAzE2Vl0V2FlrJ61vVrUFmChqnWHMB9ZR9hci3+6RlrbLd9fWksoHd0qDK0t
dLXL/ElNoWXxv5vN7GUkuuPLQnT8AfveHUeYX6t3EcLzQ4y/XcKNMVE+aZZZn90oM1RuyUt5dVOY
yallSKFy8GmDH1GCZwRHnu2LWPCeAug4mwFXLFbbrY0Boncyge10dSLtXRhVbvJrR7Bs00z9nHw3
hesUmcrjdGh6uRlfenHVs8y2NEMgbG2UquRpOHwUTV5lHLXMa4RTCLoeB7uIp7gy46l94VDDVY6F
UKE1DGGzwG62BzKVu1PCnhnwhrxT4uBoo9+pmtH+bXXNUqymTnoWz96pSXrY6pG7LnYJ/0z8ZZsD
QKJKV089GxkAtj4h/b6lJTMGwoNWCsIZgzkYjIRkxe841nOtodowaOmmJ/9dV6cRY2J1rOgp2Ctk
uyX9dJOMdUfCVSKE2pllQUinFsUeHmuD9Dvv/xIyy65z4bxFdQsQWsiWSy655NtUa1I3VDBL8Yqd
UV2wnIJgfT5MLKD/BdT7f28qw0CH/G1O9fWGY/eU1m0JNBylSYxq21Qk88N0lSGn+qpxzVA11vzT
9rMqE+eN4hKejT2FDVt7EhuL+SE7Bs49Q6bHIakUmv1eeEfDIh5jJ+Nh+COKzS3TIu2TSn0GYqBx
MCb8FLFQ4kAP2yMMsVVRbHF5oPeUTLKfFevBvil3Z7sMg9NahzUVlw61ZmQcDpKVhPeV/t1/+/3t
hQ2C+CYBCWMFo/5VwG8zEXOEB2QyJxzZQrEnY7WifGXEQqqAgaKGF5N6Rd8GPCPdNkOc8xbEtvME
Mw4FVCZ8QPCgMK86w6HqOeDgZ0QNgPpuQG51hM5y/2lKVHs1+K7Xzq1eJKfYCFlhQ5rFSm9ismEe
LdQ2tH51gSrLqMylWNrGd4LoRINUe4u0177SxCLqUM7D/qvmmJQBhzF+HwTrL/Whuyg2DhAemOMv
9MDNFPVxeXfI3QkzKRWlYfUzLn+828lPqB/zKy6dFuKdFa859WLB3LFigmllOSvqPEzqQVFBmSLx
RFQCV3VJsbK1CoyO8B0jklz3N3TFlcQfMEk1O+lo7qxaUIPzrT+U+bZzU91upI+1nLRvxE50CS5q
44klOpPpW8dbvwAkFPPNX71MYXcsjAoBt2cKKAJoKAtJQTlxdmSMEY3FHvRC4wKge9Ri+8X9XKxU
4QCsDDnZ+6x6QPhOXsx0OiLYNz4lD82WEycw5wN3wuBjM3m/0Krctti82sNP1vvcX5HfhiMOejno
747IU5AiqPR4Ge2PFUSJloS/KlFphHvxVRJafZ+EMwVUp/D8eeEXrLSfGX2dXCG4NaXbxOH2HjNE
Rpw5O9JTwYWqOc8c4BeBKSHiaiiZJmYlw8xI1e4/fZW/cDm2AKseTGDSPQ9pMRGMmhd6FPsBLrpB
ch4THMCxxTvWi5fFWtEIW39tO6rYR4sCGd3MimAkcb2Ix8GN7vO12WJAJ7eRBv9nJwpMOuJBVyCE
6gV9ZjLF+yT2+vIuGtAfHaZsLr4sth8UIEZrHhGBZiCSVLbOoKnN2Dc0ru7CtkSz6ck2NZszoy9R
l+batZkIZ5yhxJnqj1mqGqZDx0U93UHObsQKlQTbUDvHbt72idYDiEiYvNAeNNCjucH9ih4i9Yzr
05x+Oi55FnW/6gkLL9qDfVSlhEEU+7ziZ7z0PGVmyWeP8UliM4RczwM0q9VImw2MxYeZZndkrvoH
iZHsY13UbrW/C8bK9BBQiii+zIMbUfB7m3/knZY602pclZ3I5FQSl/6ma98cHEm77T1Zht3EtGZw
FYtAf2wJEMy/FZNP6VQRSmkky2G/TOPALkF0BvKP5NJpzvthMPwZ5MoxxKpfU+dsTgb2RHsyHw6K
RJX5f6PNyWa94RHSlH6coTpud1ExrQbDnwgA9G3pUVam60bCC9jsIxiNcaeGgQPjboSx7exwqEwO
s6uInmZgqB2pA/EyRjmKAMrSHYhZ1ZIQhGWG64XCplNo+DGyENOM+LzyA0CNekrErfZZyVuNuApt
Htmb46p5AejMht5O6sEHTDIkZ6wBJRoz37Z3Eag30elvY1HdHFivIB/cfgKMPPLuxG7p8kE7n7i8
ZwESsJqhlL3aVEOGuUJWcdnNy6VMBf4EsjeTz+68Z9lEZW/5iCwNdSsNrgpS6WCgi7BH1/MvIIu4
CWWhrm7IuPktivubW4OspFZXZfIGAtgXlAMLitIjBrqPYB8quITQvAp7q8kLWS+sUhD7ZQcFRiXJ
YyUcmfBrm2hznanHlqNQZK2p7RP0uzFEnRyKt0fQDqCk9LdX9XRuIVQNlHBbsC6y8a3q6AWnapDu
SXj+G941zklpJ2WDGcFSa9+69b6Vl8IS15YhFBsL7ysI0+QNZ1Pkx+DCfb50igZG46GqZKFzk45c
XcZkSQNB5wMK/NwOdJgcGZyxH3JlT9jpuOlXXiokOlJgMbB/kqPMfex6kG98gD0+C9rSkQvLqHVT
PH/hHdzVR1P58U5ltHWAUfPp8zO+oQybV4bMk7thLsgUd78SWj6QBPAjg2h6qvY5ZsxtA9B42qGA
RoLUKEwVHWhCNyvjegLMpWNFENU/X4kPViub9sjxHI+utpGg4MfSNaF8C2fTc5/gmBcejO4yQERF
L7r7uHFsZX4sp0CXa3m4bJsNl1uHEHWJrz86FdshfiIvi3Pl7/4RQG3E1Oky2thBEk9+Vq9XU+Z6
G3hEyl/mdYYRtRkOf2RaP1ydENjbw0lMovmEKB+PLG37T/gYIBvoplmZWpJr6LVVw8pAdlrMtOZu
zZQ81+7HAZJepCynYOySMCTHQJ0Lwj4fo9v+Wt75U/03IOrHMAgiGhHZAnv/7LJdFTZVCYdays8t
XxnL3NkeoFjquuljuCCKgE/tTI+gOTlVVDZOGUNd1r+4akpVsjedzr9gh1Rn2FscpJxUobthEtw9
59kiuwonCSHupIKY+rGLoee7eiytUrAq4p3WvxN4Qpl2PfTx59N5Eq6FM8u9U8XlaneKDiBj2M6C
WGK/TcJ+l0GsP71U2flqaQmgo+X9prNH+ipDLM+7gnlBJsxJSzfBMs/6/AlolaTSrU2LdzcmL8R5
U82rPC7W8LR9JEL7HyeqrrsAcuDkJVtER56dTZNJbHc8b4n6/84De8CB6BrGWQOWRsCJf69hcmHP
BTt1j9hldca3ZE6eOnvGvhocJWLLj7Z3bHL3DZhNwAsx1eZ6o62i+5pNJoe85WBgYsZSKUkqtXGz
kU2aoTFv/avKyZXbm7t0Q6Z6zv6ySNZBe+97h03bHYmwVtlpQ+3nXo0H8G1guPKaiZnuioWD3+ci
4N8PbeF2PlHl6hA//xtrL/wv1AzzxpIecgGrbEhDnWZHff7oO4pNNi4P10LxA5H9JSkOPUSO37QS
vI89ehEni6dYMr21ghvXsTPLJFlLyvyduIdVM0p5SgVLeRHo1dJSaURpxaALzHfOgipE8R+DpLxo
oIgguLMPeLMRbX2d3XoghtuIfS4OlJbFlV9QHNFqT4tLRhGzxoMkV4GSDXwcSwR/fhYG4rt5ma0I
jzwo5ycE4eAJCuVLIAtiiOc8ztkGts3ANGV51KzJ8DhLQARwkDZ7ZzS3SUkMZYVuXeRiP27KUQi6
5l8hdUfPhvbJxIfilzgJkDdXQGDrphgfzhq44BkPegurTS7XQeTjtfOWrPTSTiElE9F73fxdtnNo
AazopPHt7M6bw5fFaus+YWGFN+E4nY5Vwhyeuwyz/NCD+Rc6V4EFLNqqhSBPfdmn8BhQsrLBHH7n
BiVPmW6Xg7A5V9Vt9rT6Kx8BWTvreRftq21lA+RTxo+0gu/l813qu3wJUSSCSYax6gmnalQO2Ge3
CAr78lh+mqrVzHKInsU+fDT5IEaM8ZYvTNM9OoHawVQOeoi6HKOENzoRsjMBt7KprmLR8QBsrtGz
NJHjLfb1I7ExMG5VdgGTo3kePq/A1M/9zVvQKDKdSvJbScYvlD8Wm2kj4GbSc+1xx2qNgOIqM/Q4
N2vBXt51b6anyyORJ8jifmYMkhjeoJJkD3WzcihfmwqMkC4bqIBqu395pbtKwb3a08TAh/xG2TOA
weU+vXivRFcoEORxar+7iCf5VVcfGijxzx3TSGB+PD7paYP9UnJD62ENjpj1JhK70+QzwCORg3zt
9SJvuH5tpU0Ae7H/c+7XislO8LzhU536//SkyAh+c2yZOwyOJOkXCS5aT/Anm2rF7oYrz9rhDMqj
PHA4ZfNDgVfqRk5/5pbDXTtS5gRppbzQTeZSdQrazi9Bk4NCZVlVVDL8jtr5vrzessSCzIb6jOme
gdUtUn8YJPqBY0yJO8Mm/kU+Jnu3KAxfFmLujitaYI8sAnlMFOIsufXQJCOkKg38l9vEApUd/cfP
LP9dUHYBcZD63xkaD28tqR1uepqpwFnll3/D5P8HsSeEsKMe1K0+9aX0ejVxSi76z9NP1t9II3Kl
2Bur6DFOmeEXwVLaXqvQ+Y/s6E2s24DmZG/60meffdFCuIRjNl4nBtU0+M4v4GidoGbXwxXoJrUg
gE3eJjw/TX8UXbiCthF8ne6+fbky5D5/1j+RB0kJM6PSXM4/e3/IDoqVoplkIvTAIS/PZUfRXkF3
7SkxPTWqTfBOcu8XUX1DHwf7CNpnZg8gc+oc1fYRTcY/6Rh+v/HG3tUNRJvrRfs7o3SK40xigGp5
5ruV7gixznnsohi0H5eBo5OZRKmZuuNratRyr4wTjbdAsGQglmUU9ePiET8X4flnEQoxPZ1ROP1T
cFnP0u4U6mBk1P/Cf4lWVLy06/mxCSJTlTIGlTbtUJD+jZE/KsHsrPuFiLy0MEf1YsRQ93bqGchF
YefvfDxnjZZVOJyuHhJJ+MM7t4f6/G+cuMCGEA0cw7Q28hgA2D+2XxEh0NZHzjV6RJDYaAyDGxTn
++OWz7j1bbE5vvLSfN1tZhfK+C7Q9fWsAsXNI623rnmb0IJFCx8cYqFeec0Axz1ABBvp4jSTOIPE
+oTnssh+uR2FHsQrNkWSwpCgjrXIurg+yOcutZ8AuwBqze0O8M+53bveJQaDGusT8IhXKWsQNntA
0hpmlw37LF0IcBXUzuZcgPANBIaVZF+IE0Oaml4jA/bnkDs5G3kqHUDP0vTeZak7sW7QC6IqPn6O
y/dZnwuycUEzh0Cd0Xh+M15nHCtmrWwdzt4sDl1CEwP5VCeq5BqeXsINmfhWPFySeZDJjC+g0RNj
P6jOqsERSZr2/c3P/fa3hO0Ox84HdNNXmAjTKoa6F/Oi30aeucRZtmHOpGFKXbiX36diL75I/M17
W30TIEiNbfBLBgNn+fgb0MaNTOq4p8HL/Fk6rlf2hv4khoB4PgFR4ZLU7EacB2Mo3sUli67VKdXE
GR//sJBPgFbO/U/Dlva4xzhyDYNcnOLZL5bg2Oua94KQIgrpzqMUMFrHlSxsGmWt2bFs0p6BYuEW
6yNfwyCTsKqsLzMnMC8aMy8+OXa9+JRbc4NTbvXdD6TXF16AxTJaMS2CRPBH0n1RC3WXExakfMvy
jkjp868LsE9yfSDsvthE9Sdng5drvCcQON4dmIdW6AfFilowsE/xpHeK+HRf5i6UFqKKPNENSPSH
Yn1+mO2vJPpNoRCDvHGWLXii0wFMYz/Fbu8rta8xQ1eOLWH4Xq3zSqUEEeKliJxiZ9mlFgZUrW95
rXlugWzjXtlh3bNe9Y7N5nV0mh3B3Hhar61Ivx2hBNlglpTk0PCeDglVpbDSL5FlMHwynETltjSw
oQq/LfTbbOD5CrUunBCOHPn9BGeR9aWQQ8iGPO5UMz1/9Ql0viSUVpB4HRk8aVijjuQRUccOlFWJ
Tp9JoXuiBLNF8zCyrui5l7b6qf7F7WqqkspMvJ7zH3fnL0zC9Vg+K3sR8c8GZSQ6fVlAz0KhQ7jh
RFLp2dfWW5BhhqhO5U7NGQMy2BzLigGiO9PwN0LnVoC7pv3ddXlhlWvSdhDH+b1eqZRv2rDKvaV6
XrcZaPI5xyJOLZ5tap4SccueIWQxkV1gtLV1dJpE4rg9aPL8BM3zX2Jo5Sa/H831MqiZQtQ3QYUv
rG5CEJsIEmHm+QlfNbrRajzjMSnluro33c8XjuqQEqte+FHCqefpIzdRbApP8z/voTcgJmUeierO
tRy32bWHm+bWWvh4DyeJCIbvTvPxjS2kKDBUjG9/4finerN8774eUm0+ND3UenIQ2o0vtz6z9OZQ
q6EMctxq1zjFbSDn4ccSQ9k4y7ZKE+wTHyY0YrIxDQs3YjIgoWZHTE6Mb9XRHyO7UjvCRQSPR6Dp
jjRNhfDmZ9X68i3vmF4aGX+CQJAVBqiy6FkNttK78s9gI2xSSlRafmJBH5AfzgMueZql0kyKyF2l
mckDXAuBneoCYcvGv7FtA/Jucx/nAUvZZqLCEK20XxLKOhwP+BM8VXiX8uOkIAe6QZXmaLD0yGjO
SI2LOtf7KPRnw8sKJSkSmonueSghvYd4QqjHDyz+xCiCSIo8MGCW/8nQxNxokH3zbuH9l2mWPIrd
MP781g6yl3R6RnJ4mkU4WW+8gAJpQ+V3jAcRv1mU0/yGTMIbDweJXvO4OaJcuLb9yk3SxBvOffoI
weiszmGL39y3z1s6xozeJGSKwzJbCHcCmSC/orCbOMtrAhtkioNQBj246PVlZ3Lk/oL8V5X5TZov
jO7kmztKIe0TYDyCGM+NYJsAFfqhw7qc6X8Sjd4e/JTxNkaYPQEFiZV4MFzn4rqaifDF3a8ihdJ/
91WaKDoeSueJdMyECCYqJh5JndXNu7jbJMSB+CinvmiEt0nMTQcfoPBbI6pqZTwkIJxRzhtUxGlL
PVLdVdoptSNeQS+L4HmwrbnGbE9ZLeGVSmVgvKAGNCuJpJNrE+vpipKNGmDaowpJ5X1c5niIbYZd
jKQ4mqaG0PnbFfYI0Mf6dxp1bhMeXFAOqmhOctBiXy0l9kBXKPk/sBiKvqJzeqRZrkzVyggMacuJ
GULMMXtAlIfp00h0gctfO9JRLTQjpqEWf0VzK2ywmY7Dg8CWyAYnkA4FE6c7lW732IM4U6zMzg44
Ypr22XmX3l/J+7e7uqaK0vnEwN0abLLNwwP44gRo8/Gh03ZgiUcp7gUpapcXKebRneoYrpzNzqkz
woTj6OFH1UH/4VE4m1Hez8Q2MdNr10Jn9y7VhVCxG7CRAd1FwNl0s2whgcISfI1vbkqciJJbpYRw
VuQACOnd7LX716II2CdHh+FN7ilgx5K033c4usN1W8+REgvH72cJAZ4Bwlga0BOMfBmtG9s1AGkQ
VxquAotekvhthMf+rb55/ypGXHioUR/yA/ceqlSVk9SPFYhxFoVIQ2bjnSZWbxiji1+2uRQoMQwc
t3qOEDBKVdwt6ZC5jOp9on3wu/VgqCthW+s+qB7FWItGROqi7o8iILBlqoMfUssKTN6L7dlUS7Ag
+DM8XU/n9ux6qXhTMkYafPTApcA9JqHC9TzglBRglihPKtbSCL2k8+J04venEz2Kp8h0D09PkKDC
6crEIiIaBEx3LCtvRdxw2tJU9+Xk+eb19Jg3l1OTrDrh9PcZRQzbFOh7CTPz1aHP71+/8eV5dxx0
b4DZiBjf4gzhx+fVoyRAk9HKF5ajJnXxA9VCFlS3s17x8GpQfxKJgoduPhJ1/fAzVlt0ud+yKXgc
1noSEv7VLvp+AP6we18Tm/NSN5NdOblqwmEk+6Ig/zOjz7d+e7utmcWp4FgARTH1anRHjHqrYknH
ux0diGke1ppCAP1JTcuhXfEnMc89ZuES78pZt0twWD5DSXw6UoTuIoNwF1RkfXLbQHJ7dYJJSIB8
X67/xBzah0Adkno7uwH8qTyugEpUZx+M+YvbNRBv8k0MMbkJNXGmgqYkluLiscXpQ/APtnPHY127
8CltFYsak/4GvMDUSpzk/wo02jEgVji35RMGdllrE8jDd0uaUhC1C3EJRzk/1QTLvoM30oury1BR
lmGLhL5QWdt9xAlMgd/yl8NIdE2/oG1QBwrAyGXgm4BoohziNDF6PxKw1NIeGPTxGqESU+FsqvLj
cYsZpUihqgyiEbKIgcfF+41NixH8hQWgJ8Kh5Kb4fF1h2eMxk3khVP2jvrmKPsU1QIEMHyuJaw9s
Dhcln5uw8ZJiiJ7htDHMv9CCZ2Ob5iCQMt2Ja5jnMm0XblTtYGMerQaadV9RF9kEMeg6xk7BFreP
c+8HZ/NLG4CLudlerfpyhzAmiFbpSjXE3g4iv7niWJfvurSLRRsjHjJ0SjlNb6IvlOvUUbLGYZF4
TD2t8se4fTCEMqsoH7Ig/RvmM2GV/yzsqoC2N4JD81wR+NzOOHFtbtqensbDybEIX1rPpeRANVtI
zX+1aS3okBk1sD8FRv+bQSDORJWkOSnO/XcH3UUiu4sjzfnoB6onNpRWzv9hvgeUDRhFqjhfFF1I
L2xNbRj+SJCLLwxqE+5T4t53EGdkRr6g6a3rdH7Nad8GzOEmA95zh4j+xSywgByXA+cBYMOkUwKm
tdQM3EC2hIfBSUtz3yuWM7yzR/l9iCZkwxtKivuXae0dmxI0Th2Fk9p09Jdhk3pO4dfzJUREnI8K
aJP7LUBwV/iX20bk0qd21lt24DHLY54txWrx4bhtuqpWOg3yegmda45m0Otm4TrXMO59Y2ysFXo8
YIReaJNT2vvXA9fYjJ4qwBFHQoaeOV9pg2U2o3hschDF3j8TGfZYTMDBSLitJUZh3zmw8yDKlnoK
S4i3BdYzYRMnagu3v/NpOro4wTq1OSr+XH0l6cyZgXBFDiArTV9/TnKPLfWLyNL1YgqCaaCQqnI5
e/YZhIpQeF2TN5GstuiJdTcLIojzBFsvMxbUy0HxGUm0YvuJTil5NLIbNdQvPea7+wBJxJdGVkFc
DxO+23PjML4Ts7yHvm1vGZhotnzk2mm36cUHAoPqIGiHMri02O2MTz69UDZEV60R9NaeEbe8rCPA
gzGAHfoweEX8ojictTp9qxY04A7M5+Xei15qpa7rGl8bDyF5snVg9uS5YrdD6gE28v6HiG1CZXiy
6vtLPESO7gaUtXLwL5q126iUNzjovRLI5giNruGh7oxoepf9ExKBXSc8ZDV02jPXglqnkXCKi+8M
zmnC6v57/QNvxL/V6sHeJlcV1tW98pIRg2fSUymSmeVy34ud0JmPHDuhiuj9Ek5gvhWlKBmI7ABC
BiS2AKDcbXnzE6vPGxWHA+FZk/rr7dvOeJ3BSpjK83ESSA9owrLEJEnqEjsKBjrDf1J34tdtP/It
hK2goOTt3Vz2x1zksz0ogGV2A+N5sQFZ6jcs9lBp7AmCOhXwDGCbp/yo74x6FjOFAvv3murbk/a6
MN8Xzz8wv0kkZD4KLc3DoldLv1fKyHOrIbzDiwW9GfMXzi8OLOVI63jWb8aZECSyTeKdQThMJChu
j0MRTWn921dgzl2rIENcJzvbBeiZOSFjzPzg2sKMvdIdm3+6yyFP42CCayZHoxu/tK2MgCAwrZzu
0Pknrl9YLj1bCWIZH/wuQX7GD2B2nYBJMgD4kN0x7+ygZs3n1i8bs0C6wjLvyYqaWsPQzjsZ1n0P
tnYuD1Bhzaqf85wlq/zbPaB16B2RYE3VA+dN1MAv1jvse1Q/TFF6PL7YbRnvkAoikaSaGDKXKxhR
0GFdyJV02o2CdgUKgLAikJXVjEfMoubC3MRvDLBI3FFjKv95bWZJ1DB7In0S/b9veveVZXLFrHEQ
e7EhUIrNZ7DHEDJduz3jl+ZgCXK0l5D79wnE0tg1ioLit6Ilu5GgqEuo0+P7U/HAfE3wBqzYjvSM
fspobQq8mGBKL9prb1wMSpeLQjYm0dIaYovBjdqrAcXWEho0oMZREt3L85OJxOjzfibW4laR2r6a
1PEnOZsrjCt7zcidQAc3jFSlEpjA30MZFzUV6qaje3XHBr6TeYNPI1ZiUmKWFQWDjC2hv7TMcbFA
IbcotQL2xLmi10rIT9QmdsKn7bZORlBlCg1GdAm7juScqmbCP4Tw2ZjBdZySXPUDurKaIuxceWfZ
bIpFMxljFVYiF4RENGDBrKPtoSbK93bmohLbqYbPk85eizBTR8Ng7rlkrNoYpnMwoIgHowLZwVrG
mLNZimK+mT2ERWIKdeKuVySYqYmRXmZFOd+k/wgLCSzoImu0wiwifX9QDP8EA+m3TGPZ7BErfcbx
zrJwgQjzNfjdRv/yqD8MMYrn5gDgWae8Vm8x1WU9elXKTD3Zgd20A2uYf3cehLlJPolJKDRx6qDN
ndhCtnSCCqwl4pAfNcHdFNfaG64c4h49bkDe4yO6T0aGoENjdlbfXV+3NkHe5R57TE6VVccFbcUu
4/3cxE1Rd5hlsZwx+QfDgtA+YMRMevbjDn1557Yk5H5XcnJvZ15UNf37lA4Ju13mvgYJWhCxxpeE
RWRs5CcFxxfSMfEFVXYh/YRGwbt8BHb/eFuvnmdIL0RSpLGkY3tqssnvl9XD4HmKIj8zo6hVL36u
+KehESTaZOZM4k0nhH5vx9SgiRj6lweMB3XdU47c16Ojsi3HnGv5bYcweLIPoSwBHAJ1oo1q/U+m
3sq1iWBfgK1W7zjz6BISiEoqQESrtePemoGOGDNB/ai1gYXSr50bi8eO7OdmrETSf8Y5usyqJ5x6
GMKqrHvZ1zpFbZuQhJV7vi8Ibb0M9PsxLU5Bois9GAi6Udv9M739LFRVrZ+SpSiCZZrajuZUag5z
CCMENF7nxj/uLiAtID3w5BfjdWJkCvwYkqrJmYRl5ARrSXgNwcKiBv6NwNXAFpvSZQffznPal4nP
dUsbkOwI11Q7uE9dt0R7VNellWRsv2IQQZGOSdOGsvFLLkm6GW3hIBiuRD9DysUgPpdQ0Gr3e5bn
dxctm6Jm0j5Jo8F/fjadV2wivaS8u2WaLxML7zP9Dz6mHTAtu2sDF/fZTe6HY/q9XTAPB8wV7TEe
pZaTyAfItEkBrNkVtbTTK6kt7mdUtijrrGZqMYR5McMSDAk1nteHB8YffuSBBJX8vPBeqV27jp+f
7Q+Ct71zK9DV0XbEcHu235Pa+mHkPKF3T7Sx7X9+5aB27wzg+l2a/JMA2k9MBqg/28nS1x5KpG1n
E0IPeKB+xfmF4R/hNNk3RcflJIv5k0k/afEzV4AHfFTZqg/yi7lm3fSRx+X7e91LM1c/Bya4qJc8
1b+hPfLEyuSoREcaVmCm5aUI1h0I54j4sLJy59Hl66ClDFvaqAAWR8r4bgEzEg0eHpC9RtgYWYEc
F73u6YeXqMhgfn92Xy98vC16/izHz2qg42jqroOqbcJNYzPwSTil2HKXcZjJeVHWuQ0m4vv5j/cw
nOQk7KB6ix63M9EyBjfcfPap8varv82rCKMjJtXFN3R9MoBgEwobEVoQehkh8X5j+oB2dJZaQrqC
tkrG+VU9rKaiNYH296B7sn9EsE9PzABU9Usl/8CcfEYaNJKHcTBHxxuD6KqJO/tjcekZOfJs1Sbj
sCg2D9Lrp8/tiYwtnLrEjm2XUr8kzTKYxdLYeCrh8d7nJYvAbZr95dNWKav2QN/dnt/NFViSOdh2
4pzDaqDmZ33y/EHYwGDJ3bKmCC9UZ1TlK4aa6XTPZ8mg8Rqj//bVXi6YgBHNh9P1sl/Hcf1Iwldk
AS8WF5G9QFcNCJoz1eC04+p3KZPkx2QuF4awOEy6FBROSnA1zhWQJETjMH70tYfhf5JifP55KiIz
1wxVq10iKqVGFYEp3M7iTOb98SugIkjI0tZhv+hyu8lQRhFxLraR7BLfxZ4+6dci3yPkrRAumKQN
Dcz8SAdSdicDiJeEyMBX4btov/JKuZWHIpaiiDVRRr17FsEE6wkzYOJ/xb5m6fnso01jPRznwvJh
m0C0HTWWDZYMelzm1GDmku94uDtOO60yXgurXE/aEpujY7EVZWALWRwoP3OrVsfE/H3h9jLz9QDa
OW/1ATDEZ5NHl7XSft6ghysyOE4oLMHPVFr65P3R3NwjIJKuLwzSIoHWuwWIk3SDf9/gmAfB6Gic
Z6beD/6lSo/AsPiCff8jCXnDoakx+AKfnX0OVvAtyceOY2qIMYWCqgXOpqSrrPNDYSHB+oxnuxb8
43R2kNRQZ0Gj6Ir78o8/RIApllM6H1AK1g8NbGJVWill5pHAo2/Ebw8Wmozu2+7SucL5sMPX+yug
s0QOPieJAN1fOk11cpX8iEz3VlfXxXvIakLtOlG0gHCLFJCSgTcSG/YaXwRpx4NLJbIO6BNWwTNZ
hyfpoI6iR3VsDsp1BstG0x5xqFgB/TfjIio9wMlke0UwXKgADP6QZ++XuF6JkUz66vRHhUS6Ed11
ST0Goa/pYxkwtWE8b8rKAbsIgCSraBWaJgzHRNqHVxZ6oZ4mKwFuJj59JSRyxAbo4CTfI66kCZMW
19cGaNnrt4qV4P1TjfBRSRcWDgTfrpFouFHnKM2yLf0bZuKHnfggE3ZrbY89qQhYFMCjJ1MH7z64
nL+jOjsVFDkmF3RQWLH/7a/WkOJkFdtgaC/dM3iMvypJGISigjatSTQomYT6UB5zt1LM0yCvIrJZ
jhGTaxKrVgjBbXAXRwBpDurosdt0uwnXIXCdnflK1cPmc95SkpBc7rDtdU01RnlNKCSLmAzuoS20
I8e4OHF6Dk0jdpZHnTeQTTFAboX7zcyV+Jafk5bNHVsjgcV4g1X48tSwlh7qnMWRHqgHGLya2+tV
90PLjrbRZhOfOv8wBpgnarQ2UaKJoPysEc+ghU/4CPgKCY23WkleBRq5sJmph1xOsZabcj8wDKB4
jiWPJXvyuQiFzqZcocSxud7GycDrA2/eY/WzUR3krORCWA9vlcE+3zlHAq+d1zMWjJ80MM4hdYLX
eubZxnOHHPc7p1Q1mGugPVAWQa2pdahbID8HITyNiGagbml7Sr1f8Oi2dQPu5JwAtyf+ODHDqVal
f+8uUUgcO8+oTqw5S63rzLWyju9YXPfv8Nu2NnZLmgRCh5fjV5w2Zs10d+G4ZmfhlEldpPUaHdT0
+3YJW7jXmhpOJ50vzXcucA7RiMjR/vNplpEtMB/Qb9pspQYGd5cKqe+uunTXTkumGP5SNGqIB1am
k6VnGGJehkD1kdkgxi1BDACkKAtW5LTOvRGWBkRChJH1pMEJAYJSBwd2LkHP693SAAOUKwxs2Rqn
iqdixPSxoHw4+wkcl2/D3/8Y25f+F4VjYi8n1AkXjDmH/Wx87kyA7VJczBeMy3H053xl9hBP36s6
4RZLsthzOcDORDZXAae9klCfFK6TIqsdT+P2Uo+NHmzIGjGQ75rjLtISlsirweBrf0BvNMNJaYw6
t834f66lR4PTcqEo+EuSdVHcTEZTPwL89mb+Qm7RuA5cfp86m/FOe/U2KTZY27E5O2vawTt4JKmT
ZjaX5QJ1Wv5uuPhx/TJc8rneex48EH4IbxDvSzFzzrqyItf9/HIgCtJumPe4bQynJm86xXgHKarF
yeva6cdo3K7QmM+IqO9TRZAGYnJ2/y99vq/2ZVs/OSbIi2MzOJoxrNHej5jowDziGt0PE4HSF6YP
x5MMpEQ+xFYo2IybNSRrL/6o/YBaSvj86pylTvj+RYONnJ7Co/Y/WK3UvLiLL/Uqr1oVCeqo3eXi
I0mfe5jkPuIt4tbpRSxOq0o3YRbMy3t3zsPDVj0o8mozUQ4W7m+zzhujOUzO8NOSfatC1lFJU9NK
a/ByR8+BJYymlAtMnKWUEKHQWmjU6/VA4CAhKgFade/9r+HYKjqHqLUX9saVihcJfEzXMThyPjnR
gh722kV9Nzp6pYIO/wwJZT9bZqC8bFi7VaWhY+i/DabSoXZLozYLuz3iCRMn6U5N/+T1Q05GUvgp
soqEw+3I3B2DvmbHiU5/HO1EgyApB8TM0wWlr4fwCyrwfKnATxmX6HGqUCz2BKM8HkBsCYuFtG6l
kx6rEQik5RtTatqK4QxKC4fVuzUKWBDUZ72b3U94rXpLQ8Ax6nCNLW3DXkXzWDDIuQlrhZ960t7y
zw+GPIETXsCLKliqX32/UEQ4fI7ML+UVI6QMgUpGj9rD4t15p//83zHqG+AWGEQIh+dCkUVB2PcE
n2QA/CPlPVQwOdIPOlZ4kcPVcHBAvsrwR8BNp8rYS6G+XU0CE3e4nsFEN8SJWPwPA9SN7hZKi7MN
mFqEhebtsp3HaD0rMvQAUJ6i+xSYH9NJM+uo0MzlWYoTarX5R5qHLj5Hr4Rei010WMjz0ZpA4aBd
YtSHuLhjjxySLJDRuasq2vhHCFlPZOwpdZFSiUOpZOUxyUNAGA1ofkWTKicHaJI7ve3YpA6fWR4q
TI8tYv8wo5KirLl46lDC1zaYSfDMUwCFEaa9JRhoa63Bm4tojqS1ok4qrCAIn1Zd6Zw8hiQIy/e+
m72QNrT39CSeoeMM86066Fxg9qCeHH0G+QpDWtJnV7ttbloaWMzV4v24rri0rSqTJ5xJaJu8ko/L
cFrChgjIyoasccnwbHTDtm5+o0mGHRLxKQsZNapxs5t53u8SmB+sb8PB0ldHmpUMd1unjBfPIgD1
KWib/9LdkM0hLgQCa0Ls/WFHkC9X9QKfP3YP7BD+VTtxd1FeFQWtlTUPGl+e5GD1C8OJBRr4tvoo
NYzC9bGp4hDXlitcNSo4LCTanVdoGuHXqiXFop/UUGsxArgwA17lijqh1OeZhvsfdflYliY4Q5pF
v+1ari62PV63grC9v2bmw6kfvFJMB4XiaBRsPNpEvrx1oAKF0eiGWssReWgnZMZfY6/iakWhtwsO
Xh42bYjqFJpjGJCMZWM2VgoyzfVaiUSc7YBwm//Z54eA7mjShcMMl/JzdSQtLirFqMP+RwHiTWQW
Nx4jTIKLlWL3xh8OfsQOkKqRYjp6n9I6UUz0nTd+8m1KzJEBmtT83bp08hXm/3ekyrYvWCYOnefm
HQhg+INaS0MKJW8L1ZLUsC4YCT38Kz3HypWlGaNCxWEAJZQw1eawE9XDrPDCr8UxwEkR1DPww1kX
ahwvbksHnNu2d12cCu2yiljllJsLt3G4TuG1ZXplrkNiwf0dLT1M/M+/CgZIcVRLgpr1vcOUXeVD
vTrMeOTL++P/reRUwXmZsIi+IeWij2w9CR0jU3YEkcyCL4dLCsgh7/amT5mTGunfjpsHcGRY6+Pg
U/JcbjeGkhMEZoIYag7GIoHTRTVyrkgkezPYcZmqtpGBDQtKmerCDJ5IpqVxH6nIZfPHV1sAIA6J
D5HVhxzkqV+EK2n759JnociD+2GsTBLpYf3vy3RKMUZiU3tDugl4DCQJXIdM7y3TTJpk73eWKvho
HW9m0XjaD+pLWJB7h7T+7QmZMo14fwH7jzMJYJoNXMxfYp44hSUD21JTFW9CSf320VtuqA0ZihRZ
UweffZTNGWYPJmV7Loh8UM6+URyiU1QUABFkb3RJV3tgf86N9TNmbh+GMFJYaOo2R+z6hYEnoeg2
ZFTy1KhzTIVTiqP8n8Rbg+Bdgb70C9oTVEKY9Nv+t6zi4lBW/RJHYGJGb3aNVvyAg/IcSV+fsTKa
EtKUiUy1GV6iTEs0caoeY8K21vcO2ItmpYefStn3OQIDELnGMTNQqEEUz0yaAwJLXMRSmWvtUptH
JObWqgC4IrzzuhwjpJ43cHjb4UK+kJnfPnkPd9Dy8hLrxqA8PDpSqE2DSz2S3o6MHleVPx300BH9
Z5mIB9csREGsxVX5eCBQjRn0+7CLa0ldV1UOUmcS6J/Hy+L9XYvv0Ld7AJ99Oa3xYp46/0toatyd
EJ3/56ivbKu3GM5DCdinZaydmhQfMsfZ9T1xNOUvrNhXmO9YTv4UG7SLuV2CEIsaexKNGr4uA+36
4vIqvu1nayBEyIrZOKmjyqRTuXquB12SrhYuuemDuduTp20+X4dGTPU5f5HqPZcq9V5GV9jNnIjO
hz9KiwN/G2fAgmsIQmm2+TqGBvb7lwwReoL9KlCZn+bzL/Jw1Af0kf3Cye/RyPd7zmC8LwYyuDnC
xVGeyPVEW5zEFbS349QvzrwtZM5vzNGmbdioywDskJls3o33IM8cH6S8+yF7k8p9CX2FM8AdbxqZ
3JgZkWSkM3+1UA80PJ0hDEd6p90SwIajV9AhJfWozQnkzSjxR+RkDIIW5QPKvF0PQ/7B+amtk2E/
+6n8SOMtJ2sycIdPbhkuwAw9gf/BgByvPG9P1fmUYGzHs0G7TF0B0Urxvl4bmuM6t/fcurF1kF25
7DmJSKh0cov2xhSJkRvqd0z8UCGwYz4RNpYQHhBBQ+EdcQdmjFv8UTq7bmGupgvwSbtVdNWQS+bo
6doWPKJYLIr1Zbm+Jaji5fJ3FbiFyii6hQKXcf/wMg9izY411lhC155yhZTZ5U/OlqaNvNG1JENh
SYOtKNRsLq4nr7U2X4jxBmGtzeQ7t6somVk7TsmVPzIkSI+YPB04cIT0koonBOVmMf8hn7RNdRWv
mZt+jPEkW2FK4l3XmMu4s5o+Tbg+bHjreI8Ma/i/DrQwtorjKSahVapyxqddTVo6egKKVQEyEskF
v/4QCtyzkLkk8zqx8a97yFBEoau3SJM4Qa0jqBwsLSxl8FI9AKOQ/UYqWyb4q8fa8/Ez31VTctEM
52BjQ8sKCP0yjgXOHk00wH8MjvRpK95gLuKhsD2DLCO0hVbOe/5sNfsHXiDZtEPPGlcNZxH3o8cU
ZLmMrHFV8W9CcEh8nLkZp7/xyXYj9kvFKeDj4iCebbFi70LoQeyKY9tBIVTMDdl8Q5L03dSZr14r
Y7KTRHK+BS28XtNlsCgeT/PRVkOhmb6wfJY66jkpkReNVSjF2s455qrWQr4FQi0AQAB4VQ2RJccw
vSqP42X0a9XUKJTBaVgDrd9M+xgyXv5Ajpu1YzFtswK7e55+rIuah9IwpPHfTkHAqA05NwAnLcs1
S1wsPktqygPefaixllQwS3U0yTwLHzOAuqXxbV9pTzZ892Ta+mnblHdyLlJeuKhETk7r7jLyFUaL
ZcsHREWavoiq19alR9JO3nw+eptScbLU655GlJxdlXVnsyvdCKFa84Ffn6DUG4totgmCNX6DKAzy
zHClrVmC+iYtURpPMXakECrDs6JxPBbIPbChADZPNUlXXkNHvCLglCwoJtPmgKUXsfFgmSU2vjKo
FGTmn+91OVulmYJ1awwsPLYMdnRdlHa+xmSJ7wb8iDgycgSAZqbY+W7FnJM34piHDQMdwWiIPcSd
tbqkQ615TNALqzM9eiXiASCqCXMIe9p6ieWFI/u6jaOS7T1dlA5dwkKbVJbdqxbf+TcMKMKFiLes
y+rrqnZczUX45TJ3xb8yg+fuUDut7LkmU0Ljqal5WSW8yp09xyFUjjX9aiTeq1o0VYrZAQKhYYtf
EaQN5VIeirJEn4e9AQwVB3rNXr/qt+sX8UGafYloFqzvoUtf0pIMQzvPBxy9G6aBvlAeb82jwSkg
ydJ71acLRQ+P2TZM+p6wPxMyX86dIdpQdlNMltZPlULoqp3Vlwg286wtcytArN2vb7zgnpIUof04
+ZwWRPp7QC2kkewtOCEyyCV/NimyTfJau6jVapylgoiOEk0b3H6qcStkYqbL7D3iswAThCLxrsWG
3nLY24YhsG4KqVAxWwQi3Yo8Qvr0Q2tFcxuWJHLtqW9WMvrm+JNf3eoBL6DplcgnbMoMNATbP/ty
FsKaHrVkI9fZYBzzR4JhJweeZtCR3CyhDs60Hu5J3S2/yOxt0CfZxfBPglpFI0T4jWOL4MIlz430
IraiAmtaF72Y5+/hzTBaHZ58kFFF3UGc2XXGrf9ffvZffKgJhqka4IcZ9NXgFQxev6LP1zoFJF9d
nG+FFvUFUaqJjylaoU/4blcvtiv0wQ9QD2UfJbcNBaSRzhRtYsCjxj4crL5aYuRzbIhMAYf48p3u
cltTPW4WrJMzv1kEPstSNveU/zS8wbXAlKaERROiClC/jr+sKOfLQ2Ol87egIFif8b2YbXsoaAET
8wmeJyWScdwqS4sNsJ0f4XvV9qQ0ONIG4Wv+0RsDDiLwux8QogGzoqDbm5vW4nlenuX/v7A27khV
IqQmOFJadR+ifW2BxmELCV1xbNS22GDBH39n341nbpRwU4fjqq0uoSRG+ILzu8Fx8i5xaXBAUvcw
iUyrhG6JCiMh5aQJ5VPyigprThdPqp9AJBTtSFcPZzXlLRrTgZ24Hz0XSUPS72Cll+uc2UkJKWol
rl2VBELJ7ZWF5is/9o7iL0C5t/Rep6eBN7cu3s4NCwpGFz0PpYQcPv6NWlnQJrA6FDBJNg/ReAsX
01mXb3bY8tvUMuGaRzyR9vWK5MafB+KXiTnAQiViyq6hChOwr+0hlSDSRucDO0UXglTdhJM3g4al
VT45sFqeTdQtNoGAijS6VKYo3gboo+bkPMNteB/OAONmUsVkLLInJWY7hHZxh73uisxIZGVQ90w8
pdwzlw5E+xvL5SsBszoj8TIctNr8ejuIZkrnx2pG3g24lEweSCBL4uDp59XpG0RG7sSwR6g8EbWA
UtblUifZX62NzSkeFDReBIwVy26SdoqHEXd3/DjWeRsBeZTr/0Ly5zGH7NyXfTTadAXAK49cFUck
cskoOddx5oZMzHNIubsjLXEyV0N1dZxR7b7Ov+hiYssqXIHV8cDglth253YUhInxdHBzhprW1G5x
5jET80nGKsiinGchtzTAURgmYk3aXT5jDxuDoPuh8w0nX76GEh6fnEg6oMtFJwdVgbwc9JCTolxD
WHXfEss/swkZu6nVbAkrc8U2Dh0Ly0n+McE7+Aqx3+ejXOPmh68xA1cWrlaf7rpWNesko783lDHs
XOyRLvE0nBADsXSPAiZDNAbIEyw7NVtrgSHANzRrvrjGGh5/2wk9NhRCgTJepUTpOwpShPQl2Cfw
MVQDLYrktWdBA3vi26kdm2loiKkVzmsEpt2lXjtk8jLSN+2d+zqEzF3JW42HivZMglHinTZiqLU5
UhwDvVvblCaSEsw0Q6v/bnEKkZvb0afJgxrdfnSXjZA5MIyM4wfSkxy2IkrvSvhEWjLpEip0KhAd
c7BngcA4LpCajRGHn0sFEeKdGJTM8Nflju3NlQ9cT/7Shon5ZmKf+j15VsuNRpMq3zmMGA+rGGyz
LQRKX7nWveGmEPP3WkDw99F1dB5muE1yzt4kiEUyPsJPG2Ug/qTFt/WMJFwc9QiJMqFoFetuBzdT
oL/hfW1gh458DGAItpm0td2BUXFVkQoj4lHwFC6b4M/pVF52xMDGCFTSS5MMjHFrBRywJnsdS9Mp
AkMCIHVuvov0U3JIpL22JdW4MGIAPAQnSA0ydiSt5sdDRJsuO7NemRcUG8x0eFafPhegv/ZZmyDc
wSefpfYU8FMcJl1b1F3cYNqL0dEmDLQKhneAX4lcK+dMlTKxNZVZrVQNlPb0kxkf/W1iNecovbf/
GgLAJr3vlk9uvwDZdxwlDkwmGkCx+7dySv83S7K5Nzzhi3uIX2ffJvO9BX7DlnDsXSdUGX/4nh4l
K5Y2A8twPI9BlLEdvvhTf1GZ7mX3+waSJRGRTzGYVt3wnnBmhHs7Hx7hvVem7JYOTUWFkngtu68C
yYDmyyXKAJmSWj1j6HXTy4cRk3F+FlDxudmvBiUjF6RT/dmc0Pbcn20jS7aJOLMDPAOmPeAmeDJk
M3wzjIBvLMLILrLd8d8qBTLRbD6UGa97NbMvC1wo5Zdz4SpRR7oYviXeCSE+bFrJ2lkrfJa0MqMM
wXEvSgho0gUpF5dtkM6qJimUx4tnAqxUh5N98AfwFJeZUEoDuZZ5X6tRox2UfVF+4i0tazrZp8LW
5WgFUNeMENqxfLydnw95KYO/eWGH2LjXpqSoffLjlIIgAAL2rjt2lwY2yrhMj6ul/oaDXSBPaB9g
B1NMFhSMix043ApJQs5Jep/IWY3flSAdS1olHjftKOOeqEbb0t/3Al4XtFd35hITs3z2blC+WYga
jhS2i8gDhjH3HeuhXaSVTOLfDn0Wcp/sntCyy548Y/xpZbcZJV0SQOGWpupJqqMaxphKdqfM906x
zySSvwFg0OJceV/I3LXUL05GvijhCS8VGrJwuHgEHXYEK/ZLGmYZE5CEufF9P46aPGNq2HUddrJg
cCZ4WKLEFLq+UXo47wQXLz9n+B2BPpdiTbC9b9BTTlb0yPeJaEZawRYLBw0PjgklrI+4oKlB3q02
Mvr+r6Ldfaqb7vWxs3l4MaIX5T4+9iv4Mydh2jZTV0nFdp1KpnBdm+KPNB9QiawfXrLmRPQX0kjS
RczSIwM4oh9MDNdeo1hn5B0cNamHU7TljIYYtX0Uitw3v65sVriwKBcVvWzop09/HAjnIxbeK+FT
RR5L75/KQRLkx0Ad5a5Xbs2CL1Yeboci05Tr6jyabJbLzmQwzeZDYuUInO1UI8+WQ9CL3vchG7+O
tneu6z+lvCGAHUb/UbmuxH2jdtbQ3crybZnFFYkFH15QnPbm7eLTQXsPgeQ3HZiXSLAKgKxqPwGk
zNkg/65BgrEnMmMtfWXXoFqn5ZTgedKi2NfGPfptlE2/grnmSAtYTZFOinhLzUOfcbKqYxo/FxPq
4IaJIZZZe6LcVTAl0VMVzf3B11zHIOr6Mu1Z5jSZtTlv1qZHxm21t7THZ+kxRa1RqEf5NAPpW8of
OAru1WA5z3p+x1Ezt/GMKpzm6dDU9U7FUCaQFDrf0/XbyJ87if8WeS5CnJTYpj6mTecadRXAcv8b
wKabwQ8fPE4OTJCVxOM8XBbVCNbk464YOPD0Y9ZR3jCxfJV7evSI9u5PUuP3Vr0G0IM25wN0+jm4
BX8VRBz9CPl7uCTe5kZasvFI5p6+f8Qoclg+8ioZ5PILRNsMxh+oWqK/3M0oU5dGHmcy3tGzDJqR
UofCO2z/1Ce09Y3mPsnoVW2gwssQxOp3tE2qqK7gsntpKbnL3mxWxt8dPmSZu7bLx2YwEJAU12NQ
eVfP89uZfafPVv5/2mISJql/Qg3mziRSFoZJI7KFe8MVahJ/gxa9QsKJKnCEzyLgPjr3ygxrfjNj
MATvlrb1mdNqdRIhfTi8r36Dd9reSpHOR6Y2QYjQ0FlloGsS1s2y1NHNqJqNS8uFEvL0rOk7/xwz
JAE254HTTb9NCLXCyF+pSqfavMLjVqg+hTBUIYcgX7b+nBAb7IATRhVuBmlOR0h5e2uXjbDjPyi7
zDUc+tTwT+s5pWVOTV/zMXHEaOCyCMoovY01CfAp6RZFYFrbG+IVdtkgRsyPNZrcDVkKCeRc3yAY
+z+tq2dKYUKA4gf680jmIoCfz60Uh7QwnD9mvkyjrbwEawLCxZnjHXz2LvFZyFfNlJXFN1/FTz6S
DfLAG8hJJuzl+2B2LUdKkB6rvAGjH3Ph0e3+aggdQl30XvX9sWTgXlni7cTKMrLtRL4oM7pdHUql
3ndyWxFZJolDnTK512xU0n9jlFWUvxGXz1Cy6n0zWRl4BVzGHrSkq6ch3K/sKBBKNU1cQ5buf1E8
eRqK5350Brq4HrWArZEbbc1kLoP+XQubqxcwV0nh7DdJyTkXysFIgCVTUelH63FDb3ot3YyuH3Ih
KuSIkeIZ/cElJrCORvaHgjbQz449cez2SRyv+7XXGJLNUD4dvFTX3mlMlYScjjD4c0E5749YDssk
z/FIu3P6JBR6uOYgONqwSpfZgloGOiuiYeGbdjmDV0OV7Nsr2kybnbqdQ9Okm9Z8cN/2vfbrcsvc
PJTnZfdiaP7UwXtytZOoQU0N0factwzEoetJCUcCrWwXcRXGySDRBw4IasrbpvihAL5XNHtLkcwR
mZ4MKh7RW7p3RkpZBqtcgRGAtLQ+Dn6JhcwHCg8inJ4x4MtM515zA9wQzwZ7+G+YqsgRu3RLsiVW
5a9EGRZ6E6lWrWUdLZtBNp8D5gZkk0FBRsjNL376UzYtEQTAR6UcZw2wX6hB0xyTH4bbYo0pNTx6
g+PTio0DdJl2XSLYVJsNekzjMdoZqaa4Rx73vhk9/WRLeFwlqlSI/yUUsbJxHKnLDtv8yVfD2J68
oOsHNvayMFDEUzTN3UNms8x3OUkkaK12UroZ69JBSyyyythQbJEWnGXk+zqhJKywP7/8M8AwELj7
6M+paL+lU9IpJtKkudQu13H2rL6WwuK3YVVTf6FQxAqtbVWeHNzkYZ2oG2D+2ErI9mChfGwd7xuz
AewOklhP3Mr9XFQU+U6HKVHZbBMLtaq0X2krsNVsXgkmkD/2Ga/zhbr4hU1k0logRw62s/sn2IVM
+LEeOwfp07bjRjChUqF6fzl3IKlhMtu7uMc3Q73d+5w3pLtXRmzWkU9zvdPKi/+N5esaRn3qGQjt
kFm1NH0z74fY8iZCdkOQ9C23i1blxplagFqnocYFHaMYt/nBTKoWgCasWqSJ6nliO+VJ3fgpuCC3
wIeWExAO2N+2kTxLopbV9T9JjuBkXBZYBxOnPLzCTUoQcSfChA4NGkP6ruFCtJBMgVkTYjsazT/Y
QfjigSc6IbgFaupYOGUKI8yl/W6cdyQfsG1XoEgMzPfhpwViE21YAVOddDHlMGfvgT6Zad5RAtYX
zwlDH2PDVWIhY43z9xuR4ckG5NwX2Y84+u0giytB6+THWhIADfW/ocjQt/Syg6U7PxsAWMsiSbhJ
rrFwGtxLW3qLloKOJZ2aGyqWqkaumNRx+skmWlbVp52A5rtln763LdlUqpw5OJvFJCUD7rpSWeSy
7juuLHhyVeCjwWMqK3EXkGey12jYmp1q71QuX/W/Xu61ErW/061xXUcXe0qK3t0XeslSE75Qrp/C
gthcRjsW2nPlEzoJZooVUvoNMbxU93dMiXO8T1s2OvN4X78ngkQVf2hTAPEH8lPY+5SXZXp8Xp7D
mjoFlRF4rKYDj11kQYIqYic1adDb1sMDVOQdyhoMJBspmNT9A/FLAIrRFzpN0BFaupT+jICkqTtU
Tyerc5ZSiejCy6Twl7YroEyXetdko6/SUrRV+OtDbsTR0157xI0UHiuBnnX2GWkxR4DvYtTCROGN
ZDvbA9t/rAzhjG+CjespLJvV1QMd/nUCKCPZkdwLf3mWU9a3Ph4ShSo451ilHtXeDJeyhHzICB8K
nIlsHuwsWXF3QqQv7KQ8LXByvuJqyffyhxtiAL4G+LaYr3QTzhKPCNxgCs21G63DQwkt3tZ1Z59A
rJA4zqQ52P492n2EnLmbzP5XvABV14ProgB7hNZLsHMhBLxxTkZPnf1CpLw2MFTBcL/hCPa2Htmz
oRSi8d+SzTR0EQUx7+QjnYcDURYay3EvpAH1SrYouv6+Feul6/4yGR/sHfflcVQvnmXPmiOpCuzS
xMtQPffJpjD9YANtU6+d6P4G4+U+LAS/82k+nMWqxQUVSBEY+GyWe8mqasq/Zuthdv9clPyygntY
KAUcg1kOVJIGaWoPiYm3VjL8GWC/vg39QMc/rIaNf8AFL/8YflySXLN9KN6Q45Y9zaHfjOISSMFz
799eUTadTkRfJ9bDj/gnwjMaeMTIBCkVpZUX/aIyy5EE8DDvFxR4wkNfF6b5EtTW0c5yhzw3YyLR
xQvdrLG/0U3quWH4kGuGEb7U4Uijqk1FNWkaQCSFs07tkkSy+11A6VcAyBwypj9mJfFbVXUu63WP
I3MzysAdltfGIF3vaP4/B1LCpMpnkHoZ1iZK7f/f2KTpEHwMA2VxuYDIfLiWyv8qdoIZUPQEZQ5D
pqkHAwGS+QhWZM8ktMYFkS57mtZazaZF+fUKpUWDS69LooTag3zKpwNudPT+nTiwg+Q8G2VzadHJ
BSNjj9dhtgzEwJTUu2Nvp+R0+ACFUK2Yk8900r0W5GujtNHKij1y3GsFvCMdv/oRXESTT3FKf36H
hRhUjfCyZNX4iA4p2gHuVX88F5n2M5VIVsDNjjTFhep231mRlJzuPj3oUhX85y4FJZ5rLWpn8bcA
zr/Ip+DZddOp7HQdF5WZ964YVnenVuLTQvBGo/BROWI7eHXNzVCxxjnj8E/G07LTf44CGgLIeZ8g
j8a96IpLu0cD/2D63i06Cp1F7AbsjfXaLpztqgxo3PY8lW4A4hLna0VIlDzLiinxqBVJ2MmiYSBc
ie5pdaoAo5flPm3St9+HfeOJRQ5d2+HcgBVaxMY+RGcXmvox4MbiKId8oXlcI5aKmmv8b8rIPfKP
Jwplujxe7meFfm8MInWYqcShgjQ7cLDsm6jFFUIRMjICWx4ve3hNZDWLxw5sOTsvR6C1ivzVF1K1
Q0BeXcu/Tt1SO1Mh4U/D6rVLzebRuuxQN3Oef5cjye0Ttmjnay+xc3UmEkG6wEk2OwCZGMUQU0/s
Y1MNyqk6gvdZFmjPSiIiP7LWH78mK75op2V9PSharbHGWeYlO0qUU9k0ed1bg4T50KTvkiVbu1l2
3cpLLTsZJinI62rXjMGWtvhyCENm8/8YFtGm4Bl2pQobYZEfADnlEu4j1nDWiETDFzStoRRoc4CU
PIKk9bQmCzkBTbgvK9nkQyMH8UmvDaZFv8+zEZaQo66YwsPU3eLtOX7E90ZjI9za4bniKgOx5IBL
vN8b7+dXzIzQ4fjfBys+rjX7JPajB7uAToZ+SBJ6DAJo+vHYp2uvqsaTCoZcWNBUGYV+HHoN4QER
Z8IeSnpZLWizG+j+Cbg/Rd1oyg8Reuha2ONVNqYgi9E/HwLwtewQE1DRqkhbF29HC3PkStUFsSqy
bMvKWHOyb/lWvuyYsaeetNRge/mm1DyLp8DjBlw9E1L9Uzj1bAW4xdWqM2537P6a6wqM5lCSOJUY
TP4z7xkiOENjRqX70zAjr5K/IlAWyyDRiQVn1aAHKNbA0Wsl1I989YaVwb0jeaIF9DIEKKNM8UU4
UFep/0n/0i5MxwmCoXepjyFRvzcqrMTkLLmhKNluAYMhQh8AzSOIZJZvp6VL3A9fYhzWaVBv9seF
k4eARQHsH5OJ0BqtFSwzc+YkpUsxi3vpOch6SGDW1Q7Xw5bcooC7Hmo4tGChnTe3FmoRYqJ1AgkD
2BWnsCZsCEnvF+B6H0omkdMLdHzGbF9JgLUGEPsrVTZsxB9TwkVsRwNUJOwIecRiX56rPAA4BNaC
bsAJm7OG28yoqm6DXwyZZCOaWYw7Z70iZt492GJfJhCYilFfWsrBTXstjJfXh9/qaHCQ0k1AYunJ
U+A4GvJscxMIfuzkKK2UVMQIJsNGQLbC+jRaMhYc/0voi+hCUDbB9rdEn5H00hX5eXV8AT+nNbdR
rOwqmTsrj5rAiAHSH6Myzu65NsbxtAqU1/PZrTan4YBj/KkOXcAXzGoCGWRHOTUAUGs2FFe9nUmb
3izsOOKO7NTl8shKdAsEpAxMi69ufLLjgB46oum6F1jX716rVkZ0maPLLNlaQi5jk3Ysq0cOW157
3kI+2kI1dEnYoslrRy7qHgAhYmH7s3lEtZ9kIyO6OYG/GXpudsOKg5GLdYF3hgcoM9Qrn4pSKCYW
Ygi6aJST1wqrYwzXUiQq1nWWUChsoHv49nT9FfKIAYUkFVd2dUtmJhoXS0nu1jfOUaCpE+X02/UZ
UOYUHu7Jk/FwQPJVEMPSBEgK5S+hbELbEGsQmPfb7bP0tecGUWBGaMGgGyPp6KdlMCajIvAqL6O7
LwVKSzKsSe7jLBP2RKqG7Ct7AEYJp+MKZK5U+i79npGE9RfmP01r8KW4LkJpMMMIupK1Koq4/HSy
quV4ZVNMCCNSiZoITUe/OXmiSfeknyqpQiibglBrXZiJ855g00BPJGH6L3836UHPiSoP6xe9hvhm
9KkB+RqRe58Jtc2tvJ4qag4yhISXuSfja5pLQWPOtL/PpPgmmER5oypEg2oL219g7ptQUkGyQAR3
O2LJF9f3OEH1cbitdolUg8U80JWKr31Sws9Lv4aNwruzxbAv97jdliPGktewU2Ewj/O48Oof60Yv
eKBP9KQk9sfH/YAfsoB1x848wu6LgM+kY2RFJVVycvF7eNArDQkYy5g9mkazgBjofsD3/eSV1WDg
tCTRRif6X55YBsPQzxpxMLQozFHNwSo8omZCwujdFMeDmAExiCd7maKYg0vKTROg0MC3lvyKCgtc
QCYzBEYYhe1HPqn95sFNOTNReBebuXesJUvjnJrSG6cXZIXSAj0lPvhLG1maJd7GfWwDjA+kQD1V
mtwfAEEKVs0P4UDWc44epFqekFnJhiEvoYSHRVxZwwsOvXcwAQA4XK0Su8vx0RtfwMZq2MAhjK0q
KdE2Ch+VuDwDNzbVZcGPo2UAHpRpzzs+UJKhis+NurNzPwk1JcsbeBkWLe6ktmLLBPg6Otdg/Sye
FLdZe3mn8dZPHpUkhHgnneL76pQajWau4PkoPO7QTb4fjm9/j60P8U+M/NmlX8Jv/F6wWI4KnxHP
XmUv5i48LWryu3d5BEr3tyTlDBoEvMQNMbRabTojnptc0qPTKBNSTeKvpkOfLsfZ98Owlr8+Vaeq
t5Vhpk/khXVSWOFBZ7ZjQKz6TL1B41GVrvMqA1CQyr/lbRa7eKKSvR+RwsO9VuDSZv1CLRGuNgoA
p8GRpuHKpSEaQdL4SEdm8ZiCos1kDEd+KwWMaGWK/09xitLUMm192FYt5dfzgylwA5mLJMHRIvfM
yc5tw5PIjWFHf4kvis6CGbV7fsWFOB4/PxXJW8Nphh99dk5I7dabeet/+iSXt9CDwg6+KyY/gtZg
miF3GknIIDRmb/tMwkdkfEjbigEj9GrWKQt6A3veVw6oC4LuwZbR5a9FhL8xwHv8wyIY8VuXKB4p
+PDrwhP/DCiypHshOYZxzPfB+sesfdmf29JFnen1fJJLeCri5uBr94s3OBzqE+qkWn2obmJW59mX
sFOCk5kJL/Uc93xmbvwnyd8wD1l7ZaM/GQF2mJTd7g/y/NlGGIvt0wGVb0TK6QjdED4vR8puHwsU
5H+z36Ko57jmzAMqNctgj2gpG1x+e4zayaG5lziIgyII01l1K9ZVd4ARdDOQDSbGNJH/3UPZShIa
w651/YU0z7BsBL+i1HlhXf/5kAxjFSMWOKP3VYiIwjjiQdAsTuta8zKwl6/wcEy66aszZcHWqQlD
Pd50FctsZG/IoTeGt3j/9Y78iGt4VSON9MUg/OvTdPJwGYvbyAVgvgx4E9eYMGbUijxUkqjDh2Wy
DBV7Rk1JdXiO1yjV1bhFcnjZ0DY6nl1d5tvJpP3GrgHAm7xjZ49XbcIcPN3LOXwlQx1vGq1EbUrl
FUrRe8c7qP4rvmF1Gdv4s++ZGZTSCAo4bULQcEMR/cKa6yUwxHQoyGhn3qfGraohdNHivO2iqavx
v5W5AaADlL8GPbMd1WzBrNvyfqmmBi4zYI+u35X4CoQNHIfoRFkymsnoXXxLYonTi/kceXFOBcuy
mutpaBT/xaYBo866AJybCVhQcMiqgA7iYMGyrG3La/yD2vWNOc0NVHEL1Pn7maA51XO/mfW9SW2m
2xRGYvjrtIqJEmov6lNIFPGgQ05KqyDKkVctZ9CMl/coKNbIAtQF3z8YrsiM5S/2y0GiN7RXolPB
/kN4U0b5dsQKNaSJ36GfLKBhoPNrweZs8PQLCkc4xexS6ONJ/LXE/9bQtltWjKVkP3pVMucjBWab
fpN46ngWV45br8jUwbLMPZjB20BKzZYj6rAJNzt52DkKxzHJvOh7YgNDWdegFiqcNSLSDI7ZASeN
ceOaJrBXvx/O9Btt5kC/QjL7bHYM9l9JNvrjECom48xotY90isTxqjuOL7ptHGKDUfuCCjuwLK1b
F+9avZ6ldVQdlqYsEKdksRuhqUF1w6Mz+B6d8ughz0wSXRDX2b7AZ8f+ZVfj6/rijLDB47rEWAoc
ausV8IpqEg9y/hnkwq2M6F+PAsSRyOBNJKI9h4k6CYU0TNEE6Nsnb1LFz+hFA968UJ1sXZ0rLxtD
uQimfUZyw7lm/H/lgqhte+wN+ie4iqnFZKAYqoQS0cptV2TqNaTfczu3EHXzWQANO4yLR6c2YlF/
7/x4nRKvPslv7mqKJsoVroFjk5hQ2m5Fr5iLu1dMiaZnW5R8yB28fx3KG8717qH6mfg4W36YUPId
4Kra933p0D2YLo6mqxBuPbQIldQ/hhf3VkYZbEvlsSjGK8fWKDfKQvKWVCUVw7leH4jt41zZK9XS
KcyD7ey33OzU9sCLHNfGvZ4QxK+IlDoskZQPO8WUm4j65VcTxclcA8dhWnRy9+1vy0SgKvVh5DwU
P/+bClKHa9ynQYGbDGAQcjHnuvMLyrFMZa5LgtGm0428VyEnw7f+JJu998Fj17eMh1hC7UWlQJAv
DAqyUxgcR/LVKIBQfoPF3Vg7mlkxkEzQigH02029xKb8iE50aJT26CzUKLVAsZrfqCnL2s8Fx3DK
4Wxk6S2F28pDamnJiI8w9qpdAiqahu+zGGVSYOq6RWMufBGL6QANjF/Y5rBlj/mVXY+lbUBetELL
XHItAkfjXkqSLcXhk9nuQ4G7ipPvP++w4YncMLABq1P+6N+/2e7FAX8/78C7uuz0+uJEHob7qLDE
ddIWxcXAwSAsa8B3g9l9SKj51flwDUaWU7Voqtmwf7Jk6VI78Ak8mA15eh7Xjl+Rzkkr7vxHQDkL
gMRD+41roWIFYAb7IIgkDMqXHSik9dp1yB5c4FH+1t4bEd8KGh2MFiUbr+1JRVE0cejDQn1B2gh4
AhL0X+Ldhu6vJbMzfjpDG49jjIilLLiEoXs4kMcQPPCfH4EzYF9safuq7lxsN4lb14VIsUwUbdgA
mzGP0cYccbakexZCtB/76OVBxhrULPfded2Qc83ypoWPdKMfQwgsBBrbGcuvh2Kkv7VRiE5SIZsh
Hg/Ug6SC/Dqb7LYRXEC3+3GNXnsUSk73pPR0WWdydCPDpSpjsxoA0tmKV21Uskofr6JtR4tMqKBW
Pa/ZzUKBY84ivCeMDwFgNFJcYFiv3IE+O+4EPOmyy3K3omLkZ8PnD9SsSds+P1Oz25q0PpJ+EwPf
D6TARoRs77hwk6jVloyHxGZE/CX1l+Vyfx/CCQE/sz2Xc1Pem5XjW0XzaJT/zoVxtwge/AGxG6AS
K2IscClUK0BxxOtbjsUpHagyL62mLP/uFeggKm/bfQF6QPswyr0rKoWuqbNqU3/GceP0CvXTPQHv
h7tgz4AEme40KssVaI52pVP7argeZr4HOJUL0lUJxFzkNofR/kgpDiSdbH8jobIcfgVzMNE2tZcl
aJXcuwkDsPMVE8J3YYHTx2daFPbTS9ckQas4tk3Wnptd06Dp+Z1bD13FAOIPOA7JgdEHT5/xvpPL
nZ8CKiy+hymxgzDIXR5Kr0j+Moci/9zc7hsuG4cCRfTUnbk2pzy1CdxeGYQApbOIkkV8bbAB+xEo
x+P+BuKorH6EWnQXpoEhm9w3KBSRgN1Uo83PmnDLbVWD9hP5OGa617wWQ2wVGAW85la35kLkXmhh
MlVx0AfqlXemKxG6ANmX0coEd4yHwElllMUT0fKxjpfNQv+UcwctthMPDt5CNrxBUQE2T2XdNwmz
bJ1J/BzJBK5gRHkd2QIicVFmat8igAJgGarWYMcZksNdTn5Ti4ocYrUrFb5Lqs3PKMBWN/fiVf2x
ZsUAj/GIqKEj4RPfKb2489UL56TtoxNEM/EVncOB2XYS+B7a6Ghc4IAZnetHB31zKOAS79fskdkG
AjiMw7GPdhBXRam1SkaUeZ8+AfZ8BblTY0gWFoF3kswuuSgEvHBIlIjIZNenquJ3ukeDWvIhR2U0
RfBz7+4XTVc2+nwKenTkkFKcRH1M5HwBFYw/BOdbCt7GdcZGSXwONiU5wt/LeV3gBzAi/JpIOaLg
zz/OaGlxReNASpFH5rNQPJUOMp3lR6NShl9JmG1o07jsJm7dz1tojEZK9J7NRAQjoJgImx+hOjCZ
FUM7aPcDYtAfR2BF00E/ZphiyrRsPbC2bSvXs6fuKhS4IrE/cfaHUsFPXwJSJnztYUls4JhxAFyd
QYMx96Az5TGRyylZXWuZhSq1wOzmjkifr1Qvxu1rX/o/++5mqXcGy36CGY5mI0sk2nyYIMZ+THhK
nf8GgTJ01UWpMPB3KAOwTG71TwTUbnlclF1+XD8f1dPX+zxE/6RHV48nIv6kPAPqUv1w2K01SL7V
ElffNB78RsPFB4bWE7Nx1eo/hN3Nq1sd5CKuTuqD0Q+7/IoXYU0dSdPIn4nd+T10ob5J3ydINIJ2
tDmSlCemQaT/hJtEDuwQTcVnQ1CSOW8zVYDwyLbOuXpVNxm17X5CCxtu935FwX3JIUbnABrSC4Yh
QoPd2S9FzfJUfGYS88LWnAgrCNo1ZI+8E56VoQtH1ErJE53CGltuWYWt/rX22lr6XXZvlKf1AlsT
gbgpx4ZNq1uFTm6WpTyud+xsrua27do48xIZCtE/2rIVYdW8+y0vXfHGD8C5Xx6USnpTqKQW1N6h
0u3NPnrZD27b1v8gDvAxn/L3BBQP2JEhBrHzmTCrjgtLLoxzAPklcp2ocvKXKwGVI2BvTN0cInPI
N9UrYcxzSZzfzQPStneMCskBKBb0QUgVmTChbpaR2V5BQJn06LdU7iLzlUjUqG0XNv0ifL2tqs7N
r+LKBPKbJXYWehFLHRd6aSwi43TyQJpPA+bLLWPvDyoebjdgydj60rnglzpPzonhVocySwNPcx1g
dzorD5P5S56DZFFJ95lF/VL1E34M11foygNga+huPU5xVbOxUYEG3TxOTkoeccGZCop5xgO0SDgS
SW+ejnPzrbLfh2CkpzmGBszIXjkRAv40SzqKF6nQBfaKJPDx5t0usANPaCFDNLaLdcMNg6QFGgw4
sZjFXnFi5/Ee0C+5tCrWAILuMacPd+JeACxndoAquDl2JF4TJNBt804yzY8/8GwcI7DExsu0Ywad
H9SaWrb4L73acCT2UMdfQq/1BFC6UzH6lwvItBupxvcYsK8RJRU02obv4F9DydwED0dE+s1Bd99G
yLUpr1+ji8MdpqNdljhfMfded0pwUGl0febkiHaDfEN95kDdFN2JnDI7qN/rl81qFCs+t1peRSEA
erkYHKVXOKiaBSB/21fWABEmsZ2UCXAElviP15ToJd/dHeQ8GpNjRhAPrFpwX+ktro2AG7mQnU/o
sGOy5T5lfxixfzPBgjJ+5zIhO3hMSaOKeDuWzZSaS4yo125RZjIkEljHflT/N3V+x8btTUVK1yDx
XVsAtqRb03hFdyLHQEG8mKQrIS6iPAJm7pZi+0cQvn263c8XbnTZwtYMunTEOwwLFxDqA6aaykjd
6V7HaEcd5Vk/38d/tVMeQISLAZhkUKD5/O/uagVdOPGIklIvQnlappdFE+zX8KQOxZ8xxn5Jd5UM
MT/zcxTUKfuac/EGDDd/hpovPwvG3SXPYXWfytdSEzjlh4M3fEqc6ZpcsS9yy4NzvARR2jUXjonO
ggTyPe8nzy6XylhtplBsqUyf5AbBswpy7AF6gB6rar8Ai8FLVqj7J8CQR/EjMEdrAjxfjMEtVG3v
6XINVrO9hLuKIZWQPWehgBs/d0ZobqdeaJhacR115j3l7u/FIFGY4buT6a5SmIK+zOjsH4Urp23w
uEPn6eNhqhOLa8iFmj7vMwL7nhvDB4nYQ7LGi1HZwbK4Pswylzwqc1AnbgyyBVx5MUgsLTG3LSCh
GAtG1xOi+ZrrA8Jvtu0gYiK9Sj+PcCcCZEB624iCoKySy7v3k4SU9irJwfN10Dmm7VG9WBCzTRzl
3EwHEkT1jnJlqe62SOOBIqDhzDwcykBee8HUDGtW+hm8/64UAXBw4gOcGPxSQ3I+NxaF+2/GbAfx
NyNk1RW/g8l8qYuHGHK/Y1edQpUK5ClpbQ6AOXKalUnL//cnq6/ol6Dp5BjOKqw+nQNuITou7IoY
MTLgabOZjsa0BUGeuibQz2pB0f31bqWIeSf6pY5Cfljgwylym0Fi/GR9EOcYz/SBho08QQR2Q19K
EYUxw1DSSNNCgy3mY/vWaA4J7wwCufXxjB+s0s8W7lqYaefxdtwwJNm6KJbavPaff2w9bhyq68pD
BWSqCgcBh5O67i444bKeZX9eHI0NAasIN1YAGcHjvL6AxwhggQMuFruIETtfd9PPjqWAzTUTlq/U
o2/NSq/ahYcn8AJq3e184qSTUj8OkXs181Y3Ri5aGVl2eUt9ZvUR01+tc4HwE/eruPHo93uqSajv
6Q4D0/NKPh1VDOYYkjYp/+zb+ahPZbbUpNk7GjIhNUsJV+dTseqmP8R2RfMneVHrwsuO77JLOqKc
ZUcKprn1KXXjYcJ/tMvymDOQgdWes/fAP6CSvYlj235oaHQ4eHUJsO+ebp7rmTaCYuKENNTntUL1
cGba893nES3+qgki5IBdMwBYio93ekQG30B6LCHFUDQjOrUy0WUeXCyQy8WLvDCj7G9R83kYn5GK
cuUKEsXv8SA80CmMn7o3GwoWxrdDQ3mKvwJaCmApqFp8zERDoHPAzJg8BOAc0buUIiSHL3Dk97PK
msF+6A0WyND5qsqLvc//Rq6y8hQiYkJhBMu6mCJ1h945uST8SRDAw/gLCgVmtt/vB+XJAHlvmH+y
9RDM8JWDWQl17efCKlf8S/6DRDGobOg1E1ZCWrHxG0dJvIak/kQYLjbTJuomWTbcjQ+bSHBcw9WU
CLcJYYIrEgVg2FUadd6ZrMfV7ujXGbcKEyziP+O41DlQI+hmHlL2v9Mmebc/EMvqhsMCd37qpPK/
nRB27pJOsB6A1/IjW9jYLDbOAs6vBC1ky2I7EBl+OzD+mLVLg3mm7zSlmCZSolcitUbDgrze3bC4
a07MlKfx2+OTUlcBARrn1W3cU58Q8/U00PKj5ww7e4C5QCSOSnWBcxTszz3eM7MNL7qewNYUB5pP
8q4hJ0iFt3P9C8I96ZyzsU2/ircjjOoXTIsUtwgCKq5829MeiRZGqSqqNtQ8zVEIgmKdx3aqt88a
6jj3HPfW8qfkxuM18VBHwwmtaghya1GwODbu2RbnLEytCxxh2qr8ikBMdErRO4YE8m3cgbZBfY2V
4/PeMWH3i0bXcpk7aanq5mWehc2HuOygFmarPvbJAM2xFaGRxvWQmFgw3fqZs0dYi1IL2LT/WE7u
+EPr3/LlbpU7RLfd3aLtt0uoLjoDJMFfI46wpTHHjW2xHhKTylnNe8TMYGa1AYg5spZMDL+Jz/cX
LschwDzfPd1cSFoLryABPWubbacOLIhVF8Yx14+TJkSxNY1Wbu9dqWZYOLUc3LKDZncoy4fVt0+v
f1WNJEqqCdPBxMykJ4473S7Y3GkvgPBTD8cyF4O8DhHh3ixG3CUC9jdmfPZt+spuHxtfSWoD3LIX
5VB2UYJzdnnPK8R3kRIZNcqikr48lSUdGmI7B8QDKyM4LpZ17/69JHo5HRnZs3tV0f1m6fOu6rRe
3cG9US+0Uik0WRgbHhvgmoxNS2t+WAdFJE6mIuAGEa3NBtwJfrV9NN+EqEHoDhG7+fYfz0MWM9tN
yyDFIIRHEBaogfvDltiItwsBxbjGuYhp0wFNBpFwlG/fAuRl5P7jj9Y4TrU/1vQwMsDi0BPl/qLw
hn7v8ZkzuIsNf6jmqeOck+qyjjSxA0N8XafBXvoe2f3neY3j+XnvSFRsSa1vbavL95Yk/X3kgDLO
lUmXIGIXq0l7wSprtaX1tviI2eJbS8mvn+7dFEWcf/r24a6/iqgDK//lIcKZbHe0OgpLFWF3shHb
2nQK4WHT+Y1CcFrm6adrygmMFSCHWEKBsKgrHFIYXB2LkdnYeLW8xIR1dLCmK10KbnIiA5Zq/oIo
pQzBxhAICw4aBJEWLpShGAfkW40ML8zNagBA34x4gJrxj2/WCrDFUI8C2G1aZV+l4HqkaOaAh/J7
Su3ghJwQq/nj7YWRnUmM+Scw4CgGTuCynN8n9iD7LkjrJInz3yn6bPlXvE9pqHmhVlyFfS2XvkCF
uvSbaNjcLQQDAVqVH0LKd7uHwedmR7kzZut9kX6YrTc+GN6GNn/nYIRlmtiFusWG0LKms3f/E1KU
SoXg75expXkJrAOfTlB64z595ZFz94PJuiE+TFmgwB4geJukNNaOipDTAi269qw4rd8EqlS/zlT1
oBSavMo5osjyM73UCp/I20Xocy0+USf5i6Ma3S4Z36gvZawczYw/sUepQKo6twHuYUATRldGgOsQ
4ZSPKDgRc2u24e+dpzWNn/IW33EBCaUliwZouD43Wuiobv/0NwH/RJTDMgGWYNgjCpLhbJXNvOzy
p9arcqlJU3AVruo2N4gF9ppMzLhpck3Z3AWRDUCJjyOIIGXXoKudOIV6HZJ7DfCf+m6sWcWtnJ/D
ihAvYqwBVdWbg7lXZw9zRVHgMr7cL4yJ/X1izurZ9zRGT7ZZ/iF17lf9A7Sa9SB62pfmU1vt8rFZ
E8A3dHg9rY2cVPEsNuqw0Khxj/iALw9UVIfNSbQTYWtnLMNIuT/ora9YaXF0T4SxtAbjUqyMb1ab
bSHvoWIhzkoQ+VS7UtHoWcMp4fWRaysqU7DLD8Z2/ZpT8mRuK+eIjurIgxn54OzZAB4uU8/qZ/8k
vid8c+2rmM0/kmv/lgoxUGm8+bD/LAX/9AdvXas6jxXk9c2rHTiuiU/8oCxKPkPD6NohXf51RDGO
sN9iGWOPFWhzEm11uphnb3f4x9cvJc4oY3CsbnqWh8BaYPo6XyptlsLT1QwqHfftJrtSAGG/AuBj
leEhOrAzAm4bvK6K/puou6fM+2US73VUGCzrOKT72pynSuiAVpC8nEY6J6QrtVtz3E+SHiup0AjU
NEKOosREK93XG3XmRZRL48PPMLaR8hJDkAenKzKlKOpxNXa1g3aq218NvlaqmkWTyWy9PdvuzU92
F8wE9JJDmNxtOuWMFg9Z5nRE9VQPjR+HegIZYDHB3LOkRw0AqXe30e+imEFz32AfNH9bjRjqAURd
/A+KiM+/65BHBw5ujtA1ZJhgiqPZAZC+XrdDz/QeymWsyfffrBs5rRXH8ISVd868RtIPMiFo/zOE
r/SHR27ZF1PW5YRIR+Yee1o/YfgRRudx9VPXwgvSyDVBOa13jSfCKmlISjS+uSbqHDPYKAiL7um7
KBDlfR7iW5/X5PulMnzY6hsXtOh829TXDx4yo+koEPycwV81Yu8iXDjpU4RquP3eqhO+ax8f+fXh
Sp3NQz4wsjFpOAsBLX6ThqcDuS5NFiZ31SMTJ1v4RPJ25tnYnk9uljXX1kTAgjKQjoXtpITrEKI9
lwWtnfdj5yLyy0Z1E135bPRl6Jt7PfCLaiN1BK3sDgviZsLMt+QmoETW/KZ/tBRDT5rZ3s/0MqYM
r/BEpdqItgi5fDaLJMbgSg3+tMR+txD27yfFDuHUOOz4CvIA4L8hKkw3MloK86G3pv/DIOl2LE/6
q0sFKFw8hxIDxZHKYVvwfQKKiL0iSTeFArtzdBbWIRaVuBmoQTwjWLJ3+qt9sS1e+faBD9SdUqNQ
TQWuyAEbwAmywBwyEhxP8DEbxPuvhgZzuGoCmG30wnufP8H/8AJMsyB5ghHu2qii5cfbOWT8Ebrs
quL/PFUk7ftER7q9rvW8NOaTzHBcRtCRuXoUz8lpgE8NvdZ17Pw/SAQp8qkHkVXMoRPDLyP6fFWH
tdUXj/GlSywONc0GD7Ty6Pti8k34uZOkXLmhdBWV9Nwf/VidIhNHnbYVqTR9vJ+H+bRnDZ+2lqUE
icZ4Pa6UrYzGh1QodnbNEj2MTskYyCzZLAtuDjOhidrpm7X0QhS6j7L4wGKAFzcjX3778MRQIZk9
Mb68w960JqVtI4Lyb7nierp8bVLg8qm9xXxXOqcCSmuo1pqLikWLGfow2VAVVnG3QD/BIvrBzJ9C
pTElyz+P9x70eFKKa0afAVk97qmOdtZ5iaQo/nTzfhWG0ALd6Jyv5WJLpKsHvIQs2KyjaEBlI3v6
LMQKDrKM8ZPIdztKkh8vYRP3TFDDAkmfwFgZYZxfhjUNTsWqIfwNNvX20A+D6Un/h8gdeeal6jHH
ZguSP6WoabkW7TTNYljRP1mLSB8UXzcWipE1KJOeRJONGUFYiaVgPMaJjDDoy1eAptqd9DJC4n8R
e8KRukB6S62stIn0efGLuj8eCicErCcA53ucp8FkA2IemxfO+ZzXMkF7N1IzhPMMuwnShl58QOcn
/jhR/2NZBHwdBjJCwAYpNZ0uM92BHAJe/UKnkAq1HRkowSrBkgeV7uWxGLgJceDdAu5KYNZ+XcSh
X6aDHYkBfj8tCyfK+hntRFn7X310vtNpuVQF1bDDP0UB+ulA8kgvGm8BwUmsHbP7x6KB7/xP7i7z
inRzKPv1fpJthauqv0e34AE29wWwoYrzUKRkYpQ4WDbO+1ppyOVfsQRntB/pnAdq+gXciLMEa/0A
MJkJeYawwv1zVoQrEFr+kkbBTc/2XYL+MtIjYEMvTpS8GLFGG0/9h6G0CWb/edA0GkJ8xk5Ub3oM
gxp3XaVxIBE1eKebVKPY6mBgsWZU/cVfbAxnG65gzyVFgh2QtgGBH2NoYUQdpxOVTv1SSiv+4Tgw
Z25tog+LB/mRFyCMuoqW9ue/BT+b/1T6AP2LsMMWv/Rp5mdzKHFLqkGhKh2caGZ7nN4NpLMzYOO/
LSIRD6F3Gl86Q0fXYY/rfs//1uMjdrMHb/Rr9bNF4o+5O6cNfMp+RFUJZFpDxJrqlE7XkdBU/cUN
LYy6ubFvUTW8JgHBHBn5YMJQkUxA/K8P8WLNjqk7x/xMDX58s0sE3Dw9JWvjq5zUbCF4I9ZukioT
Z9oYVF/F3PqvigSVVmZ0KKMlI9QlRmsq8CF18ZrvKPoDVMQfQyDK0ZmwHt+EAV1ooR1yM9smCZiD
eNiGUPxXyIB1EfERzfwk3N6XkrTlMtQ7jNmCCAETHNd14OoIUbJGcCxEbELP7DriS6XmS8wxBq3h
jzEP5hDeW0/qQ6SxA34z6b2hN5Ql2o3exWeHinpbDW7CG7llLF/b4DsaRZeR7XTWJokKT1LYpIci
FkSEjI1LIJWXYZs/dMsXQxz06H/bLA/EwN3vrXQit4n1dwlmdANdfvHlXsXeQZZwB9cuLEfT3XBi
I7ajm+VcbN3Up8HkAxBIDTy+TiEtLNjAj0bD/rDq6ZOVdCalhR/kfS1ulnO4A1LjWQCZi7l7aTrS
+UHiG1R8cGCLVn/b78n+3YOZhv7GZJd+ZmLWcoTeiCACS8KlgNaM/GQ5JS07XLy82ng2W359Wqf0
puPEIzCthMKhhbSkKICE7hIa2KETvXHlkb3qFBNH8P/YPHd80INqGSkzDjB/OYoyfv496LUGb66H
rhjjevPc32qqbpJuB6Tr2riO15zNBNy8uLFA/wrBJnIqFMZxa7UZrmEeQ5x6EhCDufNjk2tWsLpz
a+XK6YALROWVNhMUmCXGtFc4NOj7Iynik8R5B01ftCfeDl2MdvQpwImUlVyySjbnrGTO8kwA1i30
hDEDueGvCezcHgDj2fiDUQxvuas2DK3zDuZ8RWh2mTX+Eviq6DGzRQWBsnzSb4ZeYTZWTSuhq+3Q
wRyaX27RSmOUGJ0+MZC6VCyDdL0dutsUx6XGqXzSAS2c9e6O0UeuKioitjeYVKmCOWrHXN4Npp/y
L0q+GDySuSXcTXARnjykneZbYWFDao92BSc24Ispek1G58NWTMzRsT28PzHoK58RtDtRHPkNO0QW
J1I7jpO6jkWjs5b0hbkFDIxa0UfC+ZXSKEcFa7gwk4qxrr2zcwZrzsN4QhaZ45Kjjk51gECBLKkm
oKcaQae3bC8TY1Zvow/FsmSxSxbJ8n3uA7CmAtN9gfNtZLe806r6xBg/Ew4mOBXnI5oXB768KyJY
0F0zkdGREAQAa9fiHVk30WW9FnQ+W5OCV58zse3UnN2CX+OjiiL3R5C9e/DPyLsWgLoeiCeWx3t0
ayWNh0dlsLlTqz4inq3srFRk4ZDNPzjdeRxiF1HS9+ppBGNY5OvCZGUt0hcf0fRKWy4u2L/kr2GC
BPVIZMAKvRutTex/syABjnsPCFk5m8KMbZfC0bvwZkM8c8jaJGdTGCpZ/jiyXVTubzkGOLRjst1N
tuVNM9RFZUn7obMcZGjWElAr5LuL6kxxJxrR1K8JAzzh4an42zS3hdqbb5IanoW4/kerbvIZGdmO
yJqverdsApci4Uz4awJYb5c3JzVBH3L+tSg5OODWtcIAdja9th85nQe/g1i7lVIM7vFK0TzovjCz
0rUbeBw07FtbIitIWR6GA0ToxgiiHhqJi1dSEXbx9Lzj9p0PqczrYzvfsteXhg+Y34qXf8rhLJ9F
SAS81SAJygocU0DcoEsFt0UjEe6yXSZQme5H4ubn2YBxLtHfKIzmLzEnDhRXe/YPIK/NxmK/0yo2
iSks67o759sY4/lR25CFpXTTCfBvCHBqFjKc+uCDeMxaHLXBM2nhWR2jgT4l849cSQRnzodur73J
QmO6NxX3LfTcAPMO5I2QJu387JUxABsivY5O/bWdfXpnRsUgiBPXnTNTkhhA8RsZ6PiuZrspbUm5
22addS8LRPVzJzUEJklpsXVC3aY9/jnntg10gkoPIJi5Z4O0KzUf6Dzx0zejxdAaZDD1QHJMU4M+
FnM9SxbNmBW7d7nF1hEh0T32DY0swBeRgBFaEu/f98VdjTdoKr6RqGtpCxDPCguqA6oXR/aFCgEi
VIT4Bdj4RmW4tOTXlpHpD5onT3f8YePzDjmHLbVY1dS9HVgmuBfcnKTn6flIbF7ioFppu6TY/WCW
P3uyLDT7N9752NIFXTxN1FxpM23cilG4uz5MDhj/LMsTYIRMpiSM7oyMENkqFwjkB4mMyROUSwDD
q14ndIT+Ck3nmePdMoJWE1GY5f36dZw5S3OuBMWZ2LwxB18TBq4ZorcqrFNCh9Fo33jeHXvtad2r
7KXO7W2ic155d6N7IUe4CbT+2lUtGUkjXdN138tyidAihvnweDapHjBhJSCNwGkerdmrUiu6tBV3
hAnCBwSplUgkuSV1MV2jjXNNvfbeeo5jlWVSYOBoE/zZ0KgYOEoQdEW+Sfz8BHenyPOUrhC/V2O+
y7k3tqP8C/1mvYDfatRB04izhINMLI5mJZgUDRR3mG9M5+3JxMFkEl5FlZjy4bwQix2GfiAZ8xjE
5eN5P7CBMlo+FvaXWGbRkOYST+qLJuy6X3Y2pZJnpuZvjZosKwWBtDKZm2BYR1GfY2UhkxJzYOTU
kMcXhquYp8Lz52Opqy7pNR/k4wN5rWmXZbZHccB7a30M18TLPwL9mLs9pxg/USKRs1jmjKZ42SeO
xW2V6e+LCXHWmIG623X9UrX0kSR3m4WxxiRrKqYBdgnf53yhI+cnaHyrGQd/VHz9cpn+wY7eXioV
gt/+ZY9Rk6r5IVVynRn4/Cln/XPmbN51vT92Mo+G15KngI6bU1QWcbLSWfpg/CwENcvC+NZJOfeM
G9xpJ7Huh32t7Pw6P5J2zJXXm5jtxPrGiIK/rEJADNb+BR73wsm0zHeVxwxZGyfTK+gAGRa3Hnmj
4QfwrU4g8r9nUQjpWDBHxx/lYmyeVlWa6LHG+LNOiSJ8x2WpO4kCdR7XSmPW339amUBRBht92NSs
CTflC5/+89dUgxfbMO/WMptMnbnlU1c3b6afO4IWqZMNgR8w+L2T+wiBXijEJkAzBYiSbodN7QgS
UNBMgprWqpK//93PczePWNwOotRXKiJukxWTTWSlyEcOrtngAkxiTdM4YH6JKJillHVz7IShyPm6
awHqrNe5JPbmpwUNIciwpRj2JsfuBMr11MQB2YMOpTtTskvWURoXPXLG/4x8kaWqOQbRJIvnuH8b
zhPVO2l0YDJSKSbg0FDhwY2LNkoqDim2Z0sS/GAoUxhocUI5ivNgZ/YzNMVlitZuOPaRfjJtTJwR
IRoFkgG1LsE1VYonTydnkvQHPxQbDysxUjzdrsQe/J06uYS2149KCJjbzypkeVO6Xncjlv1qu6Kn
BEzXepx7JcA+bFY7yO1S74LT4mYs0R0W0PDg2mG0ba8LD3scPXLfW29B9LRg0RlTFPnENq4llJeE
YRow3104qwuHidwnnpQhDlphcBxKPY05EXai072UndwBHux0ZXqyQRLYiixtQ4oEiAoMmc2/KYWq
3QcQyfZ8rBZ1ZfRDJh28ajyjFHDVSf18WKEw0E9nf6o2LxJg9zpjtik3MvtqeWqLNkpc/EZM01LQ
49KhXun/fLNcBDWphQbQKb6G5QC4j01v6M/NdIZjN21zq4xub5DVsnvnM+69u5PBNPNdcShA0SF4
xalqIdK7nt77yQPXfNwTJn/Mti3A+2YF5fT0J/2Gcpe8WQa2CYaXnXdqg0KekQrkOedZ8/leB4J9
7UdOvuXHRPIpOBJuuG/9o6Vx20ZGT6poLInaJOC0GVO53ZjpZNJjhGbQ2uU4yKK1TICyS6beWT1P
DimSM23nNdvIBGFHyhGfxanpakbBIP47/5IrnAcstncunef38guzr7iEeJcPnxLz/yD0Ffi3KJW+
xd/hUyR5Y4PTikvaIAmhi/p8uDyqZWxVyDXNGHfPrxs9J4DE1DtPJYjGHHWqxHU46ueIp7KqtYYj
Tllq/exl+nptPovFEdjXjfMHlqze/QYJYSKukyv3p0ZcodIezQjHOpfUGLBr7wj4MNYcrB9FvC37
uTtop2mkB91BSRNPzgLbTlWmGBDfMYTxETPeMcb8CL6vdU2Z00yzJDKGA5QTByrPdHlUKh34iafS
z3KxXuhdRf74py0wCyv+ikJvErVeiv01UaR3OofAEKDCDc1Tis5Xt25KRTIQW891bj3Yb7mvZfIk
9TIyc71De7wib1PaVIw9Qt403uUHuSQg3Zin2pldRR2tZ6LPjW9UCwmlzpcXKamz6S4IZytCOvob
OFdiFQlz8UkHrJ6x8l7RdljUhUkG2zXjP/Xjf9vW7wgs/ncky8XNKo3GtjQABwY5/U5I+XLzH8Vf
uY5AuGRdwOWSI5nOM0DGHgGT73HSoBN1sZFfCQt2z3DWEF+/aNgnO+2v1hL3h+ZzcpPWsQegvdTQ
5SXHgDzo5abDEb72gntAHeaqtCTlrjYZFkg5YuBKW5J7AofeMbtiZxc148/GTupoUFEwgKjZLCP/
PueiR3HWgSAdYyocwozXX3whxxSA2RSRe5fxqDL8ZaBp1HwlSB00aaoKt+lFTovR8MowdpDvSRv/
+YpPCUt5O2S5SePM/WJgSxrBrNOVpKwb0txUZjmA9H9LRPrL3knpORhQeEKmSuHI2CkYZFZ01wOZ
ntxameIwPZ7ipUv1jPRxWvNT7MGCDL3VfUsDFUNCFWPpg6GFah1XCt9FwBji/pK4ecKqLRu8rVVa
2hN4ze4bDOvG1Jp5z2elZGCjrJ95arxK4AP4BB9rs6EbZGejX2PT0H6oAAisYWfF/Wvm5FznVefh
+jSDqd2uiKafWUMcHqvRhsqtk7pKSDoO3xKsJ4DLqHgfgKXiQLs72i/xVdtzGYYF8EPDIVyBfp5/
LaIdd809bCiFrrgHL3w2tA1lMpmrB4feEDRGVt4YENKT58vIQ8gqDRWopdj7RgnQ/jWelzwkBOJE
824ylkA0X6psBjqIv2xkhHUBUvCcS+srwf06tUx0DVv9Ny4qnF9Auos3YoqwCTvTwgDXvg9CprFQ
ojVYVXGq2ZvfxCl8uLkYk4lQrdSfx07Ft48UmL5MeQekljMZCJmuOh37euPPga07PgyJWY9q9mdi
NF4l6bZOdnKaGYiJ/ES4vAJn1zS9AhHzwVTI8cb2Mua4fO3j5TD8hTrzlwgKjfLeZBWFX42aqp/Y
BfGqzy1jdsxpiEvaX8OM/auV6Kl6uWisT/vfDyQ28J1UlD9ivsYJKyITsJxOlyKuEx9bglKtyJ8n
Ud2QspoM/x7s/1SNoJl4VSXCodsM0oMhGGB/g+rn3lLQEpUaVJDpNg7yWa5T1gmpTe9HFUI6mBCf
GmSdBlMT7/FTZEUooOkgkie+0WPYeT4CrBsNCVrKNTFLWrrzkh5TvzWOL3KVcDnQXjwUTi53+EnC
ako+jxMt6XIlcb/4JL4mkNSpWH5aNSVxnhdorjhlDx6bBNn6MvZYIeBSYhg1/1m2rAYRz8tYntZr
Doq3DZNsy1U7qV7zk+9EsX2hRissz+zVKgeRl6n4EpZuzvvNy8QvjpFiLCZT5XQwEz1flZNnTQrm
zSLx67KuGdqpEbzn+k1L+NQDJhqtwwlg9Ju8qMlCox6vyy9IHW0P5izbjMGo4Wa2jSkxdVajhOUU
IZpgsBasmoGSeliq+/fb4q+KeXMaq60tsqNxN+vKgbg2/Y8MQgFTT1bR8L4GtK1em/FzBZx2y8Tr
6WfiaA1R01HqMUz3HBCxAH86kVRK44Dvn+pT2FT46jy25qPCzwDNF3Sy7/zvB0FnOiEYjM8kVWWY
hN0N8eSaF2/AwxnvKppr4UsMA8ztMNRn1TGeG6XDN7kK+h7ucuS5JcCYIn78x3d0SPvZjrwXfqh8
CxrOw9r0CimHslTfZuUVNARk+WYBu/swdkOoLZAwg/fhP1edSbfo+tEVF5I1ADWVxwlssj3wvQLD
8iGNaIMdXPXZjfW0rLD0QFSiKj9Z2Z9KegSx4pQUsnmhVNT9YbZyF9pBVp/ZNLUjh+CZ2337rlB8
gghzDg2xqo9eQXoSU6IWYDU3zVs+Uat5FJcJ/zhow06QddO9n1s26Ny2BIt4NJdpANFjvBEjA/nF
hwXnpyqIIBfsFc1Cietcg02S0+ro0UqnWp2SCFUtvZrsLpFt4IAjNx3ZR876e13EI2GjamAYiwoK
sfvR4ljIpJ8x3AYcW5t2Dr2yE7te33XMFt7jmM0xT1sIauh+P8LNB62UsRtAsjXAouoqwZg6H9+P
fdwKjPZVjS9SXbTXtGtSh42O4qwGo8m2dmoh+iecI4QwBC4PXxJBYk5UQojS9mgFRA771cED3tLv
wxPfyQzkIT9XAhgUi7srenZedZme0qDWWRbDKHBrvr5htwnl7bCavjLhmHna4r2kT1h632OoeFg9
4J197zDZZD/k243AFX9+BtKtYasAg4TdXkAConoSZT+kEEZNVfg60XNM5zbThGjPFLqqAJbBw2TD
REKhdTIiglWCk7L3Sp7Zjps6vDHvcwq+7dc1tZDsg/Qb90fUeL0lg0xTPjyTH/TjxfxXD3eNOIcM
5oeFD2vokrR5WB+WZweFmtmKbhTRy5hXyxGyfPldA67SMIv7IsUBX1vIuKVrAd6NuQqvOAcTOY0Q
Q0yhRW3Qwf1VCeIQ7Te5/7ijSJtGVRwSk7TdUk6vlNlMmaLrT8k/NZw8UxO7Lm3a1Nw61hQJtfeu
qmV2mqsxBAKCVDJwwv/uRaZ14N4nUCpz6+gXQB7GnaEebOcezAFWVtp5CmFL1pGZjRiNuG2nUWEg
CbhPYj5GCDBejh0FqM/IbZDkLlPF+1ZLcMSPyrHSRrtnqksU8LOpYmerTjtq/AMr7HeQuBGQg2uM
i6LZd4ys2gdts8DVJ+q4bpHjS5bs2C39IXrGSVDL0n7fLErqV4mBDdkygzAPmNrmG9XPYugKjPDp
wLuLb0QZcLgU6K1YJkwHQSnEJ6rfFF4W8kxqbeu0d3idK9LPcORFLcevr/ePiEwslzzh+gCV/A/G
ajjxBQRjB97iDTjFJ55kjxyeGCeW+txbXPgjO3PeR/ZAWLyEEarjq6/RTxz2nqYfYQPcgvuVtabS
ka7s6snGThJ1fXYqxOPVs6OFQZ1NjthmLLvRmSzjkljAI4ymw1PLjWSPz89ziIS69zBajd5U0ioM
UDUZWn+K2mdge/IctyBstNt/3A9VCa2X+jF8C7MBTcRfi8f7xKLMqWGqip/qY1o7iPrA0cgQ4cVd
ZLP1OM9Z8xYBvt2Xsmw75zLciFPDlLfCn7Ep9gvQGqn3dD+UoN2L7yPylK0oejLCjElYqbepURGm
frUudh04+h8dGOE0cYj+THILC0TJA+Lb1rDS5RZYquN1uHykqPLqduCtt0IJsAQRJxWw2M/h1HqP
BjhbbZ9NTswBqMc1DB4IqkXzBQZR7HoTnnUoy79PvOy+OYTXLULSmwWKpn/bbEpYrc1My03EVv/7
O8CT25rkvVeXF6pg4z8f915+septoaGISVhqmXKuTKCZ3CR1aQKj9q4jDs0V21+jOP9gfwFYhBWl
jsnTiMkc0BKj+ilk0nPP7ipJI7QMIBI7ba4jDsYZAPK46o4IN8iK50A8lMY+cFcKewfckvFduLF2
7+hYfdqZP0G9PRiF9fMp0nNDtKiVx+YUbfuXV8Di5E4XsMKCx0vXCJBKBVNFORBXWbnQ4qKs2qFC
ogdNgUd20gK9LRD/xwor28kcf0cZaL5LqqX95LZOFFTic3niEnOLM9FwoeZzIidYp5dfu1wNDOjv
Q3AwR1ptYBLC6l8j791Q0vE2r8eoGi3I+PkWw67DxS5vRnoM2kyvnhtah3N1a/mxkV133twSMSwi
kzTTtIRqXM7HPX9Khvib9+22H5sMWLLdj9NC8atQDM2NZRnccEqNCIKeV3EDi107EXCGwDvAdDJR
HwSaqITDIZOKcmFXdk4eTyD9iI5I+m8akN4vAInNMA57wwtv7w0iAX0aQpIuxCAp8NU7rEWeAean
wMePrYmgWAlf2flK5JAtb2Q3QQbyX25toAN+18Nu2h7R8Sed3TY1Y0JoGfNYANTcNBkjmTWApO5S
SO6nIY9RL6v52bam738iFSeGaAEIIkW0Er33J6YLvPuoUZTWIbS/7c/OpJ3PWZhIbqhakox8/g6g
QDJqFSJOxciodqsoA1UTiye1cTytisIt97jdTOo3C0Zt4m5xfXhKvsgc4nVAX4iIyEFYBHY3eMT1
uAULQKD/Gbzt3Nw1ky9cdNEO9WIJFLXG4wi56AJfLLr3ipvImmUudjJJBB/uHEhluY85R5ItWYZG
9BOdXLsTTdej3Dz7csa8qrTWV+xNryr+VqhZU5vquHd+WOifMliswygS/SIEX4jWvH3mUaF9gFTa
58iP7gx+EQLZP0b8tE+UIFMl/pvVs/iT6t6bIqaAv2bhhIZw9yYGNP8aOgHzwRXLSdlbev+4wvkb
gVnyj9QbtRbtph+0VTELZcydt8ZfuP/bLny/HsWEMd7MBUmp0p69L67JFnNb/cT239aOZTbpoJ2R
tSjo/T7Sin8OoWEVnzcFF8jDoVBaW0ReXWs2pOs1YRyq6cS7g75qZj9WZz3+40ZLvupt7CW5JHMD
jmSNpsE4paRUVsqUle1LfHqxPLRz66onRRyBGSJxWr1v43ITOtuEitTucx7Q4pYhBF1JVWPoD/XS
J1TdW8MW3aigkxA3mZrlXTXnyzNsysnWREcFIGg5P1dvXLTOoGQw/HYPdSzExXvQrQwuhqdo0o8J
nMQeIYYlTelfyfM8lqPssa8Vhe+Zh501Z6Z3+xYXqr5X2X19me4mHiZuc8uNP8qE1GLOdyRcRP7J
coySFMoQoawnheMXqLtKfrde9LazGVsaWOOZAs+NmOaRO7ow0rkqvWuvk9tSj1uiT/lZqD6AOIo1
bz9VD52dlIIOWnXw+HhyrzNWkg/uzYax6J7kEOM5/SOi4BUEAGzRCvBbKjfcFYwbh+ECWqt+U6/K
4MZG8IRAXAoXmEN72BvNcAbU/5qcIByy3i9VAt50zZ7gB+jZYc4TxwQtVdTB1ABxaKgStwmBvyeF
P9vN00HJdZnnW4p3qyC/9lwOHLZ4Q6UqX99zvXtC2k9l4d7LmFzcDdf+5E5AtJFcSOFRSeRyLEOT
9mLGtFaXfMa0AXDXOvZvV90AJDznLkf/8XkEaf7DbKmrPyCNZjH2p+TSXUwoGuGQYqdjlDRrTRap
KsQGBbFdLwwEjlQ10MTjYWxg6Gm++n9IPKRBYFhNOSTugsw+b/qNCXMHs7UqbaCHOKDb8kuRd0jc
zYnLthA29LqZrkNUdRGn+WYPtBLpsTCDKlkl7B2xyzWLYESM7DMUyhhkhBJWHD7K/2BOP45S10/l
2v5eJI9vwEj7+HKFIa96eylFG47rIps6gX68UhH5cSFXbcunhn/6LMwjBVmFhtv6qp9PmKrrukGe
YWFalsT1WLorMyywonMe1C2iLA4QxPq3pOxFR5h0emvW9YeoybUtgEbBjt9JRIe8Q8WpPE26Nzup
GLvcoWsQWrVbrbt17F9a94G1zopn/d8O8n65J97vv0mhD8TVb2rfLkTnGeQd0AmaQOxoEnMiFQkh
4tzla4zktnKzDOcwsZ5MWp/AB8FhYRKskp+1HPqs6eWKgVhiyBgsEnUq0i9bqQ4DG8aImQWjYQWO
yWN924GquYA2mrCqw7U5TPEIhosKhplTUlQNHn3j5SLbDJKl7Y1SEB4u+1UzMglDhGyJmq2ICexE
ZMmc95yfLMvqrO2tUoGz9ZXWrgViVxEBVzHzen8PZIVqMz3a3iztwxDZkeeSMu2Hfa3BuSlgDo7H
/rs3BnJfB8ztgt+I7ZUwZhWM8s+rttWLX9vW0/I5o6xahLyN7yeuVC6wdgJp8cAQJ3wmNS79NZXf
6b+lTAK6HTvOf5ds9jV6qlUbCkSP87C3umE+pXkdlxHWerzYM05y6zB/EnYWXgC0X+PSwQqMYmNd
75tLjN8zCdvV9qR5/or7D+hP1USdACPThRzslHU2VysJ6mX31ZVaMXRF7euEPp6CWIKx3/LmRRt5
S0VvyBYRbM2/LqzfcUmxPw59WmP2nkIs423XxGbUN5Q8PX/3kcMLjZm3Q55VXi0rdPaeRIGMloS0
ZSsJIajSXEGJ76gB/tfa0e33hDJLrnI6pE9BrJGNfkOMSyBVRsobC43KxYAsKXXGaCqZPEsjQHoq
w0phlvQ3b0GcGJwqCNFgj16vuc+efPGPBYYGFaJxRN0xftZ8fAO5LU+aNKLmAYShtRFOKUnoLIEI
seiWAft3GGdgxb0dzfMPCYkrpxB1ysOx1fdq9KdMfbUU7uXMVD3iqTUXKbEpulmA/c4KFe7eivo4
Lk9YI9dC+SGU4frAoJMPhrnKYsUA/MFVEMGl3skUG+GWrHw+JKEKrdVp1yclOVf8dbHl9pUFXpJe
bkJnCZFM5EIiVaYb2dWMVymC9wqC3hDFWhxldz1WV5uqyKK07Oj1xrYncYZ9nnEylt3Rszx67HwG
kj1xuLwqY8ZOq2Ycccien7sWEUWRz0KDIouIFkAG4c9UjQmlKCWs+7wN2QF65Q1e1OiqhVjxSUt3
sClLAwgM9bp9YIO3xE9yql3Pus+rC9DbE9YrfGTPChVq71/7FtCWDtIAIkDR+E04KSsyg/LO28VX
jysYzI64u/IeJPZiCe5mDavPN4FdF4HSsd7bYi0SNWRRNV4g5NlnUm+ELs5aRGg+LKHOMrRbshjD
/VgBJ7Fvuepxxjdgjsv3k3/qJYnIJGPPXpqlY4NGDr1Hjw9No7bbRWJItfSYxPH7wjvQmImBB8dE
WxpbEkcscu3Hy9e/6N4+L+QO7OCmUm9ra7x5FtK9GQayttQP5YUmY3aFLJidU2EVmbyFtQ8/GjfG
lMFwOfuVE4mVBufDL67yj6z19/8ulG+/YzbaLeGFqe6WEu/jaSnJa8Xi9yThyoyLTB3HIVXBEQ23
ReSl4OCWDKmGJojY2ViEqwt1iJq5MAmrqrnZsfYxB7gVk0RZZduf09XW6g22EUnEMHGsah+pACE/
HXZObp+Yk0enokqzuG1atr6lmQTOEFw9J8wDwsi6VFa3kGscALAuXdjf3XL657nl1rKh1PlUSBd5
vbiMTK6qaN1tbFbEuSBAYQ8mr45EQg6nKIdETUNy7FMnTEWOtmep3WRSlq6AwFsKjXZT5NOiV5bF
SMXErAXdwZgdDPYs2N/BXPznwknCUKFN8DzcFdpOWL/6SYUtRnEybNZl88rAqrvnyz0vr2hNwJgc
iVGRM2WfxObXVNUoHXYXqdr2K57dn+F/VSGf43UNr78bA3Xb/tnhFSNC4rl1yXv/+hYPo/VkvA8+
BP1rcigu2T165IuOHtivpXoM9isT01dxW/N4h186Qfui7ShCiEDXifvbwI6VI08FOf4dbrPNdx3j
TPHNPe9QDlEV7mZ4XpvyOcDp67mDB9W3nNaMtdYW6d1Idsit50HU8KR7dtUvUrFuNC0sJxZXm8SM
xX4dVb+xg1bfqZFU4TqmUHQWhonEbV/u3QaH5OekuGXAnyaeIZWWYhGiTm+E4wsufsuvXrz9t6a1
/dNwFTbHHsaRb7zparKvN6zz5RmZYkOtmfS55opHNbstyPbKKLBRmN03fQiKBfxR/2PK1siCSkcz
8EZf8PrDgL+U0x1hul/onOxqKtgqPCnwHxZ31POSNCJlSHd1bZBNbpgb0wOGimqGZYy7Sn9WcjYf
RuH6ydeR7Q9Pd0sWi5gSTyoRcdcZ2/b/wc60HKCo+w+MSrOHL7HxdMX+aW5vSehKF6xuPrYorUdp
1MBCGdSWuuw3cbMu4nUXz5eHMyNZIE3HF8vtYzK3JaWoEbf2HNf6Emgg3Rz7Z0AXRP8M7QY8FUIq
ur2dFLWkqrcyEOqURb9jZ6c/TdmNuarazzXpDXtY/ellPpSiwKrU2r/Dz6N0Cz1CJiqBcRPidXnN
hnSRSDFSsj0r1pxpzTSUdyKhDb6FVI+rVRJUsDiliri3r/KjgVOL3YeB7n7WXTEwVUun2Tdp60iv
CLdsSPJgob/JvD0F2xNcWTRPRaxvuqDafQBm5RpCT2lzfbWlPF34X+IYKDq1/GAIBKGQUS4qwXim
Uukbvz02AEAC+iFgYp0xSUqH3k2UAQjPB+i3uzyBi0Oryn+Sfna64KouobXA19o1e/rOf3IovlTw
1hJtcuJBYqViwDlWgtMqGQkibY/i+H0wo8hZEJggdA4/2SJojTJ/26ovTZgLXiRpF0AsHM/El0Iw
Q6xkiwMCGHh2qmdgtrLAKAnyAkEFYtotdNXnzTZIYDVoQByZ11Hw0jZeWgwV23ACoAFOeOORf+Y7
RzUP8oGs31RSHE9E0/FH3eoeWOhts63ngBo5UMEwplGcBRLhomStumAoP0r3H4ADv8yub5EN52IK
rbPISK+kmYN5CiMPU+y66GtoO2uxJAqcO1Em0OcvRVFSRzZjE1+9ow8egMEnngxa4jJ6Pv3gPiv+
9qSZr6d8YXYRs/AX/EfVY/eViJmN+NL0KvOq1DyVEOEImiVtQLAIIy/DXG5yL8zRAT3Ts39y/EDX
Xu/rHl0sSxd0WCg1oRCZ4nxRWO1MQZXUtzV0sZN6vX1NU3jhSDiXELq195ZK6jkunCBmg5Ud0K7t
xIHkPKn/nZS7aRs0KsRMBfzWsMbFOzTit9rMQFgGsw8MOt+P2nnMeRJGotkIn5jsddAlxpLmbJ8w
p3TvJ4f0wGxeAWK0g+bHUE9cXeS9cE+dUcyGWLOcxSOAdsYPUl0aBC9DzJfXF8jaxcjR4NeUuaj4
D4BGIJ9GJldurEca+usAK8NBJdiz8qB6DIn/9yjCk+V9a6RX2qAZ9di5+6okks4NvxCKR2VvIlsa
+U4c7I6zsuVlJgHJybAnDX2BpiegFh41i2J4t6P+U1yj71eW8iKTW9dtCl1vnhgrWD1daYfNDKJq
+VrqTMpBQiExY8MFllQw2TM3rtj1x8cQWIyI1Y6fP++DYXoTrKKVrGUTJVX06m5nv9IRgLyUY4GT
/WiEcKanRK+Q4+iAEji4cASZ1OCDgAic5+fdolzrXPLJ7PcpQcF/jtNZ7ndfX9re7xpVK1iabke7
XQ6lZ+mXQ341mMw+wvdfaR/FYAPsEsnvK+T+32ltWhtkH0Dr2sdIRHiKAmoqrcCe0M58Cj+bV/vc
0hF764CaCnnKFwP77OE6kn5S6rdEsShUo4j4/FI7LUKIXcV+Tp+rpCZVVGmSziZYa6SsI0YLUjSZ
HNtT6KRNoKshInePWi77VtSkYSMHSDSN8tysMpv0YyBJ2DmnEtSvfEJlRa30kDLKDHKQxCgYVXel
BuagbSzTufiGWOtCe6S4y2gylEFbzsq28RvZ10pC1+0FxUJzxsTJ9W5ewCqTJERvQzDx7BFSxEUs
f96uc6L4/kXmlNR6/X7KkwDGSs4rctLsT2v3epO0ZzoPUD2Yi2QYHhG7HsvcyaFUvTDqt8MQEo1L
CkhXFQNeeMoba7BFBo09aimFiiL5St9hdO80ixzk0ATWIL9y3c6RHo2QGJBr1Tm83RwaNNccvwkF
LCHP2v7q4WC2o4TuYcjR6vq96CiYRw3Yi/XVOy8bMOw1FP8MZQy6mxrxWsSG36fnp3qhzgBgl9xt
ZgHNQ2tstdAIAOaoPQ/W8mcE20QEcICLFA8+OzPpmm3kmFJo81BOHfuwlSkCZNlQJrVi5WDfirxq
oFnBJO7ZW0uE0u8ELpM4nsZWGcgksk1C2i5cS0SYWbm3taRz6kiofKfCTigH9TUZf6TmCwmjMtxp
nm7lL87pBzpaVt7JyN82OLeXiBdcZq1PGL8g1YO1F1yGOeZh9nnj3c+ImrohdAt3ey9eGRPUePWZ
PdVKV/pRVNo7QehxCNDS3Qsk7vV7v3KLyWBgNc2TRP1efNex8na4h690K96KdFURhOb7wZ/mP0Az
3s0IsDckugDR6p5F8dUg3FqzwmDBxOxnG6kBMU+Yilt5Ct5YYT+s/SYtur7VtzkGaFoQbLSxk8nY
e/iMb/3JFS0a3Y9OPJvjCoFH71/IyIqpoXkxHrK+vNxXQjuaxI4W+IbkxadiHtpCxsUg9Ee63RmG
viWm3WNYUa2Cbl5VJuNPDmAQPcJiZvc1zlheQUDSl3kW6xoM9tUF7XulJ7ebz2X8gtWWWJhi7ttY
kL9/xXi+kDYbuRlPbHwKQxh4na0nuCr54OcIt6swBtbTelFuqyampaYzgrMYbLWGYRb7KD+n+xyj
zkjl8k2+1589q1TcRKdyu28UYGvTX6Ian0WZhFoIbkqu7gXZyAnvmedon4nMWa0iMQzEF5YoLXqc
cY/vi5fbsjn61CnY+dUFEuE7KgaMRhQv/qosx4txsV2b/rJP/d2Mz1ZIl3SS7C4eE5nNUFPkSQF/
RNGwVJao1HCzurKbjsTKQIMXr2pMewUHiXoQ2IPxATGR5FcATEa48JE73wZWqhdHvIdsdBgKI27v
/QPG8hwASGt/sV887z3qyqRr6r+lMU1cuQ4fiARd9RZk0xFwsOwEbxyJQaxQfrwXlsVN3e5/2sFk
5KeuVOCdFPJSZcYY6uMJqBifFXMxUkwvXWvSnlGFLel/2EFBkkZOsd8TVwlPcdzvm/u7WBiWZzmE
IdgIa+67BIQZKZMpcLU9EoIbe2NxCa2yi2OCXifdFNLOeOGZAvisTeTqEuPHqxEd/DyJEHiCsLtu
KbSQjDj/9x6G5tLNQDag5Zxyho42HY+ENDZKoP4TpAtrLnXiSQQXInFNapSaJIhmm5nMut3DjNdC
KikNjyYtusJCSUQDxNBrAdKxBxL6891vNeWcDRGN9FYY8+YXbOR1iHhva0DsvPrZ6fo/9FM9AQ5a
4lVJaNdK/dTP2yftqW7IH49TT9ksFrFG3yhycUZB6I/6fWoQhws009x/zej2qm4fnG1g5ITiyFi1
EvXOcCQLRSkdt+14ojoZ3yb+IDROto7KyQOuaIlxmeygu4ELPMy/iEyl1XH3jiK0NUpTZbpw8z68
phXMG2R0uN9pOP/96x9QZm0Yb5ti6WLzbd3dw77gcEsBn80jHyXszKFKxZQFY3atU6VhqTcgII5A
6E8Yo73JVzP0CiCb3HKHfSaPDggOqg8FzCcm1och1SkTs4yANRGz33/4FKvv+e0frZZa4s5gUlFs
pb9KxCK5IbeJSiXcyzOZ/fNvqdiVw2FzMveDs6SP4kGRqjexnJq+mmueUncQ016OqtWZBaIOm2Dz
eSCWlL6pf3622RUOc/Oy2Q8aNYZ+cyUtmjYL8bqu+/laQ2dVG3wvuwMOfc5jTtRNqYUTKkxjNfXO
hdCeBuKe/SYhG0mli/NoCiSPZQyOXNT7LiH4oYQb+343FgBdgPfsEwj05qZaaUSwIKfmV5sxpvBc
Xbv9GSOSUThP4icby+VJrI5f2RtGre6vhUEeAm+4Vin3yS27sjS/FRkrFUEaYIXDXixdmMclLJXY
g1X9MXzZMHny7hNb/zk4EUNGBHcmKeGzpv0xvT0vM5hqMFiwQvPktDbKkXJ525IGzckx10BG5+au
4zcrUPsFv9ww7LFtrg7Qr3WU9ZOJ8YfgC2eVeaq4QmUvMxNBs6nRWx+XWqGlXOMcWqdYRg3w+FaM
qMWQmwBeKJ/AhVHroACD2dqMaaAnIgjPC9CcQB7to9d5r57ORgbqyul4fE6BGiNA8vcpbbwm5r7J
B1fUUBb+SIjCMCIecMyecjjFECDk4ObhDiLw9FPpKtiuOys9gWZjf5R9q+jXqV56uMWE0D3sEigU
qKo6gyIT7xgLIwuQDx/V13UjIANf/IWhHXc6N3AMHWNx2IpyopdtLpGa3wlNnx1LtVB6A40Ja3Ss
IsUIf4ibjyodT3qBFrD6PN3YSuFGwdiWF8PITP76l8JMzwd8Ia8TNL7yAGoMxWlJPh/OxvR3IhU2
MFG6vKDiSKIWWqZmLrFsww1N85hFT/wnQfPCBteESZ7k0XK3RhgZw07T499llp5xIMX2Of5y/jET
C1nfrBRQIr32kmqZgCzXzbuSQOcmBX9cr3XsDuKBkHj2oxia6InuSzC7iB1z/lnJEmgkBYHg8SdM
q3PSdi1uJ3GjFZ+sFR0fw+IqoS+oKXiDT1zFIGZHFzKiRNBL+nmMc5UAMToQZtB8Q5dngkDIaC9j
vI4j4FPjh1vM6D4/r3ysF51ASHhbJ8C//7DZ2c4cUpI4M+oJSEnEtpYV0jdAJhc2tTak7cMYrhI3
Yi+sHNDV9USfTSIIiACwBEdbTbDJesIqZKWpLIBQtX8V7JxXQ02NR02+jOmAbJ6igtNTtKFewGHA
+23Rq2K3qTHCVy0VfRx+SiszmoYqPQn5nlCPzuNTnRDBNgrYKPSNBvS9pa1zMoEAx5wukehSEU9q
INpfg/4vY7d/4FL+oABbFzHFS/rdUdufVHpUj+4Q0YWidktgcG1KxerQ62zvQ1sFrx/Sa5w3mQbQ
epmMfGaVExpNxUUkB3CCem9OfoflEOrQ3shwlKeAKrfSTptKJvXDvZEbRGh7Ic53WxlDv2vSVfIg
rT3dCnskTdrxpQrDQynygA7sp93XEPwtBPJ/CJvZcYzUl8gZ42xThadF2IlZqHiN/ZDLN42zslwP
lkuMHGOTwV89o06cfK2VCzlUOfQUz7t4/fj/yASJ7yfpDT3KH1fWAW9wGqZDnrHiE1nxhKinD0O3
AMqe1/qcqsZxuyVk4y83BogdxvUPv2jn2/IcQruw6Eez+xw6XTRXWjAPyd23UYU0lxtHgbWhVrMX
Aq7dRJK78PTWiblfKpVPF2EE3IW+t2bX1AMn2FGP4m9FODIQ/6xtUBXHVQyV5sDtP+Xdzd7mFhyH
PkKIDbgfA7hFRCjiEoAnZ4P6DJ/urG2zHIdioEpI3Q7J497DOOrxsaITE6YSA2ik+1MsODtSMbQV
LQYo3EWCQvDVdYVMzHITmv/+A3+ILHqxlfWpSTzeVUdlmBeQiLXlOitNby7AvHTCJONUcEZcERzW
rEYp3IAR2OZd2vmYcyVjBI3BovnXArlWeI0koH9c6XeQT8d94/PujC+jM0TBwZwgPYXXgxCQjg6x
CuKFGwAnS4bPlCCUwCqfiRff3NcO5EQUln/rtPaJUa8FZGwxi0ZvfLZ7g3i+ckVjVDWB3l03YPc8
9PTsPg1WWs4Esl3SnXLIVVKfQccGt5ztPz3wQ+FfmqMA96PGiX8Ftrpjdnt8K0d9+ZxwvcGB0Whq
+e81ZDjEKK6TSOhBS+nkRG8gx6M/WbSH2qsbVcPzQ3bqjIxjRtw9g61zPFqtvMBm5pVdQ1zRVCKx
UO0EZh/8CwEOWZvtZjMGy1Ryi6QOA9xkp248JJbScEslkiogq4rB3A2svm+fypM/rsafOWYLMIAt
1XZqZQ6yn+AaLlxujMLLNMaBiwlO+WW7GvB8deL93i4Gm+dmf9W4ERbtHZ0MOPlsrnOJ8B/n4uR5
9rjyEQwY59kqehrEu5to/BVsL+2MTSBNHxn6Ik03DESQTcnYjE8l9/cIFqdeY8CdXtqoFOLXLV/E
sr3yMgo8UVYIBukAqLpBR9P6w9ceL+oRcB4781Qt2ODAoSRDdPWmFa+2Nc55AXEovTeHBVltHa6O
Sm2mNp2snJ1UcmYJ6hN3KsU+KVASLzeclFT3G0+l34k6Q9/i7OSqKQ9wTdu9D5E5mp2RdQp723pI
ehOsNce95WhGlF5p8hRnjh6Q2/h4AhQG8ggr6o6bCVceB3Wr9tGfWPWSwDvKBUxPeo2pSWNPeyQu
bKIg1ngicFcvsqfobUqFPiZGF+ry28q+3wOqJUGHssqjEEiJoiQg+gGI6NNFZgsWWx3VQ6Rl5v1R
jyYpmkgpH7bnnTTJjRJGYHN9Y2g+eE0uACgnsaHjPnVXbJq10Ni0LCFcHH9emGrCXaA/w+2YOzHu
uQSdRCfb/G617XvpNXVOdUotrQ+4YWdu9WnpAOhlWJudaUgw5tumKzlmWk5ipJm0meEzioyzMZQP
5iaGa0mddw+sWuuj7y42VT6zjWc2whC3g5WmuaIAnOhJ6la/4Oxn06mYl1cq98y9TtG6p4TVdx0q
AeRcZ2B0xxthvS2FAsR9C4Y+g4ptdeweps91e6pOsFxe6xZ4O49A10II/4f6s4tyxcvWDQpY3CG0
S2N7f7OI0tyo7yhi/e0ehQpbK5pwZ5neZihnz9Bkk1V68Ke6CMJgmn8Y61+VA3zBBIg00e4DGOiy
M/mRK1AVeVenMapIzxFlmjz365zd3S5WsUaCCuu6aaC+oQtyWNJoFIevQmNEtDE8FiedfBJz/ZbV
iSGPVnkkhJgE3i3K3XOmVKNrwmVPOqQ+ty054ukxrShe9EsTRPIvEALdx4W1GB2/EWJx19eCYCX8
3guYlZZGnNZCM8S4d7W4xJlN73Uxb7BFRSDyT4tlNFahKXCG1nO2RNdar44X311O1EonE1l+6GGN
gVXoxCVXdp63BSum17fabFav8BE/9ZLmAYDzq6/bjsIQLMGfdoM1Qs3rXm9vdm1rw/uV8CWu3D0b
GoNVyEyJ118EVbpIGqnEdMl5vGDtCAi8WTSya5NERQZruO94NvE2K9QtHZSO/X2b7zeuvIk34+Td
ipDI+AWFIkQnAZLXc3JW+kwlkrG/Xf66aoR0ekkfHEOl6QVoLPNY9118dCZUyQTlvfiX7JJLgDWl
Kr59JhPJ9cGWMN5hW0wglyFhm/xEfNFZQiy+zTDUkoHFEbj1r2kNeaq7Mh1WMAHSTJRSQOjedAT6
3lmc+am1l0+e73I/R5W/JHFAKr2fFR5Es7hsebcLubMedcnDR86YtfeT3DPPb9Qvgsujud+omX8f
xfivknaerJ2pM6lMM1IdoQGIyDSjPA8Cjb1nSIMYxfTDhCDSAt1br9+L5m0T2bCT5AS2tSsx7ck5
OAmjHHGmE57N018+nimGUzw6Ju+gDUp1PxGoDofOmo78eAOFZiKHvPUWG4jrNUtaAbapYg3ZriQk
DZtgR9sLGe/YGs2R73u1DYmNVP/8gqccxJ9TNYVrdAfbX2RkbKVoAgnvYUd8AgeSzWZ2TI9U/Lw0
tQiKn1QwUOR47J1bFljdidi3OD06nS+Uf5QE3FoCJMA4MAPaWhnsmyCIFDfZqB/cOGKPYEwWe1A8
9gRWw+yPvTWcB9lQdPs8BuhcCG0z6CTPG/NvduaQcsTYReYC8S26pwiGK+6caTiBOPKr5XpGMjzT
pikId9j5d22RDqWZJlNf3TZKX0pr7SjeAdE/ATOhoVm7l18Gi0cDkzZTDcyNQmL+2UJIciJGLboI
XQ/3fyhW40SDXm1NkGjhYCP+ktSr8SLjG35/CBXuEPyQpCDD3dHP2l4HA8ikzw/ZG15ajPISm1Tn
vtuMXIPy/2RNK8PDXVH9DdCwdlrc5Hz2tK0ZnlZ1dZyRSGmzFAcviww/1xDXgJKvJ/5owu5OCawL
bSjwkktgkmyZUpvGfXDd0BAWq2MLt/KbgwbN3O5a0thUgzXtj3Pk7m8VliLSg1eK7u2eg1H/7say
BrF+E5ANLempreeDuI6128paMWWlpTzsSTMx+SiCaVXs0Mf5dWYDCxKh9yHQdIC+41UcuSvOdNNA
0NkUYo6Z6aFGcpF3V+8myorY9WIH9Qq7bLiXv/ZNsIU1U+CMWJkt7CtFgquA2JqSfb5cq61M1XZs
RFFkfItMVkB2ublEUmxGAd4+GekO/y/hfTOdpHCUQuLENlOn4SfNacBgsaj9ZRPEzYrCUVsCWrRL
8lYFkKxiGRnKCgkDa/AeXdoC1yK/GKYIukrjLnDAAbLvNFKBZMVz3PXo+Ny25JGEeNZRDK0JF7AK
XZFjMsA9WcGtKgwKVqCCbImfuhQuvH2XNbfKkuT7qvVmAClbKSst5b5ua8x6H4N7iGn56pVt8Vvf
pHAKy1M1TkRKpsJD7Sx1tsStvQ2ICkz1IapCpI4WvqAWmLFbv9Qx7jkE3VxM5oG3S38u2Kc5SWDx
IgI1gsmxNlhmjT1t1hCnUdE6H1gNUr6sPBNtEGM5dE8Kv1lpxfaonUYGQLcIVjF42jrpbx6D6DzI
ACcCUZbol8VaxX7u+BEVIL4RXifw+Ej8kKrTe1FVD9VRwJ1M3GkJvKqEbL9Jl/7RG9yAr5HCa423
fnShnFOOyyq/QkTQHzHfpMauFo3/hCiCSbntEvd557TT43xE2GSnOjGwAK76U4kjJkn2TQ2cm1z/
2qsGz8mAXFhcFieK9bgRST8Pq6uWPljz0eQXiOWlD8cblzGGS4eKPFuY4bgV8vIJxj1gVBfl/TqD
X4JZSycWzayMXldFbC/niGpeG8ZUK1hzxei69L0ps/ruVxmEsPeg1tV2vsJW1lViPt4sGhfcVTGN
GfPD05Qyy/aK9o9jHJ4faFGGaYZ+UJtdGobOrI6FJRcOt/AcSeZvdEwVPcPduT7SLVoRPM6dxBJ5
IjeLacUohVV72ZwWgV/VdDWCI7s0DnZdwxOKGdxKIFcBN310fNwmws7IJ761+02iZ1mvBzRt3jaH
zEoP1MQz1z4Hz2Eo//HkWu34cLuo8IGVtDPEVyLV/NodaR3i+K4wOzlgkudy3RIWZzT69uSG/iZD
fi0xZqmxN0xoQ1ZSndX6qmj2RGmcIPBn6TgHlDtQ+Xp5p2mZc2WBGWCfNv4vIm9l6DgPjO3K+Cgc
D1l2Wk1hcLTAJtK3mFo+uqd8Zy2/JzIwhS549233varIBYE6grjn3JsK82DATaDhLU+ehQedRG7l
VKC/6MQvOevW4bI6IUK7FZiS2YPHh+5MVdic6RiBvQ7uEj0T+qIzgs/uZyeMvwJOyBZMgy2pePmR
d26jRZNkrwdccHZDCFaCl2CpfgkBP72iJrJDa9Xi9mPbMJTgNO/GAbb/J2/+juiKm+Ku0N+gyTra
y2I19sEo2dtdNRJhYPaW/pPm6XAyUN0uw6mKtntKj9u++oV5fEsqCrZITE7k+AkSSozWW5Uf7oV2
kZVDnhHXEo+yQiPLwpfFVeLZk3QltevKf45LfW5f8DLxyX1+kKe0YXlqAbLUKxjaJSVt51EZfvLL
d8rqlTutIOGyluB8rKVxRw37W645vYweEH8AGKxKR76qUk171gooJWJBtX3W5XDSEiDvJowEoT/D
6DbCO15sgkoK8TLQCKRXDyrH0NEJj6uxel11Ltcrv8+wxn4VSQM48rUXKAqaokPnZR/GwzqSgmsU
ExqU79zdnoMvmNUtK1ZTOpmy+/ieywgt97II7s7jJytYqv+HhyYwtWZuJcP/Nye72iUaWRWz0cre
2NTO4v0tjKdiMbPcRoq8jM7QyUmLUi8MAQZiWueApUyXPLHGfTKy01lYmGwFRfUphLuvjkvCRasp
/Gh57WngWxYXqVbQxSXYTpbzbtTk+l+jmscctjYazbqqtQf3tyZ/WDnj5SPnHcLl/CCn/kSzjFO2
tigXHBCiiElHMOR6EwiUP9IeOx9eTnLOz/4etXNjyVA+7wLSWjx0F851X8IsljYKiVrzv450FsJS
6jl3IIWcOP2S656FPCqMAyyev/IyOPJ4K76jmpgJHHj8EwlJnsv0IrxypakK4VIJQKGPdhmK50b3
4cHphnQ5fprhUssN0lx6lO1M1Vb1q2rnxSSXbxzYQtiCmrHeDYiww47S0j2sYRplhN//BgXvL7x0
mjDpbsq5FygBkwIArfQK9TOSpNQKQbA4sdBi0R6riJGfpzkLJw/q2rNkpsgnxjbZ2dFZNF9htZQW
RkXP0SJ9Sjn/cOEEDPfpKXZPCQodFrb9NyHEgDD9eL382v9teC97eMMmwLflQcDP9QTeUcrw36by
LCwPG5Tuc1kXMg4d6wHq/hugJPqazTUbo6Fdu7lJQ/00hFOFn+QWrkQ1p3/ChQuZMGYxS9FNukLe
eY5bkkc1ZhSU/wbQr67HrMhODYInWxB7JL2NgsYhx4G35acvI1s54CWlcdLJzUnQYs6FlOTx4L8x
zZ+xsLtCUMyDTLhCJ8vkPym+/sbUeIF93kvyPFiKmrWYjnzTXrxgpi2/adF6srtf7B3upbfYnKON
L9ispGnmFJTKEVH7OmLWXMrRBpcpUwkT9KUHQPdUVXtwA6V4Jp908qIJEG/h8XdMVt0gjAdIVB9a
cnXJVrYYh/j99dOmDC0eqHj9755i88nUbQzpf4xwkUgNLL8JC5e7YOFVsBXf6mwEJ4dWfx47lO3E
CTphCqH/xjRwuydXqWrBGQi3uvkz/rE3J04nqQj0bd5MLniaibOIN08+ksQgqCEftZNUrv0cUIgU
8kQoV+eqLnB5+dq9jD2UefVUmJZJSI9bv1jXQm4ZEHR65DgpcaGGSQDP35xoH3nQcGYRuE6CoLlf
opEXBlBG3M2WUGUfHoD01sVAZaWrwij5KL5pdlJrSNaRoyPRY+Fa5BDL3n25XHaV8hRwkizRZ6xD
NG13PJHTx4D9zCz0SglUUssZ6EcaBkPyd5Pja3YEMJV7lvAub4ooMMcT9FODST8VmKgW2SSpho44
oMskzVj9S6EPp4n+tTbgHY7rSb+IujaVMLzmn4KX5L2xGK8h2kBai8f6yDog/1WEmhz47E9oUd8C
rlqIpQroGgfMcFH86NXclPb2Wv7NFmADJ4yfRtUEfXifWqndYSy6vLJGI6CnepStPH7ylIqyHG0M
/GFd9sD6M4I1ZqWP4tKGM6SFbNaGmEngXsiSNCeqRVotcfhjp+8VaV4vPSwzL6RL26RR7+oBIT3T
gCpF0w5TFh3XVZsvhCeNzveI1beif3UgU6B1VJTcIC6tJT1LeeK/vXpu5FIpUOngxuBRwJVjP6TV
U+CWKA7E4QZUvTGeNvjsU+fQJapQwBnqdbJUEfyvi2VOSKGOkzPpkgKYRFszBAiXI29QHVsabku0
u9F5TYgIxDwwraXxX/8dwsdLGJE4YxifnBiEmxKTgrFX7pbL0gr3zZDkb+k+BWEJubeWU3ify3en
Tnb47IVO229mA5ZT+5GkP596HDAb2YS57skiLpq9eEYvflLN97bvtW7JNZpxGir+hi5RUfTvGYL1
K+/b3OiJzTKXJgGKXPAdL8aJPlbs8Utjk4ES74z2robBLJn4AgkarAehgOkDY7h+1Rh1RUB9VXW1
09ORz0GRb16jLNQ6a/Dgt1DJUC1m32853xH2Lt6PyMjR1zOAjDpOCcRwGEBIpscK4eSuSyHPp4GI
IEQg16tacoyHjoGeehuBJOD4Mm7pi6fXcvR7RGF1vzyoPxGi0FRNv/0RAmNd9MHAOPf1QLnv5A5b
qtNLABs5HjIJhTbEibx9UmWqqNfeP7BTIcYdPmxceU8X6jQoEw9GunHzLnWfavEHm8I4+n1ezNIS
EucYNYhzl3b5Brho0hfWkyJkmCvWjAaN8TgnRfC/dt3qZjPYfzBDkyuAJ3A6dRdf/Lf9BrO8QPm6
CkdUkJs9p9cO5jfHUqp8sTb6hO3Qe6wwowWtG9OxcCWh/VIFDV5/ehxnuid+osRzgIl9ltkhGhov
mweRIRJdUOnqvsxOYH9I7SDj7FkIaUl/bVVzUcn3CBzRF767k3Lk0WpGA81lIYWS6hUUOUOcdTjx
TrEgIOAMAmksJ9uZVAdoEGBf1Lx+uLzq/b1hF9Z+vb6x9Mbfklw5TCq2fD9b3543zDp+/U6TMZv5
ADbAg5PKQKMO5AuSC+p6eFJW35QvBftV/bB0z4kQtp/u8pI5HMCDdlhB0BB5AyKNfwPiD8eNa/ez
Rk0lQ2odJGvRNovfWAIdBkd0JNItDszo2yGsWfBBFPZMkoXk1YYVMqb9VGEv+QVP0N0awL0+Y/GK
yIUrX9/godzfyfolsvNYHvCG4KnU2Og+XYLlQm7AcZtZvp4bPwSpju6zA8+5350VEDhS0jzLDfBv
md23tERi1IJ144uU0+JpaRdJDUCPUlDVICZIbo59xw5EI9Sp/2pMDiI+YhfmPHmnTIcfHUFm+6/L
S3Y+4k727qBWsSl5xzcJhMHxxYoeMuLlm6fYXkbygTeYpeo3aafKRRlC5vUAaU+8LJqobZbOUxjW
6DbYaV0RKRRb8tsgh5aoQPx8IGPqvzJFJJ7XeRhXqh/xVItMDtTyKX1SSmMYQaqncp8XhEZyj9nh
ZUCng5e9CYJ7BU4E+PinTjPo11a2Wd1nJyvFV3V9gau/BcEm43p3nPxfgeQDlkTNlzrLNIyFkNQ6
yuqw+vEeNYwItbaaRJU9Mqp4+8BTcgkcVc1CpRItO5sLpwzfe1PGevHuvGKnHZ406LEUSZq4yVtz
ohsP9hCH+uDIaeHsSgfi1cZW4b9ykDpGZpf7VPVhDzYNbmR4+znIqdAEATRM+dMvPNJ/UvbLEU62
KXo2a6MPqemZ0mpH+2RaIhOlCFVJaxZ2uO1rY8VUS0/M+LL4UK4YaeNZ/OI8K1QoEjmsh7Z0J1sK
6rMAMG2FCJAMX+naYQGp9qGkxkvBIZcmCTJ4Tou76XTB9gAnaprYR5liGrWEzwWSF0yMP0RpuMlf
MoShdp/GPeBK4nPkBT3OucFJc+elV3Wgu5/Ma74KNmQYK5uev16x4m4shY50od3FFTbojCIHlvGc
jws4EORvqwm7vPIPCa/9lFTdAy2FxTNddVBDcMDvrenWLZvbnYEypUbLksdT/fCAORka2zERt5n/
N9MR0720Km0cpKuit3E2+NlB7316z76+TpXYRYX3cR/5sbP3PoyQT8y8Po58Qzj8FMhOhg+kO09p
XHfRLaevnhO8tdEfCuTgKfFGIsqN3f5EEKiiJoT1ac5EO2mZq+9Fek9wSKFH110B2gJoH4e3Jm7K
Z9E7EEjBe68Ff/DxobCTBb/TvGsohQmelBK8La0Q4HAGgy34HfMyKKZuBj9+BIM2a5koRiT50ALo
Qtv4wRx3875GpNRIgViyvfy8z5wlRS25kEald0GRbX5Ic3XQvovY7QQ01BdYRXBAkMbp0kUS1yUS
Vb3qKJHuBIEu+M4+z/Fhd9+SuHpx0W0Hb5fpKxrb3w2N0EGQmL/J6LCn9uMAq+3U33BzkMHWHLZG
MsEfAAq0K/oWYuJdSQlDTDns+HvQ4R0AIzdIE6Oucz1EoDRdJrRUK2pX1l+PCaLvhYgmbQtliIWx
+MoBYvVLBvCwoW6mlA6g0tVuVk2eslnL5XpYAobWzZeDEX5cW0w484FWIFBSYLX+ifqswJQ7ZU4C
YmtocmfmIzXF/afwD0JTCJ8TFPnXM24lu53r2rZV8YrjjD75zOIzWo74oBFavuDVG2zf8mfGB5ig
LEvycqAGuVc27ZZGoxQ4ukNjUTUCDpjMAuwyXscd+xpzZAbXVVUgyxq1/GOn3uQ7TOxcCNEu7a3a
ilQrkTFKznr/qb4/wujFvy1GTCe8g+DYtafHYQYYqnlJ7u7hn0luZDqPP30pp7KUZTK/6XxAvv85
l5qmvOGCEuLGccLo+y2FC0ON4Oj9gJS1VchFqSjX+QDiYOBa3sQLmFKsYJ8VHW6ZVeuuUTahBdWH
8leYwFYI1N08CRUwtT6USfQZdDa45MzmDoow556mvvtRUoNo6l2xZgMKXWrfnlD/iXj9zOFVbzh2
mIQVe+3A+8HR31Bvrt/MRoJtRIHi0CHlsPw0kxin+GvqOXBHx7ha4749Kb7b1u1ckuIhwbHkpIRe
ry4fl2hIBl2bi6xbTXWYQggvwn5R24C/lwAq5pGqY0qHwzzmRxj+ytgdyq+9rAfZyyfrwDWKhWDk
1GeOl3vPX+UqsaSPoroVF+TflYk7BhKhnDKti8RNeCzu3l+kyv55DTWio0HaebV/FWTCc4SkfUyB
M5d8DTyQzcfALJKwWr29p65NzKspBjEbBxpI1mqklER13g6zwGqAXJCUfVKuGF7tTzc9S0NOvq7R
JQkkK84sSWybsn93nCRQDSlzr/880G2F/Lcqiz0gBf8hVuxkgE1WzKi02I8+j6r3x7hG3nvCxAv0
sg0PZVzPfG0cS2o/4tEf/aPbMjDnfJN/MBw0kcMX6SFcSvO78AfEphe01B2HXSWtasyU5YrolFKN
PDCsH1hED1BtgW62nMeyaRQxMCYmkbDdF4OAFVUJd38ZWBZy5XrC00VTQdqkgd//BnZkW2eITMxe
s6OyQOofZLwO7y57wNL2Joc87yZvtG8vc2emCdE5Zq4z+WO4sLR+XseUlWaekDW1EVIJnBEizonV
R0SL6yVBUQG8z4wYLdWAfo3gYGXA6TglLpgyBKKFMV0YEJQiuIq7jSvaB4keIHcG0DqBUWfK4/gQ
olXPs2Amccp8QZR3KI35afGcprGVHBVIfP7T1ooaBajHQ84Ls7M8IyuuUaRmOKqP86FQNFIvVEq9
li4sg2LQfEgLktMH+x4IYOe4CCE/u4x4sGj6Ssks40Xq0RX1KMpE6NqQAICj5wvqhxqAiv8C/oFm
9j0h8luwYeDtNhG93dwXYKGxLNp8UBlrJQdNX3AjCsyV6jgZK2hyctoM6PfV6NAop3ZokDcohb8Z
fAl8QDF96niuy68WqQeRQPsYtbtqddvka76QNirtgz+eoEVKgZNLJf53MrOMPB4rHr14B7hNU6em
kvn9BubSxhYHYU68APmr0ARayiISITnbxyrCzVOQ0X4GGcANBe3H+hWX58YcOdnvgaYzn6hCt6cv
WvdhdUo+oUTh9AYu1o3k39b7h+sqeJqRgME/R5pp6ysCsrFTFhcDkIxLgaQtnAJrBgmlEgd8ChID
RWShuq2ON1ddhYBYrwCDwG0P++FDvovU/IYNhwSKPFfoD7J46NEisvcTl81zoBocI13lhEXAQuxE
XPiltRNMXJ0kR3i4o34WZw7BTLl7eqFuy5BxrUh8dt2O1kOiorue66JsYDPwyXqGPH4I/GX/ibKF
63TiRwzb0SuLvNsn1bNzfeUqd1iGD9ii59/6+WDL5Q+EjDaTca9t8LyFpywJjIiDkpRVMTt6ErQH
zlp+c0BxabmdTL5yP2xkzc1pyhlt+oHDMarvyYz25UbOSRRO2I2ADCL7L6VDvj4P3HTUd+5SE2sO
rd98zOoF4cpLJ6pJEQ+tn1fIH9GuEoyCFSCod1uYVNftGJugMUdwkOUgEJH7AnkFzjwxR7B/H4IK
XD09UbB+7VztLOVDIUwMJLSMgZNCgGC68dv544QxepOuBrHsXpLwpTRMIl7SflJRJ/zXXHjhAHFc
7bAJOwR2paO+fnG5FO7l4Q5T6Zk0EHur9oCm9o5lsDO3EWWRJsmCdCI5k4bhNPcvWDcA6VLnaGO9
ILLaWtvkpRg7/JbnrCO53ojZN8mH7dH8DUUSnD/sQ03j9aLSk5UrUZBG4ykH0l8f8HQuMnSVbWuj
SfkM+QTurBlpVGCWJUueqQl8GXHVk2hEAAVLv5NLw2pPcOkj7TWSzBpI/qXZw5ENwn+TXxhhaBK7
tedHmIAvN6jS37zPQ9f98ssPFPahIAvlVj20jh9Vk40pJ6UwWTwoyKaRFU/534OLYuGpnXnB9QcI
xrUowsJKVcCwywhOMturzOg8Euo+GLcFv+NhgLZdf509UECA/wXbSxauGUlIxSTJOV86DzFZxgJJ
3A3VKmyz/SrCk2NJNKF0XpBvqL5HEC918GybUPVYkzYJvlFIPmTFRt+E9neCRZ1j6gFxTp4TBL6c
Nxry/4OeEY35xEcvwy3cOXTqKd5/BCcQndixL/oRiiqeml78VDPVG7Fr5jNSd5hdKm/Xqqr7XNPy
ZWnNmO58VzWRXeE152hU+UAMNo2WdHl6zhHT/9iSWTz+uEuLOnyBrEizcHul1G0PYR1+5A1vOVkM
245cDKgHOQjhT75OJ2vUuZJ5/DnYF7wlpGIC6+i6rH4XED459zD2YD4zzn+slXyCgT5pKBFwVRJL
f+QnLjNTSGqXbGXTwgeP9V6K+Ei77qrUWOJzBC155ffX3ewLgkmTcGtAaRzw4A3Bo5XIciasxrad
KfnuWyjUHACfsrVl7N5teIPgFeEcpxsPaHPcJXONU00tG21kLIP96j6nhwKf0ncLnoo9YEHezGS8
AaLUbPNaxOUsckP/0sVdlLr5yjqr9liSAYv6QMzM0ldBgSBaDM/Sn0itHtz3e4qIWWXh0AAxnAUf
Luhy0oHBWZBVWEqvOpDotZI/17hAmT6t/leFEsttA6CQy19gSZS9BOHejkO+aGTMifppmvY+dykk
ePpbhPfn/lBavYhIAotUs+F6P++jtbPR8B7/diN3R+PCV6PPSgC1GbLioWpmpGTrXE0nS6mFPLSt
PpRtrinPLffEhk5hQcLT86pRlKk4UDerpy0dlra1LaXy0/Z/YJzTkbAyZTCRmBQe2IcaID2li4rG
YtpUEoqExm+8s9KuU153K86YhQGH8vEag+TXVDoqyt4wnxDU4uhpp+sP+cWcnxnPKIIDleGZmvAT
WLQiWXGAfqig6LIee0l8etWdfInd95xw8KcoCmHZBU9+QycxYwCj1f21ECwEbxz9f6p3eJrfrvPq
ffsnVe112ABAq813k6bp3CBa594U6ZpoOKJp4AgYl03DqD7cHHCPyOMA4r1zP2o0fUX9LjEIzb18
LNplBey1Zz3pyMRIVolRky/UOj5RB52KoSJ8P5ZwuvumXsGTc1/8+qqILRuOOq6dq8ZrkAMryqWs
9/xXN73Hd62WYajcaiWBFCC7s5rrdYnVem05EsLEYnaD9XTdJvM8QWTlOCBqBTeh8PoVzaQaJSfm
Ufn4RDb/F6JpPjJSIk7ErQ5ffl+U0y1GPGdSJ/cpPY0WD8jYyR9QABvKEKmitHNR0R6n3koO+8TO
kZsGeSfVQHhFB512UTPi4wvG1J0UbisvJBuHyzpMz7vjDjMTQLF/yzWWh2wVEVlaMkaBr5d9AObj
NUaAEwBXBJVQ2HXxF3TwqEc1SxSNeL3B3eUF+XZWV+VLoc8Eie5lUmAGM7drusmqtfoSyTY1Mpcx
GvFcmQglf5mU+WF0k/glr4WGgPvxm3CtNKKZYJo4UX3ObwwzGq20gygmWiuZk3UMrBri9cvFxHWw
ShGhD/piEmtH8QbmI0/NPXq6xPuclBM4rDVXJ42TJPzo3jqvV7tzKBMNfCckXGpvayJcHuRqtTyO
/Zd3CquvHRam2V8776agZmbQT9ALHxYrZVje0e/eRAX9xUWmivmkFrISjfui1Bhvs+Tsthbv8LL9
wFf+sUHVbasivxgP4w8VQW8r2pyE8S4EEnQMk3awUBFf1TrtzOoG4dCdlT/5G/XFxJ6NHMA05EGf
nB6w13Yx5oRAmeGyw7p0QDBgSomyLYjYrfwhDhDrqnnpxeoLBxdmcVpGElnRi/4a0E6hxVLBVsXL
xWvMbDkBv4yY6IFaFgjz7TsN7SI68GWp4PAjLLjs5bwWLjp1NcQDanecEj17iJdwf+m1ot0mVOdb
Po6aU1DzA5HYBACqN+h0p+T/haZDIKvtmrPfz1spr3mqjXFMdaCxCgdPgi8Fabq+h9Fp6ZDiKx3p
mHUMpFVkgD0IWxeRyFaSawldfoehhcWL67abEnz3WEOGXOVwV/uJMBSpfmRR3+rYQy+xG7Tn+2TT
boWlUIZnzX6DRb0nbd9EuhRnWvx2wSZ9RTVp8Sl99UGWS1YkPCcl00vroByp0NPcCQNDuxUWqUQP
tbvBh+tgmC/hLYRKfhWmlR4GXXCM69eD4VgkgmyV4QQsrOR9Y01i9aYUK5BsvAoQN+NWt0Yecloi
UzNfxUXhsT4dXuhzVMH8BpBUzfTzgByE86gI74RwKnrDELEqy9pCllIg00NZWSpj9iRlsNmWhdRR
6etBIfYkbAsXMCV7bFYmEt3qDufoMQwGb/bqS06/1hhOywIIkCbyblmjwfxMo/AnDJE++cXdECDJ
7te3p1K5uXarf28Oewz0XDzZvi9v5PTWUFqrOmbyljyidCmGryuFgMBSxhrrOeKLdfoOsjtWN/iI
sOdFbYMrV/ill9XG8VLSxM9sUmWoHte0SraRsJDCEfvbl8pXx34by2fzH63DGNQNrTdDVt2TrSdb
p1vBrepO/UMpw1BMcTsvmc6MpjztUA4/IrCjMK6VU87WAoGRVsbVojiZm1Yng2e6YERM/2ytU9Ya
9jcg3KpC4ZcwZq2wUYI9wZ8W4IfddY/O/GcTS85pS1t0YVktW/kvhaGZTQ1HIlN68m3sD66adO/y
Rc2yGqYqZ6Olg5Q/AeSFO0+0nyOnT5g6t11M3j5zh5ewX/2EZJpU2riIWnnI0njEOZwuRFow88FE
5QBHUEIyBoH/50iekyhsfSVAUIRTgnD6Ui+JHBgNVm7aQ54+4ieyqB+fxcAxPuVGEScW4s99XOgz
e798z2UhXYaJa75aofLq4g0nWvsbtGUi0c+xUbWYKtreshf68sH7n2AgxDo5ZLEq0Y6y3HhO2MMm
eGhwZvXVPMqko1mOU3LQbP4g/g2oJfgU5rjWppK+vyQ9WSxIrer6XzYbFdmxpenySKuLKP1sM1bu
xRxLpw1VW/H/HQC24UAFTP4e8phgH9YZ2cRBdtGqlJqSQF6+fPdEEp938S3+cWORmonwbaKCGsv9
mZMoTHh4Tfe+lgKaLDx+krHILct8w3Bhifl4YLTqXF6inqC6mzVuKf+LPyVnjVHJXWz5nSrIKQCB
6wkQjdbwT8qLB0VsgyMGP1DtvCQLvwyJUzH/hQFLFgxpKjAlu3Ec9Ao+E2Rtf48qeNx6KBnT6k/U
zddvT6BjzKN3+M7ujGUmKjHmZv+8cfdUjE5eN/ng8myzl64N/pQQWrqvm0A+rQmNhdbwEGJlqkpZ
oBTCGS4y0Gr3itsIg2kiEFeCRk1eMsNZA0BKHNU/cFBL7GU7U7oZoi+w5Eig/Uqe49woSJzGwjrL
zU9qINqGAGGmhy2SkSLng6P6fyCp/+mZEF9BmUJf0iNROpplxaYRK/feo7tcsUYg3KE0i/xpOLLk
I4loai4cVr6NVC2GB4jdRNPDsOGWPZwcfax1KIW2iaiaYr1Ey9ajXJJCJNr5VioLAzOzCJyjqIWM
RWUQBAh4uJeu4gFPhGCeochBBUft2jKSnT+pgn5hBRi7mm/DrN/UA0NNgRXoHR2eiIfIdTK5m2Ts
/QSrMy0fD438g+7xDwoGqW1F4Qwbt0YwliZ2TXfKvlDumH1A9RDuQCMCnbZ7V+i5/AQ1OUj8fOZH
/Uq+WX5gQgsw6MwT5qYBW5FVwUNdnrvcgB9MZncU+y1xM0gpmvI5gFQopaW72XpOjbSLj0Z5kyfJ
pfNG5nZIWfT9lo2h5G0NrquKFm6Rv9c2NPI2RZeUN46UbjmWTAytrjgcmCcD36SA9/i5HwNmUkIO
Lg6WNEd+yFRH08jtFX/hEYi+qzqSSWnhNvSVw5tDktg/pUUd10hwp30Usli6iJnFALw4B0OKOV0H
e5cohyKOzFO+d6e65vg8GFf2SqMDXfoaWrjGPtrUV4SJSF/qjNGfMLemvb/YsGkm1lc4xreKXKhT
S5aNOExOslGJdZWU2yUm+CmImokfhmZlFliQMGWpTqL5yZIk/UOxgEPWFa8+EHI5xPIdUttEKcrF
hOtod08lQ6lSAlRXgDJLasDHUwnWyFI9nuS9oYGUkn4yfcCpUh3rD/Bk2zR49+U2Jv7T5WUXbHlH
ZIsicpHEZzC8Z3nxj62ADw0G3Tp6puZzDlKMnwtPSafsQGnTbfI2HWfbNOCrHAWE4ugWtJwwMFkF
Tu1rw6U9/nBpDOYJNhqq7zq5ryUYmlvq/sBozBKQUOEpuoYQFgWf2fgcqtoPYPWo+FPb2Np+z2V0
XOmRHS7/Z2fSw14s15Vm4TXxtBFNejMS1FzwSp3wx150+0p5IOJ5shxv867rr3iJx1ExWcqLTPLy
TJxr+OBaRC6MgD38aGuZvddrHIOeR7oazNIZ+w0LVFQCXhBYpwlFxG2pOzsPVYuHwTUM7EiBkQ2f
IsRDT8Vzhe7RnRcXlG4u4lPCo6mIoVz5SFO9/LslUw7KrIjJHzuiO0Yepq3ajij/vuiO/44aiZ7S
bjXKsF9aF0nyYdiw4z4CGWFtuudMZF57yNHNfP5ZGn+U0g7yNunWP3FDD9ohWG7GcvYPU7JAbfTZ
ilE9s6sEgtAgtZpu8ABooRv2lHeUjJHphbSE5ybZhCj93PBil6YcSe/ab2apmTUkcPha47uA4iE7
JyedYt1cULF6Y5ISwn8wM9VrtyCT3SdwexFbiPg+deV912L2bodnrZ+Q++iA4o3l2vfQmu4Rvptx
hFwXjRfiIwYzMs4HJhMPGhqYAnWD5S4HaFExC7DIFey3ge1ZXqhOlxUlYE638FDNmfu5aaXj49lv
CebIQo1HEq4JFL/yqC9liq1IoI3RJ/nId0quRy2UlzRaIPRyMo/UcPo8KfKc+tzgH+Eauc9h0mLv
RIALUIB62i5cLGMtOmlJweKqp0sapI3n0fEuaHi0LGbaNGGo2HqFzdms9BQGAlwvji0NqaRlGtbt
xSVvUhAK+8+zbSg86ss6tThPSG4jURj++9y065wwxBJBdmezP8nrCbj1Z8y4w7pn5C23GlCZC5Ng
1L2evUPDMD0YYUFb9x0yYIeso+QNhz4GweWmu8ZB9pPYfuvl7U5Vn2EsP+t9MQJsAI/SN7xWuUd8
DwT5NE6rPRJzpO3KOZW3qXCkZbsE4l9ZIQWTibG/6SHDrBZNaJuFUCgDvXvKVaWQMIDQWr9P8l1k
Aa6t9XTohG/hkV5ZCXn6fB5vW8uDIEuKQo2v4sEkhJeRsqe9sbBkCPXyk7eQ8R/uChHGS7fCR5vB
LWa6z9+W6qxP6Z5qd+vwhvjXlwjY6zZ1cU4QH02m29dVEAzEnwH2K+8xYqKY/VB4jvbn6jbe5qYT
xN92NQ+iPl/xCKcODmzTu4Xaw+BghvpZHrJLWQabC9AP8roHpgASVsTJKxcEO+OIGWdNpwC+yNgY
T7H6DpWLCXyo7HyQR9x3uGVs+l8WgmwqNHS3RzuRR/Lgu/5/P4f7c995zWA59uUaM4BdbWFPxIb6
EsJGeVlUE8bB7uTD4bO7MfxbtmYPojsFOwL7RGMsW3CMgx8rE+xCD7b5ufQNEENcPJVswkKV1dXB
i60BpJKyq/wN9g7sMGEGdbU7UsnL602huBblFjw61TpoZ5dKQUbL+Ft6/1sE7JaiVlzXajhjrQLB
eJHXbgCp8b/Wqqy7FB0zXiBv0EppFWctGZGHvbqtmfSpGyBEImS4tfXbtSeauUhsHtdMLI8moDdr
dbYXXPofBKOThZu9HJeE9XSjKlo8ZM1wraKd41GlzdOjYfxAbAufO9j2ItFtEvh46EWP+7hlGaFI
wKCra9cbTYeAdKeaXcyTcrulHVMHoMfKbbucoq2cnNq8/vx24+JqN+zQQH4FbLN62ROFq5t/Sgs4
oTxPjFSWb8gtqWA21xLsSo28tJsM/KfYn/dF7UhSnZxrAjfwAbsk1Y/V4ShBCaHMPA776IhvuSSy
ucjgrrJDdhkFM2T5Y1LyjH0ARrv9IXILHffBv/2i9I0aG/bzCPkxb+4Fj/41xEOUyD13IYscC13a
jw3HKKWiZRnxJ+9MtqVf45VxIdDQ6fIbom1v58iZEvWsK41Tnz3aZqgHCoqmBm0e1wxGqwSzfwfE
XnvgG4UdIUB/o/gL4aF4hZmtadZrAthbMprJVTlWevA/BNVAEj28mEOjdF+SB68/Pw+Xy3rXH9D7
PaGz90nafSPgQhrLuP9mKCwixouB6azlrWBNhwV3mY0twtKepIJtH/BrLoy8lTG8D1ZbV/Hu+FFn
VYI5U5eTEg6kpllfmvFgbiojy8+KGASicS3yVbmH8v+ZmPZvmtdYeIPurr6b7iSNZUpNa2GRMMUR
vV8wpdPSaLnyTrIIomtMW0sTEzeGqGcSRrblVNkXSDfCVrLlJLlKL0BcORrPdiUA5dXp+xzeQ641
PLGaiEv/D0WsQNReznSGK17u/L6wHsN7eNq8+4AtB7TkqkdK8nzUNABCHhgWbfVjmTSURO7Rl6Cf
L1HFOJi3eLsBiNZUzbUrBl8Y9ovdxPqxHW9l7LXr1egffvOk5RO8e52oXZW2NVyMbauLvw1QNlXa
h/VUw88yknHYIUUd1lkKXmA4cyvVB/YjUfRS1R9pSUmQt6zYWK/mFKdgdjrsB8ThW8VgtemcDXpY
Et18RT0UJXdRqefT2xRzWuI+9893u6F/ELcdEQV3j1BvFn/EYgx3e8r0y8OvB4533ywd8ZzWpLJ5
rQ+KjB+3OkAoYQfFQYjDJm7d24GcRtZM+EMwqzeRjYx9NFGdYYOGNk+F8ttJUIfkDqC5n0XtR9+z
GWSV1fJsE6XmTNq9IkFyoysbRK1o1I4Fobn6U2WgBkJm1ymv48TG/mEDVekPRuVDykhwYmiXDvpv
C+57ssPKkqQX81KuctB0p529/MGH1myVEJ35c3stjRHKLn7FmvpVNshbWmuhhh4NonLmiJlzeM3U
ngDfdcP2wesF1939gIB8Qn1MF+N4xHJLs+sKBQJoRjur4h8U3b7AsYodyFPnH6tRxWfKHPtESXZn
wlxjgbQX8okgP5IZDfCIi1jwUDflQ86r3C6WWxXyh6Ai1uKnai2OfyUm0/gDK2Ui9joKgsVnK4UI
6nDNtj2NDTYkNsQ3WtcLf3V+rz40NkR1R+nvGKfhRgycKVu4QLAEeMmwAZMV2zanwVovYjRLMcD2
BQh6OkAYfqVhLmgbefxxvAvShYswt2h1sg6Iof7yYtaJ8+HnEtRvAegz1++3T6Xr6foBfONAf69Z
uEQ9v6zITPez3rNOkl9lxODTw99g6QSkpbktlzhhYEjYEZEJRiJgOgkFR7M6vuBQjM7qY4DUXeWB
/ELqLfjAHV2J09y9ai9oy3XHMtxpT3A6MnzfNWJ4p+w3A16q3mNamBVdmAowdOLVMnwhnNfId4Kc
qlTnLdOG3Sgq7Y4W+0dum24LtXtxEo+t2/rhWc5PbWPWfylNzhMhmo6icCGVnnMHhqKvoxiDYrwJ
lxf1aH4E8P9sAG4t8BamyNnHuVOMq4/AsSy+YGir5AQ0U7+RaQZZaJsImhUyVku2esNkI2MyRLyp
9rjkl3ddW0CjBQVC1WnBiIxhQ86mrlXskkIRxojF5lLB5lrH3mfLvWqB6AOdbWNpwIbiPvWApPcF
6PE+//9QnxfmzVvcs8tvj/PmRoSXXsxbVoJ6SBL+Qi7Tm8599rP/ssoJr1duNc7T7FtV2qPdlTtY
oHOQyk4Sd3NUqutMitG4l0M91uNHaFoSasrsS5pnlBlYv/b3xPYbAyhXSUhfahNxzXYcIo1g5lBw
U87To1TqovxYyF4SoMhrZjlegWt/nvNSQhlddNbw942KLXX2EwQAz26tCzZpr6Nlkx7buO/c8ylz
IxGbSjKJFla3jkJeoqtxPs+YlBaQkUxPSK4pfhn3Hpx0x0TeeCLP6VLW/4oSkeUS3y7C6AkZaFIn
OabZVZxOe4nPHMlk7N/Mmgm/FL4Trh56gmuUVRIysN5DI1r8A228B3edruBduT3f/gBAbLaCczCM
SxURxtR3juDSU3eSqPKdVltmdEjamdR2zLA8Yx1PC/0kP8BJyiYF05QdxGDwdzQMgq1Nh4RYtQmR
vHPyIn+2ZHzYGu7soQrD/rfjxJhNhXCfb5n6b0lsHANyaGlFiUCqw2Y0GbdId9V9BV6Mblfy4mhe
yX29TLl9/TMKWTGF4SnelIQ1sHxj0vKnPKlg/3Xir1vm8Sb72DoO0as8DZsJNxE9oYRLJQx3l7js
z6Xjtq/KFGNXfjWYMh8nXeXxdpds6NFb9Sa8P96CPNmUMBW4RS1bQF7Ezq9IeKoqWJkQ8PJxCAMn
LqK/euOU1cfkn0Irl3GEH+qblRZYcrsTYlEAR+TVMX78q/Ci6iwZZruujzujHApRDp2lC8k8hIKE
nbyThv1kU0CsbqtBQlpFXvVjedlncxWEuVbypHnbxRNMoR5e+qmEFNZQELMEG5F/H9E5ITXCrwR3
9rBATQQc83l72j2ZoZWM1zj48oUiupMxk9iMK1gAS4MivwWPCNQ9npAODSJrc1875EjB6OX2PhyJ
L2U5S3Jmn2akSxv74sgk7Xd9djOcZFfKPvfq2vIR1R5T6kR89eQRUlkx/97ZxLir2ZGFltxd90Kt
ScutmEy4GIOSLzf4Hzib+QP3n2kHlqI3WKrvAgHyhVaLw2HXtadeUMzkJlsiFKbk2RXqLvVVZes/
WmgSI+bUDMySvqhu2Xg31s6fJIA5RZ8o4ysqyyKKPnqUpSWeIpQNebw6lAtd2nus2+q8vJjGNjAT
pdV+oN94Fl9puit6oEhHNyzDQoMGGX03oibfv+jV/dRMP+9jxkiuddBsdN1HwdYkcmS01u2Z49Lt
c6yOCvUD+AbTlynd5dPTh3/YDqU1WVLb58h/UFbYDJCDHxwWLYg4W/FXXq+LbaK63cCH2s5Gf5Nw
DsC5Zm4kgWyRgliNqxos4ztqkXtyl+eWp/evBrk9Vv+GhOoGRRPaiF/P9h6Wpd5DkDzqFA/1/e9i
IrSs4QOMX0omBXpGBUnZwvABAtkJWtTfyokG0uTpO7mrf7/lJXQ3u+pVJpHsYtfJcEFxqP+3PrTE
7pwaoHvkhBzyNMaPVfvGdgY4m2TSOPfMGJUtbveNZoV1dgY7HMUpzoO1NkNuxzwiIYdLfYOKSV9z
K84MNZ+/1LQTyvwogCm4Ej/fQekBa/80FwI4W2EjZrX71G7tJbxE17i8YYjw9EjAGUBxsvsQGy2J
C3xdz9ZcSCikfq1OGorrYTWBK1CxzDUOkbsVhg6PYsfOBjFyBxO1AeaQjGKPKGa+7dWw/yFgw9lY
i9WNJID+CD+TWzh9vtRFBZcY3xNoCqHAQ/E6wvHGXSNCJ+spLPUa5jRV7clYt+ZtslIYi2HcQbCD
FN5Trpy2tSyFw9DdRwcaEHViOpntoqGKcvyk+4RkHvMWcU+hCPKptrEBjHSpNlUguePFbvl49opp
eNJZybJhbwicx6FPnDMBSJpTAJOGX902rpvt+Wzem8wf9j7P920HFhtRTyXjES5FmSXtwjXsjD5Q
tk75dZE4hFpyvw3gX6nj1WxebKEJbcH7FN9XKsHb+uYMXUwR1tQ3yB6/16mfO26Ov6izF6J3XP6/
fb+J8G1faOXpk1XBBViUfQgGjx6bopvsnBR49RtWGPgpRu0uRu9YrjAxLOsUOmuVH21pd93+0zso
8r6+cSxGO9irLbm3IDFqtllU93T2Wx01o2sY5Mh+M2Su5hkRG5RsoLfmSF5PgvfrhjMLk2EtfdYp
rwld2vAXSh+d4N44nKhejJGwqHzE3mUiWQGkZESUeDvSc5B3PaXZ58FP+Qp8kXRElkdrTovtlNGY
VLSKzmmM3bIGgGpZFBJ8MLwJIYuZOC6P4TjAJDEAtBs2K55gaCmW020II5+VBGLwrLznkOGEe/Bv
aV4Yiwwe0Atv+ljUZAsK1DHE95qOz04XMQmcB5XNkaAHqyMPOMdo7xb3WOXP2HUNAU5dK1EPffYC
7jahTffLRV/fSvmb5jfvxXn3RZrkcLADslDpJif/whw/vOY/35yyRFDDvbSEs7hX39Awcpr9+anN
I+Jamw0RYrhfDNXiAcI7ZvidfBl70nY4SFIOpp9yYfq1H6vrAamIe6s4gPlfiPW3ESpb9cLu02EF
Rj817Y0x50ctEJYz1UmeSW1XsLpjg7aFgFDUOPGoSSmYDXGvtDaHC9PNILRGONlEfMIesc2GsLCU
HcbIINnzIvAwbfVawvQ8FeBzNcjJGZpy0zp+NZTyjLXh6FNuH80Z+OTZaqQOqCg6PMgZ7vz34U6l
cBEycQkwVFDAsCrlH9M36u/D37lyiy5995QeMhLjzeNkzHfJtpUSMqGh5NngPXFo8EflNV+4ppiK
NCdytUMLdUu0UsruIx4bzvWm9ycyfd2T/apBCJ61SPN5CJdx3vpKyb+fhX4pw8fnSPN5EOxEPVWA
ifBiYGXjmfRPG1MN5rToBZbl71tgLKST4qP/K2BbQSywYylmQ4AZllrjqnZ1xxs+t9JSqEmpbDwb
x9d0RhZsLsUqaV/KMH0IPmImAPkG9Bu9hgnIhe3YpnxdH7fOh2+EOl2R+b8uMsaIX27nmYJNWXK0
3SXeOD3NhbAVse+b3AL8J58FYOdhkDvR9jD+4gUfyIw1hDzCa49s4eAbZmcrHpDJ9EkfnDb5lyM9
ZfHluzoAjYNHKDT/FaTMM2o0sS718ATgu8ZAtO43XvRz6I36VflQPIVm2a9nTjzs0k4Iez63WPzg
5ZqJZHGz0d69qpqVcbzmjES7Do+bEBooSisQ2nALiXveS9gYrU3VhdH2qu7zmccFUaWLVFUVAI89
cQ4/Xf9fm4qOnnK68yF+rD4INtZPjO5wvKEhjQGB6Y/GZn7W/tRE4llEEG/s9+bsGGV9g1I8zpKZ
fvTF10TxYt+bcBDPJQw5aJDnLfGvF1Ea6y8XpGnwGYl2E0O9cbIDsrDhixg+RN0x1yY7rXUzlyxl
jNf46sPXH5mT1HOUre/T1h2xC16ya7u3qY1VIHEvShFWhjccXPuLioHUTlld4PiIbMw/LtytUK/M
9Adoks9xu/ym7QyMee7mCRHUby89/izeY05Bdy0wKuDbZHkpPc4FIx3hqrtMp+frxWZN/KdkgW+k
Dw1FjP+ejgLAuZiCxRQZYRkClWb2Z8/THNxJDoa2nPes9o3a1SOiW/XnN9AiSKqCMUFZfl0ThZiO
2bBhuQ2O6ZsJA8eEtVBQkyXGqE0dOShe4DyFPrhLgZkJAbV2COheX1/+nKcZJe8U35bH/8bt2kEd
6nTLMzU406pRNqOfPkISsvFiR7LVgXK0eBo0Kr08RsaozjNlHgxbJmnEu48x+tV+yeYgxjnaqyWU
WjO/PNhnRWG2GoQ4EH93D7G7SB1zciadcxdINcmO0x5iyCj2hNW4MsLQ8aiTzUECTiWiWEG19uUy
lYMygYolow42bFHx+GMT9BpajwMTptRsnN95uMid+BYAWLPxGvuy/qPGLRKY70W7eE5b8XyzKXgV
1FQ6dthpqB7JWxN2qAMg5dCeghdPmZUpzEUfHeuKhoMJi5noN2S5d8UEdapLmSB3F1oI0KRh0Jpi
MqwlymVC7/CoaAnnamAKL1kaViok7/0dneyUnBsIvD5U/Vxp3lmrJleF+S4Ilwvqp2yVc/gqab01
Q1IYTou865t8sezdSdyqEbxJODjQIZf4MJp/TvMMO7KFwZTRlxafhrMv26hgoI0M5xTRObucYI87
gj48LV0txNzmk9D+cH6qnlofFbuzDqpFZtAPKR+CPsCpf5AcvIE3kB2ZoT3Ga+L2yUCeViKZJy0i
0xCqPaDn+exm2GNPaJQeW5JO0rtfJ4mV5nGcPLc18BpVjVjxGTTFkzBx3NRCQN3oJ5rzE5K808/i
al859K/iX99Yu/8WHAeouXAEXc92AFSzGLbgJdV+kFpD0A2ZBC7q7kREF2BYNxnTytVHGZtEiRw4
aJ1liBRGfaBMN58EPjD8XOYtoRxyGHB9z/yPs9eflS8MxZN4PSe0hvsyUznTdFMa+/daYSp1V1j9
yNXyApBFDAbuUOJ/vT8oUKqU1UehKsHDLP5ElJbFKHk5nqaY863JeiSJbQAxQ/EUMxlUrjGHabjR
YB3ZWWQasWmcC64dN+FOV1LekVEwUhDmaaJb6ooq/7nppzODaqMnhej4nv7CtA7wzC62UZcF+1ve
dbwb0Txir6mpZoefRHd+axtEEFCJvzYUliFWB6OKZKxiDXkiFXepNoRfGkT68mugpU7YfaBZEayF
tceTJ5g8H5m+Y9VFn5dX+JkWhnLo9JuPfOuMtU4y9EWAcBznOxgYJy4I21wijGLcoj5enFh1zi1P
WhAUta9ZNpkUvndByqG/CNyg6ACJM/BbUH3ZPIhchMExwaohpe+DG9vFpEzcJ6KwmtSmMrxz0s1Y
/ZW2Llkb8AqVae74WPUwnC+q0bNJf/kARGTeGpr2RneeXRTUfP32T6DfriGEn+RZo/nFpkTC3K4g
zx28BiLDKGMgu+oBgFAooGZTwgwrmu5VrvlbyrK+zwSfsKD4kbX3Axr1burIkbPLublPaybAUHvr
usV9wEC5m+wDMeAEFesOQpBKo+hhsUs0ZK/9bOTODtS60tv2vU1pBCXAzELt9p6Vjqg/ibjMhwTP
KYUdDrT9WnpFeUjpqEtQeOi+3gtSBOf1cd3SQ9d0N7MO5M2G7ZromJvmTvYvlP//PnpwQMwoS0UH
F+GCZkG0GG12QT+rKNNhmvQKOKKenXBvpal4G4sGFYjYpZ2YwFAJjqa2ffTzCnBRP9wIUjZEp9Mk
2865j3nlfDfUDy5Ce4tMIUjyTYgkJ8TfHmmvkQTEBtKDVFtFsXVt+KvPqlYaG8IziIYiELrpbFLq
KbLDdKSs7+Bhianvf7wlSFGqIS/bqf++oXf+3q2zLDffhr2kL2az0aKycfDHTpKcMNy/tETOp/9P
c/4sp8NC5TO+TUVjGiiY2kSEBSf0D355RKY8gJiEFnVDWlwE40TK2kvznrZaReKM6LfDeRKPJv/S
UMWrvWeiT+33FI46qQYDXK+dZBchbA5ykTlnyfFXQiZKgH8W54K50Ccma/YkJDZAEl7Zdoyh622e
Fl69QDcLEBsFlmBUMAZWlpGm1uPt1jVZztOfK/5biRca5MFBzpMe40qslcnEtwzrmv9xW3UpOkIY
s3BPs/HE4Pwybc8o+b/soYXYWxrzLE8CsTf2q4hgAD4Z+jwIZGMu2WLxTGt7D42R8r/iuGEN0Psd
9XNroSr9xa35nX+2U5lpBX4G/fsiIkVzpkd3nOg9u8iRYHhDr2qjAWS/tpSlTBNdTqUot1lHaeml
UhBbwiWhCanOFVKi6B2CTWC62/trECx+NUglsPYWIyLRVzQ3iSRGTr/BuBDLs7mXbRximfgjvx4e
YcfbrUQznwJIU1krUUT9APQfi1HkZZMbAVSjPHGjbP1Yh2rxW4FHsn1bwEqYwFNd8MeXHOTBkK/i
stA67PJmTD5Zenvj/q70oR6pPLbr9Ud6U+5P2pIJQtM7TudPeGrBVvkVMoeJ6WuqOZGPgmwiLs7m
5/vPRdX0y4C+qaDVx6Ilft0/mKpX7RM4ZYjAfr+E7KGsat57gAIfe87zpesl9w8RsN73Y4A3sS7k
iDiSLro2q9XjgC8NSOJPvYHm5GbnVw8JrCwsyee8MDhKDQSPoniOY/lAZpeNhtzgPFnUX7eWdagG
X5qf7yi3w9mb8lESqDFcnot7JgQqsWD8xITpJWLQ0L66fLqk4584U+a3g/JPfYZ11KEX2KNT+SeR
jrBZ3UfbtH1ynFbKya5r0nHv9HPuGLAY095J/UTbsugxjCOG178JOzihCOtOKcvv4yxy8MJAAd1i
LcPtjpyCARKwEolDvY0u6+cFWnOeSObAEYiH1Ijvkje3gKGb6/MTYjpPpCFutjLJLxN88gt7jyWi
Etjg94vPvtNfgQ+bKyJls0KXaSVJQmRFFk7PUy1vRV1gQCdT03eCtPeO8qaqJhl4lfmDrPTSsAVQ
lsYGDefxzWj16X9ZuMhTzPa2XTgXQblefiYSNpGN89xeOG21FFuqKjEeLf+Nvj5LK37B9LKs61f4
gy2gyGtbjZfDMDHf/YAJa60me81i8v5nzuO2zMubxhd/65OlRqQ7mIqiSYpE3wE2xx998KY5BfQq
0Q1h1GJoae/wBkEFV29caVsyKlIjTBxV3m1af1wKZ3WArC6VRXVzO/6N8LPE6KI2O4X8ubuCWkxw
HlytiwPKxEJo2B9HtOkNr/0G1Zul/6kR4i0Uy/eKnNVQbg7rOnjGJ3uI/xuhCnze1vMOToBmqKaw
lq88ezjnFMHOewSPfhEs3Cz78pC3xqx2WgMmTgdTnVZwSHlLNJjKjKtNXtREHiMREljTqDvHgAVO
l6CRsjWwzoCjVlt7vVnnfYYwc5iXsBTDMxV6+YOdVcMNF7yM2XUg8m77/zVSo0v9V9Bh2g44ERQp
OHutUhrwVhNECbCOuufCcwh+H40a00APYp7XaShmCYBgO+wmP5X0wNRxeCFEkMndcWiZ6FezDnAw
L1u7nO6nFP+fS9OtzQ2gkC8DDfvW10CQmebcAJfr0oVskX04d9wN7AAoRqFpAYIHUFJRnOunvu1+
V/Had+Q34mLd2X4i8o3GJ7e+3Y1DLXmpQjKcJBjulDU97if1rfCykUD2bfrsQ3oBP3kH9O0gxjuQ
cRtur4ObQuTrmXSWAQi6oscGmSgb7b1+NGOfJKfzduktOt5c21ejX2HP/YFRYF0+25Kk5bgDSYJ3
CXqe0tA1eV80rtLrbzA56IfvOb7B6yYWrxi0q5eAp2gqGGvgcQiPlVHy0+wAhJC9+hflptKnyrV4
/kkGqPapuGPnoEaEoXHeWUpHgd/M2T+LJdjKyrJzoaLX5ui9ULKm2sCfrvWfPYxvtX8SvBczewVR
cmOMbfynmF9sT0PB8oF1ZjtZBJ1G27K0udIvzhSanmrL12AVuQVHxo8V5CohKbFBWOUEz99RzfVV
3Ns9pLKVQ+AoTXuvYbRHEz/OLboZ7qjucpKljatJGN92dG2YKWlw6gwQh1kDnZgqPW0OeJdq8Zdj
XZ7knNBf9izoSBFLtN1bWU2ksZVhY58MUs96h8eaxw0Z5RT140v/XMIZr4ZNsZ2IJ98FBH65qjaf
P5VhFJ8+da0ButClBL+f+sNDwWn8c+xR0mS6Gdjh6aE2ooNPUHELt4c/CbpcMiEAMX6gOZqfXjof
tT2sqUttqrHlQmJieviaYPY774u1a4dLXkCLqRFO0t8JBgDbyPmGrUnXuYVzbXRJkIpmGz2EtcHC
DHY/cwqvovEanGVf9pup1QXn254T8vNS/Z/TP9vEC7OGsr57P1fGTCb/Ixlf0/Dpod+5Nc1FF4pI
pMNOiNC4tzz+GoJZMEJ9Vaal7ie9peDMXj7SWeUXlnxUY52HWlExSVIchZLzE2zOHRetGT9T/DJm
zmOQUs2slBxBmDXUkUSWXzkE+6yNQMj8E/4WkHGKTq7GDgH+KVJBGIKwSrT3Y1nEUJjt54NUxWl0
f1TKDXi0ynztcS/YN/Mov4+xrXEvKbOMvu2YXZXBYUg2+MDsEjm9/duJtkh/6Ao8xNEgkC6G702m
VV7l+2eVpey/kj69FPolEzyQn7R9RTAg78DGLq7mdrg1bRc1CY1ztD/I9vblRmgfdROlUg8+94HN
5UwanKotTYOWQj2qAD88hpDPPlf2MPMKyX+uasHbFchDdROQu2McXgLI8lkA3UtGi4ozDTq51S3D
Yer3QqOMl343pr+uksZ2VAd4hRhYFE2xLY3VAWwi6nwXTU4w/kb16XiPVaK951Ss9TofeGOtkOhw
c8CSmBi6+59yNYOdayQhkYKXsbhJzh+s3fflifjayNBI6k0Ycj39jnFsvr3AzQm+go/U10NwQ5fG
v2EYgiq0ab8wJ8cW5gFPqifeGSaqrAUAi83xvcMTYI190TicYY0It85mtuUsqQq+8LVVriWm7shM
FHy3WdTX1FDPxbqYC9foNrv3+44lTup9aZc54aCc1lok9hCS2FMqFoXYieGaMpdHFICHXpRk7ZMr
gy2uRUyizQy/UNFnKcWWbB+bID2xhSfBfl3pr6qZIQEdC7YOgwMKlb1T+I6c8tiV7aEeIfRZaLia
uKktp2SsvIwLww7vh70XHwMtCKnnzH3WzvQRHJMF4EroCH5GaaPzwJnJA+GlrXGUcvG7KtBU13kT
vvJL2VSn0bEnboQcU6A6ENiDIaBOA6HDYueRLq5l0PE1VyRZcnv7ljUfTudmrGPwpsUl5yKcq/0S
eA3J9hgVficZRl7l/61EI45f8jPBlKU/Sy+9fKvq+7SvNuG1PGGopXHJ+hkd5Z/XL8GrxPGflWnA
49h9nVFT/6fIFSvOZW5uB5yEjq2dWCwFzyULNTZMJ9NDI63suYOpKLSfKgF1daaJQo4/25sGd/WK
fZDNHwJ+eet5pypkwdrwYfofDmbhNiSAcvSQxqDdMu6EAWzIapEMCH5q5THwWpAKntWh3RbCpmaq
L3RECc5LEXn24U1uNUknoLB55dojf1y+e4EkYfv9qoSam0clu+LBLy9ajouz21ex6w7IaNqsHSMc
6sboY2nxTZIFi5PLa073ZzfBxftN2ZqtVMuOkICYxGHk5oTARXGWgJSAP46rxr6WvlHF/synBuYF
AUrDpqNO8SnkB6zr++2WTRRLz+adYrLEJbk0hUI4Jncq6kk1EScdVVq3D/0TJCUnn49glkyQbYmc
35gJE4VvWU6V4Z+vNPP1IV3PN430PSCTyVkyhc2ZP98H2SWqQk/HhntxiF6KoD0yRYaNPF3BUZVJ
SWME57JL6xEbQKIur5jUguiEndkq6PUUA+APZAv1yF29UsbyM/axJFgMBwhoSHVhKd8CzLao0xH6
FWIFmUIOVeYmPJHihWWRKpryQTfZ5C+lVp4wppYpOJ5fEXIBzRf/edAMs7OOR0BuSnRiulou7cQj
rxm3cH/chpR/EYnIvPm/dU/94P9CWagRgNzYx9nXqA6eSPsgYqNQXsMhcDGzl1j/IRuibgbQ8GkY
RQ4l/egQWvAJ3pqwe0ABgzLMffjGGGS/cI86UV/BgG7egQGRsN5PNem0VLcPXaFvNnhMMi0bbUgv
mRp4kXEJH2jHJJSpmAs2VapFHgBrd02yeAqT/cOtcmzIz/Ob5Q/46uHIHQ8IoKHFrtSE6wOmIQAr
Nk/OedcXPX0Gfhb/MAAIWaY1IgI9RsNve4bmcErcU+jzUfzAjZUmowSMbEikrjDTUeYuvrS2KULK
IMLMpjrAznftrNmmJcqvnu1XPvPRtJeT0ioEgwLBevDdzuo9aeF0Y3XlMNogJiRNkyGs4vA1vw1+
88Oah5STJ1DRCJwU6cEL0TUC/1RXg0lr4izPo9TirFf9SMGi0ql87KnxNkwChAYt1K8JIAyb7YRQ
9ZOPKooPLQHxTU8HtOusanwUY66P/quhT9n4CIEz3/d/v1KIVOYI/jRAyvIw/3w7ZxZg+NtvOvkp
2gsWu9TNZvKvB1OJSCXfP8kpVZjJm+Y18C5EmjlfQWjkj3LW3lCl9MGH8XuWpMlOvoVdIn0zrSQG
vEvrAzVAZGS/DkuqC9hCrPyDu29VQig5a0/UFE2FNkfLGg3MNV3orGPjU4Wcpo4NrcYJS9zO9wme
3+GhFbNWXzuTuBWauagsQdsdjDD9MiE9pkSOn2p1boPC+lhs4kvPh1eUxwkohee2pkq+FUOfckqi
qEiURWlkFxoEwU6MtBkf9+698u6DDWvNeoC6o1ONJVdEDxHwj/8gCCvmg6SjgWG4yfjpHnQ/CgkD
Ds0CnIzZhjLOfjduBdQinyOd+pR0uVSFcNePnb/jLT2K3Jv+Rst9GQBvDwaP61SB6RzhwY51jWUf
CB74vTORDzUon0aWTsehoah3FSJFlhtFfvil9XSzFnCn7Tex9HWb/DuRZWBEhsPhu1AfGx+0bT1T
xyLnrIfudCkInkBdBdPda9f7XDruA9tCbPzhB1pU32XfKNNruIFm/mjzKPNuXs6161LpyKzkm3CN
ap8/zxHcx5feAYj48z4R/lsdPprYDmbxkELwNCIswUYXugEhoJSCL0wQg34/Yssml5ok38PpBENu
I7Ahg1IHKbDjrTBu/AdM6PwPAh8Aw9xjpaKG1Vp84w3xX0qoi9+e597WvvtI/1lgXcllY23Lpb5k
OCLW+gJcP4kcP9EWMSwzLguPJYNZ/hPKJLiVsM0l8dy4cvpirppGD+x4XZW77Ese3Qd4C1rkeq1a
t68NUlMoz5vumyspvfFyep4eFFlM+IGWIKp8G1KgTvPk0WnaF/Qt4EcXZaup1tH6H1G56zJx8H6o
rQ6UUbMJKHcBzxvIpOKjRunhxr3C466NZq9UF+fJwW43RzUmLQiK4K0tGIeEJo/LrIf8leqtL9JN
qC/5l7vUN2yOtGR+pkMq1vVt018HWG6yxxn4EPUncScTYPzHA2grj7lcWsCrzvpLQw9GVEZ2D0Ul
M/zShC0Z7RR4pyr6NdslobWnLkljO509ReGXUfzh9c1Vp97sgu1ZpU6n0/YvslTZNd5u0h3OKF3u
OBqsVBf9dCKBm5ap+/GAI+unt2D70p7EeYH63GkGRwE8VUf/yl7ik5GvTfFdBIRK0UeUwj1V/7Vy
VP8cmIgI/sJPbANC/nNiKSBgYhzb+zOFEHQ8AlMpYC1MVAobvV5PC+0U3MStO0A6jCfcgiJTAUds
l69Uxx20OR0eskMT2UlKrTcCyi0WlIq2anjng1tONRsqFESg09qqt1GwthWgpicMRIkPP4G44Utm
Vbw690YWluV4pLVxZG/1s93ebc7IkZFh62FSj7RyGrdO1DXwE9UtrhgQScF+FSpEjkO0R1ZVTER5
p5r2BI6DW+N0vdjzM/7Y89WFyBGOsmX49qcyrWZh4L7EKc8YbOIlcS1IxtLbshyaAl0MCGXEDdv8
jxzmNYov8hIlXznonxx//yzC2gp8aQ3u+hMMJqtO53QM1dVZX75VHkkxgkGM95PsRrNFGnI4qb/3
3wMevbESkR6AD4hXHRAULc1nUbHoIlg6npEcXgLyEEoIWluIWsCSKtkw/ie4R+tuWr1nwdvddPeC
K0u5qeBo7C2VnkheTGUZdYnVPn6cELs/KE6te1Ldg8hswgpIaqjCduN6sJbE6Ib8CBflFPYKb1JE
/5esUnuIE6xhMh8Mxss7eLRnhkKG2cfijE0lLt1Shkfdyid22oXpenhiqAs6AFsGgNrCI0seiCYG
O0JgS7Lq9DchKCfx1LwLJXWIKCWm2Z90kTyolUSTYceXAQPvS2+e5ZyiiES/AIRRoEVXWiyhEsHw
CRL4f4OxH3bKCIC8p2UMHz8C5pbV/MmFDiiJF9iIFkc9uDs8k/VkdbOz1T3/5U8veFsODyjaY/Rp
xsouCSntYZoJzIijTt1axJGM4KtkPns4PLRHEddLQXIMrfp9iHkHMKhf2Ppd8/+D7/PFX16Pwmgi
OTaEcROPM524CS+0OBihjCQfdK7qgRpqpYnpozIar8BhNgSU+O9R61lfxVk3hudKLWCQDZnOyPBl
iFhVAK2ZATTFuQ6ql+cBJVUO91ziPpm6V2a8NpfcX4N34TBWZiZqPN9B65mM1xQ/KAhQnOuWTbWm
tIP92D7I93GOLr6CKR7sxMAV+OseQOo/cEZPOO4XQQDkiO7wayGxub0aMRVQqVEUu3JLVHu9amSc
TMuXqLzYfy9GoESOKRYMV8uX3y3MLOAo8era7d0jk0Nrj0AFAGAkY9NbL0d6cCILO4/hSYmkn1AT
S1ujmUPVKedPTb9XsgO7H2/AKO2xG9hseOQDe3FYLAr1gUvC05/anOww7mSdRR8/X8CZxHJi24b3
hBceAuHSDcwcEBsF7j/es2t9ktkLEqS3IqKc6PGMtMNA9Np8Jc8bBiVdTwsYTo+fBeD7MAJBGGCP
Y2NDrAYMa065hjIZz2NMeieY6WdcSMWSI71/pUm5f1+i4r+Z5sdK4iqetwjTrKFV3fNhEfAXoyAg
C81d5ARh7CJ9VG13BfsJZgRoioIfi/BU8dJeD9FXxiukWHg3PqW9CrVQbZgDjJd2N+QGctUzZpI6
yVAHzhKDLSIMdH5sHtuTxHO3396rRHUjHkpLY/kMwIchR7J97hzXpOEw6H8p9oQarhXmJAitK2dC
n127fgz+Dw39vdjdA47vmBSdjAm4x7eWXxCt6PEyT8bRY5dD2V3IJQR4oOzI5jK0xawBo8SDJltX
krwhplZmMyaO6vnlnkWw1mcKEH1QDtqXGy9fFS+z8Wr1DyNFd9wJahvWHMU4nbQV0LecTRrCaQiT
mSL3tln0gevZt7+hVl2Vzpg00Hi0ZFeCGJ1By1TtL8SnQeEp5xPQN1UvuPuu87KOj/h/LfPwmG6h
x5h8PAws8YfEniJksnOyMET8S+v/FVifxdzUxd+baCllfST0jgWuR4gYa/6qmbLFu4QjOfBgLjmI
HwWLoJjXDVJlLMRRoX7kSS0z8cYGxM5CGc4QobsvWb0dmSrps/Yze8SD1w9iqYswzn/u8zJCeIYz
T0OheO079JDfzfvVYwQeCehsMm6/ozSr7MjwFXA7Akmv/FfVkxdZwYJJdvpUjncvYjohGH3G+5WR
2ptYE3fixGF3pV/xlGqjCAjv0dcpKVCGQAnWhk5In8M72XE+Voq4KXfP/TJrL0SZQRmCD7bxlb+k
y3TP2fJ1Yz5MRf89DUOnrPR+XFd5K1/+aekKkEHsHipGVzVGakgnfZUn+L5knxrXx+F96woC1GcF
8Xc/nqR368l/eRTcCti3uxonYpAY9NP5mpgsE4WKoEYVkDzxKc1VHnOzzousyUNNd7cCcLXtyE7L
xHcl+U/ra0HF59pnDMlVpUMFfLfO3l0zh5a67udgHxO/bdEJMzxO65/+goASvIAab/94vpGzVCc7
B1IlrW0YhrjylqN1OdW7RxAMrY6EUIAFDvfmVHivVoDzRtUDnoeppSHVjtV0kFUlkz7+eD+xL1o3
SMeLja0RBqf2rTgLLtEFYujemZgoFDrmUKNfaWHqRzgleuMMADlfCcNPIeJ2rPEei74vlC6XDRlc
9Sm7DbmZP73vVMyFtmlRZmPtt2+m8/gFdye0Q/VcgweDZHMWX6RM9BMA+4ZF83M2pxo0BE2nshyH
U177yeTxZLq3Q3Sx4yoqml36Pm0dAsKkqw8ktQCibSuD5lQ3jiHSW/HnNJSuYw/wLsQvLf0rr/2Z
ZBtaOUqC5U1cHyC0GR9Eyk2XN8HMGNpIJrR7ZrbXfY4IheAnGpu3BKC0gnMxwlH/Q2LfuQOb7GPw
dqSutjBshTBfXPX6RznBztTGS3JnRcpD2EZF/Xh8E5Zu/BPjo+Vv3pOuzZwkizEqAnTAzGGK3v9j
k1O884NVik5IOtpDU+YnIUjQAlJaV7P1r807G5uJdY5zrKn0Cr64AflombmQc5lDf0o+QoESBkX4
NOSSq7qRIYhpOYsiYE3u7OlW5gXIu9Cy86Etg18oSVpcvYpiE4pOtTi7U0CzReppZxP4oxIPcKml
2LY6v8hlV6PZSZmi0OxqkJqELm0aaj+TmbdWP1d2Cn00n31yhQJdd4SpspACM43f4RyzIMFDcsmH
B8zvtxrfrUBi1ntj/4fKEKp98GkT/JeQqR/guWmLkJlnmwnTpCJqx+ncEqH7nHvfo5Lc03XzZ9iQ
LyxhglEdcDiMGhGm6fgZKNPw3dlHFJ/lpY6ULvFIlRx7uzQu4HNTPqYEmtSSgSa94gK2g4W1fKDV
T079HHFHCbGCepdC6hQWLXuCBkpP9KhgjSYT9sE8SusNvkP9/7/7GxFAM2QpMkpP01TCiTN317Mu
YTc8YorBWzoWgljIkFndXCIR0viPzJfFu7Ann6v9o9DtB9ohsSRPMNlBXGBbi6JgkkkHQ5SlvhWM
G3FGZB1PkxDOAnerTyCZrqTtyIdCnbT1nGGw7fZPEEPWvabfOlsOKdaA4/Swe/U+hfYkW6LGudEb
RZlvREfKA65orcmiRdT4rxjUna27HD0aEL+mvi9IfogQCbjJiKBo5LLmfsx3emiEEvCjCXnY6IbM
xDx90gIjrIrp1mC7Ph9TN7XloPbsaQqO9VwPFlgowKZI1Q5VeI8DNrJCAg4YcVFKFAJ+WWz8S/ly
gXWYxj09B2bFx102ysmP6SuUkuyIpePPpks7Bo8DsO7m20ZmBGcxJpPCHgB0W6RDZJ6CkuArs4XY
pC6It6gHdiz03Uwc1W779AFMbyVqy3IInWzVGRgHkpOZYKKrDWQWzCWdF7UCtgw5ycw5ilDZah1L
VuV3DBKsoDyrM24dw7IW37snnTA209r74ttB/PksM1LS2pR6ewsz6MqFAmr9WRJmfCN1aJw+4wqG
m6Poqq750bPpeY48bklcnsM2N9Z0xnizTYUHCRCqQAxVVJ4fVvoB1u8WTlAFPtq10h5W/jUkkYcW
kFetiAnyrU5cEqH6YhK/gCs82gF/S8Th8MpcrGyT2S5rVDF7WHeFQxCJYThWbLxxOGDSHiTucbil
HsooccZR0LLsHKazHCnTbFNTtaS2VBDmEUod9L0Z5S1DyX3WuYmY171EXn1pPRzlS2Zs04TGY8AT
aCVMKqkZFUBTa9NCQUnPR+20ptoqYaSlGJyI0KqM5N+n7BS9+HCzayH7nWm3Nhru+EFxDt3rfOGs
No/OOm0AlaHBfVxhp/B66R8Mb1LO/ov5jxj+rRe2Mil88cFIoVueCYllbdM8PJ8xbPCH8nA95pc3
avxbQIrxr2C4gbABkadJI1N8vWLw/8abGRxFWmsuOXNm05esAGovb11PkYv02nbkAEvfayOrAp5J
S2Ss8qyYKF4bvw3CMmtlLv6FD7h1+lqk4BTqfZTIxurofMqbkPv6fkWIGPTyy1PgWIF3WTN2P5h7
wbHoAwFgJ5Fchv3TVmNIH6Kqrh+eKOHHyP+7TPcY/eRKF99T9f/t+xDkTHdIs848kZb2t5XFyt+q
DX+DSXVZoWff1yrCm7GNoqnkouBWJ+ds5wLGkdMue5aZp4BD+8Kd1ZcLyKroibBthS+btuW2jbpa
YclficGGP/FYDKIx64DF1ldj1epVN2lRsFsQWoeW8/0ZLVT0ITyXMaYcMf99U36dSomNS1up/H47
cG3Qy3XGIODFIUSI0aB8BoazOjfmm2ev6yq+V5A9RF/oIVdSzEW4n2tiYyVhg6D9vcBQir6ZkWhB
1Krksw+EhP75jLCKHxxH+kxAasL3HO8vStrNhUV6pcHWflr+ZGUtr4YB6i5WQLxAdWxBbG7KVy+P
E96MLvgHWNZtl/7pdL9T84relZ0g7QDXUXhreAsw/rZc46fvujpnPqXnXWuDk5f9Zd67LFjLKfWt
MOndiU3CIEP/4bNwrlaSQO4UNWTyUudXRHTFi8dofFNpGXpYA4X1icgWIly4/abn4yx9JV5xoJ64
gfTvC7BxIJthy3KwnZhUgelRd9RhLIY00AREN+/bvr0rWqjqgQ1bkkpyGKVqPJM3ZfX54/viYz/+
ygBSgxpkiCf+upqo4nW/EHxYplOA5ojkXAhclB+ydKYH/e2yireklReXA30u5hKqdIFtbYj1g/xa
mmCuiKMDWHYArXM1lX155Yx2mjuGYP96IKBw2MpONO9dYf4wrw8/JVx9c7Ssl/MvdprjrziPxknC
AZztZa+VlTdfOMW/stD9SzVs3i4SI/i4D6Ckr6W+Ym5WJxNdINsop6sQN5HwUw9IFVFU8vXEm8we
IXtpHjRfY0JI9QHenLzT5JLhyYHHtHuU+9pix3mTRqiSKceG0T82qDkQMdL3H8Zfr1sJCOy9zlLm
kbtOuaEyZ41snGpKyaxArhJffVGBoI2hD90W3cFsut+kG11Le89T2xSf7Cw5hy69uFG2aUTw1wRk
Gy0pDCEXE7L1Y/gu6K1lNC2KjgGo7ycYjHr98dIbpAnqgrA5a15vziLduwskEHLXna7Hepup1cd+
9IEZuodWIiD3ddZtnR2veLNtIV9zQiODqJNukU8U14FmMCNqGTKzYKtVj0AHlA2WKEmRebP6rzsg
GNYZzcRdTk+PTRRdc/tvZfBD9kRQRfBjpwTGI+zWG7XJPuJhb3E2iW5SurCP9WA8L3BtrWu3uVfi
UoP/KnjJ2h3MJehoQxk8ifUZWYOl/V3TdKWxnaBINilX1/RUFeNXd4kcrsak0eMDoufFo4Fvd65f
5vH15EY9nUTpaFE1YJ1dvRxQDhbOvlYB7lM+TtuGMObvxLSOv/b8S61b586qaAwYKjVlDUJt15sM
XfjctJhTij3MqDJOchFNQ0YvyNHDS1/ulxDiNqe5GIy0E3JifOhuEJalDSnhCCpxsaGXZIw1sIH0
itmE0bhC1K47AWz899Wyad/241i3TMyuOGl81E6MAgdMoNeBhSvo5/aCNEvZFAtKPgPG0DjnIxB3
RqXteBgqKbVD563v2LlKztqguRl0EG00SeokqrXzoE1+UsrYoGqT6EwGav0tpPLQAuI4YOT2BUtd
W2XxRndpMRtzh6BcgLnjtniOo3VymVliCG1hMLoESTJiEH6A5MJ+ukK7o6z+G+PA7bRhUMpCFeMu
RWFTa1sgWeHFxLqtZgc6VGwFBugM52Pz3+Sy64s3qmM2FsDfpeoycFOsxd70Dg44oryeQYh9K6a8
cSFcdjXP5QtKoWTfTpDSN4JfjV1aeXo6boO/vWr3TjLB1WTFNji2rBSLxEknJaePhcPbRh6NQeD+
2ZkVflBT2FEwQdr0hJbXC5E85xflnWTMpbi23cjdsVW/zvcctHSWbfy/EjfCV95eVjzz/n9+C9xQ
B+f4w62+TzdkYqSU/+olfhXZar9YEgIA8P42PFjnwSmpNqQozKNsSN0Bh5fwuJe8HTcITZK2Tz3q
MeCPyUH01aSCZgSu2wUX+m5ZWnCiqsBJxkZuv4OB+ZvGHpu2Q9hDhUDhxkws7VwHuVWSdvDBk4Gn
A6h44AgJs9MMseoUsuSxyFQ2Ppspjv60IuMr8E3FUGA0KW66oiaIYGuYaT25JnZYnctOL66wtPgc
Kfr62D9hVN890AHonZC74vYSDUe105Y/Hb2d0zahFy5eYur568pslzTLnJM0RBFgoEtYPFCvvVZX
WZh0yv1QWvFJLkH+6d+6zEWk3OeNOH4Dz5bhvWmu8MeMb+5e3kOFXkw6bFMjoF6CWEhUmBhU0uyR
Vg6EHgeYyWkFDuRMORcODx/CEAbDBZcnKT541PlL6WnxLuagfSHeCcp+7FfbJO1i9EHtvU4H1V3t
pNLCOUEk+pPpm6g3m9C/sm2bLTy4ukMdfiqIqCky5pTknWMOXBSy8+yS50jQtwsRbCwV9bDKU+6h
ebOUGHbo17m5j5bRMcHE6JiVSKjP/sYkCO3MEBT9uZUafd3tQBJeh0x+MNbAiD5SWRkVAw+PunBs
sd/d9Afsng+qDs/8fEbncL/Q4v1uHtNjvsNs/Jz8KlUZNcUJax3EM1D6S9PV6O9+6DCigKoRlp3e
qwVUg9MdRDxswQFPAsK9bHLsUT39rcLvndkbtTC9FBd3IE0b0rwHxPbaI5EwzN/iS/ckLUtYOo/1
jkH4RCD2pb8OADrR4XLPKxTgfyzOleFn8Zu9dy5rl36mvE4mCtFCU5IuEowaru/7dMZq/IlyRfZu
HHRbNDIh7H6ivvfDgA0gAxKQfHpA+U8GKwehh6qqXH322n10Thb6o/iAaH4bPq2jUt15kR+VHYmv
6VzmlK8igil4I9l1loIdfXD5OddvwupP/sjDfP2LZqmQ1DBtnvbjEtwXGxJq9Ht6j+tSgg2QAdmp
rBur4uIyDG/HSoJWRobxsWYr42dJNAY4OdoTLI/2Skqo6XsYo2HEP7/vVNam07uCwkyeINGpdThY
vr67XTFzSMIGBdBQn8TIXrwz9smFxs8SOVcQ3FXXGQ6chxW2LPDInwZxoCOlOEpHFi09UmvmXHTB
ANEB4T2NHgbTQVh+EQv0JVmNP5V8zlX5tqf1XsCW9Y0M9mh66N7nBJw2R6CorNt1v2gx29hwav58
iW5Waaq0llgfJGotb062SUQuH4AWEPzrmBpjho5W3ErRDUEo9P8I4xsMI41GsgUhYdaiKYFIu1DP
ls+NBY2oodTE+F2AO+mHLhbM8ahBS9//t7r4XA1jFdm/sRBO0TehtHnflY1xAs40InFk6e0t8ofY
L9lUk4Fy79nV0a1N2Wqg2CTlOHgLt6uj6FpAOEqGD9YA3dFRI5+W5or6WBl13IF5nOVz4j15HgJ/
2g1ZaoxosvTLHhZgYnIbEvG3An2uAkxGS4mDc/oOFx/CDpI+jY4cZnV81aarzRBCOYqf+nXGToUc
31xJR2OUThFOLi6pZtX6JL5jXTQ9k4Vg6o8CKFWn0853+Q0By0AtA37jq+/geYJcnXWb6RJy5kyX
FpCupEmcVPAcvRqfj9wgqzCVekrKeO0OjDu/8JqBuXc9BEouEdNk5X8ae1tbS478AVFfFtfzCPEN
HEaKUViNP3REPPTuAOLQx94FhqG65VwI6rVKiGCwL8l+D2TF0sYLM0PJkljXm721Hl4VCbXw77j+
zdfJOspCQDNq3CHjSGcmFhntq/2mf/CZThq/c5p1wMM3BJ/ZenY+nDx3wzUyAyT79B2XVK4kkE4A
NHDah8hpZlenBGZPgAK7MpGTS/XqUDxRmq6tvctKAvOiFmGPzqrK0KDmxCpeLZV0gLchGE922nyh
jc5cUXVlhwXi0CLenahHSmBm5W4a9f5pomJ1juY2xtd/CyXrKzjQ4klRCQt3XHFA7BbDqrdrsxVF
cXEVLTMy2DXPZjcs3UG7vEJsspWVysiQxVobDKWdRf0C2hoodXfwonRp10uHYi1Ks7XTuwF0Pfbc
JsuBwJqKQb61EgzCOPwymNc8WbrFMz6kUJQRqGL0UhX2JGFResDXEBB2F5ZkQFE3/WOE96GJaSTz
Q0pzM5jRyLtUFBjQQwTGZk3fBmvkbK2pC6NV2gf0JDdS2jcjzp+Ijv8Q5AH3a+ieZYQgTny6NM6Y
V1R0I8Jdf6NKZ7qF6WHOU3Lt8Tx3BJs9Dyh2Ze/u1g+39+1nrKvqdWAy2koPnVppFjL9NC9Z5cSH
F0XLJqQ3sErRm68hSOJLuOsgZ6488k8zbBzMqJ7TZN81Wezq7H2A0TWhIrQWgL1VL3Zb5TNIm4Dz
fLsHIGS/hA50ird8wsxlTa/PPZMjrKEwyCHxTd19u9iCWnF2Abau6YyHraSgTe//gbxXrceR99V6
Tsr3kULjMHkGyKjxBpv5WKpLIRnrf44wZiPbyjkSL4tJMhqPu3FDE9jrq93D216Nm7nF14aGckFA
b4ESztcjw6jNFFdCr+hLm8PIIrn6s+hTvSO6msoyaSajWqYzqoZFBDF7vljvB6ZHU/gbhSUiHkBe
ks/iGSRC43oWbanbBc3qrxTx7whHDejPE5WLlGbrc8diRjOqri7ChwdLqVhKbWV2B8wkEM8LzglF
gDrQss2+YiPHro5HsdyOC83iPRKBszd/H/iaNo+ujrE1myXzmGdEgnKwSEyL0Rp3BgwtvRtCaFMc
qROVQrgE6EeY3KmoEJlEkETC08aGVvcgGJr6LyWxG+Fd7eyheXoncFVfFNEHasC0limue0qxS5+P
B2xAtjYmHA1tMV5B6ILAhPx0kfRboLDFuYF06vcEMLbpgDDGaKFQ+16syhAU4QMr0x7vlgmfa5ug
63xanGOWMj1Nr1WKMbadBZeRG9Tk8PQI32ILNUTUv0WVV7t2PuxsoyRYxhw/BoHf1FxLuPVxjF4X
8EJ3xBAEhq+lae6TZgyLrzXU11+TGl8e70scOPjPYV5ijWPrhGjsNXWMZUMR76MGhhkTScPBPy9Q
8sGHmeaonwxseOXC70YI3CG6vn3T67QpsBBjoQ2wR3YFDxK3OKQZaUpc+rwdUObgpmJHHLPjBRQq
pqcBNnlNU7MQ3epDAx8VxsN1GCPwP5bwnEPwXZyDxgj+4FH5Hq/jBDiXtv8BMgfqzyW7+vNJp5dL
q5puwqrxNQ8ro2zxz0PAzCnTC67HwqdvftLXgFVmR9ynRNghLOVTFCOybwoNGtF4if1XJZK8PX3c
jBfsyoyBWYrP0SF3xCURa18o5EssDmP7uRsB8oTBYjbh+/2gamQJtyAvaJcrvaCqeq9xl0gOJJRl
LUOGUM1I0RkyaxkRQ3xDBYm7MApWBWx/geilbhNyFPdQ4SghbMfQY0ly+2D2NyNgMkgNS6+/YtJ4
yrkB6qNVfOd5uEvTfrsdaVn0FAMovrFPsSeRXzEW/nmSmtm8UgMwjY4+D8A3nEm9qLSwDpxXE43t
55AyJDpOaM1dupchNm0+RsxxKpKghLpS6GosCX5aJGwxghBfMCgytpJns2K/F/hVUkqiMzBE4zoF
7sJkqYNmTsXyg/JcKa+O86l6jfc6mVxVHgXwuzBsr8qw3QpMsuLdLGo+tBDVJfEOQbQRHSzxafyc
BAQfiUffn4jmBvZrYkdv2lr03Mq7l3XvvUQnVCK4oaes3pbdO9DIFlwnydTBHUsBJTmnYw5Yjm/0
O18nRyfhsebANnT6e5ZiBliHkIObrA18l8gF5Go8xa+LhDYJ+ieDAcFhvv1Hfk/GC2Wm6oJcYmkt
WPKsNWmmI/fzhH9IRFbBQlCGdSwQmESh9xPi1P9Ts/TW/ZZt0754cZl08Lwca7X/HX5PRY2mBU9o
wjoUCjaqau3ARRDsd7oYU/j7fEyhCGs3xQEFq0UVUQQIL8RAauHeM3ggY5oKFqBJ0wCTnM/9zunL
LZ4hfgGCjkLMfBV5a3V3snnkfFA1MHn2DnyQci2056TUt4EJ8z0M9H2fF26QFR0jFyHiiUamIqgn
JjZ3blx50QxQ7LOO2hvJxnQLvRc3tiWG/2jr0JdmF4df07BRfNoJ8XY3pV9SpyaJ1hMWHG063ZIn
1YbRIYRv8wz2FbLo79Udi0Q+DWw67nAKXhy5lPJrZAO7YoD+1qyTPzADuYLM3hNAzupefjSnkIMR
zQ8zgv5NSZi/BNtOaVMb73chiEWmdfWm/AU19zz20rfx8PfrAZZNydfAkcn1JXhNfpFCGoMyrOM0
xV5z9BWI0/rTIVCjLny/dprhipdzAoiI7XIYKOtlg+SlzsOQSrZ1Ec9PCdFXW1VOIYC5B/6I7x6o
UfUz1FRTqgyr7iOEVMVlhyTxOLhG19beihwGWU+SydK2OHvahOkPTnjGFAEVUuUfAO27v4Ps+ROw
IJIZwh4zKPsuIA1w3dISVaB+JHV/APQWCL6S6gW1xFjgCtARWiiAePO60gfZRsrdpivwilwIJ8Os
yN8drJyBD/A6/J7QWCmgV+neue5dGxgh821Ge5/iSYHAj+CjtvWYRot7D8cGKUtEV6uh88KgK284
44t5M7sEYWdvbzI8i7rKvjE1W0700/5tuisCv6iPc4KIEHtQhKWHlwSfoUScvVz/P91PViijuIfh
Mnh0CabLEe7y9XvfdQvLpPssPsWohq33TfXyaE0E01p/qGAltn6hgjL+sXLO8lnS7DjK6q7wXjLY
j50xsFbKg6gjkTvMM0ktWOLUx+Lg4vDSGQT/iGQEXqh2vlLPecSerETQllHFYJ+8uesBz11pl83O
IDjvvN8wxuuV01wbGD1HMoYzn4UxmAfc1uNuj8Ar9auEVaDMQq+S+uHchQWDzQAp2bdDTaSzXrYz
RcnwgJLmiOEjs9a/4KB5VXeC7tR5qVf2pIIKGOYhgmgqUTB5XlKNk7cL06d4JCArF8Hr0q5R5nNs
+k8EvVVVN8n7SpSCflByaboEUnlgaImp2GepEn5uPMTk5td6rEmA2KBThkla05i1Wc1SMWqZqKtK
sPzP+S420TuDRKcQ0/1h/kRJO71lFCsqVUkbx/Zd1n3WMVAm4H7OpTTxGDOHqRogQ90IvOzSQKo1
NqnEGfXEBelIo5B5OZ6tX/loi0lo/E9tE25VlgQZd+3+uNmRAUdMfSf/vTwJKGZJfORYaPEkyu0T
2u7G6IEoeznFj7DCAuGOjcV3ZW7ARnvefw2McxDTTFwHONVtfr2WvkRuczfyttRs5WVBeC7IaMgU
wxjdCpk6RZVdl2dDyzFWKvX9oocd0Rh/3isgtBGLfOIJ2473H6hvqZYolay/l8A/QRaoUniRtHGh
/0Q5xUM2GonnU1ZX05WWmgLcU3jaEnTeyUqXqsaDn8h9qL4n+Esx3SuZLuHG6QLRXTlqdXOA0eGt
MBXa6bm0FqtFzO+1FpwyP0ZHTlY31xzlagqWOhFfoIv7UIVTuGdAsVw9fP+pe12PjXIHndbiyKoG
/u+KCUTYCo7RULu6zRAL4eP7qHcBNqSvOWgzw2CMa7HlOlc6L2DrPVsy6ckCrmOzBRTFeYU3QzN4
wwIfo3Esq8nXf1i71akWhLQYnq/H7StHelSRWKlxI4BwYjTvcEG33PQUw0H6JRFAw391wLn2TXBj
sWTy/t473l8Idk4+EWmxTRCZQQGl82JN3YcCzCFo5WWzGNTBzCJ+R/kEbMWEagZYlAcSxAWRFp4F
E1oUhrxRcqd9X3qdWevNimshlg3XuEOe5ntLxgSUqBVB//67sh6maQQM4GR1U6/itRxySC9IdGHn
p8iJQNWh61zKyabQdm5ALRkZXa8A9boV3WWfkYx8x65KOcmSgBXcU5zbUQfgJ7mEC2VfeajugJxY
YfBUMwpJWHMEMRvsIKbUAQe7GAEqxOJRHVXOYp3Gm1HYPcplRCmk1ZBCHn2mMN0sv2X9aYRbEpNv
EXn6Grik1rHiQa3FqBJ/AdcrrgfLQitiiaSUCOPoa9u/zU8FXzfJqZC+Vb/i7zZSBc1MuUsmYmPx
i5stlR2rwrFSSGUs31+jSxCQw1/cWMUs68kNopOP8nbf+WAVZ2ncnk7pFBbl5keKiQ7yrkBkz2Hh
q+Gi3qLeBOwcbbpknwMrvJoXdHjJFGNEvu2l+2aaQLoTr3pIj/SbU4dMcefJVBczgtmPbi4I83hD
Ns8vosapHJzn+96gFZVA67FJr/LGFQCEIY6hRwPmV3kXD/cC6NukkTo+mXHWiAd7XFnW4XUnBVmU
+9Lpo45uJkz7S3eHuww8Oaz/XWx281BizyssqZ8Dj/jFo7Dyh4SIm9AnPMP/hJFv4QOjaqkHbXQB
AeuakXw+bRA+03/OCoGiB2YdrAPZvvcBBA+1VQMRkg0puIwvxJ0Ojqy/LZ4bvKY7qrOMyGNEzSVh
r3eywxC1OCyZKVUdShk/QVqRowK9PC1QGAJnVFG4UatkMbVz9UmhgJLU5mq5+pa9u4zvJiO1FC9p
A3xa5UFePoxzGsnNIP5A9O84TXO1xis/QoSRil1PZDby0EjAu1NKK9UL3RgVrMaQ6IA/rnxuzRPl
iHG/HBhcfl/YRLTH65IXbS6THNN9R4Zj6ZUyhNZmaLd8nOvdHrv7jg/PHU3+tnqzQaYvczJDh6gm
3t3EQE7gOgazbg1Ai7jkJCGlbVgZFRZqSGe80T4OljQUA5Cz5/uIs/F56A2NdVbgADnmH7FsxMJv
FisM2+5ybu0aUKcA+tg4UrSKPDEi5OF0Nwh1edfyGIp5Qmhzr8OcuR/Ur8csGE7oXIBi55J9iC1M
fb78qyH44JcIGzB6vd4VBRR/3fUJ8QcNi7AJR1dUavVeIdijfHy9ataaQXlsqAsd9zGHxKtYbLxL
SLZIi7H1cWq6rbNztZX1issF2GYWdebtmoO561DL0PjDFV5SiDozMXTKO3FyADSIRrj5eXbTJTFy
1Q/hSPHnpFsxLlI4TM/U99tUFcjta69JUGIbPhsK5bsxDfEQ3qnMp/p2hiEFykCr5RrsFvaBtwdJ
ORMjv0aC4fSpQmpmrEkNBD3msBLSjEL8NJhq/1RBbIPk3VK5dPrwCyDPJK3n7/MVStayg3jntXUq
L/igoewlS3Q3TsLtF7IcqIlqCEV8IVFbSIuJAiX6bWZH39b60PDlAl/tljuEhySobWx9qNpCr3OZ
lkd+5OesTkpG6g6o1F7KKE4K5ojKzg6vU40MMNN09lmz+pfpSC0Abpv5XGu/8WSLqd8y0JQLdb5y
8MwampVsQwrSyM3mme0e8DlR/I3PjQVyNSte8WQGUO9ijFsRCTvCryWoJ1e9X5XqenfFYzyzgYMu
HEKRJP0LlVK1jsuhFxbE+0x+29xL04bMOSsXMEPdFyU7p7cS2gY8VmKPoa6R9CXqItGE6/qgvj+D
4XNTrQrrjEvV/izP2HgQAqIUwY022waoxnJyaDhJI8buvjvCBcsGE4lWuKQTooCaIXg6eD8t+5Sf
nN/3x12jny3OI4Zl0GP+H+9xU24NXtC0W5H+DwZkaAHy9tXwoC7IJ8ZZjso8AgQcaxXA43grRQj/
lOnCut7vFwEiX0bMlX0HT4ArvSCLtoC7/sShgZkuCGixGGpCKAwqhYyWIs1L67PcISnfDxWG+iyq
f0yjt4KrFKkYmNW+9VipMtg6Y1OpdTPrC7jgWuF+ZLhb6JpfzNG64nEfpOSKSYzDC+vQnwvaPfMf
TjZ2jGNhnbfwnDVTFgfD8Ud9L2dJuPwD7TiUp97TNscfk0QRsQGJ46OohDR1sqpweLfzEdFtvTNR
sh4TKIypSDwJv3tcIoKe4E2QuTA1K2exQwgJY+oXx3NM0+Q18zYMcK8zmaQ5speSLgYj9ZHKwfRi
mNCWOgZjVBhGbk51tKsyRxVuVH/7Tpv6Kv+uKHWd8uJpesN9xvLfMZJy1JBWuuAB7B0HYRBJI5Jr
yyrb60A36TTw0HYBR109CceZyjZQt+ixkD5cCkgUKDAx9841rmwfDSj4ZhU/C3P3+D0EaTrdQg1j
a1Z1bzeIYKLNT7SJRGCkmW19FMi/fNH+jbUKeDKvQ1azLnuESl8mNgTlA4jPXB+heMoosOK8Nib/
j1/B79phqB+xeTTb2/rzMWBYQ25/OYxU68v0ZEsVnoO2fhg98FbVnzeSO+HPFnC1XfzPW12LglkR
/oWYJNgrgMdI65u3iIUvvynlqVfn6edJ7qTmF+w2d68iPpLEI6D2MHkCny0+yprJUbBJE0EYqmrs
nUjULzcqHPppw8oKXXx6bfYxndmnvMIsPhWoH+DTvTbdGMKlhYc1pQSbEjUod0Dg8jqE00G6gZOp
TW3DsNReRUlgdfnarHOs+ibtSIn3xB1EzmWxWfgjjvl+GiSPfseFwhx+FlsJv6o+9UuG3w4GoMZF
uZXdNqklW845YIcl/TYePUeD/KQRXCrDAm8V8Z3VJv9vreLL7/Ej+E7/qfItfxdPpPRue8bH0v5N
GK+ool3WZpP5y6kaLrFG6bpl6Ea2CssCuC5R38zE7tUClFcakhXjQ3pskMwuRyqJQlU2ti9+nmGV
lKQhyMQ5w2XPmNNQVqn/R1aHeRovZyIQeOTWIqzE8LaQ4bQd5lD8D3LI7bteVkrTiM2pm8Ckd8uw
k5NDI9BeMD3A1eXvoCDPdKmGujJLGNELOUh/67prVKrdl8voRbmLHiaknRrpqH9p5/QwZh4rpZH5
kbSXD345TlEYseXFCA7Al8B4VEOkns6rBJ1Z5eNPqIMIMzqRlFUOySdGnOZ1c7+Ew27VuW6kh2LY
5U7d6QFD0DXFsphHFYJMBOa4qqizB/6ycAU4D4MNB0Oi/5nNBsAir1IpX0OVv8eFsEXgpfblro/5
ScW5H7HMnPWi3JeqWvJ6MCaku3gU+2VNI8rlLBS8KZ1+2VvIifU2X+cmZzipDHAYdRDrgBwmnoc6
erNmwDPWrx2absfS9MROYfq+qR4BwnK29mAI+qI+vhs0LOXXO9aUahgjvTWdfFzhAQ0a2ucIEUvv
9TaWMQghOqK9K7t4+ld/JpwxSrEYVNRiZJnVbA09F1YtkOT5J9PlmwD+x5a0vUMCLDRiKuV/WcJB
AzpNAge+mUdEzI3G94tInwg3VDWZMnqnDwS2FfpnVlfx7b5iDgs5I3wgZk2vG7j9K+sc50TFWv20
ECvvRbx2zCWUYQsTXeGjop4WyQp/iaIye6ZIoOr5/QEUGB9UNO0ZStwCrS/mLUPYBR36pZ5fn38c
GPl6irpEWrS42R7AAjX7ejrjW5QmhhE/ZH+SVyCian3uHO6lyUhqxE5+sG89tfwhIgoM0HiGKGec
j+LLOKWwbAZc7tvgih38fGF2S7r+5rlCgQycD5+XhJOudj9+NMZ7L7UPzD5OJ8LgTs3a4ZGGhE7d
khl2zV3lfGmb0DS5YMDu9x8JasbzzbNz+0GFG4TmC+olqkJ/idFpGsnQcFcvv0FvzG9UinG+sh3v
Stor26JCABqGtnwqxNYCfd1PBaNOPSqDPgZan9ePGeNMU0XbwZ3KjXQajAofqI4ikjAHbYXXsgZl
ygATEvqw5whfnL2y0Sv1RjuDGGSQajM2+uqHQdTVcqyIcHKGcj36WNXWjNMpTQvTschGlxLRcu8L
9MwzFUEWv0DUsmE1csOgU1NZtx6jdymG69Yy4H8jfHkhVFlftasTYApsZNpbNS97UD0QLCffRrRG
hZcDk3Eg9XpKeb3luAUJhiGUoaoZzSop8vykBbBFz+kqvnGTPmJRCVvJeX7Oo9k2gddWOzVaFlip
6Zw5qfQYAjhn90jPuoqZIxNlDKa7Z6poQZAoQZbmEHBRDkmOrtI81+XFL6TiiBAR+JeFLSH3xPsR
URRyGsE9z4GE3vTx1oynk2TEyLbAtfC0l3kQrIgX2FoqfGok7ekP+eqHHszFziyuGlbKoxgByV6w
XWA68Z3QKZveWi07WSXOxdNSoGNu/VLaC+98vuhX1gy3jkq0ZXaKGxy2dNSzI/KQM8bv0GhIacNe
q9BR5JHIy0OoygBDXLJ1t65k+fHVU/WpvMTKj+s446HL3OR3pqkbn4SPCYRVEyswV7MwH3liDOB1
1/AAsTdYz8iz+CpZkKVA7E9uJ5oZGN42RkuKQrfd/0Y+3WKvqNGAf0C3An6OcGzI4VfZ5Epbw9Rs
UR8i2eQ+u3eQNv2lHkdy4Ac47uK3eCo+TnAUhFVXBlQSPyZGd/xMclcyfgIums6lIpg8wldK7hIv
SaSH41GxSWk0khleba7axPZnRfed6S4k1VIKg1U2y01B0uLCiw+j4gjYfvAen3FUCGlwjTPsAPvM
oi81m6mOmyWYC89zuA9UjMRqQnTPmYD5IjxKGum6UfSc3rqrQXz6h3PoC7RD8hJpfZJcmaZCYshF
FReiWfbOpaXRO3zjwh/Euq7ChUIGdfBAb2wCS7vleilkjCvtUGr13N+sQpsry93gXzYnJs6npV/c
BmatESUXOw6E5jq/L8SYdcv3W7TZIAWeMYvWZR5bj4CVl3Wu/BjIrE4twhbm5p8wclvG0lPfRybJ
QBHN/P4QYeBx31QiGMLWMh78Qv8j7PxNrXHDH8zL3+7O6dLMDtxNN+0TDwQPD78f8udNQ7RrtYlZ
OQWSAMGM0n13hiwFGCxgCkon0jkGpCAZWgE6Klp0oUjt24OKF7KaTG08Mm35te8MQHT3fll8JcHr
EgVW30CGNUvg/oNvLEPSia3W8+TNyPaHvZrNqZwom2RtC9LAcw8WCaRtje7gIOISo+Fe006niSH4
sTpXUsVgFYrCDwfdd80FT7maV1bumS3lHIThM47ovcJZoGgKt1I1c6jUbrgNlSykJOJ9ov33tG9c
6t396Ky0XauWorrumH+u+gNhF/qxhxj3X1SXVOnIl9Ygvzkf0CDVS8ubZeiuYcnMXhj1bnDVkKhR
/p6ngiFUKSgAb5qgvvQmzEA4a33zVjLhLSNCTF6vLwaEePDNgl5pdjuiIOcyuEQUynUO9a/AA2xS
GRg5uyUfCoSVXFEk8H16NdK/CAIE9SyqQu9dNiJt763xcG1ywFSHA/DJtDLadiyhLnOZZPdbx2Wi
H5VUVQ8zmgzgNuMZmzDx0Nqz2lDesMEaMoNmX49959pqYPNSNPSeTV5L5D8nqusjVqAn39XtSWNF
8D8coWnms2jjfBdHf/4yaCUtILh5qzcViKq/wMO73l5CIXHGnSpn6pjNGMhpgdZC1WXUdW/9wW5q
1g9BB9gLXw4QT2ho567zd4gm5SvPMB3mBxZyAKGGlyeE2C/XnokbegLDNJ5EPE2ufF+iXxxEoNmz
dPYJ+kIW6JQW6gKpyQI+fgtVWMS2N+Q4hJ3o5umD8sg0Q+mVPUQXBKFxM7TgWbPulmWMCRnMgZ7j
NmNZbND3/xDezozfzwfYELzJapY4o3bUxLu7OhCUw3p+4y/41iCBKSo6g1iC/aXRLd1ebIpQY4kU
TNXaPrGpFN1Ujeqa4pF7lF2j5TtadPtpOzA0fsCFTJ77B94FH/g4Ji2KhZPM2ujKQqUdd3tp8Gs+
esbyDlvOFgwqEOELiphewOiosJBjXp7Tl6wR+MTlSiyj9xLKOISCeTXE305w5nd6DfrS0a8sEMjW
OW8BSSTk56YitHZkrR9d4EhjoOqbJleaTDeDwpiMloc5gH5HmjEbPaWze20a25NP8BTYPHwCJZxD
Ak6nD2DdFkN1fT2U0psnk9GOAqK3ZrEhQLc9DXOV9OMS7PPFa3gItFyPqe/3w2k5Ro5MvnndF4kd
1mS5f4vKDS+T867EO+jwMt01GIL11u3Mb/Hgu5M/8vENMGKYGqbaT3Q8b3r1ThyCfnEn5TsLEwGT
+EOMPQC3FlAUxw+jURwrYbi08YXHVxobuqYLrpAzRF1BEtfkGQSxWHZteslbKplrK43wW+B8C264
oOB87+zkRQJFlTky/+MSzwx/yJO6axSy52+jHy44E8P4oSkS516VggjPxd4LqdFU1LvSoDAtAdTd
kSJu87Ler25aAD1U/lSEdDnyVaB9ssPB8M71cs1f8nq2/tuelDr27FXItd5HpFmV4ojeUcMqcGbx
ltlHTrj+pxDB+olpfbMQyRXzlaFeUjq0MSZSZPW23efHPptfQMN9TNn0Ts9eijb84q4TFAOUfTAM
h9jKfXHDZfxjFZfu/XYYgRvScEMwStCat/2ymFcC/I/VLWFUnTqsR3X/D8gnqGevTWcd0nXh3WBF
TuCoHplkw9xneetlftLyiQtkxXaou5eOjP8VfLlquLfCqTF4xVsKd9HhySY//YubCcrHV3tkQF0o
YY82HvTL2elCZTkQQjOe2mhWFzuEOj3kB4svYpnwm41dvNYQpKakb44cOoJcHnSSUZcdGWVDTqZq
y3Utidb3ORhYnA/avC9+SILAzhA1SQzptjXkdcyMtmcYOUgQmiJKZBWhCKQS6cIs7ypi/D3+P5Ew
x5t/ff011DJUGW1y6/EHSHPf3tYJFm3o9ZRQdJQg9pnYy4zwCkjbkhleJvqmm0esk41MdjZcog91
clpywguZUFbbowmhvgCL7PodSw9RcywZ4SoN5/RMPEMa4WNXpxYu88vZIVouYhtsa87AC39H+H7s
kPn9M/hL885pom8y3eYCAn7iojg7kxRuwqUp7PKU/H4pGmxdVcAtwP4bDcFZoOcZkMfgwRfC1eAR
K9m2YVJq/l7PlNkv0hBwIbx+4EzwW7oVPI0CKq1YwFcCV/QINiEpG6KP0Z0hpzHsIaaSSo/BeL9M
OMzD57M2Xg324FLTqsfU1pz3oIwrXMApD4CfhacBU41beAgE6e3hLGuKUbJhTqZmd+O+Pn1iBXNR
DTjmJ6QAbi+bXz86njYZeSDdb+CtrGKtNiKs0wL7sxH0/JRj0nCbIIR19qSLR2xbMqU63mFWB5tr
ukTPMR97r/ADOpdffZRkF0tu3asaXGzsNyGWIr6Xnwmvrid5fwOoR7SrQMIYbbheOd9cIyNZkDMw
cg5TpEsh70F9ksDSer4qJD2myyqiMf6cFV1DqB/73lYaPulB70NSIQq9IB8jUNhzO+hxSwaYkQ/o
Q6AidXoegZy9x+6ksaEQJkgQfmF+7ijC+md35iP1ygUyH0X5gdKR5AxzUSCmmaeMfNnxIThKI5oQ
qD5r7HN6wdIrBM7p5Z6uOXOaKD3Gmrke8BFwsiobnNQC/zjABqqGNjhmzjkbkBGtg1I/7BwsnLhd
jBIZsGb4cJPRr51VMwSwW4o5GYKYZBuVHNjhkkfwS3rvjDdhj1bgr9XA1AqlQgorqIxfJ/wDthQM
3lBnYeuRMSw6l8XpZH2vJLdcaZFbzQKZ51eqV+/eOW96wgIs08RHKCYnN3bh0TGKtzCpGlJoGa5O
/jH6vQA5aVSkzwMO2dXQbFM+4ZeI2drSJ1VjPPr7pcEzBy+NghiUqbTTs9nhz9OJx4/y+I41fySR
1nRAd1SXEKQfzTOOMb8PkfZVtKd4OkTbMlW90CHYCyFBXWAb6U884YhLBhoKeBNqOja9JY7BELEH
PlnXbikRDpkQboS78igyBXyMOiUQd5wK/RhKCDZ8rjQ3qVsRf1OEr3ypDmOH7DbQcEvUmioq9muF
LXNC8Yfv7QWmw5gtSajMpE85AERH6TJcEOFixEAL2ErZbTP+HqEY+Nd2yzUX9AyhLHdiOvyINftR
xCLK3d4Z5pe9vn4pOEUvydKlFk3twkQUPjmLbckhobX0Y16OZqqGQRmoyaCx0PXrC8A9PLWUoDGj
qWa0mqkEVGa7SnJ/JBulCO4Ko3MBDkgSxSPp0Rgvhy47+GDWIUMYpfNVhwZ6b6Sp5Nq7V4PoKVZE
oX/9KcOyiEnyQDiU8QXKp4RLGvu4Q+WoZtiZqWgd+g9+w41LO/teV6jf2UM3rUVBTmIF7SE5qPHP
SKlwJdcPJqrrEt3GX4CrPYmRr2UtrrH89ILHMhowH65XmKirgL2c1KyyKBYe/ZjX93kHE21O8b9s
mbKgR29BVpjM4vP7JfPIM1M+QMZnP8cD+h/T/M1A+Pa2ZHrEsECwDbHI1ZubObdUKFaepS7ruyiy
UAQ3F0bkpTDDmOMKFpJc3Ntv2QQhVKKY54VS6f1NmiRuVQ+bk8YiMVjXcXCiJwxF9T47X+wVXg+J
HxI37P1K+EGnGXyis23PUdhLhiOzzXACh0sjscbmTpSmEnOvwaNRlTX3AEDquZ5oi19CaUMRyq5Y
XpooXiY4FJ48rLbnZkx7sjQbRKzeGQrnuxX1rlm1pSnXB18hgP0xAPwxxmPpjCZo+D9Gv1ny4BqP
TgMEQjgGWx6kWgpwr1SLiF68YAiU5QDbdQ1MC3wKvVdqE44R79V7YI6mT6nT8ZECmUxIwvFBilBV
LXayDkyAWUuOtYA1EwFgwORPW75J/g3qt94Hzjei/LXFTEXh5qL5+2rll1hUVRV9HqCO6lETm2xp
WYAOnE4uK5Rss7PPAEApJjaMuGnFwj5QGUDNLs9zp+V9e+eOIcciZURTtsfh9s4Lei/gVW+Z/NNG
3xAx/JoAj0Vsw0kWNaQvyOcYRuDS5SNHBEBMMIgXjMFYvBbC3L2p/aGai1KPpuG2+TJxbFVFw4au
p8WRj9gi3WZce9ysC4X9dbBzQWSy8ltjyN6RL8uXXVe5ZNewi29CevNrWXx6UDODTVhe6af4ZYyX
6i+nqBRRC63oz6Kg/4Q0GlaPD6BnZlAapEsM9ZZ5FLkjKd3/zinf3wNEVaPzEndbP81pkroN++bc
Ejrno2omTWJeNqcPXMToia9exkb6mvbJHy7evxkUNWGLux9QcCHrsrxwkeBRabmoFqStXgcVJ9p8
kxuxznZbZQADhRcM+k/Jf7usGSWaoVt4z19oDNvq5VtO/GtqnYEbrvkPrftW7eT/8+/kkoBbK/I/
W9h9LMdN/SdfHhrP5aFzYB30tKMmq0T23HmO2qxzMqnhsbKkxVwdRC4hT5HkhV616A13jTeZMc08
IhQwHYJ27ukyt0ySeJtrlF0anlGVYc14uTiy3dp5HdUtUuIPcIiSF0+mNkDRRUk5w9aEDN8iT+R1
tlzPqOQtfBH2d3zNZfmqs07YePH4yGmgv6/s3KOEnnwJ5i3hioxa6zBXWYzZzT2NM/3nMTYBpBCy
+2i3vyI6nvp+1Zjr2iikNTp1ZSydFi8/AnezDwe2YTvxuzXfocYoXFBOr0vbpqMP9FIGajcNEWyO
fmm3EYoQ2HcjBzk63+GDyEVoSjYJJI7bbfYUUcJyq5YrGpLYAd2W9caKkeXCB0P58GnAg9ZAGvBc
iXb/0aqyiv2h0W3xc/kPIHMK3p3EEByt5yXCmiF5OU+8OshaGboiLoc7D7UXsWcu7+dI3aL+fHuQ
ERZtn5Eobj79YDE7MWO6P57Odyby+DZmfaLhre3KmPCD5tEP2xKWAaH8ItGWbD46oNZpTCtoDQsw
yRYJppbpdR7bBy5rRBx7REV0/nmKYCDnaM1OWmXh/63o1wh6c3SRMhITTBqOF2GL8Wt356Gz9Gzl
aF7YfZKPGHjWRRAqgM8uQBP/+jXeuYc0+8iDLN/EsRF3/xgiOaJKL9MI9N+EREAzdEZ/5hyjzMuw
qhxT25s+H2u2aWHmJ3WWO9YwHD4FYA80I5r14WB5a76i7KWIzu2Kn2mUqyS1XJJQAeMlIcXWNBe6
upIP9pK8Evqs2hPqB6rgw673rwv/alc6SMfaaEYc+tuAzT8Bhq2cGdBEy5zr2wuVPgNpvXYn3U1M
fiNEPXDDx/KsFtt/5ERlnLIeGR/7QhhDKChdzEPwtILHEK4goKY5vBgHZqYeMLm2HOStSOwPcmgA
S91EX1g5UHiZcnk1Y3K8AtaTKbL+JJv30+vFqiYF+EhPO7bvw6/UC4Zrz9kucDXWcuV8VV35PFS+
9GiThXkoKbxboqi+NbkOra7KCz4E6an8C1Wxt1h0ai12D56pCKdJo67F6iPU2b9KgdMWSExZHGlc
QJIfYl1Q91ZbFpXluAZaE0PMSsRoVs8pzT01DM88AnGxyNG+kO5WN5bGNnGrG+kpqaIV+03z7jNK
AuHM3FWvxWbeDWDNWTQWbuGNzP/6BQN7mA11RivGMCCp1CUREBuaTS80Z1eW4tmFPsogYzUU0GV9
DSTHFOUhoopti2ximJ8wPJBjx4haMVy4/M3rnXR4vHOA8OPidvDfNsk8n0NDhmQGgVuw/iOUExuu
abim1ECOIn5FXSoZ5ZJuGbCnTb1d/ctUphe+XeD9CO/zZShJVzDArPSlu9epLsSZyPqprJWLkQQ9
SbPeruC24AmGShYGQbrq63kz5YsSxe+sjVJJPJWAkp5KvANKCf4aFkqz6t2rdeq4qzXXlS/hNTiz
YkYp/rBeC/hvMECOOBkIxSdmZEFOabd7ZGRrIZq9Qvp2ebWKeykpkRXvEb0m06pWzU0WD/VrVaL1
2F0uPpWcBrH4vLTsnlLCquRUAjxDtQQjInyJzTrCLT4qEmufwBaxIPs1XsgyYicgjZIT5e+/gHdg
3Tj8hFYVFSYgtG/Dceo4oBqM3osHbYV+FvZ6qEhG6rjCWHmKmQ1k6DgLZ/hUEJCrJ7nowhnfDHjk
/nyEVagJBAS287ZkCI/5Ylr2qd2NwMzzvqFP8nRs/9qCqMK1K4G+oA0SppGyCwZxqG3X5G93x1Iv
FSEk0qvTtAwLSliIOcepkBnXEwSZyIDgQbLyShbonWSvRpKVNnuQ9ki9G7/QWxbeafiLG4owEeFi
V+V1aWsPMyjoG1zb0AIhkDa23DAxxfSkMSbbsjp9hM3Zc9gsDTuXSWXePd+WetPKwscabaaW5Imx
n0kwIlnlr+zY74e1hK5DgD2FTp/lfVAzaWhKL7PcRTNi2zew6UOnM10dEp4rpgmZDwLDd9nUr5EY
aKD280iUVR3Ox/Ko7mQuLO8EmeFWBvFO+VXnyn3ktHDhRwQh3VIVQGTOBEkkVB0NIAc+KrhnWds6
slfTgd8d1F1/7p0U4CYdzhtaeZlgJOhTEGOLga9DJiNopiFCq7XvPUAjRNRRdG2ssEKBjeDnCqc8
p4RFcj1vivEl51Z6WzJUAN1aOfQ2qMas4pnqcgtqqRb21SolAq+wJxSJcMagBAK5VZOrkBKKZq3P
+ivck+q/ijZLPr5PV+EyzVCcsxNqM7oELxUEtld+E8UWEtw9cyIGBtB1E6wVv5WT/7jt2bPyC9dN
Y4SdLQFrwAFe68WPUol2gXpBhCqNe1QJI1e+sXyVdste4vNgGjQbQBtAHoO1htlmYn9cNyU10xRN
3zI5ULV0Cr3FciehM8w7R1QQHVApdM7Qzb1hkzQZBnSWUZWTgkgOZAn23kx3ijijzEdLnM+8SMZm
KVN2c71JMRGXpdMRNRPQjp3YQDT8Ct986XE8HjRjk+bIMXPklMMSCP83JZpeqsy6ZdJSxCztpkBy
TgQNXrsOIUXL2XSVR0yrqD9niIyrl7hmgID9LZ7pw7iiWRMNcfDQ9aI98F6hpiRlE2i2dHLOOUTN
LB3EsC1cf5WIZu7N9wvy/J8ynESLQfg/sSbP1qh0FdeVw0qF4ae/g7CyKFgWDYXyeEqAB2wrZCAY
Mo2MQ3xaSrfIyuGTy8I8Jd41v9UeCVTYefyaYghMV4skkUZAPXRWiZ4+aWenYeuk077QD8OTCqJv
4Xk4fbP7OX2Nu/sCtjWHPab6bNbegWu9bkWj8faVMwwn8cj/zqZl9LY6r78PNWKG7Th7NDpaNLWg
jqB3ZLqsK4LmkVTPm9eLH9Jt2YFw+vZvZMxffpATvxMlE/icnSJikQcpIyhjYsXkYdQ9p8LgYIMm
Yh2rr5HYH8CO6weXBXW2lVZRN82QUxV8VPqlX6bYRylplWiDPKqxJhKn4gWzJCx0mCRmtC+77nuT
Lc4hm1IpF3jI4+yD+xOJixNiKfVxge8WVPJGHupQKHvLThJN8IBg+LEn1vtp0owRipx4BvLlQm9V
JDRzOgEaShH2HFJlBsp9ZPDn/epCmsy0hjrdqByrTh8qT0MAF31kYak4A6pA61sPq+u+JdqR6Fw1
dPEXcQPP8wHz0hajg5Qqoyry8t1ZylmYpsty8oyZw4t7OWHhC8fG2pyvHH16AlokBaCXAlSWPv3I
YreDxLBmddzPoCwKQ434McjeK+obTPITXh7kLD8zE+xbG7ka5upyT9SyedqVp3pvuMUd4SYQ5Bj3
NgIkl31INQkdgspO0o6086pMNWDBRADmYcPfROxjxkfy4d74R7jyVR7KeZ9XQfm4Sp/PMYN1hlul
GFjSgQ33VcStflNrUjtek8Sd0ley2s3JahFvAavefvS5eMltZDq7K4d6xHtLjDFte/fuhXm27wNk
YYFlaJ6xuyjvviIW+3uMaGXpluP9aD8QVqz7vLQc/jgH/XCBj0vJGqKwnBuUkoplg34AMtXuNZOr
qFP3rs0PTenrRSXtNkGJcGYHmvbVDbEuTKT4bC/4PfmcWM200zmgsa14wJ2+URynHydjJ8PG1DSd
wO/SRvk2dGr0yOflwveZ4D7DOz+B3MykB1AkJV+xV7Cbq3Kl6HW6U1N2C5cQ3r+5+Uhpqh1D1Ljg
lOcroduuviANlmQQvB4d3lDmZMLsnNT9EgdCDwlffoA3RZWSDS+d5FlZKPRhn+6PslBG/1VKq9J0
0NijIF6+vO9Le+by2Spk1K9KPsvCGCMcPAkDTsbGBSwjxIA7VQWRslLYEsKgPCaaSt7LsVn958IC
9t0xvCXV1PCBPG5Ku0TcXHoYoipvpcOnoNdZuyPvURequs3PGgsXRfx/0yuz4GSBUxN/CqmNtILk
9bEMSuJiqY3d7LhXGj2txjXIhQ2cw3QUxszr1cfPUI9OYdMQkah1kfb+MyOCzy84xkihPxTQuuUK
NRpxAdeCxYwt61Qe9VXxFR8Ts7PdOE1YToPW8H3Qo/IefevJtZJcNP9ZHD4lEHX8w+opInTGMSZq
IuI1xHJ41uWrFGkYCgzvxPcqjtQboEk7N+DNegiSldBfiTf92nwdTSbxHZN3N5rNFpWgcAxBEBew
Yy1jT1BMy8VU8iNSouhkFRqv84hZLqNQ1xffAxzsllHhFD52Uuc93sdbEFk1ethRT0nB8LprjV9d
aOG1xrH9L3b1Dl2XxUDL97oD5PA6jjcGkupqjqQPPMUiYzIKGKuck6/xpEJBaEwJxkAIc2eSJyrV
AqPDgZ+3YU7TPXE+Oc6C5G1KPsWhIwSUNo1yPt8WWO9NTVZRt6ja2jAVWs/6yTDMJDxxk34zt74+
uhFZHp5ae3XwU1NUoiWhXzzqq+PitvpCzyF6JZHlYJfxNA2LEXCABqbTMSUeO4O3Vni07PKoYYA4
RegDPTTIeRS6xlpMOFnb0/C0UDvzgTcqGQYskUWtSib1tdMQmsd44Q4SFlQk+YTeRZO7UCkr6xEC
+xDLrQGy07n+jvKI2tb22KMlg4KVbmV7sFDRqFSCEPUNezg1QqVX5B0HW9f1Hb7j+5HnwlB3zfOS
g/jzV8cStSQe1xiGz9G67+1n+vZj2oIEO1ciEAoWNUQn8oWpImQsdc040szKWPmPtYc+/Cx56Oxg
tQeNas/VjHqrvxzocNo626UPbXONwEoWRxfZGRSsGWuGCFHqvv/axtyw3AJuZAdXM7ndcMmxkBPT
qFY3I0U33SchYarQGaxXQk8RoBHWO9JCTxWkgw+hsUXNjVscsfQ3FOY6GV0c6zgBcMqjuc+cwoRw
0FodTShZPPOU8Oq1rlODveNmsGkrRiJkIKSVKVpmk26aDQiugROvQ/DU9UrfYlXOS+TQfd5kSCjN
pp44U+VyVBQqay0GTKvjLIiIvP1I5rJcvSKbyp0vgSzV/6sXMSEd2hqFH890B8ydhMajnHxj7CSh
olJybba1a4wRyQaWr85ZXF+qn4kN0njFioPPUtXyb1Fc9/XifwpYRKODnerjIlXKLlOPhGTBHYd7
5B9e5+lERDk/grKzGjmixckNc3cl2wFANnz1TvcQnm6BNxkAba0oYzqO3jywX63s0wuJ6miRcSUJ
bRqA/jg83WYo3yVqdLGLQOBVh3ytpEPqqq9fAhI3427PIJmiFX9SIFxoJHsKS4leolTIlcI36Omy
EQ47HvTShX2391yLd7Uz3th+AYrzgXPVglgXGjo1ivQEBXiw3Eufrx6ihoHiwA/AEqJuNJVWzNQZ
ASpUZyZr/iZjaIeKyKgGd09MvKATvlt7MGcQKD91u5NXcgMUzzhycepOFpMjGXyyaOrkykAGZzot
959cTuto/qs8ltP9auzMh3EDmbpm4fLS8njjqYis45fzXQMWlyqmQxKgldIOiKLdwuERoIj15UST
xtoEqZSmQ5pWgZnESX9ObDFWuzYmmyf7Mzw9y2hwIvwYU942p702pJFFt8KPyNw7y/SMDvmBgQ6E
1YAL0zt7YNg9Bu9WcATDwtnpw+DPqeTDaOLEkFJ8xV2gENtmCFvcSjfbjfQvgSdoFec0h3XJn4+Z
tBErnXpUlhPLSGnWXKG2VN7QB7k4HRKf/V46dMYxMJyj5UsJGxo9mdXGvuFdZJ1OR0U4QbRu8WbG
RPFAseCcfIpu8U7ubKsGWMj+/k8DGiUETXA5KMGt5vOjxTSMcYHMQEXuv6UbbUtkR0zS2RtouJWL
/OhSRc7f04BrpH1NGG1OY/he5o75YFymuljMVm/hPJ8+WAayrjYDCZQgLRXSCo9kdmNSBKNmoqrk
0PYIgoxjFNtuOkfm8oGB0oinS7EBebXghLFttd9zvdAj88LFI2JGFoKeEtGuAkI7QK3og1wSzP1P
5/MkG/4lHZOKigt2DJ/Uytp7ryEAXcXs6/ynliD6p83dOtAlHbPk0XAh2pgYb9ygSSRe9/AhZwNF
FUnvS4GlLYtWgLCE6l1lP8ajkfKGA71IUc5wxbBUPr8mi9bTWuu+RAwtm/t1tCad76WRM0VSjzc6
THyKfATC+OvM+scwIMBhD4bUJjTDaXhk3+5C1ILAxVvx7uvfS3OBUirYe6AmkOUEP63GNZ92aowH
GmkUdJS95djCqXEjpHUSYnSRrBy/cuXJKs1uGao6riG14sa9yWEfIgtyMXs4U4Mn81hO4hoTsB4H
i9IfOMDJ9yXkaJQxSft7n94NHL5DyTke0HX4shcieMXEsqPJaRwS/1gk3Yp5FdD/D2YMWFdVbLzo
SHDz6+hkwexXKZg0zhTBVJYnZIbCBXBA8pjISlQ1BIBTrSvcuqj6Z6sUFvJQsPL0Jl9A3+fsDzz6
QNVQFJzt6cZ1j76gjRa9/4B4IJs6Ydp2gYvC7BTYolQAVVCt7vUKz9WLFLXStvZOvb6qInY1u0AV
Xn8Ge/1Lxoy+lRhc9v6XXQPkA5QHJJb1N850UUkKC2CWzBEAU2bDl8cnoUKi4bz4fS9ojYjdcCs2
nBePtLEg3nkew4EogI7S5IqWIqZ7Ik4WzGlcRmpS7Wxvc0krk/vgAEpkCV22qoA0h9yB2TPz6Fps
lALRDLIltG1SYGEpwds1kel+jttxnb0ItEaOeFAQvw7MvecC370tVpBxFox1i7d75QL3ATFl0dYO
K+MPiixg5H/SSCFuwrPC8VVgS8i3oWwJ/kP29X9t7QFtD3VOnIfaCAzroZHKugrrRowtSKC53/nR
yGMTXIgE1YffJlG1MLsTpkp189rYHJRcZfnkyq7N2SoU7Iln7IsttDTWx5Pztdt/LbRLlFWm2jIs
x3KTt+MA3ggT1fozLP5ueOfYDHS56OjWbG8ppi2XPss2vI3kxTplYn/ZQlweojpUUhfImtD47Rnt
usR3UxPPCcYzxsFvbLMnfNw9p0vacw2WW9T7NiGFn9Km/v+UebPPX5MK72QDVQnkFh80XD3nShJ/
TY/K6I4c6/PtY7vmwJbq/dz6+23aJd3UyPJCbsaK/fQ7YNEdh+ohaL0Fahs9s/g+s/Xgh7bL6+4V
wnSlBpUnkyHzXa9Lo6Kila1cj8SV7kMcG4tJWWIwvyEHkHpHzZHtNOvJZQF3xzr3EMNDs1v3x2Oz
AogVJa4/PBoz1K8GdvpRbBsw+hkCMsOfR67pZLqmgSOe5YZjUBaLy9QgF/qll3EWjrFRKFSBy/Vb
UdGaFJ2EdpD5sPIoqE/VI0pHz34uan1Xf0VNb6/M165YDxLLj4WiZJGOv4NbyHdlx+dsIUiYzqxI
yCIwb256pCnYpIEcCTxe6Y6gkgwOUp2TpdWcOspis6B76nFGtL612XVkN/45l6WQObHk407iou8l
iNJxd/oy6oZQUWVHg+6XPNWvPdYq2AAXHw8V8fkgtmJTzTpctB40yA7SWFQOwa7fQUwzi4lvVugD
heShNcRzNcKcFjqknUq/HUfkP8qu3qyrlYhC24UXhcQdMdAclK3Rn6CX/Usxl9A2EKPXcxj/5oYg
Ec4Ixw7OfpinSW+i6QCLiZt1Ur7JS3zY+pBpa9xBCwe2nEMWGLda3J2CdgGxr1lTlUEW0tAoK7QX
wIkgz5leaGWepmgVKksu88ISne9gCR6oSBdZxzFnLStoLMzmSP9dh2VWyEkcQrBCdoikIepImAQ8
AL8xyWIrsPlwE6r0KHktbqdT5iMcioNHjBfADSUJzDM97DG4/0n68AXM1Bs5Aq34BZBsN1kvToos
ofdRbWvCwBdKvPWLJsBgD3AY2aC2c2qYhi09OlV9WgPtQYAiAckCiU6k2mKVvCR00gE+h+c/4369
ugvsASp3wqJ/e+kJWBYTs24gP5QlQAW59uAetXcZyNnnXmBLREr+PqAqurSWTUsNwd+GvjFjF3dD
3opnywo9LONcqjadpAnFVaxLT8Sw9VsEEyYReZQvY62s5kpv2v8rvDPYJ7h4sb2AYj3/zlOkfIF7
J6G8M3rSZCRmfD/SrK3kxDVLunUn5h9fQ9LFdpolsS7QLNmwjsa7KMsKyQtczFiaSYrra1y0dAGQ
9v5As2Lvc+q77vflyqYr+TMphRn3tsDmM/zUSMPLNRlgD4nNfeEswhAZQ1xOERkBGqwKYuQGY9N2
qwbFLVT+Etqd+6QFlCopN626ndf8KakNNV3YpRYQV79G5tHE01GswyegjkhR/RJJ6ngFsS4el6+z
11Tk5zgEi9RhhQ94z2TWHvytj3pgCJZYK1rExgQxTBJweWPXJzSE3b7ltxn/2tA+HRZOC+q7M2Js
iCtEZLmC8WTV+T0mmnK457A3xaNpHsRQumw6iYz7+cCO8dJPLftASXXn329f2jhAX73pZZIplX8k
qcsKNlbVxbypXMcOb9GwwxMdp8Qor8ttDiNCzm80IVlerVijY8EQZYP+DakNEZ1jyc8N+RJjvhTC
Q8lLN0Y1tg2fVNi8VFm4sjl2Fm6i8h9VTIrhI0+iMZtXQCFsuXIZU5YpH4Me/Xoe7ChaNoDPwNUx
/uZt0bJtTiH6h//c0WJyDlzNqJj4x8WJdCZtSYoXqqHZbRx63Q2/kZTO08zLuxMBCfMPx5gXL6Uh
G7Bm8okTlrSQSIkAh7uKzMq/H0cN3aMRMTZPR05rPWxc43SBsx4BZyrPw96SdlgB25Ix5rRx0JPz
6qxqy7tnOIK30flSJcJCHJPx6eyxEpTKgiZAsxn6U9/wjBTmGNbmZYfZSZB7MgMvPlRt5z3SSXqm
KP9LQkDajv6/Ypx7dXVEelbvTfqhgxn8rar2lC3mM1kyxeh53QD5eDuzTtynKgugoag/Vp6Sto+S
6GbosFozqURxfa4ftnojB3uDomRnVnY0jDzGh4IXyoAG9IBKSNcU7CCPaj22th9+0qgPx/mq1f80
qFxct0eaToSX0AV5p8VgLdWf3ec8FQElMU3Gqj5LWGBb7YM7+yIg2E+a7GTzSZlHx7ESoIvw4YVe
PSzi+urL+RGgHKJJTx0s/zzb5HoXqwAQWazq1+UhK9XahVk7maqCZo2RJGtfTdcaL8xF1T/OFkSN
tmp2vhm7pJQaZ45CPIyPakHF16m1eug3mzko5B7qSNPfOlkVHrp6liOS/ZDd/yG/Xfbl97slnLPA
7HiEaB353iGWtjvLfeeEggFr63DLdB16pQzSpVdj7QXXDu6Ik8/GvroSgPXYCw3+GplXYbF6aQzy
EvqEzEDIBCABbmi2MTRtOcNyvWcH+Yl498lHxduf93w/8un7n0wVptKkIVwosvatsjM2DVEBLJ0L
32CZLZrJ+ECftsYhHj9t8YDlBjnXLvGToEmD7BFrjwv3CAH2v7HFHqU++ZRwmjUTNM5glF89Wjok
5hpVBjF5VuAyYvN46CWuGD8uMhZX47ZD0hYzJZruj0UmQVrlNoHESuf/6jYt85Z3jmZ42XV/2bJF
DrMxZlW/HJJn3wUtfd5mNo/bpw05/L610YzZ0M7wgJQHFuUFS5c0PqopatKHNJZhxPWkx/TpHXaF
rlewGvsJvmaM0tYadX/+0Rb5b5/OlWHV3k9+C2IiACoFZG5aEzkmkAsQVRLPbGLnIkwMUzrRH+Nx
IGUNze+6rIv3Si/ooLUxhOv2u/nOUFVVV2i+N4Z4Td3Zcde5xlb2yvGGviLm/Kuu4SGkSiOpzcfJ
efB/QefD1mcnqraV/TRTgq0XgQfrLTXbj5cmqVjTUCU3yG6jEV07IXUwAKs1IzQSYVGz8T2PDRgL
G/ksF0X3RSNSM0eoO4BiBBJw1OdT9Y5z2QUX4FvMmy08v+rYtaH7SNJamb1g2+HLfc4wBO76mheU
UrryANLhmtG3mEa28PMM1wzk+kbtDTH9sv7oydQ+1pLfcrzWtITkeAzI8C7z0WOkJ/1CQtfq8DIt
cC8KMYmftAqabNZbyZDgVdPC8pYg9y8jmHWN7bdbCxw1InboA6G4a0aqTvw9SGsO7h9oDhtVL8oQ
JkhquenEH94XN/lmVR4vf1I0wR0+yWrCP5jwpNpdxSxzqsgjwHxhUTPGkqNHR1lQQTQ/+7+fppB8
XSL15n5Rav9kmQ4QDAfRKm6KFnEHSaInDzVUT7dfpPzDk19Aio4ZPybTSXyeN5jilgTaT+apYGYA
rpDz2bsJAbPieFQwrnF42ui7z1KtnXfhZ9D8jPYF2zOVwwmuC0lKVnPXeJ2bmvCRovldmXN0iKfE
MwVbpUgh6Pzod8HiV3xedD7ZllxgYvqMRQGr9dnZ45Yl/ZSbebHEAx1t6RgQOzWY6g8BeVZlbLas
383uiUc6fN50/1ggV7LJATkT+mTOxJ7xb01+ReU7z79NBVzfDyxRlRDJuNwJ8PFij2mL1gXEAV9q
uAXZh7qKXrg37AofDEBUkieOrBRMKQ0lB5WT9heePs6ZiCXssLLJRCLl9nZiIV4CGc5P8DaT6GmH
KojdUkWJNg28xCiadQbmvJZIQ/uEFqhsFUbvuf1R9XB6+kf8ZIegLoLbIUKJFWXAGjC5SmELlciI
KQwZvpMPBdbLjt50f6bwI01KE5G3WB2RRtTdyNrq2uk767DXisW9uMezsrdluZ2X/oznsvjs7DRG
Y7W3eWSKWuY3r2jxaiP0ImVV0em2FynSzJ/YWwIMl4eNYxELBYEZ2waZRl0/gd2wg3hvgWzbdXGH
wOXRe4CrxLjUyGcbab4KiZi0wfpuAdwwNdkyGOK9apvopdZ2yIMW1aYtJf0g14y4hznUxPevx7M/
HbZipdMzc3YbbdBueAHi8xL4TEVa8kwQMNWmoRDC9fHzJ5c5bXwIg61/WaBTj92U8tG1YYJPSGVh
8rra9ZyhEz4HhiFFynDs7BtN2NVJyZSgDuX3P1oVqGJDBtB9+e3P1Lr9FRTr2vNU/LVWsxXma/Dg
TdP66MHDus/NEM8zKmlQrtU9lNwkR5c3eGMGe4O/MdtbhYbI+nOB27MEnDI6zjZlvr+i9eRPX9tP
nIypJMdCvvKGhKRkTZ5mtkhVkTu4/2CQ5a00mFKWGGQXs2F8+vYX+Jg9WBoXEuBtsGEJp32hzOdN
6AYMTPC8pfL8w2H0vzaRQsX4h/E3WkCpbtxyW9yjbax09LgIsTNlvUkaD1X45wCiic0NG2UOQIbv
sxLt829WmjDb+5ARN8xlUt3qNf94IAdVaJ9DI+ZYioq14PXBbk09n934oxkGAgnR7OlD/V18rhfq
ifXRt2U+cBcHThEYVVS2r1P0cgfJ7FPOv2446t8XrrN9NxVIpa3VhGOgr2GP//8kg5kLMNB22tEC
Yrk7GwV0x/LKNEomvTbnI9B3nUKyY+bV0zTlJRt3ZjPwSniozRxRdmbHcReVmBu9OWOlaxe/RBBW
7OyRdNoLbXbMOTXG6EPLdmv/CKQqi4mLuhXtARbLoMyoEPPFuSmvTAtDBsISY9Bsl/uO6+xlgui7
7tKB5TNYr+I2VqFRCzoWVvenF24zxC++N9e9a58JeLm3wINt+BFKlKNOrMaEeZqPrWFs+d/FSWTe
g0Hv+7HnyloP7CRJeTL6oU9+VTdPAYAkisFNRzyeGRYuyI8/Ad/JB84WztAYtfaFfVMyW/TqB86P
fxR1K21nJ1dWo65LzvFJuw35R74wg9PT0CIHn1R91tQbynpQCexIqKEo0Ttb6bfrxlAp4KDaaUNH
ReGM/HhErUpbEDgd81QaTlph2Q+9imAxnEBRDyJkneXNmQ+APJ3UuduNvxg3ZY6Dfd9yc6JR57BG
9adXs0beZpMemr9wp66sxTRq+/e+8/S7zzCl0YDQJRpwZmvioMqylvAkxNQnrPND6+FDivMjga99
yKSnhNCiLXBylNSCuDtOs7TTndNE2O62h81/1nB1tLUsLZxN5GZeA3mapIPk7aXKxWUS44BCfT4/
0O/dO7SxdD3iiJIrAAdpp17HVZZ2sJBVn8mhb3/PGjwXtXAiP7kiQf0Eoh0v1ACdfA3r7TLMG91W
bvYz4XCletjfRJq0Bf6zOctLQnvR/tiKV4LL6r4mD4HYuBfJoxGiL9dQS5CXwwaHLXx9UAkqJV42
p2H7Q18fwg2H7KjvkNII2RvWCG+o3P2quN3N4y4XMQsX8+sia//j2PA0/oYIsi0IeAr04tjz7EIp
eBbFtgRrsscKH/2da14rgxwVM4voikAT/RDkHkr+f1KjOF7rTTVZhdakbcXJkBsoeq0RrW4m3zyc
p40+Um65+1J2y/JSjapQxnBEBtZ20Xn/8nvkZlQHxJeayohZgXUJDkERPaXq4UUoKt4PQnofd4m0
InFAnjbA8Tl901Ve1kb6v+8b42CsBTWVBMjSTHohWA8/O4FETFRxw8U9GFAuXzhLrFXD0+A3PZzC
3M+viIioCUeTu0r6uYrevC5Jzmev8aBNWj+EDt6vi7FyoxDkjr7u1juF1nKM46TCbP084dOEjKmV
psrClZ/w431shZmN1Y9JgOfv9hL8DmMc1tApp6VLVLVfqB5QMUX7ytM8g+5/LLUKcufV+AZIqsXf
Op1s3l2K++Xi+/WIt6KNxOZxh7LX9wYLTC3Cfl0W1NsNp7kW8cFuC2r6Ud1GwCSdS7tKm4Wt4Mff
E/Afjj/m4yaB3pEwbYeWZshf+IPFTQJMnT086BjacvGd4Oo+iq70BWKiSjVuiJ/emQC7Dgoz5ZWT
LbwBTtyLXzEZVDWZ4/5hAOrnNCf0jXRu3c1E9ezKfOS2wR5bx34qdr5cOnvGG6mmqQ0ZG2WZMTBq
R+84C/oIXJ+IowZjUFMvUrOFP0RDLTpNTeNSIcdqEUnodrrmydZPMCFe6Y1jkqD9qiTw696p/qYC
QchOTGL/dT3seKyUzYPC9TRfc16knNx1PQDCYFCyFLzz4/UG+9c/VW/mWcBJHapsAW44C1AtOiD+
wpKaBAmvwQph7lDuGR3DuvJjLCFMnuliPJHaE+cFTRnkF8VuSNCth+XRTCsEftijO+tPU8yNpEz/
GLryR00DThC5t7nUtTij0f4nKsIxAu6pGueCqKiz/dh1xSu9Gc/wJpUHBOsVQhYiDae7VR8IpBkH
FWcGxxTQ0fyz5TCIQjMWcA47B7Gr4vZeceb8Jp45+vMZ/Z1KWvvgTmjcbyPbbjWh0bbSOkVc05m3
QirZb5LUt7/6ioFQW35NkIXbkOX4b4NaqVFFZ+JF+C0mGzoKS1awegF1nr+gHQNoDjrS03arseWI
ytMzkUWzEjxcUyhtWs/yhYHSNbyyre2fw2Dzcf90/n5cv0yXEzHY8y4rGNJUSZHrjn/f69Ubrjhq
Xa7zAOwIsPlPQ8DVPSEg7jBl2uo+89ZgLcxVRrMD+bGkUv3ux4VJaRyYc8AgApMcTdWZ49oQDpf/
bCyLwB7FJcFPp524cPcFIhYWbnUT8Whi3G+0vED1oQJ3uL6/VonXryD7fiIR/1+IFUFMSzdMYZqA
Rn053i84uTDk5u2PztXQ6sbC6TSF2B8q4vRto5YE4B/MdmETpXtYNLhMeKBgeX27Z3BWCzqzJ4gX
abYCfnPDoA8nbtthLoUgHLKkKESd0MMz9uS9E0OKoTDEOhAg8CLdsw49TbfJ5NM3EbLJrYgTxOeZ
JZuGSmFteaDgXhY8iRtGs4BfG2MJ7AXVmaay3H4Etr557cNpSBJmAYKd36fzJ/T9qS/SvFSmMnCI
fhcoF5fSXFfNg3kQvjhea1mA7kviEnBROJiOs8CNNWYwKpXKsyJ2AcFfQT5BeBCfowmwN9+A/IRH
qqyXTj7lg90LGmfr6GAVugNM262T87tmCs2JOkn5Oip4wboL72raRBj4Jg+ro0b+fe9t3VBUCs87
8QrlCFjWt6xL5HzXYK19OIBu4ideD5qAEuCnInsdVUHBhUZnM7yFBkz2uHQE2JSpFCbTAXO1nj/9
T3RdWI1M9/ypjiU2heocGWYaJC5C4iBXUPrTZMinXVmAVI3TxAJ4woW6KwHdO3gGejbfiODcV2Fy
YfC1QuKeqvQ1ThtWK3jymM0d8w3PswDAqQm8kQGZr95QjAkRaR57oMQQZuU83ALOil8NJSaUgXFy
RFTqNxcZO9YHyILYEdDVrQVGhSwbEBhKf558Wzu6aK5u65djF+Gj3ZEJBGzQqIQOAodZwz3iXFb7
KZeSS/oK4bOjQoKjfXix2E7NYoSyAQ4ikP1kijFFUieu3/m8Jk/xtnEJs3VCELx3Rr0TBi7ks7Us
gfWNmLkW3BmErymLZAjM3+3i/q04h/j8pDuEzmZAHl0N6Nu1OHOj/sY/5CD8P8C67Vr95rxotpOh
tuc4Gp+aVaZS3jlrDn1c+vxrynGcPTiqf+w1rZEfzT3zVkOF8DP53+Vif8lpAMnxzQvcenVf6j6T
yOul7n4UyLNA6qSSpHZvZQw5yh8wugvDubVwpm+ThtqjiS3WW0DhBJ2Z7b54dmrca+yHXLcJfX2v
LP3iBZq9iqjTPRZpj9PfR6gIU9iq6Wg3SmBDKxmc2/ZwaDWIHlVZhz1hXUa2JGtjpKxxUdacjxpO
WnoGCpezAakVN4G1YYld2gyfLwTXCyU4sp489KhQJl1+yRFNR4bbXLsy9IRrIuYi8EWR3cjTGxPB
BHTEmRB5+ihNUvKQKpKL/xIujYtWXZulD1tvTkt5IkcDX5mSl+6Q0Py/KLxM5SVDylgizLGQn5LR
AYdy7wGiussb3DsvOds4BLhrKmSCt1nrh0+N9h0Ms4c22KMCoPlb0hjthB/yROaLNevdSntp2kHH
3vQE2sz/IKilFEXWQTlQU6pKrjPjhHjlOIF3NVo/e7gNsK+H3uF6FPpVJkLd4SduFEC9EBZrEKz4
WFCkiU67wqO+BtmB/Hva0b8yQafY0EgxkwWpKogWzEg2YGe5pj22/VOdy51P1YIQcJxyvd7QEGza
ZCMX68cbU9ZHW6tkl1WB5CWWMEQA1OR1ZMnD4wW2D7LJ/bKez+HsgHlCA6pd+p0zUddKXf0mSRWy
X3IdqDwz6JO0awBUVFwQdwfCFbHOMjGeSqHJX1j9tWRWkHSC5XpD4+KVRKxexZTbPur5NEuIerGg
Fd9kW6X3vQOIPTEN3Q8V2N8jWK6n7Yoz0dJPsDIcLG4LyObI8ChzNZ0NUEkSrarikSJY6QYqlTBA
FGmfA3rRdRM2xcc9GPuYU4QwcI+snZ91uoFarw4NalVbxa+cJlaxjK6UKOt2JC2e5ya3KE0WceZQ
P3p2fhjRL4v5NEKcvKAgSdfAvXbJnnNZ5HFYnKVHbzjsqfUh8PMWuT66sJM5gfzweGQU0oT5F8ji
czrhBFlORd1p6HiuEMjySoDrt2dTrgO8ZxFErNjefYxsRLor0cmO7I9HApjD0zZAGVF4ESsXQffz
NMdmizbqlDbNqj0cnXF0dC1wxLxYsDJKgaBuxEwuYsY6D1LGYhXeHfdrPaVnfbcBWdEZgtz5k9bl
mhxegLfhc+CB0DC1pdWNbvZGi3pJoE0Mh+Fv/K77Jk9vXbmMAvHsaXO5GtRDPxZRLbZAfHeKlBaz
Gg/tS+FDdVvXTzeGfuTeLHbQxYuiAGyD4dN9hfPIwdv5BYkALtCyi4YzncUtx88HlWL00W0DTOWa
MQj93lU4bfgJdCE2msGbhM8hhcFge7fxvu006XJ3B7GMMNRaTBla4COdIq9HdRhCQHUPu24vhMDh
qmOtuDkDkkakdHSn7zOnTmSePqGxyjjRysI+ytcf7hrXVsg6vGBycE3PWhcpOBKdvqdKubi9uVc9
9I8s1CuFgLIqnGVWQqVbPpKPfz5HBobuyZZ3Ihgbs8wS6PrDdZFGsns3+FJdq0v5KVRymCGWTEXp
xfKpxSeflW12HZ3bemkFA8EsYSB7qDAE2rF77JEIHIsQr930m+pNrGXvBBRHkpz4+f1jppEJqFck
VNbUvG1lfR7fFdOniaQxQglo+ZUGwjmpD84lQa/4tzRcdSePQ8neI0bH5BZqCJJKXIv6xDoW8oSB
DGHWAhB9kLlxxetuzR95VnyMMFxdYZALkup+GosvzibooGcBcsA1fXr821WCSTozacDHIkhomdvF
/bECpXPCb2VO+3sUlDk2dp5+LDRbNBjeMFaxzHul1SBrSpZzzfXfd2Gel485HKL7Kiy4X9cRDgYN
Nv2/hr02EisuMh1xibEGx99gpPpyFmU5ZxC6j+vyKkWNU+TbfjRqb/798x8IWt36LwcY86F2OVOm
gzSoSquBCoJSrw/NFeT3H/7T4cVQFJq4/YJLn9Uw6Y+dlWXwtwAcO0+G7VpHekhYWFMK5ZarFfAR
S0vrUvN8ubpIN99oK5MXjcTmlnmrPUcpZOhSRmAhP7btNCZppKNNNXQGiUgtTSzbUq+qd6bcpbdy
GiXCh+Xq+8yGvWSnqSNI+VdTmPkQZDXVBUD9579NcGSTc5k6mR2X8MJDxuoqVzS22NgeYdkvqEc4
HlmE6PFagjsOWzV2B5hWCnHAh18jMLTe/z7MYxPHkL0Y1Vmb4XvWYIY8nUrz/17YouDSN+FdxkJ4
5NQ4OFR5MYeWaZ92W1uqXXKmdG//XiaBDtNFY366DTHSCxSb5AegtDGlzTiee/XegRoatbUKZxfB
sNuM3xTUBML8BU4oY8GBl9xhJ5FNq+RvBPwqlAgce6SiMUyvgko2puoL7MtDIRk1lEFgV7POs4y/
5Kd4a3NctcUI66ikCgqd3KIU5rsU8Lv/6I81uxqNx3iHkqUnT6EM5zMkOqAY7ZnktvkHv/8oZt2P
WZ5Ygjp6jY3R5wwaDZWstKN55I2LvjZCabWMq2zU4h/PtYdO0ophq1CuR1/pC9vDgEimbFDJp9sQ
YbWV00MGf9kByV+y4K7Q2ZL6iBRvzAfvhnQk0+1UPK1YqA5T7Cl4tbwcCy18ibyODaDdmT1n+Mdm
LJyhb7bzJcwKaKnYJT7bhLbYAPpxwCK1I2HPkRHeiAK43qLrSwJqaGg7/ZIoEvzS43G+CtFh6N7c
BPs3iycdHliSJS/uLDMF++SjpL5Rr5noCilarORpqiLho7x2Vq7AAehvl2KeLdlfkd84RzQgyC0Y
8bZ7Lo6E3OKZwGB8B3EhE4cP+N4mDWW9MXwP020YX4PUPGMCjTYcpU2k7XI5vNnFqGR+3jVwLbeP
PYYdIieknDhcaQpexXD7nvP8puazPRy2UL7dnMJRRzclk69+sLx+HqSc2Bc3cLCDncRxY5xmfjAI
wQy+DyeD6VSYdS6e0WhzSBnP+tgObpLRlDRDKorwQl46meuxXr/zQnI/mnhaAHwqbqHIeJvasGvJ
gEU0lHi4TgzYWaaqJU6MnFEVmmIfA3+MHrt4Y/5rEa6A8ykgSo0IiW0GL4634Y2e1WIP5lykI7ZL
OzXzldwzrePrA/nHEbS0SZg/+tqk6VGwSuu8M8pYSe9fFEyTdKORDueG/Kvlkd3FNSvgavB7lWiH
3EoRlKmENxgS7zhwA4qDHcZuchViyBflDNCXdCtkYpynyJ+CeRh2oqGZCnHJvadZLJMjekVUXXDQ
YvwLZuqqOOfzLuyUnTdk3vxsqxXoa05Fn/CxMHh5WYA6XkWsOQ7JfxdcXrKn7XiTQTgKVveMuUEg
9HkItQ1SCETt33hbGrggCdQNvivJ/l2kcM+7VzkKNGHN2xgYVwr3m0D9hGGe1xSxNkxjA6SXSk6+
WCAmPmEdWt0Zk63Twbj3lVI1E+iZosQQWZXCfB+YqBbvtsAMjSFtQhGBC2idbVe9mk8RedRyM8PW
ZXUqi7QTzh3EFKkLWk3r2xT49dKn19wIqv9Z6mb6MPIApGGTNmhXb951nLHE+xMLAHmuz2wbEDhb
Dh7ZkgVKRyln63IfeJv1VHN61dmpE+Mb6yo4C80GsU1sHP8KzWblEmOXo+hgulrZ71gbYIWO9T0E
VwnEgs7adPTsv5V7XmFY3/6Hg/P8Y3VB7GpHp6GSXvLP9OgXg3mULj9OKYvJnBhbqWLgYhcZByDA
CO1sWFR+opxUtxp6K+L6IGW+1YNsnTFQ2p475DUPNc6BErCODn0vbJ2jP208lMP3t9MivFUVqFpS
EKBi2bD0VhzyNuqRr8OHJJDd56QvYpzZnFsJSyY1kf8v4axzt02dHmbDcs/RIlMJzS5mfBGOG2BR
JNxmTEht3hieBRjXL9+V0LmgixxugF6oPas24FZZGXN8UCpe20iYlBr7H2HFAkr0ol/NcUPI4k1C
tUipcXfQg99bIBL8QgU5V+pqHvhYTIXCXPkncKoBFuk+NxTB59fK+HS3Zs/eMpn+WvFAls8rCFGV
foVFXpySZbTGKYSTGJVclAq6ui+1OUvvSy6Vwcrm3UXdDbfnOsBg5GGTEsSOzWe41PKIsbikZf+9
fLG/gUGtG80pszKa4jG2vRdmW5vFYvl9ny63yfrewzrJmjwrffOPIjO/J7sa3Rb4e/oPQzbOpZXK
Div3neDlZOckkUTXfRPyMbLkfbXRPjsPQQiT8K1OXKE2w3h08GScpdg/XdfXj4auQtFMEP82UChH
DtEx8pGuo1ZWeXERS0HdMsPuul2bu6UaoxVE7GtdlYunjCOCBcRtnexGu8sE+ZmakeaJ2MbrfmlT
7o0pI3cmGpCUa6ZCpW3iFD/n7KPnaXC4XhvzUbQj4RhzSQ4zgMsav1d9F8hEsuSjxL1onmGaxyif
qayLXsSuTgNKFWeD6WFFS/DU2trUQs36Tqi5JP3XEMPRr0Al5Fm9jd3b6H0n2wc7DDew1tinkkfx
/Dz+YAFgZ/lPGvF7FdNKqJPd7Kjx6Y5Ffz1ZiRRF5aZU5x9Yu9Y0TgbT4aHhlTHTbvohd9+m5pZf
aoxEInw1Yuds+/kPSz2FTiw55j34H3zKt7OXpn6wiG4acDKJPXuhQUdlq/X10za1PF8j8emvrU7e
9QwfQ0ivj6saqUliXCb1qda6sI38QVXINXgvpCKOo3Dj/pimaGMqZUMAZnIWu3WmJRoPcPOspwSJ
slPGlLRKn94sJOA9GmC69oI8XPDQS4iySvIN42N16XUzxzpWpgiaalt5JKCdwXvT34OxuOS/bFyt
KlNsbeOWPLJu35AACc0iYu2esJWefe/I7k1HbdeJkoMcNGKiWwbbuW1XIuzbr6JCaf6xiwdrsBjQ
SXogZ7EVBfbehCV22P/yJzZBcNu2s2QGTnnzPSEc3vTLZaWaK/EK2+p8flFjjmlLWFR2/uYUM8Qv
qodUVRhjcs10UKuvefoj9L9dhqcGsJQGbyzB+QQl+4Aerh0CBPiQoOVO/0wzrUgIzNjrQ/Iy4zGW
QeGkM5ER0RwcX+YxBHpLv879XQhjT8ctQWZUsZwm1ZB63thWNAxlz86of05EpLuSelum00UFePCv
hu9BgxgHHI93n9Nr3Oqg6zVmAhRAwkAyAPm3iPy8Jvy+hz5/sWOTlSoM/mjlAjV8NCGVBWmE8zYq
io3mTMi6FFcP8L/ENeaFuCF2H+bneE6/1hqo/dKd5+1faM0EQeHzNYM2HN09waE8oOO54a1sNvBK
QBE0DnHrOPEBA+fPu5/FDz54jNUtOokauUwu6R61GxPx4edHYFwaUnSxHPBKKudTctWT9DWi+hEL
dZNKBmmphS9jENdt85FqxjDl9NmoZ7HIXZjboRc21WRxmsEK60mjGgxOTgHPxdDxubg9XI6oNpcH
5SJ60kTEEEQWu94lLD3czpjLpA0shn0d4BG7l1Pdch/3GvmSBPM669CZJrrr4oKxM99O0wavZ09/
so5A+mH6Q1XZUu5Kh447H/XqcQ+LbMcuC4NuF8xrYxzg/vYvFdO0LwxsySPGBoStphBYd8EAZJtI
To4N6dYCWqvtEbIi2KOuDUkSq/0qK6HXeQmDk81G3RJc5f99YQY5m3K+QCha/mKAoNfVzHGygtU1
IEbWS4Kqb73DPuL4VR4w9HeOkyk8ENuVKDC/HKs2W8OgJKathJ9bow++kaVYPRsztu1jk/9MadvB
xxtTFYphsLzSibQqO4bm9cvGDsi3/lzwHyfeizmDidjCmiChLs6Fn8FuB9q2dvV2FONFI3nRZooK
iLlAacPx5LhssJJXfm1NdQw9EdJj/c3dYsakaWtWLqZk/KymvNu8fToMv8BBeh6YMFlIV0tRsqdS
AdvQVOmRZpBCY55SpAWNiuwXz2HUGWCYeJhHcbxwiBlqoqKMripnBlvU3aQ6vLC2faUYiCFnDrEm
uv5wbhAnqsEt2UTlt1TxNPrqBTpdIUrB2yrImTb4RdQUrKnBoDXroZ46DFfaVTK1dZL2DmtP54jf
pPHU1J01Ic/ory/q5mZezAx+dYkUazu8Yb9sQVLy1qbDeg81b3/UAL8fJCx9rnPi6Caq+L9J5bns
3xDv8oJuG9l0+NypZPHH+LT1Wl1Q9IlptM6f3af6DX/nwKJXfKzsL/UNNi1whmEpR012wqvSuMYX
abT18dcbLaF1twD/SrYOSkhVqT6X9v7Ord4CSeNtgPiU4n8G2O3C8KSYh42AouFMrupxPkzwCDtf
bHCeBJ66wKZWZqYhfnEmfLNafc7KwqgFw6WkSMYU71NLKs/TMNdCeLU/+VxWZiLma2KtZA2LsiAT
eH0/gQ/lEYpxIgQpor/026yXBBHCmgh8Unida4fdb9B6apRQEP7ajydPsmZ4THs6ZNlS48uviRXB
yIishSiVzzsF3Y/FGIkmcHGJYwXgNSeyh9v5g2K8i0AQkmQNdc2/aSB5vzZ7zxzzihskqHwoDall
oIaxPgMi6scJ1Rv8LL0aVgJ7Odtc6UR2FpHiLrbexG5JTHCjFrTanSLiY2GKs+XQDBjfICLTsl6a
4drRsPUkJ8J6/c/kMxy2Plw9ATNTuh0x9u01ISdJcfBjYdR8jNELeguhx5F04/bEMq8tGwYZ2i3e
8k/6V3X7nNOPu9fZgRTLiVE9tHOQBwZa7kHVusTDrRqKL39fMeGyzfuBjQ8OrYPjxj5+4J1iJakT
baz0FCNMjElbe9edN9DyDFSxLUoGUUbIW0Jy+EBQ1BRH+VSKG53STlNe9qDvk0JI8uJQ8N3E4al9
Ye8l3OwWffPS4NYitnq2RsUcZja4fAZmAjhaIsGUK9GGM+Z+9oN73BiGrHhY0ZvgwXaVrhevDM7s
4gBSLQtT2G/BmErbNRSZzR8or7lMjVNZ1yO9wbXX7odqf9bwVci5kdy9h5CBHJievHjRbyk8bO5A
CgLY8fRiD/A+372epNi2lWF8nHAADKSR8+4pG9CU85jhrALc2Qh3+sUUQd7bTP6nXRFRsFF4wUbh
bfeATCsQSOWcoaO7cb6irbbKzBr+6WunwdC+yhob2kCh+TDBuBPVcOO2gcaXQnAMtBp1o+6uf53V
ZL0HC2a3T/xrDDovkEPLvMYiIdiCf55EEFxHyzCq9w1EC84hLZKAQLfZ/r2gEkQ0jOUieJ1j3nlj
s9MHdoqczqtvZPyiCuIxTI2aw4uTj/QUBel0RNzO7KjSbmP+v6GRQp5yG0V0rw2y6sU2lainNnn6
w+cyrCCQWduoksBJc/c3LuqE5U6vgqKt5DY9Ws0Kvc3SezVgrLJS3pFETFPhpqTT7vCoUSk7rzLg
9T1I+PepL/eOmzlgnLUe9DGAVptWJsFlnqY12A/628wwmms/w307lY1A76/mEo8C5ygUwpVFuryx
loLeMH2LHFkjwAYAO6PjZPKOjuUU8jmYYw34vTFbf/yS4xsy2RgL+vJHAF9XWMlszDNFdfqTPrL2
251IVdUgjbU/6ASgWDGhPB1iRH2CGg7teFJ65/LeGX4Mqj+ywcSbuhbm5bcaU3LKnHQpG69atGIM
iSqxh3uVHkq+J+8V5yoyJvhOlnTws03IZT3UIBiOzzLQkX4T4daVT6/usmTuNEu0dJzx0Z1hRHwg
G6RpaCXwsUybbwpRjWis9cglgul/Fus7HntEJzaOmlnFYyuGzlfl53wup9c0DWFxWXKluB/R1Syu
LAf5jGckW9SSc9/nOACiOjhNc0uyJd3jRiHkqN9pXp3P8N8yDIL50O6AEjrct/jUYPH/srufbvUP
gp6WvdZdVZVzdA7iCWq01guca2EeHFIkCPp8e/R5lheDlziGjM+tqFz5Kn4XyLPaZHABGx/XkF6Z
dk/XphpYqjYP6Vvy9vdhzRak7Q4Ttqu9hdD0t6GMC1H4c1KEDrYT/I4e/wpVknBrXeHjCKJLtdia
9U1FFBrGMWZEr4B6FmzjPV6MlxAyWZNFq0msEV9GWRilF27NYnCQsyrDU9exyvUpoMt3pvaClqu7
CYitTXbPMt3CtdBAM9rgdeUIHbgU1xSCZdsrLBdBs68wwtiyUgtEU46WGWW8jfhGmJUJjjsv2swp
w1ntdkNXMYRP9UrRpbyjd8bbt0jw+ihktoT5s08keyJVimGTuBaafB4+ScULlOtgoVjX7fsyQOgh
6tjs1XlN4xipSJK2tWRyO8OCEfeVkg3uGUkT6X0VRQtuKjEC/gMz80cnbw0QkSm6vHEMGClDsFGf
pV02jd6Taw08lqFBqgwExd8gyeGHGP8y/FAtbzl0L81zWWciS2dRqLkkPsghX5PJJyhOJ9S9LPN0
7MThd72qPJojlkvE7WrZnvQubc/FEn6q86Uhb8x47LG4E5Vls6BkGB6aOkrdu9lppgAkOgnWur1b
0IuV6cY3P6GoAyctzgklv03VakBx9s7jEf8k+BvkUst03p5Zws/XnABz3zl45BqZuUxbT9Rxboyg
RwuO8/bXF2hYhj51WcF7136bbOLVHhsdySCPDDEC5JpCzBbpkVaQrRYefgm0bmHflKZGvD8S0/vS
I2UUpMcWnh2clmvRWZGdPCz9RERJvoBVqlc8f5NNJMpZBYyyBA59MD5j0f33HclBisOIk9SVLaRr
uMGI4Ygy+xjtam3EAA4k5Vm58DDd+bmfxbaJrFif80QZx2227SpI//nFLPX6YgKxLUjbQAyhGiY3
ZYAxLX+s5S6hxCvwgdn2vbEnEPw9yxH4Erhv1BeqtWKa32tq8SV3F6ZPAXnxN/iyLIUyXEP/6f24
tC+b56XhuhkR4/h1Dx3V/AIGJhIqrfjggORVZg9Rs1NfZ/IuhLDXjSCgxiIHjisgN4p5FljQLBvT
VaJsgMEoFSf/67Q9GQ7wAKdbiUK47lX83ZbJkuK0Pz9V/pT0YXey1VNBN5y149hn3TL+OSwEHEIb
fKnn9nRrsf2hYJj0OFftfWgFXsQzfaXxcbU5DaGbl6pLH+IQqr4I29fhKGxdzsyTDU/w0Vc7Rvmk
qwGt5pQ7/HH4P5+h7TdAuuE8ckQxsBbcXENHYs+7L/1oRsA/HhzULE3oLbvD8sDX4ZnCFQynmYAo
7ekIjg4+Q+ZW6Py7WQvAku/XzvAfhdaDULSGtzOOKCKaWEdYcbgxvGimsy/O1a6PqpTDNYx1Y7Ta
RhOq56W4DfhxoESASHIh1cR64UL+vSLXvTfv53IloMwKmLNnoVN/29HoZyo0Ki1pCwrdd0JoXrxX
+CDSmgBfsbysParrg7/IkUPJfu4wi7pUcCHRYlFqd5fWFgptRsI6miBiArZdHPdEaVc/rQBKGfvD
JcUGECl8uVR2m/fAStRhqpmlfCJNdjEwJLojGDO/utHBO/0Acb2EDRJ8/xml/+U1cbO+K5F4rzFQ
X1MNBbNrvuXHmQ50A6xZcSHL4aFJs5/IW04FhMRc5E0srvet2U4adMntw5zEqojbrBrfi8WEIhwc
kD7xEOSVbWy+aj1hRP+1LWOK2Yyby3nlhfY3WtFPmaUn2KfoXVcYztmKjg3u3hKjlvKUXNSQcg5I
07ECHREAQrbF5Df5ukYFkgf32o422mafsGnamQ2a5cLIfFN8JJwQuMqCb6ZvkIwjr6p0heh8oy07
ph6kPiE1Ygx9ijiK7dH+44cPPKwEMp+CVWK5QWAFhb1IFrj2iny82+hVHDo/d4XkHWnAeta1cz8w
Zcc+gWt/JvdZfv+oCjL60yt/0PWkJ0VIyUusdpddGEnc8msVLjd6cOiCaV4n2z11/jPmlEMLLyWs
hxAS/ZCLOpbuPctakL/PTj58H9utqVJOaEs3cmLF1lzD2kZi9bVndgj6gVWQ6YXx/CNfPd0f22HO
CvumyiDI2wb5tGH26dkSs8G0wCeobaudJTc6TomJC6ZUxGbZz7ARBDjve6vEVwWNbGVe+hjJ7yBa
/TGWx2W2PFEDAsdOvhQ266jJ2NdmBqjGMB6uV+CplKvLO/eQqMhqC9qUZf4oYN3KeYg/+WMwA2do
nN3rzQu7QA05EbBVykZdD8QaecRTsEFIV21hJ8Zvv2tkM/RPgxq84ZUy6sd9AOFIehTv/6uOCSpA
5YEMPvfdePyFSempUtjr29XwW+ycNJXFmrU7lFWlPvkoD564cK7U7hMtCBNaPOipHIuIThtESP/y
LGSd/KE1qPpvGsvD4xHo8ZSgkgQ5AgC46/24hBPK8qAB2BwBGB+AIrRmjicGKekueoUCrejTq/R6
WqRqSpyjEcVizqiiMYsDg0QkPgozgXcoA1DxC+z87x9FMVCaUKMh65MRpTb4CM1/exVtLgZBS6DF
JTdI5KhsvLKHAj4Ubs0T+Dwt6+3wB8gXANweOXL5XHV3jVFntm9q0sAG7+FLm/0/nMe8HlNVteH0
mUC+A8ELX3Qh4LhUCmuBBV1xMFIfdbuAoAh6LYj/SMbwbMvD+h12A1ol5G/aA6w/y3Rsu+zOuZya
/eEBVfVgINr4nhuUZ+GjXiUoEakUpYW3ejXyjd9vWiq3+CG7JYlIt5nF1pS0kUSRo2FbH5PuosHp
9Rh3k5zUlAWh8HnOEjcVbFLqem4dCxP61rFHtwevo7xV6EjzuSSzRj6uBV/Vk9BUQ1/NkIwm5c7V
iYk6d/HD30iz1qFZfhjDqqn2+uUDzUwGhdqB27c004obxWXhR5bnmXHQ9bmXzA2c/TC8md+/Zi/M
/aEEl+UWTWqJFwE0vWofYHM6GkXNJd7i2cylJ0t0dCLxZltW78AsztIbn+ug50inLQ3PEyeAUHa1
pHYKt4RjBFhGjDrHzXCLqeh2g20LPZdTAmxwYoMiAkyQyhdmp3RrnDW3Sy1DDXfYWIL4I/GiC7B9
3b6tzsIbocR4I+dBLBGRHav1wLtVD4mPwGwS18YXajqIxqEpe0bss6u+ajSBTQfaK6ykZAn9Ycc3
mKbc5aZUSLwMjZUEn1cIcjxawzsRFgV3I0hp4AptXUYKobJSP3rh6qrkvFQoNP5HJOPVDF6GS7/0
2tyqQldK3coxWS1jLKE1XfdVdxf3HJS8KbUYyoJJ7s+eKnbtPqunK/pD+9lkmnGzkOqZQj07TxYX
tzRxJfgGSVW1IETlQcbzcTQASgk8Nm75fLe4hjC+JKv/ZmZHRC+HyUbAWuqmrHvebKxBG6/n5MO5
WlIxA/493IEOQ6HMuLe1Y3JPvt3rEV766KIsch7faGDdesvZjTwEarNp/5IRpGmS9pgwnZOtYPVX
YjOBiz4wttMdIqtkpnzGWvIwDBLAms9lA7z4dqAE9ybgiydhRRKWXzBJYIytBKrlVtgYyivmsIkE
JTS8tdbRRC6si05t1B2tz8LSSdzJF/lCkRCRFLZmfPzwvT6NqqDUzzqpwJh0fJPFwPtoMTYV3dH7
qT/jB8re2CEyewdjE3kuCjR4eSiZ7ozPQDGRnzK/fjQHrsXcqH625q3C6RvWVj9Nc+DYAXHenJA+
ZriQSTMOt3iF/VQJ3DhdAmKSSiKsixV5qyfUN0vm6W/v5P/J0wLc8fdEeYm5Xcn6cMMnAN//WvdF
kXpct5d8OeiGDH9wkyBxYvOcG2UmayaEXCq1R6r2I1BuatJqKrqJQvamMvv9VaqUbgJh0J/LgmOD
4/OVpZxzAubBUbq8sEjET7EnYudP2wx+h9+gtNfK5x2GGo7K12bNTeRc5UHNOstVN+z3tsuRL9p0
drk4nwdDWYD5PgHJY/h6/IPS27KLrsRHl2B++BCRONebMHFTac5v1oJVZpE3cR/4dHy00cPSWnip
vpNTJq1NyICMYImuolRuKUuKKQ9PWFpEW6JGw44X+HDzt1it6vNfxr0yOhdlOEjFnUZYMjPFbhwT
pgrrWbVEh7Hk28650l8bBBa2+oGYrA8Pb8bZJjomWVq2hrSHbFhAQi9aqvrjH90GpcunN8calp/w
sy55fasAJjTz6Ekv0bTyUDR++SJldtuObiI2fMLAbB3p4asLWctim284v5LvgEuNud/KogFxaM7k
GigXauQE4RECTYbLoepKeNyTnJBH2BLn0+LL9WF+TAZpp37uBQNCvghdwjslwDTEbOgg89mBt+xl
oM8rVkWCyaeSdsIk60owdOIqHjk+lE2sI69ksYXYfc4HQdjpA93rpjd7QHdoxNkREJ84EEuxtl+p
W0C2I7fzkrCBis2JXj5DSldWelr8n3hl6XSZBRWCf4eQ/CF9u9quPYGh8jx60etWruGgWy6vz6mT
I8iH/50nT7CKn7vG6meUSbEKsJeRLJ418zXr1hOLBRDoCXfmkFxM+Qki+hSEAU3KQl22CfSrgIpj
h+MRYiQ1GLVCdFOn5ka+06BmqBIDA9Zm1NCcnU3siX8b26m0wx0M71+PyfdXDpnBekoX3c/9vg1G
++Apxp0DEefH8AQ6ZGPHAinPk7BeKTTlqVBr+mmj6Nut4vhj/62ZGshnuUYVBKfhpBW1KKsK3V4P
GUkPyDa5RRHr3RGOJaV/zSVPCDoqqXr7YibWL9OjmIoqerOR6eY/q1bl34PoyRB8NjTWCOm/SDYn
5MGXlmOti6JtUec1+2FxgX+bfoglvM1Swp+Lx6I2nmgOd3+S9c0OCGbsKZl4ZtzHzELJVM+eHqoU
58L8AZubAq5tUwoFMDLrH5iqYDhG0zClZaO2yR56zvqByiZ5P6t8OtdhDG4mBX70BcJmsN4F6lae
/nhK6gZWJ89sdmtRmrCbyn4/NlcTPLFE5plS1oASw+5gFDGFjWJ4t+wCkYxGCNhJCG+V7O6gOv93
W9WBgmQ5PQ4AiKO2PemfOrtHC6T54wTM+Ehhdh3TDWXIW56GxGtfqjoJQh5vcqd+8XdzC6z9a0JQ
GW+vuv+jOi6cmf0m8FQTKDyKpl/RIXAwhOWZnp7/4MUbQ781WaLcgkmOQngaDtA6eR0vgAxPBExi
6Acsds4F/5AKvDiCApbXGEFIVZWizxw5PmUwOZMT2Nq/Jgt+VkCV0Jt1XlCIffRgdP43hm1cEucm
+X47j4nnYOiWciFq011tPiWsBlfjKrgcIQecmdRb7RKIpSbJKv8Fvgd33/OjoMp3R80K4DZaFpPH
WiUQTLT/SOlWmtOTvt6s+iWnSXQ/lQLj7nprSUEJjEVz+lM9XzQ5ht9hWK2G6pAc9FoV8YpLy5C7
aF9FOUa9feGfq8FS6amvJqsvaWpwSmzmFAW9CeZR5LVLgJ46pD1ReJ/lGm7osQpUwfOx0IgIYu46
l+IPpyZK65/R7oicTraZF/m+SFNWyQQGqbi4zqvHf0i4qjNmSb06BLwVBxquSm3o2hXovMppuV2l
Dz9N4qVnvJQp22ILEcxvQI1jVY2BJSokfqJx9Iku44JvTmx2MUOZgkDtASxGU6/ORej2gvVY+SIf
qGjkUaHGex2O+iTnYkWrRzgm28psuN/7IfL0kiOcaO/74UP337UlgJQbtWbBS7UiPtHRph6Ya72C
QqWMzYFpdJDwzB7zO5Z9hK5Br11YXlKBpTv8JzCs2wfV0Kq5ct916G0b6KgQllJ8xmG0tYwssCi8
3tMQs5JwQcypuyHFUL0Ga1TeDccWlG4qs3gWSiiHC/yqTdC4KW8y9S0jWi7AEXI+mk+ifH9PCVPp
L1Dnz/4/0fEhAFms0GAYeggeqB2PL+yNW2i5IPteQlEMwNSGXltlLJVIP2iZlB07X+evq46DdMTx
SNmrqdwZXjrPfECAL7oL/arkZtpTYVLfOjyljQ85WuY+hYjgqDh2TmMs53A0AV3Cj+n0c5hWKpvY
oC3omyoMZL1sE1LLWSktfCrKcUjRUssGyJvbcIp9rLhrVfRAoTm/4LoU9eNIeDmNT3OLbDPePSoT
upaqxNjcC+XlM4xOPNZt8HNI5wBUgHe3LuXNE4reBC5Vrjc8yKAb+xLwzhXfgPYfr4ZjAS7NC5OB
rby2BFh3TRcjQ/gI9mz3Gzbip+UPIQ/5zRo3digEbqNV5TqFBmk+0l3mWYO5zHTA2+TKETrra7ma
jZGqaQgEp/TisqD1dp3iuLnzGx8s2YvSK3wQD8cxqdjNgmnMTb3Xj54bXBcfl3aT9mq7HpGFxuJS
JRN8tzi2tL2DLm5qyav0Q2E8mYaCKV4IAiTSHsRHFdKNfyVJpkViPrv0U1Bny/uylItPun2JmmVy
R54xxJ3e43Yz2bHOKVxdEVtxydZml5v0yMLegXioVed8MNKLCjrVm5nNS9bojyuz7TCOmFEVjgGy
Qq0k3qx4YF3ZyA6SlY1nlnAl+xm6/6oJrmQlf0aJ68P75n68GBD+8HesVy88rphLk75e/SYbeA7K
D49Xey294ay7LGssVASC8hwPvpGonvJ0Q/hhxhhVDaghiidZigR3ikok4NvaDysROAoVLqFMXU5u
HFW4QZBRkPXxIEF5HaZfyHPud+xw4N+Sjxy6TTEKcHVJtAJbQ/x8DnIfMIA2CguP3IOs/GuOQtfy
j93EtLySoExQq2g/5x8gEO1p/ELg+HV/8NtshTZInTecL8irsy9Tm7jRFUENUHOO6+xEkNxkrL8F
x7R2aDfkieUyfeEKnHJocsdf3aovRu1BTf2eF+ubcoMkJs9KvOpa8h/ncnjyBSR63eQXQ0rrNVb4
h66AwqFMS9+25eKnghsonbz3XUSseuP1dI5OS+/HpLDGChGELJi+XEIy0yfryYmAHLmzKu79aMX+
3mj31JpKqXSiptOszy24XqNFV6BqjeGRgjTh7Ap9zoj1FBNZ/VANbF/yvUMmamlNdRgTO0rCKbU7
i7DBR2dwgEhIo2J/pdzWXt9QRkYP7HE7OW9eazLiQs8caUJbpfUUWsyF2HTfk7g2VW2u+swT6djQ
RGudTcjTbgeqFvdS8+oEQN62pkmqMfUYgGMczbCc3q2m4SRCVGtLMnuaTIcaewNi+C8wZCXmqnWB
qq6AzD9YGutWhdu0jkv/ZP6iJQAidQpboNpNWA8ttz94Tu67Lci7Sl44VJujqOGWaN70o39/q2/e
6TcggVWD+Ep+oTMGSF4OMsuG2O44y/DF2NF2glqAu2NAuX03LoAWUs8CY1lyIhpwP+2DSCg+ria/
VmbbdAu4fVDVdXmEEH2ehONUPTeQbDEFQsa5e/rJ1/Z8SA3LnA2s0e8VmjR7c6AMqzbC5LWnphs3
GQG/9++8dNKuAP0F7j4dC/MphyupV1Cu2L7oPs/QDgHCPOf9HfoA4pxzCxj3+4guSQj3lQ0vnEsm
9cnkc77PXTQikd9LYggPQH1SxCy/VWFptKweOOC7vpsyFxLlnPv42qi7XgWdIbwQxyNfBnAkyDwr
fEDZyv0/719fai8dlVbUZ3Opw3TozAbTGO6oniSbyC6JRg7ozwSoSbXXMlsEA1D0WLdpjeiSbBWQ
5Y1uyw1Mavwh+ZHWpQQN0Q5fi5LdZxelTW0ddgcnQv4+QoaDAvEZ6lw3R+pHpFF6ATDbmnD/JnhS
soMmkkRv2+LBzvjwtbFe/FFjvDcZoi+h8Pn0TkEy6RuHjO7VIVIUnE76BwzBphQYfn++ywqxF+qo
huhmMa9+NedZX/GdS58OJvE2exDY54YKIVkD2Hdx1sPO2WYuKJ/+HxLOuo2pmgBEkU1bsZTrX/hd
WJviXjEgxQZns+HMaFLU8ze38/t9m1fTzIQoZDcW5ORmqlZzv55EAbMNJFMDxSeBmd1gkfuyyLEb
0yoGfVQRrHmPutGFAJyn9nxvVTX2RPgeKGrsZa21S2cpgVbb6Z5fogVphUv63BM8rffUNp5c2WVq
7JDES4BBK+SxJeIKInfJqeUc1QJpTU8ZTi1u9igKVmPE79RYQxkcTxjeOY0oAiKsV3qxqghxWEcQ
Nu94ZSZT+8EJRm5e1L+9dx0kX/hT37PkAThT/UMYMtzW9ILzXV762jlEXcheDWPuYyLl7DrZLB5o
wTgrAjOPlYiZ5wo64M9ySD/cMYZDatw3nHjem9sEmZVwBbqJmVn2LdvaL/VHPRi7wSD8qAZdUERU
hlu4IBr3rJX6woONxrm7l4M5Lc+P8JpiGo3nxfLcPyKk+0R0co3nSnkQK4XombyI4iCAdQd0/Zau
RMblqVNbHA64eSzpgdi5KcUROFehHrP+DrSjc2Uq8wrjtneHlAvrZUZQDLnEI3Olmfa5jJwqadHn
vwrTIi556iuLoKV00DJjYYJ8mQozwU+YPseqKMvrQjivlTTDKW4PRbZVReuSevfs82CzpYXyccKU
K5MlftfV99mu45vQ/qotWOoU6Q3+3744SlT7DvfKHAbJoIZi3FbyPqRMYuSeecBM9IYXp2Ln0IaL
wsw59Vtprcdl22/tdIsp44NegQYx96WU9EP5eOOMqPsErbTo0U+Tcs0yEW9lxysrBo6Uz2Q2dhUU
3r76iU1SX++NcOEivW3+v/KB08rrKBmTiggpeC67qd4EAyOK9kvfriyAs1T4DL4xIDAfUMJZlrET
M7FbUhRM3vAsbNnZj724V0cxGNgxXG3/RUzf28bPzGHGVjSb5zGZ1AD6VHs+YdNoc+faHRPkPH6i
u2KG+/BQHLU8aOZV9z5hI/eK6TJ64dtz3IHsdvfVbYRrgGFHd0l4SWyTBtIS51XAOb8Bns5bsKK3
K7KC/CdPn1MG7D6I4ITs9vmh+HTh8gq/TPWucqRMLD/zezZp9uM/gF3+gt8s425HfB+bkgy48FPo
9fz3weN9NpmYaPx+8FKaQMIXbQ6TIl612RxYJQdCGvWN0yygGZCTPse17BpyBbx9hzfVujR019xs
qFiCPe8ibnOsAt2rjPKg0eqjSo9/4ZiAkOdrqI5wuAToO+fdC1S2vwiYPTx9qsQlfDTjBhSK6PuQ
rjAGiNikK9++TwwDjHR4p9o/24kcmr6LVZz2wbjsWFq5aeXpJ+jUdynha8lpduuO2vHiGeTvqvRh
8NXP3gPJraj4tJqkLccffcbcJ83fS3/yqGFa4nmgZD1MJfQLVAKLG/S+qRco91wc0gDxI/I8AnDe
U6F++Ni8Gd5x6C20Q/8bDnRP3WcvfVxLUQIQJySmqlbtt4E17VCayDE1cnCqfCmetgySuiG01h5t
Ou+H75LYo9BUQuUH1ow7oUkIjC9m4/ihbHDkYXOZomgyBaMT4kIkBsMr5GZDssJW9z8natZ3MviW
RmgE+thkjv4hOzgxtCn/LBoqlKMO6VwBmzRp+6fIIHrJrnnY7kDa4McIUGv+mieymj52RK7ctp58
701yoswe0lCdQ/vgT6obtVSDnVbybTHv5SH1grWKR8LmZz7V1UsSKZtT9ETxTgPyQlt6VmkTelys
s1pSWa660+rAwLZBiQmhIoFfsjb4QFdu8J3lS+sX0j5U0ztrqwvoN5/YAr7OsO1WQyn/dQvGSgIl
YaMjNCC49a8/4PiUpKX2d0vezEm51mrKmaN1LXnZM3OnbQ9DJWWWzD41Ini8A9dm2K752M6lkRGV
aVFr9ZeI4snDwuVCdo4qiImeeyo6NpuCETc1BWSzTms+VcVwanJCYQj+DT7IRkpNfZebMB5s7g9e
6D6YkRytVYK5bR/MyT10wmelbBPa9Y3wlfLj6LVjdKq2gu7vFkpS29fxKuzcjhJ98Cf8ir2gdNqs
Zw0BSRRnqZAp0eqHpnSxjyIeIpg41pl88kAR6LApjx8hqeTz1NTpwdpw0KszT5qTMGm9dzR/vio5
dYMdTtaWIO6mAzI0ICThkRRXSDNBh9l01pBD+TBjhN5HxhDNjkSCSq0MPAn3M89dBeYkA0RD2mqU
7qpL1suQSLwLYT1mMLnx0SQUxKregRcWNMrEacA8dYzV6schEVhjQbE6RukEa+BWDZ2xzVlekKKq
sOLbRPt5VB9TT+IuukVN8s7jlLX16yvAD55l4YuqGQtvtfPjADNY2eniepQHDLl+HOSo9d4y5kgo
jMcBtj3/VeeLmRs+jTK3ZZP+lmtQp6noSwDJRM3STaVVgeCmpgKhgrCYylmjeM8So7ZNOQZKiV6o
QYPlS3msvF/67VbFzWTqxeD/OX5nHfSPN+5yThn3ucDqGRgfsyxQZgsQ1OX4//F5P5eZg+kmLntW
zwEcHWGYr0eYCGCuZdjW37wRUvRuYxuOvsfaynaK4T9sbQ5gUKR1BOL5rdA92YEvLeB9z6MCfQB8
UrlRCassygyYefbqq6Jegb/jdgKu1e1VrvzItSS3oOKAxIClQCMqD/2tNJOtizZnbAAK0sAYA2fi
Fwthx3U4DnCVghjvDJg71n15RGiizDR0NsD8Vog0fsccVh62e/kZgyCKu6Se3Qxc4usR4ewjWJ31
qDDLjVfet9Tp2c36ppQu3yLb94BX74Sr1d1wuyEzRg4DYZDS7axpB6jjezyLdSZy/4yRt9ziIW5Y
J0XAY/JDvHblE65PNpDVXZxcrmG/HLF2tMGQmS699q5hRYkwfF8UySfh1kb2+Fbo+6Z5HWtsfzmj
WCTYoADJtp5BVaz+syhKPDCXRUm55X4VeIab+LXvUMX/pqX8YAwwWYS+YvDf1xihxeiJBIgyXICA
yjC+MKWNhnA6XTsL0krFno/D23mBCifzVPy9zPdgw3usCJCHjhLdcAj9UEPsUTBKdn1gdcnWhLoo
fNI9A9ObE6Gbvz+jumsNFyJ3UmAxIIPQeYFjTNwH17bgzI9PFinc240/C2wd7FAFKcDUcM5dQ9Ha
Zg2OslbaB4xYRqlfp6nGM0QcMmtz0GZ7Xj237ZVB/mW3RBZrW6VtDN7cVTgNiWh0/3o2Kf/diD5k
J2HOhuaD113ZlinSSJxYBlJbAbqxnuGVa7V/vddnmgTbe9Iopg82CpgcEfaoTK/Ybdcz24EYD9Ds
XYEVWRVpT4tkT1jGbqCniW323GxBky/gfSYqy3TpsXizrqxxHCAWoncUXN8IYb3B72gxJnYol6rO
dzxobbVBtcGKQBmyCs6amFuarY3lFVUrwIxHHrRHo2MD6NRDwZzYe4Ktigk+1o3M7vzrgebvsr8/
XBKJFoNnQ/c823cqjS0AZpiC4plnub80ZlATBzM9CeMgQqo/NunydSYZDjllfTu2uXuh+R+zcYAO
fA/muJuWPvhhzU99QZYN+KPFJlKDlVJp3kUHsMvm+Ut8fpzP5m89p+OMH9KpUOMJHvCxnB1XaQqB
siUZ1CewDW86sLipxh7uP6JjIKaqEArDXxCPMt8ozJIG5kTeiyRSXQ3jtMNzlKS5hEmsh8XDWH1K
VX7GQV/iBNnAIJYez/YzHm78MRTrNtwnA3KLO8g09HdSqhCBzPt6eJkgkDGfiyw0slTuQbRSxKBU
uVofnC5nldOp0yCQ7jw5ltcYxHfXgHxhgpNMdo1Bh9E3yQoumDpfva0Ji4t2q8wBTAPfdS2R0Owo
RMFjyo7Y3SznVoJRBBUfnHO0L4UfWbGuERmuzPShmv2J8j2iMYCotQED4b89hfCCRL9prSzdH8QN
wVUbLlyjH+ThMf1Lb0PPeEylQBGXDlwkkS3jcIw5+susYjWrzq6YOGRsjdmau+M65Mj/TlQc9+Oc
m73x6GYBJR1VMEj5Sm/NiZT6EwOE1Ih9z8mmWpdFi0/yXdM8AuqR2U7by32qvHqAhwkSik+EvaT7
Jaxj/eyomE61tWn8YNv+zHYoaMtTMFdhNpPCRR8f0pTanawiEVzokAzopgtKHh/AXodTTNOeP5kw
Bs2zgrWdbCm+7+7D1u47L47/Eqg3FkkqWJRAN0eF0XOA31lYufRLqW4p1p2IfEqizhLAyEj9wF3r
OdkdhAn/4PVSsdMJh09Qb320MGRwZgyaUKFsjxM1lum7gGXyn01ecFYRVLrGjGA0qhgu04WVJ1W5
65aijR8A4I8nVRkvagDSFSKY4GavM3cn/wpDXBQunAP+LLxRMa8ZbTw9AEXvVLqXNyW50pmqt0wP
WvlZPogJKbLfZKzgvORfKd/aIjdGsfkqsUECNPptfHCFwKnU5UDXrSBA4t/fXzvLa9xTt5wkXzMa
ulIgZR33VYcd0Yf+K98t/HfbqGxu01l2YnXBLosFKbt8bGfnl46V7jIMQDJagRQMxE5TYaNTpO9j
5+TvfV3nPckSpIVnRZw+fjqr8wQmpUW8t8RlgIt6KnHr2Lwq7uEOFZqp7oEKstCdaryKkIInHxXC
KApOOnHS15f8c3cHUbzV30om7A6gnPjVz0Ib7Y/1FW41xt57x79smlRsXBdb44XOGHWkEPMmwknn
tipMF+qH9lvDPE3ZxEb866CKEqeP+t2skaO7PkZjhYvuFdPnwaaLnIF5gmU+pkUtqpq4Vc9PHLat
ZbR7KDFXjhn4jh0RQX9MCWVLpZiy6y/ttIazn0oADReDVnMtXFHya2eLZz2azBz1xEGqu/m0R0gW
fzxqCFMjSFBugwL1q5LQUJvcTtV9bvhP6rm14UdQ4RGLAryuLGHGES6iDXwpbH+p+50/QxMGJQoZ
kZfzbP5b18lopHbjzqelB9pdcq168elhdEEgWOOoxUriYRs/SG6adHE4NAW0hU60SIDU8SI7rv2d
RZiBJCcmBDsRXdD4azfxZ7R89n4JW6sWOpEmnjCQ4AJXLz9y8oNm0DGGLfEqulkOMlQysjCUpWTK
tohE01SAwbHPGE1G7atLhginEAe02chXBlo8NwL+MRktNdEuRZto4l24k0HcPgUa1njR3rfroKzg
3jWqvVb04nfLtL4dW0McvrkMB1Xk0pABZkIepCSmK1F1ThBGQ6h96/0TEFGcRZal82DoSh3CeQed
jiO3grFqxV2vAhYFHqpn7y3V3fxqZZNhBiNhffPPSt18S+fXB/dXzt2FKOT/iBHku+bgJaLfRUp7
nFk0ByujjsIAgw2CCSpYv6GndA2V5QlwsH3dQIHdUrnm2rfVZG/CLAaf2byn64Tw1siqkK49MIqq
uVhgwB7G+qvfdAerv8O8OsXecgA1KHsrMZBIq0KkHk/4ans/Zm/WmDlLwrVWPD1G+QfS/K0qkv+M
0D8MLPBGSdtEtRp7DiUpXEuhplVMIfQoKdlENh4fui2xWMynbrMPVrY4LiQGxg+eyvr5bUImjWbn
K/5SGYWQ/cRQzEq/zxPdcHvu+11Hvt3zCk07brnLOB3K8AundZrVr2fZKHGdQxcmDS77BIrMVd8u
4M2KN2RYwYg/pGFTSznjeloPJHcOHH8hUwMuyhzmY6ukvgDO/VCI3wxpdvXLuGbchvdiMU8fSJB8
1+xS0johuinteOrpdsWbZRSnIlPpkP2TmVBCWPeOLNWCZ3mAwRT9oDA6RfdBGhBB3jL4VLx2mbpT
K+Wm0J792zx7YaPHxD9DQ5pwjsne+PI2KrvRcBhC6mG/yMiWHRcknW5SBuh6oSl57Lmd4ygwuY2e
OAIY3Om1GjWZ0WesR2V3lVFCz6ud+icIHrduDLnXkfhG1OpGXVN+CNIVuHVb1D2jr/vQ7BfPxtmh
X9H2shZDhO+kd9sDGaHMffYK5FWE6np9gP4HYBZ3e+1zAKonSqC39fl6SWjUb1vlLk5nsHrSUCYe
1Sq02azjOS5uoP6qNnVexfh8L64i/1IYaFENXHEWFJj5PFIluYI3340QTD49qjSjy2iMKHOEY4IQ
tfe5+LMnlwuAxRFjOZhtNvoaSRILc+rxY2ROnCWSqMkpbGl8suUe7chn5MZ7kO+1q5oppxcwcf2X
7K3i2PFcqud4T/9ZL/bqAC+mPx13yeHj6cCzaKBe/4dYpxUSQzK2YwkGxrlYRCB6GZqGlrvfkhug
SZK6bfT4sIbxbzmIkw87h1NTiT9L/2XADwsVElmp5jnhyxdzrisq8noL4ek64Oq1WljxVKsIunw8
WZmT1wfe3M/33rRgH4Uogoyzt0HBVBKJcz1qXVpF3MNFU3RAe9fKHO1JVdEjhmLpba70SfBgwIyN
oDbuVjfERrdGI4GIeJ3Q9BwmbfXn3UTkXQVaBhxZ9zXnAz/hrGdyYTbEAKyFRe9DL03uXzlmJd10
WQTdk5rnE3DsIg9VfBV+yvsCXuoZ4bkB5PLrWdKxQEPSTgLC/aMPXeMF/gVvM/++6FGJI/HsEYzh
zX8WbSGZ2+Mc91L4cKQ2lsuGO0/bMEaaAWBpuSHfhUiMphZoIia+7ZdzFMIIRrBcX/fd/jA7fieK
W0dCln8cfRU0YA+po/NPYcNltql532gKtPvAZxKhqBPiQcFjYYThc8nuYGlL8qxfe4OeJS2qfsDu
kpeZgtuKLAJkINqvNtTY486TPSlckmgbuDyXVXyzCKP7q2VM8tk7xsiu6uT7t7h3t6hGoxHs/O0b
RdThkAp+4MtPbZpM4kCkRayi9plRhYGtjBhe6B1BSegYCtiEaXAf2B4sDTv/YYyBrkF4eM/EZaQX
VjIz1vhr32IkDk2xxjQpMolsw4c5kj/j+HaorH5TissfY8nJLagoj0V8OKJou14Mef4gCnQJdiBH
D7YN4YNy5fvc0iB3gFCsbItLG5gEWQiB2+7pMCMpOXSlJOOFPs3uF6aztnqQTTMFQUYRYFE3jUlm
+KweI9M8RCmDGZO3LI+YRk68+1N5VgY3mfLtZsq0c4x0OTnXl4on1D4RbbgoBo53KubTPre8lBTu
R+DKZtr73cDxoUcNZPEgDCl2wVq6X0sFKT4wyPc0+Kbi9liYDikjCFz0MiRRuJdT/uS2bp8lLtE1
UzoqRGGh12u8UZzAgMDITPdH9gsM5aK/OV9DKHEA+yyYNMfMNu4BY3B3Dh1fnXFcucdFh7TqWW4z
yi4i7StzpNDkAhkoSSI/cSN8zr3TYPv3tQQK9ZKlIUXzG+QIszP7bzjZT5FrGU9x6b++DfTfGRKc
fcvIhrOPKufseQysduUImQurZKXs25HMNFaoWp6f9aQ+Q+m/pDagDis9WNg1aIFHqKhhjBSYrgEf
YtLlEKqMT6xqzDelhI6V3/Jr/rP8Ye1pbOK4FnS9DY57qWiYLhffeawWBME8xXh1+WcCv0uglzB8
wXGbY1Bd9ctOsMtD7Ws6hBWMzvvCTG0yrU+atRUInLAnKgNQojEB7CxoKKAJOW5v0Td/usRjvhZj
z5zqbuUtzddnJz3Qp62t7xyJb2IcQCxKaAYXW0jzRRbw/xqRPbqIspr8AaCzCczJSAyYpIXs8u33
QKT4OWNbO7h/YCAGPylxvhGXJRqpvmIjBGv5jWeuLd0XEVHIq81Oh2JgiegdVsPBDnA8HdM76SFF
xfEmqwj47FDBevi5MtxqmgqMb0RgEtX8+FfdoDKzpwFq/cWCj44QuR+cQwSMuyXm1iWQ8HFWGMAn
nlXJJCHoHhOUTHVlPMXfaCBGAbPtEaaLsDLW1IA3TK/Zmc15w0332uffFkRSvyCvJndRA+Oewfna
D5tO4fm0wraNfd+pFNLCC0ti9gJuKmvgDDZKxX2vUH92Kfzq4mvHwDCE9QPiN+bYyEpl5zPB/YGt
bMd81gO2EfNuyHHK+1aH0NqliUtVue0TwDlYCqmZT46mv7Y+Fxmtxfs2iftM7LojAdznUi15/piw
4Izgm6l1U/xl+JU7AABfJP+Gk4ISA8jHwEJvC5JI3EZgEkppja3pKdinXGzZMU+uJIDcUYLkbdmG
4wOOZpWlRQ+33jVTSi2Nb8bw3xt1ozpwwBpvm2SAs7uKN2s3gfaKO+J5Fq1fq6SoFQehpXVHBo4s
h19X6m9QHH49vNuk1X6kYmlSSAENqLPl7PYbOIlkeXlNJyxBQ2GicqPZxeVNGurwqpg6uYtP1fFN
w9WvBY6JIuX1QvQeOGnxPMbkkyThSfAE0DB3nbgHzYZ63Vz0AI1AhAnvXaOcaGusRe/W818HioWq
aH02YsjkXZb4WttZXK/sGcrbgZenmb9kqUEjy1jenqmH4fmm5AzzGF6AhIETqpZuH7/UiK0o3CqN
JUDeDSBmBNNULVujlHmbkVcDC4wVwR/ZdFfJ8KeH1lh0mdSolmWgCZ2dUUtCX/Eu3gHdC9EKMyT6
LMJhid6l8NeBa9tSuBsr3nw42sksdMH7pW+o69+2J3VummCez+B1IOVxRq9jZHnNRnyO3ggpWa32
6NizmYmp6gOX5PzKLlsJaqdzF3TD3R/zIYyf+bgYRE2iPpae2vEooRGU5kH51KaYRpIYJsoUEXh/
e5d+UeJCpRGfRwjelBZ5ZgngPFtuY2+OLb5yajiF/v7z2ct1yyDm07sipwNSnH+dNLHmUFbfgAZF
yU6TowWw4ID2DDOFnbhwRmyErgxEhgBwLGAkePuduKl55iijfLu2rdGnTs1QoPOgd6T6jD9gallm
chCyGtNEJDB8U5lFQkYz7Amhy9ysGjYHDT3SmsunBDMcGnbGkUg0jmn1IAx8ALB77f8K1tJS6TfK
vkQwxVLsbIZFl4Rj0RVPVPv8BPVsoKDyJZAWI4xsvbSx6HjilsNtnNNSvu7dOcQ7pH5bQ/f/OKKn
VRKB3W6SB7/gvmWhvxnixCyZ2DZ98Jbk1RereYKszqBXwhZp6gA25y9enLIjrVQhU6h/OmoRJR8F
Sq9d20P5tibDALrlNgE8ku4bV1IEYCI/g4zAb79z23ZZa0XsAnFKg4DomV8dbFAsCKkn/Ex2Lu4w
lY8mUNE+L5CH063NVuFbXgh96X01WsLnTsyNvx2pCE6Kiqkjeg746Hw+q9swq/C57AiCGPFj75a0
bd8CbmC5heGMs/3/+9TH2g857sDo6IFYIvfS2pBP5kV3kizdHg99ks3ptaXQ9ai2s4coJNBYo1Lt
7gtW0SVOjKIf9yTctHrU1U32iSt9CDLna6Aewf4puxaEuFcbnIuV3Ag8zCgPiMPf0ywjBjL8P+V3
p6appPvOHiH5h218RIGi9XDqEqrEdli9dUOOH9FcNkhbbN9p6AE6Syb4zNd7RzsFC1DAEYLplD2t
QNfEWuqEWPEHUujNTnbHui+suPGEWQtdKnw1KvLTdHAAZ99ku6t1p1cCoj7aJIEXYuwhOH89GbD5
SaNTT/Lul0nsdGVWRyteBFkwn9enSsRUmXNyWY0dD7MJrQwfjKJ+dVzSsZYzZyQ75Y475pvxlXo0
0nWan39jjrZGEpmq1M6dlJ7d4LJKUQG/wLFghJfHTtCERapkb+VZqafN8OLXspg3bV8YRzMF4FjB
OQi1qnc39cEdnI5EACil9Z7FKwkvC5TJw2Fo5dAcm7MvOdQ3fasKdc62/I/yITYS+PiIETNGMuIT
wLacQd5HI/UcKhK7WQJzY82LizLlmROk+p0mAkjzUuAz8xiuRJlTkjtoIFtVVyXX7vD1eWjswDik
KNqV4CZKn7hcZYaxe1WaoXUsCGQAwUwIoAH2BVJbvyn6sW/k2Krb5jfYdLD6Hhpw2MstYDmNc3Ct
7nod82NcBUSeQcMWaa+jLYiJRQ58IzcUZ7teXNGYv6f03tHmkqGQ6Gd/ixBjyw1MHExwSxm7fkQI
9pHtV5oAVqJPQABRFdIASF3FobK7B6M0L1ejBEo2QEvDpcEN3UmVhleFKXF341T1NzpGWgDmKauE
/u/K26T9KMq5vVBN59moP28rVqz+N3E+vfxIOdHWuJApYyV/b+cPCxQOzC/rx919JEjP760xTbWI
s4n7fZdIvj2zo3Fl8S/RF1GqaEX3dcPAlSqf1ns2Le1BD+gTE3YKSEoQ855Ccr/ndXmjNffzRMFl
rGZdKVIqW5D8VfXT9OqHHSSPq9f8zCpDm228fP2qkh9XbsZdds0VxtbwzoxbDmzwJjQMIWjazco9
Ua1oL9fQBM1QiAjtAKQkWoTaVhsIQT0nV1yl5cOKjKG/BXlpVJs7c6OfDMB+QggB+D2ClphAyqVe
GQ9FccpTR3XltIw2yFkJnGhSaWhq+pHV73KK8eabXCFc4FY2H9q/qw4ZIhjFletzxZ/FSvRofXQC
iZPiGIuy+yQEI2gJdCfOFP8/+fVAc+qbAk9ubsDrd7m25q23iSVvbArKLft9Q2sCI2zPKvAfnGAt
04vBcO2DPlP6aHItvInSI+ue1yc4L1x+QOckO+RTAGVtp7HsndD/SdSrJzopRuJ5PfHodBDeX4J9
iJ16s1RvaDLbuUH2fOhk99gmlkuayxnver3S5E+NTt9qvAtjLk1Q8RZHy/yqhy32CwMEV81sfe2t
FueeDP5+EXw41UwgVc5yZOIgH8E2yw0oDoBNzuCLNxweddHtNufa4i+U8PUqPKev/Ekaon6NUHuC
E3hCmmvv7wgC/PxVbBafzPYPc/Pdb6LaKwSRw5L/pzRdLAq4/CdrysGjqCP7V2BApi2nPhJmOQ5T
mCCi6tSK2c03xZyP2ZNkZttKhk+sNn1yNxF3koC86DMXdrL69PvqCmJxL1L2na+Yty2Yx+vfEBBo
INFCyJs9D9NwCIKThZQ0RdtgHkPoId/PTLLa3CgMrvfh8VA4FNFrTbl9svPRKgIaftqJRHQnGF/G
PmMDA/bIMNwj/MzPfZSSdHeeK7SlMBeEM+d8f7nu2ZmvZ2379WlVl3Qy1n5iL0larEJMNPBg9b+a
BsSoovfnrsX9AG3M353D65lQZpdi6p84l2rnDUazHdlzf3W/EmfzQAiSJWrhQDZZW4Rpft+227UF
x/3QswPnLE30Wk7XZemWD7MV/I79oEW6tA+n0X1bbTQEKZf65jyRiLE3thiVJ6tG37Pnjf7DYi8p
ObHA1NglMRZBG4QaQpsMxxlXCHwkb87BGZoIyc7L+LPoqowXL7I85X8rpzDUMaSoqGqAt/UX8x7x
pgIEGJJL1fsSwzath7a5TTeKe9HreEgysmKR2b33QlrBpNaFj8Iv+v5og+gEXe67ifjvSWiF4Vzo
WuhpNiRkm6aHDceLeFLpW4TQq94dpfBAE3jnom8PLLtgUOIDJXuDGzfNL6CumIhwxXbdifGDWNhT
lzjm6R3eAyJLVh3lOT4zAEito/qPH8oibqBnFB5MSkeCc8D3ACb60AdnRXYFaiwWfuxF5XC9QFZ6
TDdpvwdGhwFmQle+iiiOFgzbCVn4UDWRXHzOrsNEqmOop1bz9TiVoOG+NNQwfQOz5dLPdhcPzfPf
JDU7+g36t6mSY8mPNgY0oiw5Y1u/4JsY50yCT3ofD8swFKYgJB8o6voGSagf4f8lBTkP3RCcSSEf
GSYhBd2PUcjzGzNUgzlRQROFVVlNQTFzLcc3nqpaCW3dc0R3xyzVHI5ZqdT0G9te6+8YTaQt561a
jcICcawOjipiwungd/M//d+BdOS+Oo80a9PevY+Wu682lTusgcr1fLVLgVI2LR2HsLLC+41X9raz
hy3BIbEYZ4JhjzQXK7IR+i0vBRKzzX1WVYTUgFiY/RV44d1YkDTP8NPZZz6c+VScFggMAxfgAcLE
uIYYxu1L72BIQPzBzufPHAhjdPO/v3nyEOZ8Qc5NuKw2Eqfa2/SsAqT3/cODtobLHLjL7Pjsxt+K
Tk+xbE8o0P4O0KMA4VsAwsV7iLPIeVkibPWWmbZj1yGCKeMdifoNjITHoEkXno4Lw1TqGzrBShZI
HnVwyuz7XYx3ZvWDbE6BwtekWY8Ss0PGB6NKZ2tTlYht1q1xY3RjGatrv70vv2CShi1KbjVxULOD
yk+H1kzKqXeNS8SHiErSQUwFf8RQLJqKoCPGkdyvE4entj+Xrx6KMvAtW3H130IQ3Ri6WPqgyn6r
ojuFPwIaEn6OWTtnWZ171+jxGltPL5AviD8BWy5cdcGxGAdK3aThz0XdipCnJAF9/1NdpE/3GBRh
LFsFadzb1BfVBbmwkJWIuzRMYj9Xy9xsvng+u2p0na44/ebVXO7Gte1gxFKcVweyAuKloctDV7su
vcLP9yzo36Xh6C7XgFDGHQ6rbFRHdIlouAh2dAaiovwZVRac/B4aBnzfkkEp7LCQvePoI4r8iQU2
iwPNQLEp/Ixz/dvPUPOShQFl2GPyySI9xpCR1yFHmBMVMfrqTAKNwYNhaq7aOhne/ClxlTXxfTTO
tGldhKOlEeviA3mVWOu4k9OeCu3do4l/oQ4z8oPkT3JQwCZUa56LiyEMoBnIgqjVnFaCI/0A6TIC
Xm5tA1YVUWJOdSZe5bGk2/C8TH9h+yN1isSxLlfNPOMXhS0YUT+71y5V+5Y3BaddQ1lvqa5Xxmx3
eOyUP4tFbmUo+MWQFcJF0Ux7V1OW+eTUorAjFnsSGtyfydK0qylcQ94y1cH4YdIlzXr2BJU11ncC
1RQhhwvIbuMNjlZ7B+rw/as4LvhYdUP3HN8GYMB7X1esdupc+7U4onZAhcXokSueL1cFqan4gWqb
zQl1Ur4Q3kzuHg4UHkLexRnqquIQ6bZ+os2RzvXR0/TmCpCkR+r7WgPJd1SIIZOwopHWqhZuBnCc
24k9Paq0JK8WdQnc4D3DjwPU6kxTtLFt5ztwKxT+tR8aKDEMq5l3XrrH3VuY2qfxh35SUzRru4ga
f+cLVIuBnD+tRbwircr1XWAOtPeOZzU6aOOeL8JtqWVmmPSFFMwevf7p5mesFF3bD7Fatcdlfuiw
R1nuK+YO/sWd3EmQNT+FzsEMHJ+MYM6+CORvj1mTyn1iht/ztFOJgPNm+e5rBUFauoTLj3z6THSK
anrs7dohXuPQWTKxVXG1I14Lj8kkXAQ4ZHEyMRiQFPEkquKuu56OsfvSNsBqYimadHIN14dof9Uc
qZPnzadJYvBbVo22eurknB3YYpJp05rJ3AyfDz2e0+qv01CCtM0KVMPMIYm4Faxplwtyq6Z2JLs8
ghiwnYMb8xfSIjgakwvfy1nogxkPEnxgjsBV9IHZVVR9xjupgZw6PAB63Guf18wTUL9oz8yXI1Pn
NmYEcGzGi5J3M1j9+CSPmW5j5CeuLaf1QvWaTBk1dt1xur/gpzOEso4h/M4X9ZmsgrGgPQaaJ9tj
lizwy5pssAvt6I/JVcylok4R1tsLQiXbP0U21Xwy2CyjuiFICMePyZ0p7zPqIgq6hDV/ll1AgJFp
obYsWKmreOyObW3zLjkxWcyRIuNdtohDTzIWjhaqKXYxmit17Up10PI3/knmBFaGyiv9GLE7C17R
CyUGhdB9absWDfF+XIiZs7ielsH6x8IKTxc6NI8C+r3R2AmYc/S8Nzpdg7lf9q5u47+wBzGiJisT
xLeEWPDYUqRmwMSmpQvq/9Z9a5geWF33utnC9qx0MRCeeJyef/cnTAAam3wFyRRdtN+vkTbRygLZ
YSFaf/bHfoKIK20rEkCxIaSbRaWkOyx2yg7OIaySkQpMLwfYP6FYxeegICT4x/OjCZGM6shBSaPa
D0rsaJwo48tuNTMoq7UcZeyWyAgYEjONyLKzXtEBh2++543eahYvwF2noTJRwNs/ulWuJCm/tEs9
B2yE5Eff+MGdWzWcLFnR+iARVuotRyS1mDZxEsjfSsJYLdJ0Bv6aWu2FYlzaCA1DWj49KxfPuTwL
4LrRHyey0VvdpUs2XAD3B4/bDw1cf4FkzshWwokIVnmuuV1P/mC9oqua6QOu4qjafO8XqZqb404D
nWfBnYqIsGABYhZe+asj4cpNJfD0V6if6/rvDfutdM4Irz1IlbZOEeIEYvpur6X2HOZ3pwOuY8w5
Ak9q5T29mQ1q1ella6bbotaS3t67O+GkZ7fd0CCpQ4gWAY/enO2zdh+AjAx0hfMqJnDMA8PEEp9e
wMQr9fnE0lLCGZ3vwYbb6leHYi5TFJOh+cpTUXRjM5wXPynzDUcoU0EqOmvliBTR+ufpnqMwVXG0
ckUd+cRV5hfkJdRVD/HBuOaShREambGyG5G9gPYrZVRafAcfDjv7mT4IYIEgVdyTJf2obuh3Lz6i
MrPbOalk1QHlCv5nu9QF/ScwJuBkfdLWDWuoarxcXZZ3/EKj0/YBIv7TiCt2HWCZ4cuRFLmvZZR2
mW3m8Tso46xBvQWH3yZhPLUb32ZpmwjwJksajayPPqqeEpFPW/7ItjzxeqvZLeyavS0OBsd6qd5B
Oolg0NgdPWC72Lg9/PsmteIBHEf0UZBYPMd9xrQEn3CZu0DwFZbi0OVyDdeF+63uRA2I9TeSnD1E
QgLv5gYtb2we9HrjCg9KDs3Q41oEPiGfVzIkiemt+q1kIwns6TmsHKzHNHeSAPhkYhWHoWgSnmFH
ssaiXzktN39nmhIU39tRKdKOvK/uviyY0DWOhnj4qhQVgpvj7QEsJNdAO3IExdlEZ5++HECUxGRo
agVPBe51Qw+RCJiDRRqwZGQsk0dNtIFG70Ko8ldV4dvhyGc/XGIxMPsD9ZtPmGps3eSkgKdHB4nR
janJOIrIrO371BQZnzjH17CBffWI8Cch7/cHk7fjJA1CIUtPXwD/XXeehJHGvM0GJjAr4KGAoF7F
tpioN4WIoTlWtvJEz1eh4L7BIzR6ICmGLoRI7Qtv/3zMaF+pe4OB4nfdHIT2k5JDg6yEqzn64hox
2IHQ3RMCTN/dsvKbQy6gtiOdhoTjKUC5JH9bjScw3UjhRgrQ9eczgj+YmJgdjhVP2xhk8bqFu63K
a2P/oZWCqx/weTMDJHiaLbjdtfttSJS5VVhZXzkCroNvoqVqWggn+Ev+gFPXiEGUtnvbWidq6Y3G
qOv5HK8uQMfD348UL2aCeeKOoPM8BjnfnLp3Tb8bL3IDMOW9vPkbNn+wuVvHI7HeWUhO9DJn+Pkf
B8fB1YSsHn5zQ+G7fo6f5ghXCiWiGFmzKK3VQAFHdvO+BOLH1MrK3B5BjVtidvzcHTl02+NuutKM
9ioMlZC941aHqbXtoOZxTxg52z0Kij04ZHaIhXD89xm4rGWoIk5X6/xTCABrljp7Rc9C6sKDhLC3
AjvF/3w3I1h5KNkP6PLL/aMZV74hHhKe+o9+Ykvfhdzb8Xu24+KHraAc86VUy7ZUkvQrGvjqOWlT
RwYKqzIkpGHJDP4Ny9zPInCQvHfE/G1egAEO4iwiRxMUdLVuKo0XnsbCFw6DzqeYLKpP2c/q436+
7wcSaItKWpgKgVKj0sTB/D4WYEDSzcf1xsLniSa/NaxClg4aWGob68Kr0A/tudrLpDEHaMknMGdR
cr4b+QepCEo2p5UKIegI0bGhp8S4Nn2g8EZhbzw2po4Do1tJXYyS3KzbMyObLut010Ovu79bKcpp
xnjaTMMkiYcRGVvYbPU/TZ3+j3wQ7e3R0uN0QSPR78ZO1aYliSMOm5rPF2zLaWDeqrvo9qjdtR2d
kobpn/AKbLFfuNggWvVUomhBLVMn/KcRWJLavUFambyIHNPExayhNT7d0SAtzd4EVStLj9kMlZkR
Dije0jH5VD0slRD1b8/bz5NapaqpRYUcjqEqyHXen3s1ZgkgWc8/n1k+VtzO51MpzTg6p7oqO4tS
a8FipTAfVTygyOGvYHUocPahxBVLyB8gS9O9xZ5PnjP2kWUK6Ieewv9Y6XXn+Bhfi+6VdyQ+WagH
5MY9lxBPfnSzR59jKIyJ8sKjfGHgiUFT/lK/kq5TIilqfUuSjbvawHmk3VtLIBkYbVYVsGQsrAJG
KkyCKc/i6VTqyqB5lLYzQAFxUUkWbViJkHUpcCxygqAACmEhrHFeA8zEBXO0PD4jUI660K1/3S0W
tv7NO8Kr7aPqaTwpK7wCKyJVGcsYsoQdWEc0vkMo0HHpStY9MG3IGu5V7Hx95uiIGhFOuq+y5uEk
oiPvSidAKscsmrDTODRM5tAnKdBkMak4vjzbjfznGwzdQ8AaNBVYo0gfzIhwGG9rO25lSmz//cl0
NHIalscLqMdthGrlLUAeMcupfdPpbRoYmnfsRHMdy+DqYj1vjaQUck6EtVufe5dY43OxSNecG9Yj
ccKeo67R5sFFoakYpLBJQq0c+6cCp5e6uiMZarqsrvIETcoKt6jRs3jCMhKBEJPhkzSIPp6lntwZ
bIW2XNUBIIj+thluRJ1BzJ/tLRtFEX4he0uFEn6eBh0J7Pe1aXdh5nkFNKn9kqI25CJwSsc/kaIB
44UaSDzIYKtW8g08WhBPmoASSy4nYkJ1Ci1skuAYg0BPQlWpFlmHWz3cs+MV0fvLR+BfqJgzCOH7
fWj6kzVgGulYbAKwPGYzpGp80xCJLXUoSqye6L2aGpncC1DS4yhX97JuAx9GP0CsUrHVqFodvgcF
mLvlC2MNUjg+iooXwxbwsH8r3JhZwc7akCnS0DmeW5DFt/8/dJqCgDk4TK/EivnpIbkfOYZbxXiA
sUZEZoEqQZt0cgE6HuoE9k1PHk7MHMqN1LCZDqOracIv40k3t1tqJv+R8ibhRtwliz3CK+qFzijW
wMdaU0Y1C/Uh0mrbxbfgQkMHVqjHBFZpuzIyYNyKjRFjSxsXqpWFKluIgbLWPR25H4QNkEw59fe1
H/dKTBHZW84tBTp8x9dcyosDBzckS4CIzvmqOgVlAjOps2Rusa8lLR19VEXnJMzmB8tsrmnwPJQS
3OuQWjJeFIVjB4kcqMzmLMA6iDAIISe/JY6V4oGboK41dKtDLkYPBx3sCyYQaJvLtCORTdrpNLUr
8al4zDPTkCz+1reMgi8YNvmsOyTo5UZVSC5Qlbl5IK4QAnFBep0PRSOWBB19WlvCj1dJRrw6ZxP2
i0SZLR7uN379W4EUyBiNYgaXpqXLYanVilLF0XV6gmHFm0p0MFtY2OA/oxBIyxGxXzmjK8zpe9U0
OJQvGPsY8qyWE5dKP15QgiSrm7xTMw/HFWPAgXDt/eMNvIvvduT/iyTWNW194t8Dn4UjXXvRpX2R
YWMIl2lnI3brNdNitZwg79zvjMQuIUX+oJkPoVPgpzaOYkSC44kOJ/fLZ0V4+sLGDKOikuaAjK4g
6BQJa4Ctimpz40XhNPArt4VJGvtVZ7IicH4iVkhOgxs1AOMU8o09XMbQsHST213zljRGAF2dFIBA
sR2kV5gUKl1y0nISJdCHSjMVEOTRg/SYaZY/hqrZBz7q57dZbWB8Q5W8phRhisaUq3+mCJyZfNV6
9AqxsKE9oGelvb6/hZFxSW4dUjG6jDLAda8OOwsIN6Z52eLNSOtl/JGmO5/dW/WXnwfJn/0VipWB
C4p1aFlOoY18KfE6bH0nADBwFTdb+W2XNbJTI4Is+BsxdIbCx4TU92R2ZAuH/p1i148LF9EdR90j
LHfj4g7SyqBmfjzpDVmOu8jTvCIUP3y2G9iljP+3EOLlqFb5OyajFSKTJWZKxavKAUGNvbRNgEEG
WGMwqFB/ibVkBlt9sqgpWorrAfAyti5z9RMa1fROtjgLbiVHO9pm3dLWE4AMcJEKoG0TM9pIfOsd
Fj5fUyjYyCXQeXTlGm8IWcsfh0jDP5BzzmKcignNnYbU3SYR5+DeV7PLXfUrRn29tD5aQy6ikwwD
O89W5+jExMsaVsDb7eWEFg3HXo0K8/A3XlVlZSVijk4NXFfc6w/7vAwMVG9DwBeEHb/6NVRFUg3i
nqCmFAaifEjgkBi8gAc4rExX/7RkPITIY4x1sxlsbX+OMfL7ns7vuh/uv3aywpdnPZzEtes+euiP
6VYzfiI3brh+1t9Bg7u1z8/DSPbiWkJ2XxM6gFlZ6osKGQHEQSGe/fAxF7oECoD+X1ulcTQtuBxw
YyDlPek5GMGs7gDn8Ndd/l8KKTXLoGYYwwOtCvM+rmq27LJhOHrY5Ov4Iq/XUSdEFhtdD1m+DXxP
rpsSEZHCPh2eRLvzZEYSuGlQP2dYVC9VPm/JbUCU31X3aOZ4FnB32pVJWB4KsNnrmw5oahPJoh3c
EZdK+GG2pqNd5HPnp3YXO44+eXzvnYgIRm0WbAXR/GqNxWb7BnmXcQ15djEk9nVRKCKEZIhd2X/J
NXnx9lfcibL3Y3eC3A7tLDJAjNqybvq7xcSlZZfJGumV/PlQcyBnfPDDcXf9zsrShgtTZTau06Bs
gHdeksiotA08vzx+iOmcVtVQz4+1NM3HPXNE3tnjxdRvVauYIBCR4KD7HkOeEixH/5S367Q3idry
1nVhc6y70qHa6pCOebsG2ONNg7BfabLWY30n2FCyE9AByYw9NlekAwZJ1unBxzaLSuJoyNtjceJD
58wKoYS61zWqjt+TZ3Je7nNPgukR0yZBR9xaqPskIWNtvoYVERuvSw1SyjmNE/8ZGNmWUMlMiaaG
boCCp2nOlvLNJOoSUwk59Xbrx1R0FybKIQorhJ4mnJvdbS9p2KQOuoJxIHG24CV+Xucsx8kLIDsw
ry2K0whL0YzEqMJcqdTPnjvU445Xpxtng4im9XDnQeEfq59N4rsdwEO9ho/pPq6aRn9KaXODLrfR
/3mzc44rSkjJuh7LOh3cNk5F5exyCWgCiqDeyonF/szFdZbEMOwrbQxVdKboYVBxcpmDCTxnluUB
PZ2t2fKHxWTic13agqWwjmBkiYMxkbrkBP/ggBblL+eH5TW86Nvb2kZN+RVhlGfhpCYMERPJ8t+B
1kwCvehsUkAoddM3FLt516OVWJ3f2fUpwuLIYE0YgsTFaygmgKvcoRe7uZAfvh3/rT6h3R0Bi9ZM
xXew8u9YQOiKMOReTbbZJzQGvqSN2G03469YFLle1PjRCEEBXCGXCpmCieD9AOp8g26ShNUqXlSD
U55vI5i8pbEyFp4eBHgfnGpBahlnKsRBKv01Qq99bGvzEjyCl3tUsf8mZli6PgMUR5K8BoQlS7Qj
CZmHFt2ajTKD5/vfIgAZNpOJljNAWpTUNyhtVpplzYl6HZMlPozugF2BGHJMj3WgVcHyYiRPOkmW
ee94TaQLF2DpNCTcr68YQn+GNSChdKJKdDLfz9GiW+LskJxkjvwF9/lj5djVtKvWcLLVsxef2QUz
KEbK/b88vtsTrYszhj3hbxND5c3Jdjy1sGM/lTBf7FmNnIgvNurlOA6YOCiy80fLKdaL2tO0nK1d
pAYdkQl67hIrSqO5JJ0tAApGBlnSVnq4NaNBOVWHNYRGHDqa+5BHX/lSW51DMk0C/gAW6APxbrrC
YYD9spWR6+u1RkZdngW0nRBjBvY2cKaylnXHZ245DD7eGZeduna9bnEh7StdCNeMMnhg483QTjrx
bgRnvsEXjcWSdHT7ambB+RYU5TrGRePjAKJBBy1cAE4a0wB3/6DlpmAKNTbUcOA/OVkr7hV4YAqY
89hYkyyDa80t+00x9mBBhG7xL91C2wuVztR3O4wt+T+6Wa6fguV0tYNhHqPqAuL9F+39EJ3BHte4
5kLOmkiW5EEKe+4TsYleUghYupddSbf9IAalexI9o96d6xPP8cnbEKqWaUc19LRXaUo9bi1K7cjb
sGZ110lwV2T/0gW++iyE/QabrahVlp6IlbpL4Ha/RRJ21clEMePxLrqd66/Pfmy0P+4TCNIrrsqI
hqzyv8uOxdH5qArbP6ogu9AHyUTCt6HXEeWp9FaH5Ai7G0yl066KFcIfAshFfTXYK0oIymz36JJK
5lHgLTL8i6WBOl2LbzQ72V7rwL1uJr7TZ/NGia7/vW4pgI/ttCSwFHUb8kUHhwopJ23rxKmRsdzl
wTT2/3C4P/0Cq59hx7UVA3F4qofQg6QBYkzkL2d9qvFO+lZm4lI8TwA60Qn4mC+mXjv8Ndw4a1j0
XNiZMDNdKlaRzo+QAAjvtt3mh4fvUBmFucScdAr7NJsmndIC2I+8Biq9tfCTWZg5ncZxH8ITYjZ2
uwYPy5nZS/QtcFv8kUcJLx348m7trIPe1COJqKR+mSOfYe+gIlqnsUr/N8wTt0vppOFVSSBsk/bV
k+INJ/UIVo6XbcxccNIn6nxbfFU/HXOggpYHNp1SFTMroPXfhvu4sZYx1bEDoRNNNk1n/Ew9yHBK
9ZFIoM1f8ugNQpoy77PP75XzrJL2wo888nqX545G3sDMusn8aYX6ylckawJfzHMVS4I9ewy5mYBT
SJFGXX+qdpYh4rXis0gMwEewdylFUl7EnzjZZ64sWTSyajkJYN2tHzOtdGTt1bVnhAkEhndghP+i
rv2gWNwTp4FmZm0AdUZoHocqAd9/JBT/c+5ZDMphi1ImrBFZirtEmH4cS2GGy/wb+ughFyI7OXRg
9bwM2VfxXgQYdhanS6/DPxKkgfVcoVzi+kRVo2VXMBG8/Dx9tGK4tK96lOA7/k7bQlKCOfvcboWS
JKfuv/YbjIoyQysESZTIY10LzDqm94MCvICk4p5q4fLMMO4gHohm8e77JQSKhSylIv/c9EfRmzbC
juCfCW27NoPBPfe+Qpm6ZamwtkVEesKF8e9qGO1AARK5sRDcARLd4JZQRTG5t3dlDsYQdr++vIfb
PKV6fC7rFfGZ7x9XN3KTk2G4dsN8ABxhKkfC0BOOrGHU1147YsgkCGm3jhXGZvAjwKb4BMzPkk+2
xhweHyF7nZlYRL3ZXMpdgdIQIfQdcsRCDvnio98xThC8T/kMwR4krvghR+6BVFbpGxx0ZIoBYyDd
DC7BN9OrajhLkBrJTyxDj4U5I0roiCwkD4N2q8RvozWO3aWW7/2u8O9nBqi4PivI2Ghm0ujWZ3E5
3JsFHSpDL29TRRLw+4Us/o1g4wdv/JTfvibuwPIO5p3Jb0TRRmxyCTyEeLSEsqqGH16BtcsRyGl3
rukSUjNe0R4RqjhMYreHCxteLEhzWxeOmgGnRbN5arZubB6IN/AywyMCzswFTt8o6eaVL+/daziO
c6zvSpZRo53RSP2YDMNHEWQQmmvstFbxnobZC0wMRS4cRvPhwue3iqdJk24qLnvK7v5NbW4MYeh4
ce9ZH0eAoRbAqUf15s/PgxH9tGmpaXTBQHKqm5+RBQ+0VR9WTXJubtpMGagpQL86cY9afjk/aMgP
lFDRN20Q7XjtnTOBOsoGNhEPVTZ1HjM/T1Nx+EeUgC7Wev1ESodJrZj3gZv0Z992lm3ulkLJSONe
7H8l8ZAVuBTQdhxpOCzTMSQntURiZU3DrkoAJPb1iCbTLKV4bx8bg7QpYfUpUOmmqjFKgUEbh8+h
4Dy6tRy/bceGwZaN875fkfxv1NIIavtW12/2xfsDpsCrdfPZyZAl0BxXcnXmYyhKiEieLlZZfkWD
NzT9V7rwRoRTOtC2IONEgIsCkk+mgdFCnX6O/uz/XciYv498k7kT4T3P5wnujB7nUsHhWm1t8hEP
6lhVmA2vpuAectf6LYji+3gu7krdKIWUFedGC0cB55X6hz5vw8I6SnohqSzk8e9upAJ+B82IchyJ
zUjGh97ONDa0hcqXBFKNAf8khlQI3xdN3BGIKmGin7Kgu7IyukMgFqJlw3Grx3zOpJK6/xY8EPxa
bGJDAORny8hWrRRmA+8CpqwXWueQQec2/7+cQoP6viSQAmeOIz9IxLrQ70zMalw94aRUQOCVgpVJ
XowfkMJwiIK0opPXyqHqcZ0uWCYDLu9wl2BYTq7pP10pTRe144YH1iHY6rLzehtf3oTifXLI3Eim
4ieQandwJOGwc9RubK7FhvhVssCERA67URbVZRIUcYoiemOWA3c/tJSbBFpAp+StvOPCwKB36k8M
C4mLB8nc5OBrvDnpjhr4+VRHKBnEU4cGmOteChZlz+oS7Za4thMgmarvtookEMpSAkLSncz3lzOk
flbryRYioHG6dq2VGDC6hI7eVdGL7IhQL5dMkgwpioAneQVatb9WFCJbFOn3tN7h7rAtR7mMa5Hd
hX0gVaQNQQTULsMZXMClONQ6g/AtViO+l4RnOASKu6UbQlI9MAu6eswhodJiJ3JKYf4rsY760BeF
UaJpfUxy4uw9LqSLkRYc00UB5CvIpCLuQlYLSfVR2Z2UhuVzWILV/NxQc5XrKM4tWpsAfmH0P7fC
GYvteS+Fgnu/HzyFKvpWsWjd4fPhNG76HJ28UU8ym7va6jRhaywXn4UnoxUxS2PmGnSApx5C78RF
8XhRF+PtK/j/PXkyGm76WRngjerSfCgJuW1EEpcH0SfVvsf0nfMcNyUOTODQJRjAI1zViSYwlUkk
OgME5Pne+Zw5xk2xroCWvW89Qhhrb9mPfaMEOX3RQpMAVIyc4hr747RaIyNHADIk79uKUmvrjxfi
zmz49llAUzEP2y28esLqsMdNV9bDD0iMGe/RGrc13g3pZuEkftn22T44+4EPkYKiJaIMNOTEeZvU
OhSuwlSsav8NPK6d3RPtXHhNmdGbT7BNQvkcP3aMcuPlYMpRSvgqrIS0DX1+lKVbOEra62tk0Dg7
FnPcbH2drzIUo918bV5BqP2V/cuOiXBxwtDSXwQgdBiwl5y3wkuUFk5G6BSeXSI49/mfTPJQL803
TudNEhOzac1GLB35qet+lvGHi+/4UWiaF7Cz3TCRt2uKywoFNXKBNthTd+dAQZ8OBrOhK+g1hwOY
Q5Q0n2dYXcwStc2MpyQ0gFLNZ7DfhnuHxGtpzFPDPwu5ygmXAGylA2PaAnvDldygE/+ylvgnFzs0
TH2wK4Rgacqv106GizLdib616EPPOeGXENmlcN42zLFbQapNDvRW2OQPLwLSqRKe7hiIpT/IiPEQ
Tt6dNDnnK4o4PoB6U75Qt/xbVAjQ47/Fip31QWVqdZCUs+MxTTlOqSv+Er0LSXA2v2wYmb/lIpep
22tbA+xZw5xJslimzqVZ1Azp1i66gHXXT+1XJpOojbQ02MbfvViytMZWsnVqbaPliAxBwP9vN36h
XAPOJXeAti4uOWrMGzjWDTffLLhODmiSzgrCMkxFmHMwm0u4DaWjtlNViovV/L2biyf9bERS8kku
wba/Ep4WyuzF27/cAIU1JSKI30xBHcicIUUDfTDYuRIvRYDf1VMDcXO2ePsPrRcLHKVs22Izz74p
tpRt8MU8BoYCZ+PC3Me3a3qYvaV0RRRKh6r5v2MwRaHUJjAfkBFQdvS5Mgw9PMBWJA5bnlkodjDt
y/P0KWZfmIGIwb4VnRMz9leTx8c9BKc3X0tpIkYcZT3QsTQgTo0JbMGPgQvF27JSbN6FhTJVOMDc
xaEZ/jjf4MsQwBOV/TkUq52Ev2hRiFR5ZY502ftWPZ7bHIziLevDgNwwIUc8olhqIg9zkNnwfMkP
2WbJiAwXcCIBQB2dxHheZpJtWZiIaKJyxLzZPIFb1b/jYnBG8HvqEGwyToW6O2tOp7VmkuaqWbiP
v6QC7qIgZmv9ef8Z4P7e6tKKKnIQKnUpLugEjkD59/tX07UKOraFXc8iuwj9r62jKgGLBFs6Y1Ns
lEJUTWVCVDJsfmLNM1GUPDJowv8ec1F32FzO3We3rZh6HV5sPWQBORW+MeNPrYHan62IedKdsMtW
HytpRrYu+uk+088burwmEXedCWp975ZfHM5Yk+PBIqYooottIbf8lCJH5pgwNb4JBGnfjqMpcrbf
qtuP2IB7aFsrJ+34daMTB+VmLxSB485HGWvDwHEn3i/CxmFKnjAoyS4Yjrvj4oGgw4g9MODgdSSG
ncQmqWe6KXTbguY9f/lIkDOFvn1Kmxk+JIc4x8A0VZf4qejug68SOOZLE/I7ZRR5RLACgqUkSsnN
/lL4xYmDh+Fqrgc0BV87yML/57X6j56emCfckTnM/0QWvMqkRkSPQVNPCCT70Q81V6LQqjgto4sX
KB0F4uA9NRxfQN+zZlP0J5+YWgcUsD1iUwyw+6FCVeLtDRDRiXvJ2QaU9jkv8iYBc1VuP75XXlPE
kcXUxX6PooqskWbeQ2tHnI2ARympb/54Gkk60B6Djo8Sf98ZgQjCwMaHvZHoSzkUQKAX7i1/Kj2G
Fi2Gk9RRwuXGjTqnAoPjYVQLLQA7/4auLr9X/B5zsda5FqjmScnOUgyIvjFZXjNc1k3HIFJ6C1L4
t1BZj4zeb8WlRnvLypYDWGUqigTRC9nafC33BoKlOs1AAbr8Ut2VQdmM5Pv5jNuWXh49SUOU9YXR
euqDYyndHyh9HNpFanf2/s58Nn79nNFGmvHhLV4OcYSwebHKACqtbuwTWn33UjRjBwxKYdO7SY0m
kIQMlMQ3en+GktLlgPaAT7/8Igpp76PeXdGYmsEDsEJhajhWZDOeAuaBhOABjMqd1cT9Ou3gllV8
pf+HltdPpz6bEfYZVay3qTYnNf2SY6iBz2xpkvFun+TIPiF4RjLFNMlU5vcvHmo2s4p1Zq5e9ACa
BK6h89nhNwbVhqKhFFfpUMHc7Gx+W72zRLucCXmNWGImV+Lnjeq7F7IyOVNP+iWQV0JqTiDcJMIu
X42/FcgjLbxPQku1B3zTS/Q9JhkFOqAyhlM4lfJ7n10LidEYto+jIANxatEatVAWgeVEipqiRDB8
Dkl0bD+oTHAZnuhgHSiEFeYCw/u3dC5mNEZh74u0XOrdk1n6leaTTjpgb+exg3aLt0fZkZoJ6ZrF
EV2JXbh3NS6ERtOfQt9Nkbmbw3z2OgyS8my7px8Ogq25YY16tieyUb3A3fStLZyxii68t3g17La6
fSW112KdQtaKa6oSX/qT5G1fFwf0OItm24yTVy7K6pR2usGhTYLdc91fQ9jMXtZ6HSrqoHo7WpOo
pSs5IxD/22SSD21G/Qkq2teePyzwZE0bu+AvNMJ8yl5i8rxTAHYEXTyvYAwy0H6LOwfR855Fu+ha
cPrvhKejhpDtvpFdyUPr8Q6rsmrZgmKkBc3czOoQ8zdIxqmelWvFv/MrMI6eMjNdcSqvgoMh4xSG
Vprt6QKgxZwJnfiaWtwvx1KM/aQSyWxjTz7G9x8Y/i7bwN3Q7BnqArwS9F+rLbbx3x+nrr21MFuF
1a8TnAxFkq+P0gvjr6EydZS/BwKcXFMz6mDFxQ58VoDPlEKK/TN69YJcZpOLwqY05eEf3MunXdBc
8yk/KEeeaVjdVvQIN7FMp6eYg6iA/PoZXh57lb2XapWfbUfz5SobrkvyRdnXt9xwvkWTWoRb15i2
oh/GieBnUsTn8ruDJorG441dn9oeWbCMoAb3efTYMqGh376N4alWXn7+RE4DK4dj70xrZKHqiCeX
OQ3sh5vHxOpJSPhWaZd2q3MH94ZEv+l8z9l1BvLzohnyChEmg6MNNjXiRlOAkOJn6rRbl2mzG9FA
riSJPFShkwddWvCADIDZc+pHXWJuvHo7JU3oZAv4bfJ3XV8S7CtrtZHoS28wd+h3563IHcPsKMz0
fxe4b8HKfGsfekq/jeKUUqQJNroBbu8zOZPWOgQZL0bVOZTudcdFX+ABKsqjZvnIeiPSHi7gGd1G
zni034lFYOg5ak5EJsn8MQfMrwGEakPsbUVy41tkdoxRyyw1vGlUTjyF6p/39EFs5s6mcwvSagtD
+Hi+uGzqbZXz/iHGaOXx32A80f549r0MjJt9ILXsFs0cgLelCEa/BnVRmCVsRzAX+U2eA9vu2Psp
G9RcWhz+ofxDDAq21aBUGuh15jTjOjjvsjy544T0gFBJgpV6C+SOjOMKCgvSBFXKp6oJrkNYF+Ql
fr9e7SOnor1xQFCjxrrdqd66UZXbRVhJ54Fj5QeqV/BQE6xxky+6EwFzSsgeWnwbB+umSWWPLve3
u1fbTMc9bpevvePOTGGXYiaJY7203a1wX2yXSHETJnqrbyh5cwPbcyQtWF0pKGR0dEJ0lGI5xIty
N7v4xVhLurepucnMOphZeHaSc+XyaSVLWaT3uAYE+mhQz/aIXJGc32pJDHrYs2BNaTkoXg69+V9Y
3spBWaZvLkuSN66yIIemQneObqYgWZmLTIOOFDi3z/JGK8KIUtDueTnLPdSpfm4zcGwaxFgTOKxe
/0cUXzEl2rb6tLutHWkJacJW/vmChRbCZrgN2R2U8NbC6thQkFYtQBp0X5fGSa98jTfGE2JPsPph
wtsHJ1Dw+jXyDIm30tkKnPMJjGfF32GHDAtT9cn805bFn8Y8+aK7K1DEUHX/14nlAiPxezuCI/NZ
cyjh5fluL2nnH30yv8RqxsCZlMxqf1dfzLJaBMdBbNHKp05BXNH0msRed60mYW9eFbwNDkBzqM5X
Ggfiwkw9cU95gtDuW8oazhZsAWZN4FQ9hLAgNLUJm68zbrlanQsFgfkjyG2rkZDHHWWcOwtG8ntK
zD9LX4qlS5Ts0nXl6dMtJqQfhlz63fwt4gTjS96AGjfJghWyu2mtRqwgs/Y+sLfNu/Dku4Cy9YDp
eTg31EMUnwqNVkfOpyYaXlhKSaC6xgEXLh9RQLPBYbvSd3eI2bKYaJjq6pAXI1c/cPcbbyk+7Y6c
D9Iso38sVugcIgk+CKaAfYLDH1YI9pO6160+Rr+yYV7ZdU0uySgmGoB1xIxr/F/NOVkZe1n77dtu
NGzLzfARwL1s6R25sqdm/r4K0P6RJgQccwUny4e7Psu9WtVuzVkdXTC6Rr6cHcxn0KSELQryhWik
H4uBfOz0QfMpCRk/KOIG2qkNwZJBLXXcfVl/v/36VbMXg2dlARys1c//mGlE3PcPrHFzMmFm8u3N
9Ka3VRilQeGdW3FCBdMLh6uCuT1T2jRugB7t82x/foGK3uNo3cN5SNS8tpj+ggaWGy7j/g2njV+g
ZpLdtFFQEdRXt3ZC+VsmmTGOorSMAqJZRimqCZiHKlCrWgszNGuMnwks8Mq9pte3/8JnvpwBWC+B
33QSdijcMcTNVu4rGUApnuAKE0Q6YVihtXf/BS6FaPd+7crgonPaUbC9ipaOfSzgCTPx9IoW2f0K
+vOoJs/E1JFk5XP/tXy+tlTCIAdbaU3P+xJA26lMHQXq+NP/VqL5LZXN21/r1VC0ql7Bz4M1Jtbe
5J9WgTNXORCJ2W+0ajl5k5MIyjvvL8XqS9xOn7I4+hDGgiLdOkB9WgatA5+oqkdr1kaVB6iL32yA
PpzFQnlAgmnD27jwpSCZDLGl5KlzK3/q2CnwKRNY0M05prebKkU/i+yth+0z9BrHuPYIi/N5B418
ZwO/RCD603kgHrJvcI0lo/+snOGnBtX+VDPPN0e1NYt8fv8+tkWTGyqEtI85aHMHLPRpTOZaVxoN
valHwqveD2fSMJ8pefrw4diD8b4wJNzHFJ3Wj+N1XyqlRs+cEa3Loiq6uFCAVyF+O/LOoVHJCYib
39Yj+DpLrbIX2SxwSe1Yq+iutozmQJzcwH0cVemANv4iwbSmhO3QGUsqqEfiKldCZXvGsbL6PrGy
ZNBBay3gzEHvP5OPaAGWpG37tOooHm6NBWbndZZ1jCFCdpXW7OGotHOvpYTotydSU7DY+miII8sT
XKAz+CkIjdVNy4Ax4jxFWU6CZk4U2LkoBY4tH8FKy/CciVOGX+PSzaaPUOWVzBFYHvWvDmecsDjr
+Rn7Mp5gPsMS27FhWBxeLkk9dTbPC1EVuA4G0gVUNr8rNHj5LjUS25M1Z4UqZ2FUgYkTVoVsa+rv
eKzAQVa344dUBJB1RZZ7H/uxzoynAt7Z7wT5NPl1v2qsveZuEN8dp+oFHdPzjrI/Frmr7buGVbOD
D4BLEjftBBgzdtNNztaFyROB+8dyzPBXysg4o7tonu9/Xki/sqqkyzjqNOa8WGvmDCvIzoyADMb4
V9+TKRSa4t+CbAwy3tkjonF2ozdi7strq4+xfIYdiuF9qQKTM1D6jhzlmAGwaoDPoM9C+etlF5+y
oDuNisPJQIzUu6825hEUTNJCO7LIfkxgZGgMA6gOYh7b2Ht4fa7AMPT77tCNRSb0gtFraikK+Tqn
PfuPo6+T+OnwRMHNlOh3LRRezycJ9PkB/QMBkPhN8U3labWzAGb5F/jtOJO9CtNTqGCN+maZWcDf
AVIW1P7MW/3Ndcpk/d9p/aqvhD++iCU1qMTh9cPY4K7izFv/FIPJWxYbR6cr6XKOVhxv4LFCpPKd
g5u9U1QZT2SMaYaKPH9sDQc3vBiJ7lAmTnT0r6ii+052B9NDUaecfIQ9UFTS782WiK6UEGZgLhub
36Inffb4GdeLkbriIJvJUVzlwbASLye5v/No7Wyu4w135+eaMFBh9dxVL1I3ecFCZUcqi3CXmKsN
AaBWfxv+PnHAHIir+kB+BoF8CHnGwFKnktYceBWw1uqCic9/Mb6zPFwMShoeaeSHOgF4cCqooC5p
lfZ7nuGWKkmnP5APC/CAynzzrKBZ4KKXdyLpqQ3ZoHSyhKafD1XUDwOapc81q56P6JQYpBlxX18N
s5c4uvkyyiaEoVlWIL5/NqP1OJPx9x4eJf4SLJy3NwE6X+jbU1NaZO0CN7pkVJaJG2zNmDbVPDYO
kH44bg7XtGleZd6pjOo7OSpzsAOoMrgx+b/EBZs8V3B1zvhIj9lvgbZbudFPFOyl3r+4vcPdi6pE
9Qa5m4fZsLsUtuBbxzO+ch1umJ8YPkdsjtq2RcTHDCOArElvxf939To1ZRS9H51u5hmrouSoDWjX
xPkyk/eXScz12Bw+eq+5UfdNzeNZg/wB+AT0s3rcR5p+6+ojFBPYhvZVLs6ChYOapL4YQdor6zAb
X0X/mPNaJ2f+WyhXAGLwAC7dPIsLPM4ru6tWEI2bFanSd3aBTK4g08UkTyz3N43Kib9LGHlHSSwU
JV58I4G8SqtyhtZjGZdxxiP1J+XPn01rv7Sa8fQEZeHOiON/iDS4GlQmynkhRb/EVuXWhjTJwKBp
cTDAsCEnXNKkhI0x8h3KvMZ+3phP7kW6vloc2jlriqvLHtHnV2wwQhhIRFGZCRKAudVfRJnCUeIO
V1XCEWxJmABGcg8308EOork3vG/rV9xjlkdujUqPFXerf8VXYVFUZgUbHpb9CM+lZ35cl53xbmRT
szEL8z30CxiesTThM3JeEr2XylEUs+avzkWyozwB83dpb45dHlXPkfhw8+LCPlmMpibFQ616h4HH
fafA3oNOpRrZSC0bupGl4Mpu29imBXeGZfdLNCU9OEcC6SqL/K43qnmU0iUKnxk3vNR9OrU0w6Oc
oI2QXhtNzDTjqrcYBTpMljw8Zg+CzhvmP7yCSQbn1EQOghWogr/VggqVc+LWAe3Ss7cjKDboEXEl
tcEJIJFSdq3qrix7ZeX28rlrP4v6QxQ4NlxxzQFexuYf+TkgZef1s7S47REj+B7yFdO4WEyZb8pv
hqZq9wjrWKbYkG2nbo8UP+o+ERrUTfulXW2naxI0wXB+C28VFiKpc8NXr94sYHVcRn/tteJdlCz6
ER5ZNVJHIjbxibX65fuq5OiIHSbq8vayuPYv5bl2ht3Mc0mdJq93N0vuZ4YtmhDJnjTFkWZbdAXy
ra4HbRFZRGxC4Lso54ywA+3h3b/WmVfRAE0qoGzrsp/KTb3+kzOFw+a9PBZ9kAKLqd7qzDPKngKF
NJHKWwI36g7ODZCU8fEx1TKwGwmpvg/dPAKieTWG2MtmW67u7qjpmXXgc6nYkYv6rlFPQ/793i2A
z3FnnmKw0D8WG7uE0yhoM6mbq11XBul9b/FunPjpntFaAshouR/zOz9arJJlLaTPuLrdawE94fBj
by4UBde9UYTFdJgxKDB0+LMNM29ZnNyMpxNh2CA7KF8c25WEq+FnOXx1/sjzRvhzfIAxzFpHybT7
Cs/2tUf4ML7CDyS9jZhwXsyuUEbCRIeLwQzIWbepW/vIy55hEGMXA16+1kksyeSqDtM2KJFD3KoT
28R2rvxN3yPmh7DXMjzlJdqtuEqnvanMn1ovGnaaeP5RXNDPZei+CMHFI/GMtHoMMcSheXbAQbGH
ffrpnGkV0/nVTklPB2e0hhiEmucAoD9HOfm3NJDqIX7Gxch/iV90W7avFytLFOvPY4QqWyb/fvZN
7C1J5WaLnaFABdTmE+bt1Tjl1l9JFjFgjUvG8SZyePQA+fNm11c5rQcziUxQ+RuNLyLKzaj3BLgq
qt9c3VZJb8ufdGNP5ayMo6vUx4ZFqvaHlCz6V4ObQNDwq4+dVUwM3PpN+BwJplYax7iffZJkk6iW
weyYWTKAJ2IINzmIpDZEGnXM6cfzlfQBdHYFqzTgRQuoJ+Xws4PZR1SrwwaUhp9/o22S9nlPS7RC
mi3UGKnIdYIeM3jpg2TEDteBd/+/TNtMoVVBhC3FuweR1s0NW+1NCJJIx3grpuyn8ic5KISP65Fm
Cgl+fWnOavBuIW41vhykQvHbUyTikjQM5drceJxRTgw1TO/4bL+oNDraOhd4vbF+nBCAgUtcFuEC
2DGP7zpvvU4OBEWs6jY8NlOTOVy83L0ECS9DWe2pDwNHe1Ti+wtqK5IZ8l9523N/VyvfF18Ddupy
G3tXhcVXMYljFSVHO79UDr85eTKKzcw09aWhulMO9UEJuHnuf2Rq64syhpFfi2ivnS5Rku7S/jl/
yDmxsLNmdO+xRtnNUu3LVZYuMOdA+ulnnWEoPJrrqJoI9eMf0pV8G/WlN4AvmPlXMb9nCZGp4lmJ
XKS//3ZX9ifjxQ5BmbVdgv5dkqqXnDawOLz8K1/bytVAM2VHmbHY/r5jnC/n9nYT6xYKwHkGdvdH
04SCOofUKhEqn9XaKP+VCKkck935C5hCgvgqA6xiQc0gX7gw5tsSoT4Gk1hZzCbn1o/Q3sTii70u
HkkS2TR4f9U0JkShMWIf9ThS51ruTU3/riPsJmjJUxdFFjm6d+tqtEK76XSwPvyrGKD7LkClXe1M
e/lCwTgDHWtsafhZrKt6uyjHjkkRILrGa0Xj6Une+87owT0qOz/3E043rXGJ5wxYwDs+IYcaLvWM
Z63s9M7KcxGSEI3nvCInBYBN0u+ivZf9uPTe8z5RUv+Gphh+9HoE6kGmKbjQ8+G7P4LCwsac8gwL
mPryhXYxut1L+bS47dfc0UVFilUjabvYSsTqg/+VUuyqgqq3SP1S4KA1RoMJw8D2tSML4rXVlwtA
PjuYXcU7eG5Gv36vKXyDFLYhmrpFWObFSbDoCJEBeB7UGIR2WR24wLoWKOZycdIBYDsCokYbn1n7
ZmrwHq7c4IEv+o0XY3QMcN20GYeMcxW35SYxiP+eQHzq8obwYAXxTBzgHNZt1fD2iMVYrLmvwZ8U
uHQU+hmdSuKBmhY7ZPNbdB/EndUZ19FRUtIb1KFBWng/CCLLx8OSO6WJicOhZBHK4+Rvvx9SXHH6
8Jmyq0ovWiyWIimS34aCyI+QevDdaehlZKF9f9jdPmgkUeFKga8FEZCuGfEQxaElooi2wNi4pZ2O
5fZ3jYSd8FcQ9L7rjcvpzxW0ZQQ05sUekqgnGhcIihoYqohPNFye6yBGwqj8gvIsc8OoxyTustPi
lz1kupZTklRNg7FePrHNyOOfhusxiqM2c5Xb/hTAAP+sFpVk5JPi1W+4xFWAm8XiWlf8TH0lY6G/
RtPQWF9mfnDqdjnf609OoGucrSCxwn8VNYMDauKe8YjI8woF+yxzR3l8LAZGYgRONPjIZt4HMUW2
gtD/klWWCStgEfPesgfRkuQ9VBQXs4AjPHpP3eGLoCJfDdp5c9cxSobLr/bVauB66UiQDlrjS8Sq
Khdotd3FsvXUew4lJvplKNi4M5a6UWzNtCjJDNq2FgCJ8FU9PRsZwrq8HHDxBZbPgOyunX70+KMC
NJSiYBUZBwRCMecm665g0pFfzbcTLFb9mVSBqcj4X6VFVetJP0BG1/niLDNW/bwsrgtspbF85agr
e+1BYTkqly0c4AvsYOBCXEAs0MDWyypq5gcrn9YID4L0v0liRdwsbrPV60EjINjopz9x9GSqAXAE
YXqFCpCeQP8P7TG/jKL3GSSC/PLANiwC6EVsD/RXK0/BXd7kNIsfYoko7/ILoNmwcLpAPo6asjGz
Yh+PLX566eICYODiu32ra3zQqXb+YMiNZ5FxvdFpQyCiMB+VMsV9PlC95+XT7hezReAKm5aYwS3Q
tDzzqMHxyDQNhU39ix3Cb+lpta4Ilr1KyuxMTuRtbkvD1J9bq5eKYI3V2wOsZgZtq64kFIS8voBx
muAyMSDgxZD43F8cVKnua5pqbzRK7OfHOmdy7ihLTu6zpK2YWLXTAm84j9PIdDUTGYwdPoQyh9pm
6t8/eHmz8mhRdFcD/tWvuIB0SF6ioI3Fw9HTUWi/CqLglpMc6HEUs4eOZozh9GH5L4YaLiwYWPvK
duVrxpPQYWefebQdmrhLI3UkFTxuwDQ3knKwjPfroo80z2rT1aqepdKVh7ndxUcGkBwMVozOnJtd
QH5cfkmCTE1NjNykBtzoAslq6wSRcoNgr7Gp8t8lCYOFMz8Wyrofv9nURkjudDtkFw/roZ816Tlz
NODJE/Zwqn6n8XRfX3/1uM8OXO49uT4ZAPQpSvBLv91tAAPUJdWxj/rS/aM0yHCDqThcBlrvvteS
YKHk02qaMjdRrTcpdfmhGttJnfIIc7RdLEnqFlrymHilvvcsDVqDPVcmDb+T2lGzzMWQHNputmbp
u3+mjA+MWuvbIC46b8qGvT2FNdkLybUfpMlW4aGJGKMFS+fnlLEInGhhHum6o9QspmJWn9bG2oiH
JHb6T79qUqJR5h/too6OaK5Wxc95lwGuDMtmDliXO3RmHv14jN9ahKpn8vvPlDRJlArNKKME1+8y
3DCkdRt9toojAedxSKLwLIYNtMxfjvbCA276v/FqC2XpiKzYnqvR59FOsyP0BTk3MavvR2Qt19ec
kqOkuf5pqmkF21REP4BbFnHjfXAKz72DXYOWU7SDjgPwdvIa0/3ed7eNs5fPVQhCvPV8x+8hsFzM
Dyd1urd4LbdAJQF/XgrygdyHwMTVSBC7Hqc9MdF0G0r3H/w6vfj3e/xJ3S841wIGQWUwztmhn5z6
zAD69UiLEyhBX6yQQg3DJDM4GRjb02gEjMhLUa9obV41q32CNcRhHuIZo5veLcCC+5xstV5c+/Aw
Bzlzsp2S53M5y7fQ9uYudt0rmZ9bAPa7gYg9XUFoiB4KODfoqlIJ4HhdDx8SO2rOYpAz7kdAwO02
dl6xThwYAXyGrhpugIOy8ZYXZT7rlokisIya4g6wQvqowU9AeMZZUzUcwgD7PW3/sEFvV7gkioT1
ZkMIhiKntT7W7W/dvPMAQ3N8Vt/6E7Wf+KF/1/QcE/smR90w+1gEcgmjqnr2+qOddSoFi/wovPmJ
oVflKR4M24F9Hz9VCgZG0lM20GluM+m7PxguMyTx5otuS8IE2kBwkJvStDWHnN4WiMnKlSbjAY8b
qBsp/5qXFskzZE0NiOVIEmc/A8MOrzrGcf+9H249wC3h6Nc6/Dfd+SJ523T2jsNV69g5JtvR+rFk
HdePMn5UbgYg1vIcJk6T2uxJ4T5u669U+8TxqRV2w4yOABLCv5zxEBIz1q3B/TZ8B9YwCyRoql9n
j2VZ4G6/enx4tFJ/i9pn9K3RqZIvJdP8zf/hm7doSH1QehBYyYRJLXTZ3YvaFdhPc8I0TxTSgVEJ
2ZAL9K5a51hrCFMbYSMIAGTS7MmtOu+9DrNoE9lDaXHnJCJbXMzvsr7y97nFnfHUdqTEsshVTwiL
rOOC9RkihHNsSUGlKtyxuL42aTh6ApQBEzKOIeTKvicpwLrCKI40Wk8hU1nh2wupGDwcWLmHiG1P
oup1Xs1X9KBx1M/jkT9RVr0S3hvSJfA2VklGdMrv9X5C4y7IBCBeG0Sw82eU//9zvmrhvOJYVJVe
fX0VbPXs3+/3JI82xMgrGEViMyUYd6gtbv4akIVyOS5Qie9HJseX2Jv34m0OSw7+vmwGjvEoZPCO
yHMHjwj29tEee92b+SokcOF8Gt0izO1rT/OWlSguJ4FGGMCu152OlYmJLwTftpzOSOsfzAGOq7Zj
R6pyrP69yWeZq8kBEsdXkFondYkiMCiR55k+x6/1vYuHE6OXsEOYsNnbGQvum/9u0FbpcLlTRJva
2w5/tB/9G7iF14CTgMKoG3OAksU2+pz37jlwYZ3fX7zUSQJuCyL/0/XL8cqdsBSbDLuq0Ir9SFqe
/v6wmKerfQf3TSbKUbNWqPjSAemA7ERH7lgyK2baje6UGeTs2wWk7OeyUJGG1l7hut4h/6/cphgO
asXsDut6QkbA1Po5fOHj0cSjn+k53MhHOsa4I5FKCA7Lf+UbAimBqZVVo3hs35MaYH+bZ7kFdtmn
nGHrtSmlNVmDvigVxzOa7gLEHtzNAuItwI2i0NLp+DugENlmBS3/gxQDCH/xjhdVjjP6gtn5/MsN
44RoAsKdO9TJuhmpQBT8XYx42GYI3Shw256dc0NrXdDoCthlr5c8NQoNcbqlYDjwu8nBVNoiEiWa
gMuMtay/fmSsYtAYCFH5RIF2YRq2GtIBUbjQvUZCZDtqA11etFSgZhHilTC20cJGowBSGSU8RXXZ
cFXQT+RJntBj3nAkxIYYJLj6tKoY527KRie+ODm39+3L2YQwPdDw5O7cxzYkfMuQNvLH5AOnTl2H
sEM5G8NfZAiFstphgjY6W5OsBaQGqwDfpYt4R83NiksI6d0YbFp953+m4ru+1kdspHVVxnGHePk8
heBfApNEck/QKohwnC0aOGkFMH93z31gl60HHvn1fSJhtT7V+1uETOEOLq6KJiRZntgbetZ68BQk
7XqzEDNGU9dDrIVFEAHmMaMUQf5xfnwsH/9V3ZDI0pjCT707Cq7r1cgbdiTyY05YsEz1q9RdErOv
Y1hYPGys3RXbDuOFEf9SCExTKs54lgRf1kJCPARC+P/lnARFny4dyBt/xQP+rqzTJuusO3i+i9m+
obuK5HB8XOw92hV1uXx7DFiyAGg7X0AUuPLKR+o0FSCRJcWz9nqqcpxSkdGqTNPkB37dnh3fu1c5
CT1xv882IC4TMrIaXFmabOqn2Wcs3VMgEBs8dxqr5JFDawfkiG3O6QVJAeYOqylXQ9PYHTup8o5V
UU6ckcYAPH2uT/ccrQHqPwMPGnLoe3bTifM491auP3YJrcSD80MEW1wgH5JpUo5u5QAivmSjyuUy
JpgnDPKJAaXm9jIqtSGNAPzvdIMFvNo13KF4mQQuhKmtTChaKK5zpp7ZLxwUOSfdywGXBbYvTSlg
OTuiFnUMiWlW9Pa4AMCHi9w1uC6pmZ5U+Mw4USuIWxvk2oP+9Dj5Q2e820zWmWEqJCsfw6yIcjCx
LE3qkfxnz90o33BOYpXLf+YASR+7Fd/3nkgo58YWVPpQkgG6n3f2XQfA5eJkU7vbOhidcHGMic/b
K/vhlqm5dsY37L6yiZUyFygbjQnYYHzhXE0w2JAZbAOxJBzqXPNjKpEfJldWUMvFEjb0LDqbgVr7
WKVvLZbBKsvw3laoCxdysQ1APJlpByn41UvmMKKTMgK2NL+CFKjf4WPshVl09RX+oY+IeqDcc3xt
xQ668pm+ImiwLYxKfQaU56do7mrbbYZ4gqZ7HnFc7n1wkdL6VRDuuWGHXqP1gQDkJKNkLL0s2Go+
2nyUDdeAhLNs2K1FH3BWCMCShglMd/s4OL3l4wwUM0hnfyOLflPLJQ/P9grYCht5/j697d27rc/a
7i76ITRRdNAYdknG0XFLYuLg/iGapET7heYg12SbLi2NOQsJs0SGL8+nFJ4OTBWuuPKHGJxSl7FR
/BUwf71RY0AKX6jGCfzFLq+HWt9PKssGu2dw+0R/N/1Qs77RhT4dr/c7EZFC+seU+duUtPjwq0NS
P2JMG4oF4cNxB6s8o1kcwbfA8jRc2/BhRJ3x5VLIvYHX4hV5PhpYQ+PY77IlWDTIQ/C5FjmnIFYz
wdFjVXHW9+XdedLCBSbcDHWmleBnfvphdpcJLz4NoBBbjKRET+iSlco3RQ5HXxsXMiir+jwLMXe2
WIg0NGK9OJ35k5IR6lUA7ciCAxVx398V13bDhFTlTPfyGLlPE9KzVB+RNWiHIDF2UDTN8j/Dcm0i
DDYGncdHnjn/6XRBp/szW1cCps7mTcpzxq01pczwEZ8ArG1a2KdFLL87X41ovWil1aK226iyHPm7
t8Pw/YLX3lOWRCaTOFfTqU4iCrAVE/PxwgkBLXdKdopE2As/kS1FfcqYp9NNKvCbwN3FRPJHmqoC
E69lrUtxccRtCxYnFueK+yqeunDvMP+1X4XqfHLSyIECXllhJSXWUDDDYij41uX9uKRVUME8pbVH
WvVp+o4fnwlM4b79QCxiFbNfMhChgL8t9tRQhMr7gww+twPxZMcbi4oFwnDSO+SX3pZhIyTHWrcp
4IztgF3L9HbN1P6G1ENV+PGfR99kVBQLoLvW/EBeoR7cgThqkkSyyp2wnDxCpw/4XrjRY3vvy4pJ
ggoAGwZNFYXjExYZnxzi+u9KzKBvtCA2sObWhkbqBjB9L480IHQFC79OLyZysz4Q3k5aBw/EOqB6
spYcuP+taptD6/+DZdHURLAe0FvdwqFu8sW6ha6FKvc0w/5Izqas0cEBdXcAw/YEBgrlNMDcqtB9
ST7T/NjWKtju4lI6m85u8w8MU82B2MDGnQ22J6BxJCXiJdr23e9drqnGrhrzrPkUJqnnwpIdQ9WY
tLJBo+Ef+pRFykC5Fi5sZIqOwmQETV9LJEaU2RRwy5FEa66UDRr12F33kLFjViD+nsrjvUkHsXz6
xa9YrOJTQXy14gGhGhD8hm4j9YQkECBRSnF5FwnwgqPg1kDZgYd2YhYwzQUpAY48cK4liJOwU7QV
rHVSofhkM1SLLhRsW+eDnGXxDU22nulIZcp5ImegRTPY61DguoLrgEU58yMG4d11DDvRcuUkpCh6
2fMbv+FEHCcn1AyCBCEDNF5UGPeU7VDraZeEKlUxxPhJQeXi7NaD2psgZReHJvHOSqTSKDPDM8Gz
/Af+0avN5a1+/dOR0x2hqYer73UQOvd+lQJDOifpe7wGKFth1Fx+4HjMf6+nghRYw0++DU5qNFhz
w7tCVyqRM/r6RQ0qRFva6OTIxmzHD+22Sekm7tuLsarjRidm6ONRAJKruVLTRqiTh9krPmptN/cK
yYYil6Sp+yWBSabJMXNdIIFCK9dYM9BLsT1sgpPDueArOVEtcwJNBwkP5XZOVJyZ/mLKpjvfFBjq
UPTk0R4zCHYslf6/x/86TPkq7b6oFAX4RloCqZR1/AqtGUunMHSb9deBWcKpAgy4J1sxH47iNmrB
FJj36/RK9HOK00XJyChPRoYN3jfAI3IbyD/rpcij1GOfB3MxaYyGxThHQFBqd+oNQoV+Av4GDpQL
/JW7Fm/I8V/YvWhi9i9rPJMM9NdpwPFLtfUnNm+OX7vPb2v7PbuIvsAGdozOaum7Ba+qcCTjc0xx
2XAmz+XZCR6BfgU8ye+xYzPcDPShThRxrEwwbUorUWAV6eSpsgL04Auoz2+rb9UfeZI5MMeQTf4A
pn30+ReTq3OMCau45YN8h6mIdaXRL8Xv03/ww0JRk49uuwsElQXAJRIzYmcBuvWtfrVU3etgcnxD
H0702IOG1PXTf/k7vX8QrrS7SVmNPxg7Z5LIJTOI9zqfZlFvti5/B3lX8rrRLQ6K1Af1mzKfEsLZ
SOe2eSJQjWCPY/T9tT/OTAZEzsX5SYVvnzLDKkQ49AJIFbqUcD2Y2OuC/MOt9/5ARNSnigaO86Fs
x2YPxcjiNmTmbWLF86YV2gkTXw/QJ+X1RizNn3nRofBJS+h4n/QJqHepPqYDfr7Y4IoWTdRmbnMT
zCrKZLiLv6Nhf7Uk9KNnHWtJxzIMwK1od3X/f8gbPiBqIqKbKZ3DC43oY55No2b30RY9oojhwGvv
mfkq9x1kNApq4jkO4vcnK2qJ0iCS1BNhCgNbab00YCAhe2RyPaSLc55u9MjIpITqFXjqTzO4jK8o
NgH/YeoXqYU2F9TGQAzwC5nQBdRs+a1amjYt3twgM5ssaxN2edl4YiYp6Cx7IQciYWfY9NYzMDhQ
kqyInaDuELsa7ivI+hT0Qc0B3zsrO/Ti9xEJPi260tj78d/7WqafcRBhrLJeE7C//CeAJOCjJULG
iS3I0tihsoQK93BVB7PvV2NuTNgOQqFtD3T9oRQGSxmLGd9Je8IQK5PHxoSLNg+YtbRhFwVw3/f7
0RAeasZtgLqQ1i13+TOsPc+Wt9lXP14c3C9vHJ2XEj4uPdGNh/sBNkYmtBDO7IN2DB6KK7O7FLP2
KeKk1PqN50c+HH8hCKkAluWwJXz8yTem6Jr5RwGfhX1gPDZFKiNSr9Nlw/+bRUFwMgftKozgO9GB
IybWTgrhurWlC4wHbjneie+VF1SJXNc+lMhGjS+cE8fEdnd/X8jqorrKUI/EdQtW+IueGBZO2ohJ
YoUtaq4VEmpT0LJ/T7ksctb9joN89UaOMOsa/3RDFoJxGbtr63SCEF4pCgX2z5hrKR2ATacVBPDb
6JhPhlFLMSUWDBMRV17bEwq4XAk0RuXyH7oAriqWTSRQTD8/a1fHqCz2JqrZS0isz1aPm5PvT7th
8xoxDedV0ik9CQjpykDhZtC+/Vv2rRo1gFV5aR79vFfsDEGvLAu54z0ujJ3v8B9xR4pOunxqrRoN
lLZZjLkcqnt4LGi0cvCPkbwRGsjFT/y6ElLKEbBC01D21j6Nq5ALs2bpMovX4Kt31i0Xb1znYSMz
dMIXCh/Pw/HQNF/ViT24md0VhM5e4QaSuDXaUE86/hl9mi0zjCMf28/bCrdMk0aawz8xbfJSYoQ5
X7/yto8rLoues2+AiiB/fY4zuEa8rj365J5LYyZyuB9MDCBEHmshm16e3MlCU7j9HLUDcrEZIVHf
6x1UC34oqT8nqi8vyqNtA/BX0R34qp+aelakWRuNbug4uY4uoB0A4BpXWNKjR+n5bYVv6dzGAl9W
051WM3TWRbobN0lBjKNYmZw3fN9E99rQ7jTTTr8pFkM8uybmZ64NnAxAlMGg6WxoYS4ilAFvBOSn
YC6T8lP5JmlTeRVcq1Vu/TdJBql2PcnymopvzOZ4au8dYFWo/YCZWqCWcJ0oDNivZ9OD3XIXUoxA
7ZJJsRutgD/DyZ8fEa20r4EXbBsth6uJ09E5C3glTZaM0WqPzwLJ+o2BImbjShehaQ0qJPwq586i
XfGnttqnTjdUUgYN+ISHxGWXa+6PrB5ERXLefX5DNDo8Oq8TRzL9MbwKYsXrYCPADKE33zpgZRre
qB8Y6V3YT2IkLx9Vg62xkXnYcwoslTw9Icxy0202sWATJazK+9+ABJT/4JAt4/ktFRsoph08FoIe
ZYhhnGrQk79nixfgBvj6/a7vcGK/FhRASF6psk7V1o2nad193JfJo35k39ZREOwlpBY9XWDxOLvO
jrUltHcVAYcmdzwuhoqnrUaLiPW1IYImT1VQUidqOk2gwEPCfRAszlrDoe+/J5wEYYtLAgwSeQle
05BM6n/YNBQcAFXvHhJvOTwABAVQKB4A0krXArK95+dGUzFBXen8csjRWIO+qqythX/oKyube+Ub
gi3xRQyarQ62TePIr29kWRH8Loz+3etQWlrj3nxXOrgrIilUNb3JDcs0HMk62P0ORr+2X8qC9CKC
plheiASVwueZLEu74Kw0MBzFJzhmqhkxP3Xmk9cYTmDN3/C79jB4MlFVZ7jpnIF+6hmPUU//uC40
ufKABPDxVUn0Vc6g8rEG6DzNTNeggmAlCfGjf4javx/wjHtbLmdg0qSHsPHDRoQHXpE4g61AcKzb
e1GbovDe8snXjPGtBYsspowaeV6sQCeKdnPHhHKZkDh7hMqo4rjB4ZPBTly/+UParOlbZ57Cj4Z0
Ouy6DumZ/l23Jnm4WEfjrhFgd4TWFolZ5fbZSAipwb0pFHZQNMhBYGUy5azXw2g+FUECD7jBUhIw
kJHWqjxbIhLrZNrS5Lu48BrQxNZP02HOCRJlWlFdFqqYfBYt7e/t+eQ3AdNcCt73560v2D3zEVAP
g8rqrrZwbNv9pA7qWPbh7LsbWOq5jPYm8kMGmwvRxhz/TJW8j2at43KdaabPGwq8Q31J31RtDinX
Me94wh5tGKL7B9N7qupdTh45QeTP/6/hCou2OAugpq4YEC3SI9F79hs7vDGEv9EK7Xmy0ny7o+ej
4gjdBsiVaNKQwNQm2tVLr66f7kzi+xuxrvNDnQ09zXFzloP8gvRyG1oIBujf429ILZeG1H6OAcPw
eIMrGMeRUCrbyMUVeJ5spXEi8rsZ8nk327Wp5yirq/Q6P9F5784R8Pe5wtgOC8IsrPyfA8hIgfZ0
FFV8tlkLea25PTz3jgOQJnwrfE3j55WzKqJUk6FmyGANMmOAjkwC62HK/LBle4JXibqQhC5NVz0W
rtDV8ALIfjy71uHffF86MqIQLJSLzB2Z5SVIfhRotFIUQhuECJq28ea7aPZ4d6GZDOYY7C8FISXx
/UVA2Oxa3MPATOEWOucmCZkaQLbx1YHJrkxRPT9PIetRfRgBkmHY6uHGxQPlRlG83mzCxa6uDr/P
o4i3ipFtVHrhza6BtEbdkLPxXQXjy6reA/rLU4JL0K3SKSHP0qLRTtE5pz1QAx3IYFm+qReO1AN0
JFm2se0uYCebPagoSfZJSMwn+ORL3guTSZ70DAggpnc9dIJi+cDufUpKuuKt2EeV+4sfO9L3tEmQ
aDC6fTVgFjQWQ3WNkb2JZYeiNIbtzUsutXzVZLO2XyydAcU5ArzOXKVU1nDl2TxSMQAfh/tsEQ3m
ujtBF66rYVgvc7b9GC/G50iMnU9wJDTS8d4KbP9er4UCnBLPEFc+H/HmS7sktnBZjWQ0/cznPxzF
4jQMbQ7Hs9hJqPTLT55zYhOAUz3BaomICwIQEQuDQj1e45q+DJjDqpUBzWGoK/jMi+jhLPTfgKm5
iwM+8tlU+BeKd+JwDImqzTMNunA7L6w3Ru/9Bg6ZIb7eLCujyj/sIl9N3osYh9dYk81gBVC4jfRp
9s7mIwkZI5VKD/jtXE227NrjJEQ2OXxGQiQ2oDgrJv42hJ1uFsSD2ea3JNmgaYXftilc9Dujv5X9
dAfCdmPok6fvLeqzYHhil6wyae7MC/xI45q1PJKdbZfFH3wa0RWmqnI8MnCdvkNTa1OoqamqJjz7
kZIiETia2YxtDLbcqB+OG1EzqarWlJBLccm1AXqwf0j4RKxg41o4VP1hgwN3q+NrN5OcS5NaDaD+
eV+/zdp5WbJ1Q4WTMBhAYhT/AhsCZslDCQw11touYhnxQabrRCP6PjWavyUsERpRVNUKPI9X6Hg6
KJYzuml9tlCFnUqna3sT6eIDWb40eUigUxV2v/tQZxhIrRbvqHHFzaqcaxvaa/5MUH9zDzOJeq+0
6n5coU/o0BWFRGUoCL2PgLzIt2b71BIetu57fCDRrHXvgzdLGaaUYFXhcX7n38LF+AQIvP6sPNrz
9eK3ESaJDdBu5V6fLfD99cOcaD2uSMbQ956MDJhQ54nxsap+sQK6Z/EP3bsUgMLHXEprF9+QNrFl
ZA4yTB+aE98+OziHjDCtZwt2VNZOKvzk5yNgJLzzwOpmFCeXT7fmeXN3nFyxyrHbC3VXAvzxLR+0
xXTjcFleMkF48+q1aW/DAYuoBQE0yITfqGhAPH/xCWwjbDu6CFpDla4LOIKLRocjPCTuV6rQ6Sq4
9TdFLUpAvR8MupEpWf1KQ4KlXuG9knAz4uVI+cYCbFdvR0FbdVXioXcp0cH1j3bJZAdqOqRKtzqY
DAcbFP5VZ4OdLXoW16FnR37eeg6inJtLFf45dbTVBPPlt0OjPHjLSy5uQL2mmcP6wA8WYQGOUlGy
JSYAZ767FlOsCmqFxIN8ni0abhYw5EYoFBawfP+t4stw9FKDJWbA/mchHHVFc8Td2YymcdubOHi+
jM5WViwouoe70EGmiqtSsuAlF0SWWODdRqJCK54T2PQ3FulYsycZEFM9iLLXQtijLg2Sdsb/ku+e
+0GoHtcm73+GrxfFdB4Q1DCYeLCzaPME1nbSCSOAPRd/DJe8sozg3hJSEdY3M+2cJL0rrD3gJeXE
6Dpge3mcuEks+0wsxog7aI2y11V9An94DFtuZoKGepiiTfT6s8Hphny/HVhxqWeL8C9fnc8yvB9D
fPCUJV0UyIVR//TZD7DWBS9ZsspR6GaM0HG3IrVB9OkWyvZvxaMRnQRBohfUOh/9Ra9ikO4oH5L9
S9tHEqoFTjpB9NIDYfECe+abxl3SZZOIfvSbxo3qscg2GcwZkq0gy80Nv54pCm2rSiv4V6oplX9L
tsG0FYLaTIkUdVAyQzsTI5/lVTciySPC256ljQEvnChlZDsiO5wYP7HoIMWyqUg9YsMDRrnNzQ6Q
LTWcbq+NGG24nz1UZSEF218WiTNkGLBaBQMhrwYK2qIN9am+X84fOZTOEj6aAffjRR/feRdXonF9
qO3qTsxxBgyYjneZl/d/K154lG4z4KRWTaSLuGq6nhGqraye4P5UHPnVcdp+tWaHChXK3HvOq3D9
BpeyhFGp+FCKI38Yu1YYJEbnEXrzVKFPvcIXtXGFTLhNUxjPk2Mj71u6aPEELzxZLPXuKM3ONb1T
/9CG/J4rzVX1t/6p24crcA8Y6c7Ph/gNFSg0jBol5SS2biojGPpK3W33BXJSJCQgPv8R46/29DPQ
Rw16Qaa9TZyu/uLdV1O5F/fzpzmVR/7V3lYs2qbSnvUWGSVvYe3SiJuRfFxhguLFYMn33FR1Rxf2
13ZDyql/iQN1eavUNfJlEFZ9AYd36z4CFTnXocunfLCblEOWuz3pfwtXb2IWhQoPslfsntfUipgd
JWyIyupUPSwipCxRRDl2Fm21lHe4L5o+nJeFNatpXNZyuCmOCgkmH7hdSsscraDS8eXeJfjfqxph
h5N5hyNkmgdhlAVmVvOZXs1hvRdiL+iWqWlAt9te0dSjup0jAfFV8k9SJkfLrV2LJauza8uHaOz6
0JhDWMLgVb+n/4InNxne8a5DLVGCE4W2BIKbG/Vm9rBkDHpwwpuNVnKUPkRl0Qkhm1DJPrlAguYD
jNLNzQgn1CAWtjt+qEQhHL0ZHAvZDThgZ+WdhW1OB2dlskWubbVosIPLJvaROpQpgaHCqryjLaf6
3WhOlBySEDx14gNW2C79GykpJdDDkVjDSdgQysKImAvRRz7yNFYpaRzkIQVYq1ZZ0RAzsZaoAVxY
n3yuYFHndB6KxbXBZfA62d2jUc2XkKnH6c29OmlrAu0yqudDGRA3nIksNqXcSjRgMK5qVfjiXjzO
VCoCXkH6hujFMUbPzLq0uYD2FRW6K7ZTpdpzgWT4mO7mKJuNt1EoPXMXJiIQDscLT6xoqE9JtBFm
EsKd4TSisFL14kxU6M32ZAD6LTYgV4yUjvtY6SuiJqYJF4Yo+ZNKGa89RCln1dvpCiMhgLAvDS5P
tL9iB2MDURJb8MvD1ekOa/UicaWqm+2fnPsU9oLyaaGopFJXsCW/RXtigDvsFLz3UaMVIeILSc3u
lsOFFfe06m3F19NamF4p1vJflst7tZCQCDiN8KmBmNiHXxiMYQdVS9OT6a/CuymOvvt/qHTPI6iG
Yh0ahR+SII9D936+IkIqt3GD2vMk4/9oiT9j8RzbtMzilzU8JXVc4JylawV5ovqol7aie4P2dPgz
7rvIt8bikUe9epDHT5GL2zXdJmX0DgnNrS0Q2ziNXLiEDP39mrrR0bTudgybIkDLLPZRoZAJL1rC
SXaXnFKD9k4SVU5JBgAxGGw9gxq4h85D8IOsPQ5ZyNcq40T+xAzBid58OK0eRgG+GKcrsixZVAl4
6gWsQTEQOwWzz0SQMjHh8BAkw0JwN4kGhYj4jcot4dvmdAWcip2QSG834LNfPY+Ilj4I3fgd/cgy
/OPP14isXJ1DZ9/FsyO4sLz6q+/aQD/yLMH5Jj1LDvqX3TXQjdou21V2+rPnC4gnwNY7Pfq+zN4r
P+LLGnOS69/Qrj97NP12hCEVnON2D+MWnG7qJ4OIpoFnS7EWDe+UUGmi62csoM3ctb+tDZQJU3je
pmNu+Z9rYyHsx+BLCpoyO+y4w0H1O8JftaH0X0A6KglUwIxY1vKOoUenyM8ZhJ6HdQKuEKY0vdEU
MTIrEuDuGL1ehvD5/hgpWwg9pT/0hNUfkpwj869Hkr9k9C9jkOpa93bDrm/yRRv0ZmEH9/Wfx3t7
rVCXmew1lke7AjZAVRI6ZNVxO/OIvscVJaFFTBCoeWkO17JSIQTVSi1dDo3Lmbqidrzl8I2Dy5IH
6o6OhCsep7Uh9bQ4pavlN1LbD8Dd/nCZBVb6S6s2V14VaU+zwdGnf3gWDsewvUkwBsypXX5oBELp
0PCvG3A90zylWmqOEdxvDJ4EwlkvFGCrKAhBlW5OG/X3EB3wDhUalkR+hqeTaTt3exQLmlhSU1Qe
bGifo9Q8698v9TmGV0sHyUM78ZOipD9leMGvc73+53csriKnup6WW/xOwke7ikSz7vayAQGEMxmA
PHhqtHSqatBVSLsgTSCKyBsjbbEbqibBFAaDZPv9EnQxu5AM0syvj735wmilvuUlikMFM1ZGkiEk
9R5s86dZF1E1iXj9/bnzaetuLgrTWDySMZBYfs2bEfelTfLD2bXz1hTAqHQp6hdJ2mi8X3FVGXGj
mYhc5LvaKOJhCV1J7Loqgok6b1GwotYSXFtt+kjXgItthJdo8kEvMnzWgpQeFqOUqPIDPPdKkUOW
l9+nLDz6s0HieNVPmyffsULHiGg1++QCGd+JJws0Vvst9WVApczfGUEKaOYwKCsVFAQKg82ZeZkj
2GAEkZ80dnhwaMniZIdXiVpEbGs+YDKQXFLlHmreG2/CXoUuJFX/VKbNGVflSEH1msVreMwBoBKn
q5OXnYKcvQQ0kPyQt3OCtPuxzs+QgIFjq/zfRVNGI7NHPSYQB+i9myYkXQmN3OxPUVoCc3uE8aFA
eSwzi2fSZQz3p6A2tgG8cY0vLI+jujcI8qoLXy2BMf3VzhPB9ViPmh54Dyflub1Kb3hxM27nhOjW
tKXC4LesC0Rxd7eod6uS3Fgj3jIOrmaRnDJUNofQ9O3msbZV4g8oRB6rok00eC6QlXCWuM7FpyYz
z8OIU40gj4nEku6WgxI3R6Rv9xmoVXYOi/rCVmjImmg3BtSk90VZNozfEuqBE6/0j0bkYu/e3y9Y
VVrj3vIguSbC9pXAlm/IqmqOp9g+zoVWz48Bj8OureWDjMZCLXD2iCe7yU6VU9PURrvDlBd8Ggw/
s79l/QQGIr80lJLTWW5cnSuyRlLAgrY7/3DE5vypMOdUfO4jr1ohI53QxnS6sMmXcDckPxI7NfEV
oysKlhf3ao1WhlVNklHZHejS1dZBCzr93YzdGLSqnyE/ziGN0CfTvnwHj2O/+MSlcYQokkzYn7ds
ZwJBHPK+cZFXClTMImnCp6Xaz+QlV/xjPB8p9HtHlovJQJ0yO2CMljuYHQsBhzdHBIC1NMx59Y91
tIxA+28H6LDtAnUXZJcWo4bpHCeFEQeUrRQ59QJnYXzUlX+3GniqOdXRdBZZWSWZcx7nSlqdOJpu
w1/0Ou04dveTWGhljlrBG2Jz1CzECdEFzC0+qjmClQ9vr8F2ESKUnbbz4V3hPijqm8ork805qZJe
gfF1PwXmwt27sgHCp+rZcTxgsvTX9VB7KnNDutj772lzR4J4nZnJS7xMoqZFYi90T+B4+7oeoPIM
VcLAcwvolL9TiObcyRBPbIvYMKQX6Swu8P3vRMVH+DxWtP+825SgH7X1dSMxRIhrxizsNfSMUgXT
hc169w/ZtHQooIm1RuWioWiXtaGsf08jRuzaKoPlmNVZwe1te1LJSbivFIXk7s/y+facchD8nCUa
lelkxIOt88VsD4KgqWy7v+IBIi15ZXh6p16NZpZrkdt12zG6sxhVeeinNMBBIsTMcOzL42bMkY9V
5okVrS8h7lPD3NXL6AXM3O6i6PHOnFKi3N+Qar7UNlj7QW8Ut4l6T6T03OIy6L/YoxrY0YOLPukG
o8tip4k0slN4+fBxEVNeDy3Pqn69wY+h+jJsJw2PsC8cN9f4bPfsKsVz+sphPYd5x+94kuA65EOz
CwNZoRx5BB1e8NdMhQS4vhk6eOG1cZ2b438ae7+QYro5nZ4knVR0159A4IOxjj1Vv1vfmL8GBPcO
L6rH5iRJY8JyL5z/I8ErfxBvbVM6x3Q5dOanGV7iWy+fLUbJg4ZYTMTkMu/cCpexQfx+nm1HLIHA
j6ep29MU+nFTd28VIMKiLi5uCuY7389A0u8aCSP6zQg/6ODnlA5n0c3jbGl3AJkfVFzMN4bA9QUy
LCZD3qKRlAM24GmbLhHQc9gMQmQ/ANJc9apq5M+6nWksw/k2ByKN3lLbUz2Br+IbUQb/+cW12scq
WvzmwxYBS3Swha1TwooGSYXz2KKH+RMzXr+a3x24sW/wIWlpjhh5jt7M0FWxvrqOD6iJJBegYpH+
9qrgirqS6IyLVh8jv3VDUXq2V5XCLnvUBSsS/aL0LZPlBRHqmnwaWiGndGfTcv5AmUYO+hNJOzpe
OfUoVoJvurgHzYORlcO38UD9P5F+PccD6Uzz4EcwC8UqieMwqoqGjfJ+zhoYVilCgVFQGEHKU8Hh
rvbvvYHD+N0uPp9gPtXONbscEz01pEIg3wKtjsWpZZJuVSOvoXR3BhKN5y/MrRYZUv1NPzTnAPk6
awXWBNs5cQh86PV1eHNXA8dTxkKZSRvAgXdbiyPm5aS7YhVjHDv3iCVOzoPMazRjPQaemL5ak3Mw
69tqxFq3RX0+04fbmBX+j8g4QQLZSWI7xq3S7KVI//COTAOdgPZ7lJI5FiYDzGUSYXrY1c40r7nQ
t5SC5D0WpDDPb59xoOGBLJe+dmXlR7gEG1qdP2JBEgRJ3tbJ5z6/sS4v5JvTtf5u/pGdFfFt7GZg
R31Cq8Yoq4O65KkdtdowROa3UZl3T0Ty9bnRV9NaqQfOngcmuEtS5jrf+/VRCwqVCHe45szgnChM
o70u3j5wkVWHh9p7sTt7KB+ZgToBJdLsGDIuMt7z52Hg+d/ROBhDLzNaKyzpZ0nNBNG3FCo3Zhcg
Z5j4NeSBFtHoJxkMaqmAGrLG/pHupY0QC0Y/iSarZGn4bEVgQ+Hl7L8nbLFVOR8S1BOk00Y5/mfh
zRcOumfBM9XJdgYR3Xs4zsgRRzqcDddrMpT9yvjglx//vIAeyyfPzyLTftQJHvhV4XJtJj2GChzf
9u78YSxMkNa0X48n5njKCsKXbbbgkYX0Xa3Z2xytLOPWszI+tTX75SJ+dR5JHlhpwh8bDPobvMS/
CdgcKWYk27MPIdU/aBAf/XaNcg26j+7F2EzWb7K7MmbuVxNYIe9307kXsTlVIlyr3OFdFSR0VGQN
audmMj7XTaE08AoE3I+u0lHforJmobPXNUU39O3v6WJ98SztTs1r+DPOmA7U3KdhNhWAHXPj8E0h
YtRSjlVP2Mr8CEAOWpIZul9egaBQiLfK27salIVZqLdcNziJmTqDqaNGbqkEIsdFcf3rl6E6M0YT
keBW+D/YY7Dt8ZtfsCAx5ZTOg8L/K70n74zTfWB/5a1RJRtSpCrg
`protect end_protected
