`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S3wuAQVf0c6ewTjhunBLGDWe3c8uav9LYhciZ8trhISeFDgFrV0eX6oQV18TUKLPoujiF2ZUTq/B
UFhz7cB6ew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BEPJFXuExFJxxlXdzpJQE2Xiim7Humfjq54CS7NYTa7d2kYdwTptTGBwYxkABeG2Pxmqz0FXmPRo
U2aVyJqLdz49llbAxquNDjw1vwKjkr+pRKD4hSmTq4xdT0ZetYil2gRbaiquoc4ZrOQbIHgmKlpT
G0tj5GxgJD3O8NSVsjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXRD6Ywo8NDNXFhH/k26ToCsbFXBAW4kpIyxdfgioF3tiAOAaK6s39dK9YZiChZOut1kwxLDXW9d
StHAqZQaJBAYREZKhcTGuOvygECctoIqfoEYgMaIavURDe16tZ7f10LQnqmOdzkF5Rn3XJJX19by
ty9mYWmINjxAKFIGTEGydFApjI++ewgDl0rMQ/KM3pQJmBvRj4vKhiEnh+gFBVHxy6ny4BRzAAVO
e+33G4qJUEb7Q9FaCBfwbeWVCr6epc2x1/CTGSgdxZ3c3nHPiTpNXx4HaTmZ58pJEdz4adNPUedW
Uu4JjEU/+JEBbwtAhGPX3dy2DdO+aHV8Tg+xIg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JvCzHYOTM8rQKapKnyISF4GqpH2zgU0EanTk/PD5MWwGW3oAN52QOFjNz9dzBiBv73AyCeGHpAn0
PLyq67DcY1ESq0iOR7JBVlzpc5R1ldmUcqVcSviprAaAoFU4q0zmmcd/zt25Pco1scQE51gVSY5F
EoTN1F6VI7Oo32rPWdo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rIFqjA79EIE7C5luYZpPzZADzj5c2UGGCKXia1Az9C8oN+8wkUkOR1XNYKZKo9oMckNk1Me4Sd7p
45Hm3OHYdHaqC5r9MDoi/mAsX2O8w1DHFsOKaWT56IUVcQyBTAiH+pjx0hk6A9bSTh0naR4N8m9d
CrWeZKabfO68CLxfBHmq6bPi2DhgtBacVGjB8+rS8c2j2zcTau+Te930e+mPXmU4p3NCxo+bKoMO
NkpCx04zGb3e3SOwCjQQOH2pVxxVgzYbLi5dngof1aNKhJcNUzlkk720VjWDbkZgPGS7sdSE8/u3
nLw5pJdZti+D3MDDpb6fHgz0mEFCf685Be968A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62880)
`protect data_block
0eB40Voek3XE4QOCP93RnfOevygMkOlWp4qDGT43GoBRWVFG0GUihH/E7CvXCZVwlI9ksA0HQEf4
XkNK0jopDU51DeHPUZGR2Wm1+jR3kAziMNHpntJpglYAtfZFhcT/aDAzpJ6kkkYsCrstGU1Uf/Y3
LeD+qw2K3LM++tksXDWlRgF/znF+Jw9c2JQAPXKM9TKRvOl/czmCOhE3aNSoCh1FUwlKG7QK7XW5
1i+Y/6fuS/CW01hotPrez34/+2hYr87se6GBDorysLqVAXMsLY/YV9B7HhDUSw8jyNyknIEmI3U7
WudHo8vhLWlCkMQkDcMf+Ivoy8TEGZRjbwDtOXoE24Tpyh0y7Szqp8vQqEDariMqKoVn6oTmJYLq
2DpWhIEswln6tRI/+zBSleCqwfAdmXyYA/Icw782kOJqC1rm3rVrW/fPVK8K9QJVLjxlLtCOUsdW
MXHfW8zBcf+OJ6M5Ps5WfxcGaSo9F93JhZJwtp16qQc943Z5uL5S7F6uhx2/2/JNEiZKR4nwO6YF
9lApKneiqiV4lMknv2GfPf3Z0yt/epCJ1D6rwzHUxOS1WE+QGHCe4rtK8iJJPU8gdqWBAV0E38zX
DrRSC8OcTDpaHRsM4h45UtUZ7QHuncOnjyjfle45UXlGJHuJmqtQtKoBHlkWLaWs8IxPTRJdashu
kUk0S37b7qinz8QPzVNDizIo7tt1mrqBCLYTAlFjqwSpg+Q2GoQNpEbhhjJSmvYKPuGddRJZO7Wl
OSphxyLgZzVvmxDSH/t87kHgGHsFgjp9dviohojl/U/zWNmgRey6ALjcz02ZkQE6vzh/zBsU36oI
1XLzZdPOsmsFTW+hi0YtW4QXrws+XJn0lDvqAm7a/4zSUan/YXPqgWJAp0UJnu6AAEQbDjLTTbka
rmLtzTc+KBM7Qh/MrR0nLXOt+vB6+4vpyFW6VF57FxmXcsdwTMv34b7IGNAHXV19xTd61xcwO0FS
hYiDkPuuZYyI4HEIp4JXLUgW5zvyHVNvmOFASRRNUBRiTkDYHnHp7Z/O4tBKX1n17fF6v/fg3mwS
2JeiK4If3PXvktkxXJaPGyiZmPmt5A4Bthy7HLbet//JHNLV38xyJ74gKq7QU9oEASiPXGEAhbM/
x9I7SkQ7MIJFc8uqyxac3MnFNurIiDEeYdHyaMERPao3PN6xhb/2oFOdOfTFP1ukLGNEUsk0hPd1
LgkUtfW5A20Gbm2UqEhuCsZlhhN713pRuj/0GuH8RmIBQvAjd/LXyOWfuP01wImCTKOjz7332xEc
vYTB2ZLyx0dZNiESt3YthzquQ30BRv2JZ/yMS2L3RICN8EY6volLZIQ9J/ZWNZnto43SN9PZ1A4d
KcVhHcitoNxEjWlorIlUHZeWcgjrKzRKTms/5Qvq+XK9VFq4xnGh7Oac9iup4UOYCOq/mhqKA4j2
JlpoYNdiV2q/qk1GYiR9lF2o5Ecimhm4F6Qr/f/9tQ8wUUD6qfkiHSEpOGq0Z+43W/6hQ3pmdtRH
CP6CKYahbYpyAC5P664kR3KSyU3BSn/mcTnKBa/6NWGyfV/dwudwQZYVTSGWPphViyNhg4NXBZdW
VpNjfiNyjHV/WD/NL12VW2Cc1vUJznM7Ohc7WOPoxL3rTVqMbdkgPi1PL7rVXfy3t8gZU9LEOkRW
PzJtI3ekd0GtH6hpTLnCd4KmXpUwUPsqehrqFsbkKH7YNuki4EFBpsExEHrPqDWOzpH/kcA6Kdrc
YH3a3yqe7rPGOTbbq8kMXtkWN+YItZVlgy9BxRaEYkXkPwPE5k9IeceOrVP1c98Iv+echFZLGGt9
j0QBJm/V8zqFl/WSHqF+eE2suXsp689eqNMH9JYhg2llYDoxhhS7WHFNPfDyoEWMj1/FlOG8ECsl
8hbPn81Rxh9ZGPDmnWU1rLYxp70uYzLoDW9knjjlU7YCZd0swAJvYRhXsXf3VpO1kz3iv6W+nZMX
Brg1+/LfOSXBphl/YIzzMLzLBGrPVYuVX6U60QduJlfeyJj/jsupLa0YCq10Y7+A2WSQXESFHfnp
Oo1bNau5NhQE2DlB0tGBKT9+EPIslfIrUiX61m6Dkfx7lrqNHGsqror8LWJv4D6YsANdMsKop3y8
ywyUOABWxCDeC4c0Mvj7ZXbQ7mSXzmcBcrunwbWP74A7PloqWvI7iteJV7lKc7ctjR9u2w96DihV
W/DwvdUVHlOVlxCx01PJRop9W1LKbTZpY/0ZzTe7UocPsy/89bc9AcwM4aV8BP8oa3Tq0MJrZOMO
mP8yNtdJbBItrltMSYPKOFrGF8h5Z9v2p0WPw/sstYnkE2z48Rw+6hSemnVMd0wzek9T/E1AS1oE
ZrA3f8QL4jIonmJyBqQNSc2KVR9ezwV6djyk6MGEmqbDiHCADFai9EZ365ggEep82nSHyOwH7e7k
WAk5TUhv+Z/kHNdp52dLfVakxOtEHSbneCdm8hkeGJ7HytHDkfG0EsgZqwM5A1W/2scrmPjhfeMq
Z5gZil+FLHuqDgpnlqk6GwlHJoOLR6TnOa32UQ4VybJP9TMmBagp/su2C8/eaMBKHBuRVk39v7FX
8dhO0ZLg26Y43Dp/r3gPiA1p/bUv+HokNtQflnLHrnfgcNwAFuo4ChGQr1suF+/6MEZ39+YYcLQX
aZIHry63MB6k2POVKN1jUp6i5HvsZkxmE+SYqfeSDdTzqzoy3kdlF3NsS9UON2EiPWysa2Qu1opo
tMApEFghS37Yp1yaPg80jFeZRC2laiYChE9ZVjVUsteBxyUf277ypkGtcghPr72TPqQ1zQtbODEV
01nBZ4KzeBhaYwC0n8+Xh271Ug+NcvgaVLmitcZexDBHRfooei8SXKptlrX0Oj+5f74mAi29Jmga
Yl+J4Ze7y68N+bzIJgr5GmTFfbhcQWOQtM+BOeiDagj3eW0qeSPaLziyW5Otu/hbEIob2UQETk1p
onrFt1MwZK1hw3fcZGOjClWT219Jhfuyy3lsb9z/1Y0t7kkhyoXH0NKDKRuDurkJ0bKhY+0GCyGQ
H38L1GYASu7gN5ku/Zk7VkFeHIldz1l6oisOIKm7UGg0hicb5B93f2Pf12QemWqxMQgJ63mSrLMV
boU5NveNGoLsYDtDnaV2YNF+CNcyA/sJMBZrLAgN/9Y9uAUXs3U4HPLd5x0+voXUhAbX4JvYJBIt
lCVF1LiQZRVoZ0CoPFcTPy0oqZf5t/B0waoz6o3QOXzVHLjS+SJmInj4IqzXOmBxM6t77U7iJ0L8
DqPYSIzZg6xsFDs91WviLUP4T311QrZ5LerwdtK3Hk+uLWzb0bPkHyvvFAYOd0NOT/j2UcC1GbM3
1i/7nsYc4o5C04OSProKpPCFZ95VD9tiWD/bMYTA4fStiKgpG/mNKps4FVKJyEpUpF/F9lMeHK5h
VhhcrPozoTummlVlNe9Vvj9dPIQsA1gxnvLW9t4VkxX//GhFrj2GBmLS3o34UxMZaED8vODd+il6
qDmoKi0uKhKDjY+vHeO9zVnGAuhOFFJjgbT9M8pnz1DBrbNcZrdIigRY5CkGFdDO34KRb1mBDfZc
8SlwXW59J3UVLzm27HqCLovEuLH0Fub7d+4UsIbqTnRafX66FSgrUvoVswLPQcTNtqLWVgwvv93x
VlNoALu/dhBlcXrdEQSafLhZo/CYe5UdXYzo3890nosYIQlXck4n8Bp6bTGyaNGVHdskkhocokKq
Jf3zXj73pTosZkJTHQjBPPRAj/QRiNrRsKIyHLdkB4oiSkSg1P57tgzIPJ2P8FDCoEuy743RykFN
iMPj7w91PZJyw/0FAimVUpapCaduTHAb/6ku6PVq31f4bN+VgX7cdQF44ydABJHM5eaEBolM+0BN
ON8y7T+IJ/pjO8E2X+0c21BJZSx3v+qXosjCuIZi7yf4af+iTGreMQ7n0QlaL5R1k1QRVhNt/2En
oaD1qq9+mQ0By+bASF+1FfwJ4+Q6+xJHp+TYCE6AVyUcDh5DFwI7o+alR23741zPLwnnNcOPxoD6
HeaPDBWyT9Mg4rOjgUyIiiEMeC/awOci63aJQ5wviwMVtI8TuIBKN6s6vnNvQrkm963Ap/5zWHqO
5VTUM0pZFY1sk9SwX7GhihXC/g9cigdGLl4j2Afn1RjQ9Cr7jqS6EaYpOVhaW487XImYOz5KXKf7
MTIRKvt89GpH5/OkCXRbpGSVWHqKPbxxNEroYHWrKdu1SFk0qBsKXJxUKUMajD/uSN1AgDu5+vF7
vqL4Qmoe16JgtgxpkOzVDXLLX3oh7vkeUcXdo7e9Ao9YCUu5sL8xOIisKGBXaeLxm54HURlBn7Qx
tW8+v11vZ4lqTnB7xMl8kMF+A4oXgVHR8OrCfaMCudzlYGHm47fMuZ67NFkU5bbxXrWHtzOcJKQs
Eag41SzqZw8wIh56dzh4oeAMKy7mwieQ+K0jgupihxV07IqN3fczIEP6V65etleBIEyv5tyw5ZPI
Qun3em27EFqqhmWuIZhmPM2qGdzZEL8jPrkDxnPwfifbHwUy7/oon8E7RwYbMhBv3q3P98bV2bbY
8oyBx8IigugsUlobHJN9LLoMBJn90kyDFaNu/Vc4IuR9L/K6eajDzzbwNGeGjaH16HMjtoezKN7m
+6VQM6qkJnQNDcvDDu3vzNA8QiZOpgEbxgsLNvrEEDouuu+ljgA4iejiFmj/6TzodPQw8v3+OI+1
N2vWyjKmGt3ezZN/1Fb1rSQRXuZGY38lSXSVJPxQ94iphR6AI2Yi1Rgr9HInvAcGROeX7aMgbwZD
D/eCfXXE+ERF6n/NHpFy2z0f4zpQi2YWwcYPb2he1SHQC66MWSPlrhY+GqJyPzLvuuDPAf/OYXZ6
AON/+Z5dN+Wr6QmaC/8AxMz3uiNCQLPh635RZuSgHSeyt/F3ZT98JrjVPPugXm8JBia6BiNv/q/y
PWAIOUPm3EwetwMbdW/lOGEHM4wsr7Uj85qGHPbHywWL0Tk2ovRRh800OVUdfrADg4S8ZS5q6DY5
vivTU3RKqhBIRkb7hcsy3FfFNYPk/OoDnHddHtwnxlq0J+uwPbSpdEZN2mOUvHwlPp7npW2TKEHZ
HspTzjqG+51QhxymXX0JhFF+znYkNO4dh4GNJpVLyAaD8lJ45njyhMqMdh+97847VbQD4OogQeuM
KUAcfQj9I2Da/wIpQmztHn+PHELIuNuv/zH83dBAUInUsTct6aYA1Ghd46T02Uu24qgBcUZyitDY
mq6E/xIimU64X4hHo5w8RYiTsGoRjTlmPpIfkrDagBtIixlRLgZdZrevFrOA46bjl9Z/uIJ1gVtw
BH1LkHG9ODgQ1Mh69V9PnNqMyLXxK8uMUfPKUoAax8lOPaNwuxgQ2IGQGM5BlGVAyP5pdKKVl+Q7
F5u5HGpawjP47ZmiR/G85NYPc35Oh7nxGRHMr2bcGmDmuv1MlKaRKosOrg+wXIfiXsjbDOHxgQYX
AbK+jRFNAgwkvESpwAIazTVVsqwmI/0V3iBi2bJmy4CHNsa/JWSO4HytVbTDrlOLlFCQt+JnoKpw
yJ4H1RCcH49V5nvgCW2zMBOi9lw2uByhUgHnvWSwPp8GeVjCXA4RRotjtMlsoyV1LULmUxWWuSnw
zQoEnr+GksNmGGDENA3OMn6OqT5TRSinxxwGklsvYSW+qy6NWkqLF0w87qgBQZnF/+0oy86/Oty7
v3I3XwsaRtQRKJ0tDAXpowY9EWkv5EDBmsovW06cMJB0KqOCgMR8ZDRyOmbhk0qF6QpW87E0XTkP
lcJYB+a1jPzzc/0QQnp0UOePk8H4A/uQMEedXZLdV4ALViwRyP23C+aNDr1r3IZN77nQ3dULsBBV
gE+DUR2pYzluPXeeaMkkKVx9Hfn2neU5RPCKcd0kmqrdy3KquR016HVb7yKJISgWYnqqcoEtLRZg
TsziKFE/seSVVI+H3seMs7UIwHFGB1cw/8/E6ufsdZqPMhai3JJeZwaKgF4TRY1lZQGw478ZFPX+
+zS5zpn5BI3jmw65ewQA3r8k+xLD0T6jRH7vdJSQ2z+MRoOyme4sNsOvPdp587jMLzG3zeBdbEYo
B33exuZ/pK/qTKMPwo38YIpZEP2FqUG7oebVBgT5LYYUW9wuc0MtgP1PAKLNd2iwAnqXmxsCMRH7
yuTwvq4gPzdkCfJwCaNw6nHvdun93Gh12nrlyE1OnFxO/k2fLeBtnnYTi/ylNWUpWQrDeqLh7SOC
SyVg/wfREChT8BHG8xVRYBE3rvzQ9ajb8qKOBUl0Eu5RsoB1kYLkB2JmevfcWOeiaiR5nf0Vppid
iMxliuupSo+Ukt39pHw1zMTX0MqqLP6ZlUKcVVu55pZjZl0ynHXaa02+yd824WJy1Le5AhM/87J8
EqArAvboolVDxzcsnWg+dyDKVWMmgQmyLz8NUzpiWMhO1BvyjDbj6YXv8fDJDu1DvkDQbsn3bNpj
bVVyWqbqER/sree2VmcPyaxaeHUibN0GGYF1Um4uiEqF9q6cdl7QDGD7SDpdd/40M0dStPP85FF7
7qKSG+GvByoHp7aaUcdGxKAABXx4x/474HDEnrRtFvxOfRsKv87z/5VS7sz0a9nudPafGWhmL/JF
RuBfeHHn+OhXCctMdlR1ONyBVe/VSGIvNzNAx7Ryls6t8vr9zyWsw0A9e1A8QRjepGdckpI3ysiH
jDiliwH/M9mFwMxeZ7mIv/MjXX5RFiORr6fYh0myoNYmmytzE4O881XB1FI2J46H3qpb2o9z4zoG
xgy7emO7hQ8NhnZaw3XOFchyAeiJQI+BLe4IAeYyiYM7S4ClkekIrHE1pGvywDRe2Zr4JvMgGGt2
8v0eL+scCkZ9xWGSKp4vNCEZmjvjoNa5ggSFM0AgxjCXv77uKNDss7WFkPVKkVtZIpc+4rHc2rvU
0AFIae7hKwFZK9ioeeThjcZzTFxpZ4njw6C0dZpI24mqBUo69moX/4KfKTfO8YEIG2VqeChitZ4J
WnvNS2LdjW7A6l8ciW36BgHs7CNWUOdx5Jv2uxpxQtexxhwXwUWNAjexDOCO2AuoKt3hzPa/HJQo
VHTeKp1Vro3PvG86SoLxZEVMdjCmVnQMz5ST03Lm/VqAxbnWWCaqAwufA00/zup4t+jjPddBCFMD
UbA8lH9soN1jCQe0U1sfjnEj+C+Ng+YggssP9NWNdKXbsp/uyVDVBXBlJeSZd/MMBR60H0VewV6t
X0tpgzDeVFDufzW3KJC3R9Kswt3CoXicXtcWUxasjAShwMqtGyIQdTZpaqTHV/OFF7cz/aSJ5xyf
VV/Vavn6tKqpvcA7NwEnnSQDX9sw2i7mAp/bfnnG73Ib2H8pzylIdHuRO1jhAXkLYFrwqummADE6
ZLPInrqlIfviJP7XwVVACyYWJJGvj9LsIa0/RaoJAXHdjZP6YlQJ3g7AYQu1zlYnh3T8ZyOF+7xV
sh7+xjz7BvzWumSgi6UbDlh+lhdOAea5qq0L6onK1/kqKoOujXVkaO58pBW691jhWLL5Zp94vBmw
F3VlcQ/hXyJNJtFtTcq744YPBmdbFh7QJHN8ovSSAQHBT03v6YVeZIa2nQ30Pi0dGNbZTapDN+7t
hfB+MWnu7K90Kg3+9lZbmSNGv+MRQMl7SvCT7gKbAI4KEqyBz7a3AYQ/Uk2opl+v5WUjWzTe1zFl
82r3g0r+GeT8JKffZTsV7BSRW4sEFBb1MPNGzab8V2rzkVbIl/U7vwEy8RQfP/8eicKYvsOitdiB
6BGLg/6aNSJwMBbORGahimnt0PDh3i7izJpkvxyJiz+iS7TafsyqZDCycXAC2w9oOxQk43bmLm+N
XETBgvXGwQqDyBQ5Ido0RxCfESaWaPetZjzvDpZjPm9trVnq8T6ksE/1DVw6HYuhSqU/Wq0NxoTP
XC8WQxAosDUGnOn8tdpmnP+aeYwxMY8zxiySrFnPSTZ8GyBYIORJ1hRW2o+xCxI5+yFh+NOxsCGy
XWYrB9pNKKva5d8ULV/JXubxPUhIlTnGsNjfuarmJojKcAcZzHQH2NxcKO9OYMwLyEa3v+8zXBij
HWmoR8hAqZs/LYnnQAz2wK7A0zysT18PRpfD17Y0tPG88TX11Zf3mo6XRMVf17VcIlAVVIp0M91a
/AwtwlzQLHDVTQN0RvAH7vAxYV8sV2UTnP8glWut0YqKxbIC8kWEybjBJtXqnKBhl4fcMuz8UOx0
cLH5Rc1hf4w5CqjW3gkgpEP+Jxf78VBO/9MfCNpYPuaf6NAPXyj54vB8/K3723XlJAmyvVu7d5TA
3Jp6SrbZiKUG2sRDtfnrD1keVFcLinAC6ty4KD0652TxWA91cqJIAalYFbpEW0XP3SehEFfxvb17
jA+BuDSxHPAt/WuHStuzRtXaLIB228+sgX8tF1w7KCgX6HRHMTPqmnBesNbmWTS95n5p+Jv7T0vp
gaqkILEdd0J83gX/hGzUqe8kP9NNlwowRcylHSIPDwX2GKU3CAfbP48lvsxJMuX6i7oKP2mFWsiq
X1vaCZol3IqV9GYPUiDinQKpHVpJ4LTdmKEwj4cLyrp53R7uZH3XBgaT5vko9je2w53H9A6tMBUa
mFiuKWb0ArXX7/Wh2Afl9vQ4Akhxid8aOVSm1wy4XeWm3WdDRPfmVBqD/N84jkentCa87y98XXao
rcpYvMFgy5adIzpg80N7APvSwWzmbZAyLkI1HB8I+RAc8qoFx9Bn2pvkA9WCDArWWPVcMvP3QuT6
V/sKm5anje2FH/anpwSFk7zMdQysdO9NEezr20nfELgnSNmC+4sHGRevh6Kta4sRKghFeNtwHehX
mQBRGusNEuORIOxDMfAo3BSaNwM4U7MmNv5UIPc/eM8xl9W2c+2rBDWC2W2VkUSEO2vUuf/q6ixJ
GWoEKWkSsVFF7f9BEkhpOWAENi4GlwTk2AMUl7m8+NTm4+V/os/1jYfsOyL95e5kOGEYQtbq9Z82
3fVTTc5vOuJiA4FeMCkkKEQfWed9PRYU1mLqaaugDTnpryNAAY0LlTnoJ/WcV/sGUQG9HSEhE5Rj
O9C91an9TwyeSuIz5jxb9SMYB3ikHSgAkCYDCvFfCKzlUnuCr6SU6jgtUYUCX6VzGNIiFifv52Jh
LWmt7MY72AqUkHBiWR5K4+OFtt1jVtjQLLw3BvDYrhqGVc9uxe7MBZ7CLf5cDqvC7Vv4H2UDIpzE
i244BtrpYwxQ2Y8F0YykJvCSO1RDrJn/YYaCwlJbVui+GQdQzW3akuST+oLsRSIh8yjB8/qXE6nx
dkXwYgK7dvEv6TFdB9GQW7osvNATs4tuLSRMpz7tfn55pATIoyvGoy1B+FDVaMFVpsngCnS5szsv
U3JUYasHFQQ+xlT1j2VchQpee65C260nX5/QjMImgD8fNc32ip7KCXviSWc+Dwuv/nIK87MXjGGZ
R8hPYdBj7nnRsZXUQqumrXs0cS6dUwwcQt1E2dhyJR0z69VwDjy5n9zf+WyU6NMF9O0PVRk6TP6o
vLtz+XvpeAMggqBBB7snSd2UFgBas61N21ZJXFegA1HDRsAMaTQgXwIrRsqh8pgDvaEbWGto47ia
11C48PRcru1PfD07+quIzVBNIRsezQMR+DDGvLOaoV/AEAlTU7aSGQ9ogaq3ZF9iyaID1uB6WXPr
f8k1p5XLhqryFmb5I/dNdEY5iTE49Fgdy9hCBGI1WCTK8w0JfLKMs1+gJCz/LuVLJlrBfpsPN4WD
8KT2JsbikY0OfGzsgdKj3/LX6Obbqe6aWyEfVxqpwTs2wlF88Lv+Y/fzFLphv4NpiJEFU6uaI9Cn
ntQiyOIm9JjpBfVDlpC2/1L5hp6s+5D+c/nyZIlU1g0/gBEIPcAhD03iq81C8pRQpwgwTzIBdf5m
z/4GuIdPI5o1ZCIleohKcq/bPpBD3sIqmeamsZbL5F+qGddnxnNDfwgsKDPD8mzK5fmm7vS0PXTS
elFzfvt8S+w+l1vs7ThmIT5bbQvtXGDfDD2KYfLCuA5lnkrf5laPhzk9B/rlj7cNtU/d9rpY2aIe
Ee1vCaqyiQrInSATAWU6VQe1ACQj/HADcgFMTvhKiGCYxPVpqbIKiiPoKG4sOBIOlQu/hQivd7iN
nLQbIw5XBJzkUEcedo/8WJNCUNJHQBjrfXh/q+Dmx3BKwReLoP1z4kKh/GBr/HmzCYZkETzHmHQd
mdxWTyxgSo2sGS0/3BGhigZd7FfyfsahS7Ot9WtmyewlpQOI420/kl0vWrdEGmvu6jFah2B3fE72
daLk3uX5KWXgkeLeIGAph+kkoNBUP+nS4qnDhz5cD5h0uKkoc37IcMkqenvG2tFWnGFeqm1qxqr0
ov/vMJ/ckPQc70aI3PCS6m2xCv8XiPPqoFkxp3nqy/t2nAqSS24Lgg/tGyAiqydDtFRFa+4Q/v+T
kov89uJYU9MADW74UkGk7CqriqnZVKdgYtryDFX0SchZD4ZDh4wWZtPgMW3aOGTIOCmr3r/vDpaj
NhB7WBdPnY5nkPncO13MRhqfirO8axCoa6ud2oMCUx5xqlMKYOFXNLfKriOt5tWBWJH8QpgU7Ubg
hvq2nt7xaLwK3Z8MB/gHiUs34iZXHpoZDpPtizuzlA3+cKOJqyac9aLa9TIgjrqK++v9uFGB7vE8
/Vh59sPaE/EgOtlgXg87pdSj2yj5RCPu/QMePV6UYOQIwBOP1niFtlPi5e5XToLXLouJq8zQmk96
QvoAvuStrQm9118+1fw07vZWg9v23OCXi0AiNAJ4mfGvOi/7HvhNPG8KuyJQG7Tep9TEs9CGBx6v
sylc0y7zpVUVJHVj6fEJ04M2KCJqO6k1P+aUQCYAm6NBv/3myGtOoXaH9YXEaO36OZ52p8xaZAJH
3p17/OUpKboOBsOiXofhKtK+uRHb7vpyvdyzTO3QBgr4EmvFKTQKGEP7nvnb4ZLaexSm/EVkX9g0
DjyMCUKlkhfnXovv98oaGLAEpapJCeVFDmPtXt4ibvA481PU4rd/GYBnhjhEJdigINVSQ1p0Bcn+
Bn6uRNvNmOYXAt/cZQzhaqEJRBYcK/GLcV3uztULla1tUCZlbXTDMxBlHFwRyuOxcEA8UgzVGKuY
vJnl3+5QKKOLN3Ku6APUtE36eHVBzvVi6Mog101ybQ5HHDKuhfhXhLBoHThUmUJcfasYwPoevcgE
ihpSWgpuTF/wRnxqjD/VLYojtkye0rG2iWsnCWkNBc5nH+qLJBpGbV6m4EFSXwhAiqwerj9Thevp
LNK3a+LX5zaBarkJTgAz64z+o7Zr0Amg806fjfzFPpuflateupsx+0Qwk81w4051/J3gOS2te/4d
/a2MUQ9Xp/Ock+psnJV65A29nvxMLm8CEhKglkKc7Y3y3n2C9qlSGwqXdqQRSGjJHw62tsaSML8K
NhHB7lC1ZPXHkxPEM1ofy7WmFa0lEL8vI5b2fE4NUjJjGt2XWXj4/jfeAjDqQePEy+g3XZyuCGYl
sas7wrQFomenJz8E0M/YDZ9pP80xsxunwmCsbOmQzbOEiHo9VzXXJwon6juwu4rHgRsj43fvvgGc
J1ZkBOV1Fj74Jp0zrETXVPH1pP7prVpjDs6Ai8Aqesw6XcE3lxo8Cpk018UMyS+wVrqNrp7K2hn0
5BYjKNFrwZ8nHe0kBqDBglg3ckbdKiZQyQT3go8SYeIiyL6VdUG/YnPxQNRmMTDQVY42uUwXjSgy
ey8m4tdTTOck4t1SIlGioVRWRjRh0lYEB18x07+PeEzFdPll6gfFWEs3P87PMJtQI6NSwuRJ9Q+c
QZsZJ4TCdFXS7y11eWIwHUO0xCAvK5sDywBgvAwKgtVXIJe9XO5nYzlJMuZcJfrx4afSuMpXfmSF
rzkcL6KMkJnbxCsdO7MZryHrxyb6hSgToksPE4vSa0isOgMCzHRngCLg1h62Np6hEnCW3yLXCeDn
OC97yUcpyMtyFhi1r1ObnB+iDLaSPZBS3sS1MoA5qLptYdEHhuv/LgMahEGD5rMmBrJ0bizk1s7d
Sb9PdM4QGOuxiIBzETaRQj7RYiE+3syIrwkYZeQP9LBtTeWhs0gR2goP32qxyI7IesfOxc1uBBsa
P4I6hY1W073GUKRgvoNgH98RP7TdRXaJAq+GVgwPzF5BBWZc+UuLDXX7uT29a01WH3lyM+DDtr/S
ao70FFSkzeYieg4fqZQ7llBocCP8YL04ghaZ3kDtCzIAbJSKHKHoFKZ8isW9U8xxegbIL2/P3Km6
MOJhSkaJ+JpEYETH3xZ2mRsDjjoBbhZ5ASgI5YoRIhb1SvxLvWfSwo8s5B52/oH69Rw56WQ2e9Hw
8higZiuHjIWzrGflc1+wr0hLL1IIbiaBl9nmWbL08Tr3BVznkIQ3gapnkfLuL9i8ccOiF0WW/N4P
jcSfrVRgsUL18wKE0DnjzMhULKaLM1DwWWBS/JYCoveUzelH/U5QijFAfVxrRXlo70Mj7DF3mFZ4
x1mvBoRfSq4iigJMFSQK4w+G78dgoKB3McD/SYwDHvDyhZmGBx7raxqvvQlA+9iWeggTE6pKDvwo
6HjsOrB4Ac3qDY8kDnnIZfAIBN5nS+WKMGhpWdIg0/50bms7rz+Doyb1fKIkEnk+Bm7ChpiVqVNm
IssikOdn6vIMPrv14R+W/MrYwk2aVjYo7bPTqcZjHnZwxgDVUqpBX93LNeQf7GWI4g6UdGn5863U
GeOjMv7bcS76jQCA3MjJqeqDbUNOYfrEEKlU77y6JhFyqMYOkMsx2v48xDKrd7u457dc1Yu/tkd0
d6DCZXWJOiriUeT1NwGrmSyQ4q9jsHjPdSJn7sv4GAMO68cxDjn6qioJ49TF9ZXq8cFUYMYUrgl0
2ArHsTpjld3JAkSXbqAQrhZsTbcsbrVdhXIcKAk9L1MaPFgLx49s9pLMgIPv0ogv1+9cJ8QLz3Zf
1I8xUet0oLcaxLN2klVvnGqfqLTku/dJqD/8XMTQmBDU1VVd0Vke6fJmpAevco5Be50bZvR0KsB2
BEVXEme4GnvDp5vTjVkkbAz9+sRtXpU4rZ/eAi53UO6MFP8Untwz7JprDcUacC1xg8ZF1bEujPRr
OuO9DnFwoIvbM/MZ7dMKRTk886bbwVtFG1f9wzs2XVpht4gVJAxnoGvzYQnl+LOnlgwRkVTzcPHl
A03WtUA1r4PnEWn438K0YO8UBB4J2sN3b8Xkya+p73K1eET8bbr1Owz75RVPguhVGh2Hnt0rfNTB
znGgXRkq03RTOA7DJEmJSuwtLyDSLFMRU+sw+61xLW5p3Mr6EJhGDrVjTGBLgYQzvn4kwa4qRLej
ldvI42dRsfb1VBL8WIPjuFzmURrNMj3lxKLh0qgZQ5n8WRopdNd4mKy/AFfCzfNZF/M4Wpn7P2PY
NecnJe1sFCU0AeeVtkTTo1NI7HoffKUhcUebKHUN9q4Sn2mP6Ob6QP4LXUi32IiQvBXuYgUYJNRL
yBFncZC0aRn5s6m2i8febpsuq+bldstWAWEnrxiJ4dvxm+l+/zZsPpfqd5zZPkhV2HirpSWkYCgQ
CglKzxR5lKynxd+0bPNCPPRYMqLyXCsv+d9F7xO00JobEl5b47qrNPMb14k39q+xDLXLHQxVjv71
/5oHjvZ3ktzhaumAnp9DnRKIuor2g0fL0maeOfGSW61goeLW9Aa7H/+ZVo8u8vAllPbQJXEfl+7r
1qV2JnlfT/7o/5itkRX7e7WwbvDI4H1q1bc1uowt0uqaomNXyYVzoTQUn0Ic9ZDENxm5OZccBUzA
WFhPE171d1jZrLiPAzBHEhkGryCjT4O8n1XqR7HphK07kW8kLFcjrpD+glXzhPpn9F90VU6gFHLT
svmGCpBMpBF7SeQ6tAXAy6SFuRGVqlbDWhsXrFabGCytO8sD6qqNSCLVTKsRygc5PWCDPeucWQhl
x7vtvhnYEx807xpm3sukG8bZDB/PrH6SshBqE7akFAZkEAxGK6iPfCvYqWZt9H3ifZGAE24cLAGp
J5tpoIrBIIz/4d7r572wQgNgbcwpyxeQ0gYLWjYepMGaGUBt986pyYZjb0q9VNk2E1ERuKub+/MX
b2kPhzrrLj+VSbwYZffx33qpRH7fKu4f9dkDsYflvbtznI/5eQqpdIP2iVZNI4EcPByBz0f0tRMc
M+HyPMSgmFOqRLaSv5J75SJNl/mdMf3t08g57G1zVR2z7gUxeX8xo8pPkyNDwowjPf9fzd5BwigD
iGoh1Rg70qgc43qBYbYCmTQqJf2/T9pk6/6BKuikJJy/y3zAECx2IrHwJjeeRej/QNMzVKE3pySO
SYjOMeDfEBblFbhiHkv79h239PMpHZejNRDtfOvu5+ZEUk1ptYSes2WpEH46qX2FfZX4weVgotiR
FwEXnhdd1Q/StjuK4doKz8+c5RHB+XOfJMmYmGmejbihoiO0gSO733IgTsrN8tn4Bj+SvdduS/pI
tUYnScz+XR3qjoOk1pP4vAZI+Xloer2ymaAkC8nHjSlV1Yvl7EVqZknXUgSYxUtFTwW4doQOBIH8
fj1pE+Za+Pp2KiBiTsFYXPZZ173DJtikM2InT0sobuRtHjLy7BnNwwHW7p6XhdEnBdrEGPAfVQBF
NYcWpfEeIHOCohhL0UVSvz6nKiwN2qCaJDyc4tNr/eWIen4XwZkhiCXw9G9r+r22iclw3of3vjWK
0a3sQQW9rUkboHJaZuAr5WJ+yugSohKY8xbwtkJX54ZA0CuibLWkfKAgC+Dax04ARChcgTNowFma
7qggjyS4/hs5RiMISdztynD+p8S9EzQGRgIJKmA58Xe2fBU2YOcsG3of3Jz4C0ccriuNsXw9J9sm
Siq0JQfP9whbHfFKguvBNFlkvVFSyQRuuGDG3/4d61Wtr4GbbG+iujSlEk0LN649JtEBSq4mozpO
5iQ0yL4IudY0ZIwTnJmgW5B9l+ZtXZNv8rQj2BaEwMIpYobFrS74S2CUaOSBg9POODzSM5IpJde1
RrH/KZ1t6Yz6C5ZIDNyFF+5pnwgnex/dX1kBKfAhVJAPWY8X6ELhggwhZH1jxwCSCzNgj29NLbQg
pO9lPsMIE+yDf7s+gTXA5D0Na4K+SPltBrhoa8phozShNKgkk71rgzdYah3FfKxE5EcteqMdTa6z
uK+ZxKGF2Y8bABFMSpNat+ZIPN3xHDeReF9t496yKHoUR/54nfkAgjj3gkaeBGjR4r7yW1+D9rtO
VFim/XhwOm4udG2jjekAaLMq9OrZvlNb9lVmfsJShCgytKP5JdPDAmt0u0Kxogvt+B6s8iU0CXa4
6nEkh4QsoBcQmb8RUZvn5imTass2aJbN6sWs2nViRtLqKz4VbPQWcRb9LPDkom1tAuvnCBflVN69
Ih7zISHr225l2tCAeJb5cBoajkd94J1yLvO+NVAiOej+jd9B1oV6lVsxIgcWnI8jdtq4J4/Y72S4
YxOn96pF6HeiVQ7g0YiU7bhiZ/WWYTL3MtVoO7QlEXeX5jrZh2lHlpIdBg+zKsNwlZgyUGyvvFrb
IL+8E4R+k5Q8t9WtJpJW2rARrgli9AvHiGHylNsIC2lQFRe28iJTWK9c2asMP1NU49PGjNXvv0J3
v3Lhew4qAnzIUX9GWPMTOkBdmc9ZD9bPkBPLylfdR5+pScTBXn90lQ7XhxJc2CX3CSra8JhubYzZ
dYOtn4cneKMHgWTPvs5tJm7sWBscVsxUgyqcLAubIOUYOaWKO/CI69TFlrY2JrvbfVDDhk05B7RN
OzrCzBpn5Xj8+d8gtA57NNaUocTAIGPqdlo9pImuuXdJJ3pijEhIY1sfhTjmtWp5fCFHWzWI0lXn
P8Zpz/e3Rou2uQ97yH+sw0RWk5M7D5VtNG3isTXuYDL4XJc4L52xe2xIAyjNNGPC/WxBEYm+1/fy
Je9zA72aEfdQOLHvu5QTgOQqxoAxbvV7JAdG6JU8tfmvRNzbt4RIjGgQT37pKuxTCIvr3vIV4yo2
eNbdwvKWnCP/ZGi8AYH5UjDkXCyxhwpxj0sK36P39x/ikxbVLi2oYewe0I9IN0jzA6ZP2NAOJHCj
Pr3wExXdDyysHK577GzhXNcgj9v7g9i0ivdSsnhDlwKy3pPGP082TA+ZCm2I9K89HjBtHBbKgIkK
NJ1TqlA8Wk/x1kBiH+4EWjDWkyePtMa14REEA7WU1OuvmRGPIeo7vijT7xvA/j0UwPjbH9zCBJ96
E8Qqox4gWXxXFv1sez1g0nqFAaKhlU9RDUcJ5+fI+yELdiWcpNZ+Bj2acFrupI2r2n0xz0/PKVL9
aJPHcHxVoiQPodGzGBAB18jduQUTCvN81iYICDeWfb3P1g0O1sUdTkCMbx6L3uLMafNj0v4K9i5p
H7lueZqIezSKme8OkpuNQU4Ua4YAJgrcee8J2hHVHrYnQ82gJ/HjKwZT/4R2b2HAsB77xdKIroNK
FPIZ58lwBXZ4beJ/5Bz4sS9E/ivyTcUL7L2Cj3ymuHfOFS8kETepsG+BiY6B6iVLDIYUmKX0i5Nc
A1scw7N0W3Ic2uTxesbshtiEcozAM1FlazdRrTf7UzAtj/nIUGkHOGz2v1HBSB4qy7iFyNJHjQsQ
MniqnQcFUqoCsmQHpqtTJc0ukknvauaEnT+752nQjOEqOzRIKNenWOQoiOWaG31ht9GUEdfT5Sh0
45OIPGsqMgImILIzf1GOiqlKdfgzYaRzUwk1SjgPkM5e6E8BRIxlnINDAMg33yHtRbBkeCsFb5Tz
UdVyGpt1CZNTihdlh4soaL6qhKTXAJGj4ttxImpn1LZC6SICnDHuE8XozHNlGcNh/2CuGOPoYubF
bf8YpqOW2REF0xpS2AUBzOYAkaPriY/pmn44G7i0FNtBqH5k0ximPne5SAyYWEMPn7DmkW99t1OA
7THr/W8zOjqvwedj+sJXk8iyGn2j/sgOqA68f0L6QMZx2nvM+tLZ0QxRvcekMKDocjpHCIneOYZK
ZyB53WcOsj79kQ9Vq/T4BaJfRpQ1RH00oUjK7eHqpD8YCoyZ8jIM2U3UGrSYKtAVOg5ep5hA/elB
DG9JR53bIqTWenJEFHfxGO7xd0v/T/Ss6fKtEMgI533NA9+GHW6UD6h1MQtOlnR+0L2KfLzp0KJz
XAOLaUrJ5azGTzFKUwL9fVR9jCJhyArSAn0ciZyntZ4trg2Ck3x2eQMpQTOeBGJRzk1SYWB+WRpd
ig+iL0FEupy2ZHatJmKGfo44rabrEg+lNKkW1hQkDm9QXF7oN9YRTL88ftuISFJEjAFe07QyaIWD
oR9bQ+Qsj05y8nqupVcwQVMkksiKIqBQ1+4t8q2CxhtO3wwa5YSUHQO6di56mVWeLY0EEtQYYvFk
JnfDZdRI65ILH9b8PzIj3QiobZe+R7sPYeu13fcl+PSTnBxcrnWcxYGb1y9ofSrjygByLeW2z7A1
iyXk2sKq8Mi60VkHS14Xx/SkqQDGoSohP9y4gE432m5PWMFlE4/E7aoh29ja0l1p76YQEeQEHB6h
PpLFxrQnSnyttZ7eaxS8HSf/FL0//hxeRwSwLKGgLhsVMUkIkZf1N06Sw9INRVXldDyoR95NU8xx
+5HFOHp6sNyQssX0HwuF3WTyDwOdp0O5GTmAQi1b9H2yLnOI/UpvZVcQSZToDO84YMymTk9wKsEQ
HdThQWqsRT/QyD4//wDQsRizsPuZoTjT1AEaaTEXn2lxcCuuyz/ovQwhSisTmLoVt517xXjENX8W
FIjJrEDfn0SBMoe2rn531I2Pza7aI+B6lH45WB/BvUbb5PENyUrd5Abco3+Fyoj6yqzwI7u5SZoT
G15v+u+33BXkZeKg9so2G5Y1zQ5RontKPj7INlGESWVbMQlygmUhAAKllgWr9CL+EsXEFEHSG+4X
7p/JN+rCZ+E3UGaLzAoxUgU3Qbqlt0xEmieD2s5/STMtaXyL/7+cYdgBrs9e9VIjOWqRZvvIohqC
WEgh86JBZWi5nlMBCahOC+SvrZq9FF+bN+AEk72hwkQa0t7AEbOr542yYLwI1GChefRWa3W+vtie
h2sGWhkOmKbDyzTqH/3EF29UH2izEkKZ01NmnFPPHk7NPySquH5TUBmOSkfjqtayDbLE+RaY24JJ
+2vjVSWQiO5Y4Cuv3eWRGX2DyF80kdbmmSH8c7opBtj9o5CfFjaA0sTajxXnI5El0AYNH9KkF2bE
QzdGc33hMma+QxIcpa4wJIub1M6ZF4zOgpzyhTYUsOXQv94UFQKpVflc0njH7Gog1pWXWB52+YlT
PIdakReAbSox44eTiHOojgNy1Br9jpE1ZrtLczeoy3oK/VMu0YUX+2R+6+O6eXuG7xwElSFxP+Z4
xwBWOhMglUfbn0fxBOs6jc1Z5r2A/ywLkix6yjpoETsEARGGLcK6SoGLHIbqgRKDpCx2nYt24YiU
ki9dMkKzLKhqRNFWWrkp3g6uD+STvDn7B3UQVgJnnoMfBkhxEmf9XWBwK6mzGbsg9SY4yJohzp2K
Pdz/oLcTfF/XHoMuX96xz+Dle4MiM44vZUqf/w90tyJi1mGvdC044gxEmH3fs6Sx67iNzvxLnaRZ
VDBOcOQZ0yEoyUZBC9NaMwKdGP4xSPLOKv6G0svUj2Gwu50YEtPnq2WAIDFZWIb2dg0gNpnykpO6
JErIJMZ0yr1R/kQR/p96bH6LiOBw0L4ejl7OStzG8NNlDIu5zXylhbt8A5xJFj+d9nUVHaD+oVlg
FnUivjf3OulBv4nRMFfTWRcZcugDlukD+R2+NrmBHilm1+DpABQc4oRc5pqK5r4tcE8eXyeR6w8+
3lWqlnwlAP5xhu+iK1abgSBKhpMJ8Jr4f42Xnm/RZXC1PzkE6OWXWNCq28MeizwoMewOieUrR1gB
pPIyXMJKjoDCM5V/cPvKhsXGlwiJHI1/ZC1rhsm+bO69+hRrT+DPFhYBep8jZKrruMImJZ9zPR7J
vMF2F+kfouat1Qyy8uKfmAiaOainoIlxo+kt3By/ywVlfwaizJ3fBQI8bkIjDa7c9zoTb62ovWet
/iiyY3otkW1f6+Ne1+etUW9FKgO6/ckB1tNjpTXuQwe2p9mOXB7CX7/5tmC5bigUEzDVoVRdbRQo
YGtgTfNz+t1svrGM8BIcdpo3IbFj3pmeICw5Yw7KJ8ou19Xm+TmaUrtXkxm6wRoy3JFve8GRlJdP
RVR4RJANC1E2oxLIisxRjEPdRJfWqS5Y3X9eCNENVwnbf0f+OTVklVezr+GaCuCS86hXRyIyHxbo
rLadIZvwmWZaVaj3LnrPJdNoxb78VWzsspIJu+d1fZCJs1CmAJoKhwMEKOzWzsV1l1Dq9GJCpRiV
CMjLCdczLOXQkIQXOABXNB7c+6A1fm8aiSl1trsMsj7L1t+Ex2dmR8QEUZj51Rd3trnpQ5PcpR6H
PX7wVjfG7wqzSV3jYRVu/q/kYB7PvE7ptW47LlAdEEIVoDf57MSu+kcg7xR0902CoazJbDCjnysl
j9A8QVCgv7vxqeKpjB8F3KHVw1mUImTyxSiJjVhx7YeJCL2oQYrMS5eKwG3QzCdUyHg8Qx2110CX
ygbF3eqDL9KZy+MyXtxlGd7kzvJ2ooKKgX+wqpeXk/YMcJfGprROALd1SN667YFfOi7so+ZMBaYo
OXKzHNoBCY6PA43cmtvDUyGX8TipE4o9x+O7hU7R/Xq9omHmnoL32BQF+DlkYXjYQXW8F/0+sjBR
jT9kxzkJPTXEe7yxLkZEbZ6uihO1LSWfTkaLrLlRJ+QazjHcIBD+IFzEs4ysWWwgcIPZgtAtr+O1
bB/NmXbZYc8s1SPAGDSQ1bxhtizBP+ixEhkBAtqTDg8p890EtTqTjMezwn4W4wIFyknW3Qg3ckon
COL1sdtoy91mCOfz011xojXl1xymKrCrJ3RIGv4iFCWEEr9r+FrUAj6s4SBL+0zDZIgauymMKbAL
dG9PpgIrda/VO2bN5dWtWg9wLUEfQxdYvMwH0xoUFVr1/UBiI4Gcv8CF5UvMyXX6PD2/26aTG/j4
hJIzsjdjIQyb4NotRFbqrn2cElHUtJ/IPcjwAj4lzV48HoHe2TzLiGEsFVsZYsLi/umwWTF+RXdf
y5dcykuZ7l1DmLL2gk0tTrNKM3BDRJrSCFSFSElOnTkmQNpqBzJJGreolgkhmsoBoxpQd6/fHj1D
GU5xnZk4SBFK4KuZo7wXRqmS778yzPPT0CsvF+h4VMiwX38tEJD8mjapzD8+CrZtCL42lbA7POYz
iRsOTH/SLedOSUm3/ycsJlpnxGxCK/zAUgREG7q0TfdDmH5GJDMZRN4FYC5h9kBUcZmsca/VV7CM
zafiq0VK+kAD0+PHqX/KZskLtOTPviJqjDg966dwKTRDK9Neen7yCoALwofhZjqeQ5InoyldXdzM
dNXlffM6yyzDMVsvMOrmO9MEpfSH2R5jYZe3YU6Nn22hHTLtP8j0wLVPkpFD8GlyoR9bdcgFh+aq
pAlZ2/H+osKb1L46iQKmlI7doAhHFt4tfrmToMB6NNDNF7vF3b6871mXKwW+t4pgqMSzC6UCn+mW
QGqNqULvctRGKLcafdTJOcfMCWIRXs2D4WEmaka/aVfsexXA9ZJtivdH0Lwd/F9wvR76vBnRgOc7
I5le1tCYsF/dMqdwxJPrwqJACDQTIO/wRk3JBwHRySzSyfzEU0oMtVTs9ci5U3s5+54xJzfzrwgm
ksKQS7Uwa5szSdMmmSDMNT+fhOE6aD/u8oGcq7be5HZLhV79K2Jp8cMxv4RWqBI8wS1XvM8LAFkb
DOnOl2MDSFUdQwnJhXSNCTZaeSAFCLztkiwmhKa+6N0AVVrsg75cQlNOFPLWnTjWXTDk/WDwGdfG
Gpc+Lblo28HyXKsd73gs+1SIPCtCD8nnp5sT52e95o9zoYzzhV4FZVIL/gEeMfl78SXVJjf35D0H
uPo0DxAmaF432Set9sHwt3lZI//IrJGZjrByHo2lATm9oa48n3KzihcLNKewSTSklbWPN9lvhXMt
3iQLw2CEYBj2g+YKZek/pxPjo+63lCVn/3TobirgnnDV8riuvNttAWXlsYH9MjfKd4WS6emIml66
/g6fMz+XTAR/dEUnxEV3NkkM9ZonuJdCS6MNsIDQNxdeUMMHNzJqxcbhcogenwFr4MwQzSMlo5yl
9zbly3lUPlxe369Z84KnPqexCaQcba9rB8Y/hGK0fhSn45xv7qFImShS+JxI75KXG1c1glbV+rdk
Pi8BYcYz2TfBPtVlJRLFo/y1TbuxwzFfQ6f5mQWEca5cy6D4z+AAAStRrY9ypdUD7hn1zqzupFjB
PkctPaID5n25aFPWVbMdJXb3WfH+Acg5a9apYcCPkRyOIyVuDnKSxY27ePjy5KtAAHhX9gE6p8Pt
OonZXGBLL+oYkLtwoP6lE3a9GDwnMHejATIeQ8KwFU+WjhvxXss7JnK6S2rVbYnVvsO5lNnaaoIj
jRDt9XF9qPHXjfIzqhywUKhWm34APbMhGfkov0gl8W0YLl7xJhiQDuGa36nr7QPyyEbIhsVlQCGF
wcgzMoD9nGKUgOYsbqjTELdGd88kvYVAEuWQm4cJZzuCv5B9OWPDtLjc5nCqkjgre8BJDDywfXGr
Tq4U68nCebzuYsUd/i9qszaEphfO58jNDe8vKXZF8GwHOJaTG1mrdQ6ZJnv8UvnnyfP6+4mJbqon
a3WRBkvlNvvBHDtNyJZqRvuSFupvl21xl/9e1jkMKtYc+xqs+1FCjG3IdumqYEEwHTi/8jQl/RtR
91opFK3pC8Qw0fY77farNv/+yWFORFDF2j+1b4P7xGaaExcclVfQk2HngbbHB/pk2bTNacWeadPf
Vh88Qxhyc+6YEagTuGOn33uaBeDqLxC1Er1dKq5NhdnZ4CZ901elB8Gk/UY3kM2NHGBl9wWactAK
5b9KOhfjRzl/OZxdP1cCL30luYVZBy+oOZJbhm4hhYvSN8yVglFPnH7zlNjE5lfcqRo4q5kUzNeu
qcCmTAmV883a0Tr3ZSsC4ANFkMgIGwv5z6D7r3HtmxOGB23VNZ1k1tmdDCllTQihb56pzt3R4anY
ypoFvuymiFTNY9SvQJYR+1N5Q9covTLWZWsi9YguzfKiHClqQ1ZOMDytIQdr7ixZlue/4TxMmzTY
kwN9F1vWs6tfWzOr4Cd2DbwHJ7qNNClHW6LUIuuGXx5wWYiAJojfxDRmvYI5O2u38B61dQrK9g5e
UqLoJf8nCQWn1GowI9mzEQiPv9yFz7AdI1/R4zJl5YSOSftKHWegnjygpEfhC/CSo+ywaBpCYgTI
pQlsq3PdGykO2uK0nXcmxO3V3XJRINZQBYUVoMzex2wOVIVXdbe3BfsP7KORBjruhnKr5Y1yDA1K
lEZGfRSiTc4fkhO0kUM+tUw06T72qDia6UXYD3gHho6pphN5Wc5sur/fPfKzOw16Idn3o4NwJwdF
8NWpFnBrt0PETqRYU3iC2ebdADEA1coQvZXLm8fb2iulbszlcN+AEPHE+TW3LcMTjPIlY8wnWwCw
KIFD4Idl/sN6IcISYu4fZE93lAfwRJaIgZMrBtjdJGKXeEuMAAcSUzXqF5vG1l1oEmTcq19+8sIl
8WpUA4L8ffnbY2fUTTvIOPngM309obTsDOEfVuzOU66ard64YQjbc9qzVsDuoggEovcnuXmb74bO
ISVMFMfJ/N8ZxpeltmobRBUHgy8Z+TbsVos5MLM+2Bk4ajzY70/nljgI8g/JyI3EZgqwOKxvL9IP
fx1+EmI9KRuYwU7rcFjx9f9yaFtGG6G2B8p4tJtXmKh/5x1Cddkq/PGs1ZwQkKnHcmvIt1iumJ6o
6fjZHI3d0dl566Qtlfnskpya2yUnoe+HUMjBlg6PSe6ZaMKVtBXUllxb0mBRyz0eZ2lqVg74DI35
XHH/OGtBexRxDpjVoSAfCoQsz0LOiqrOaoWMNYfOQsHPXOulAh6GLhT36deS04Eg4hjZfqW9prb1
UOO+QEX0AFzgiD56Hm22Z9lLiWZZu/P9saYZPoY/GqBpgAka+FMQ3zPJtc7ueu38DutdHa2+QBED
sj1htyBHQoa0/TrcD52ttCHFVy5OlH93BF6DVl3wioZCC0xKAluXo0qNuzSGbdmVnz3+WrYfhE+w
m/+Oy+oKgWR8M6RAaTE+vTP9OVBqtbJBK0VH4K6kmwrY9Mo+L/GIJ9NGg6aRbRdaVIjc2DNnBlb1
ZYmq7r7ZwHag687elWmwzPxOd36dBrmU3C34zVlnCpYTZrwr+4cUSW5XtA9yzNEeAggVYzxM7Mcw
BiOgJg6lR4lDPaU8RkJDB8x87okH12XMAeJ9hu8kvpBi+JPveVMKHLbJX9gmrTIw/Cqna/dEUgvP
w/pdZAUNzrbVVGwq/6fwWCUbMMZOgiNBmUb0VacIHi5M0sRMGmSq6e9EdbtoPtpaDyPAOmIgixeD
sPoLgK1YeFGygVkIQ7m7Nuv5xA7Gm/LZVrI+1uZ0xvjd0HiK4e0/x4+K2YPWLq8pBmzZf+9LlQv4
xcDYBA7eyerUZW7kAt1Dhqe0IpqVRM6SMxTrvWhU6/Xkr8hk8pmvi1GORD71dboWKSnREgDfru7/
QxjskcFlj3YYVKHr4RqyrPcu0P78AcvAGdy9sxbXMIkVNxgl5XL2TsNNXOjJTpTyE5Jt5xcJP5qd
T3v9pg4P1iniaxMnDryd0PyAwQoDRkvme72cb7urJHmdYgP0BH6Je+J8M3km5xa+MC2vOT16+/Lu
D6bFH/v1nj16zZNrkAAfmXn4/G0tvXjhbXardzgx3AzHuutX8AlDMt0H+EEstpiuz8tcbam9qFks
S+ARN6l+5MqM4gsaGp68AzX8fmv281lSRnNHucD7NZNBhaCjLYU0LewmClA2PITO8DiDwDihImMD
oNEkxWXyURx53Dd9+9nRAR9h5jvZ17rVPLBnhwTO7+We9DjseHFlmRGRQozDJkCvOQC9OQF40bPh
zq5gQ47mAdq9+/RHuJ+GxnJZ5Wd46tfpt1Nb7RseltVxU5hUsffnmfwBsY/ovWy3QfNGDHzOexVR
mtrFjAJSbp9HyKdfKKnBSl1ik8ueDiMsiq3Pw/2YD/Keh7y0Z1PgwDcoa920/i7NTlNAO0YbgeSU
f+aZkraXUdFi2vMDmFyXqgt10xIYBKkSFeOd68IR7wutxwrYAyoZwJI8HIFXMQ+9QIsJ6nY1PJVd
92h7slwgW+05z3LUkHArSdVxN7bQPiX19juTuDV2hZHTbjjQ7blx9RnnhB9kmu8GTsnDFzgPdhNc
dJYXToce384gdgxObCWMd889jaRhqophtw3K5hULcek6H7GaJgjqBV9SnBau1X0RxGRqXh7OHoWL
yDTtfPSLZXz3YkgUgi8PjtkrfeXJR0rmm3frcB+oe2Io641UBV2YRUhBRwI0ypZt0oj0DLARPSao
zwI47RRAK/LS8wjqjvdS8T57S7B/yqJIHqkV6X5Nw7FY7v7OUiqcIZ+g1uk5E1a/QEA7tDuf1y6o
6hvrgp2HpVZbOqCySyXKCnnmXTlR8o/JwEmVz74PF3B/Z2TmT9uL5qkVIH0YmF7Kvo7vrQDKvfQK
oUdR/s4wuW7P9bPrgEsKB8Ewur6FirLcSsaO4vDfSGMT6kufK8A2AnLd62kgEOzhvHDelEMGOXjj
8CgaJl8E1U8u9VZVH6LUW5+92CmkNGxgdKhSGGxO6purLPG1LydqY/CIYmI2vJIMz7ZycnNch9JY
r+J8UBIQxYYGWG3cMPuMFyhyasWEsH2flvI0o8HjJubISZvQvxpWhniTHv/VtZT1ohkW00s+Tr8n
sHh1S6BoMwV1lA2MTm5agH0yQGmc59oezvrBAoZW42Iaq4WMPZUzrnyBaaUAN1pxxfNBFxr+twU3
3ocNv9Ha66TpsooJXPSCzZEwPgXIj581J8vHjYT6VDWO66FUaCIMR5jggVPf+Rl+nZpZYEhGX0Zn
dWJYTg/b8BGZmNgpREV9oV5wdfSp+GFnbrnkVp4iv5MqggAnPD44viOELAoT/dFbcu7ZqUdizN2C
nVhJV5HsKObJPThQo4/UJHDFLDI7AdbtFSZoTmp2Ve1IBSKD89AsByai6/idxS5/B4yHIb75BFZ2
rInPEpGaP+olXQ75h5GAkakmVMVBD35KwZJmRTXQirAoZCCkLFyTuvOM2/WCzi1Z+UzgiUlBhcRp
b+Yar6spoOpN/cKKup3bj5J7d2FaNlO1cMkCu/0Hxl0YCzP0bwQLqGkI80qNGSGmxMPxELsMTVZH
obpn5q9BC/1dzgGx8tVqcB0T5XraX90457DqANlIbAcR8ArVHCSPZ5wkwvzS55Y3NOl87D2CDP/J
wZZOb44B5g2WwvM2dt0XayJBhRQdKip8Fb4bO5d7Of6Yam6q7WMMEqVGqbr9K/0cJjptIBKlFcJj
25TkjzNT2wyBJ10z7vmCiHDN/BoqYRkTvmj978q3R8VZ4p6OJf4pVvlZWQOGa10nvwzcuFFDbBTk
yNZb20mRJQPU1kgYxYfy8Sr0MO8BNQHF+wc2FJc+10nCZrY1VkvfafEsSfqFXTIpgOD1AzXWenIk
ZHgZ6ii7J98VltoeJvEVpBx5jK1jXPqmEUFach0j8BvMuIbKg4PYphyVgsYLl12tUb2JFdNQIlbC
IcK3dqZlHl2aj79yMtMocss16Bi+nbu9veGhBwUqHEroEh6LvaIrJXL7nFM9YEo9CAfYZaOm//f8
jCEoGyEwFQPEBr7rE0t8PiDWxpzWgtq/1/PCONoR1rK3d/tysElIc/D5BOqB8f56ixvI/QMIeMbu
iCXGZOU0P+854OvV9IwQpNPstn7/2Mih9dzIFF4ytq1HOkgMyHOGS0GLWBIu0j5/YvWHt+1Hio5H
hSamJYJv1HXSk5yOBiIaXhokU6tw/n0Hrcf9+NFugUbqLWwSXyLxpt75p+auARbAkwG9ygLXwilC
FyrDon95QB3vhV5LSh+T4X62cDJaXnSoK6lqgcBHW5Qz1KvdBaBjKxPgRnreIk/Wzu3N6Fug1KvX
G9RsWMAk6wtfi+dTPDv/CidwvzE9jAdQecNwmRAIRzJ424B8Epp1Fu1eFX1r4z+ufonunkZe8KPu
2Y62lgLVecUxBSgmBoYF1dP+iLrgqynUVwlaUYei/C6H3CeFg9fwIKIq7OA60hhU2PlPeratYZ57
YlQgmrR8nJ64FF90I9uCJbMm4zmJcF1G/dbWAybPrLTD+to3ZU6E5qtoKaPXfZo452WMsCfJoDuD
g87iHa80zD51D3akBi/hppqHa4dLAHPzvQJK5205lCSwsq91nZfE091WBTCEbzpIpOQpU5wbAdje
SfwUs+gnJPuUrBvv9u7HbgA7RLxoJIcxleoaL1V/2RXD9Qudx+Beblxl5/2WFTj08shoVDUIAqIf
1mSg06Y0wsn92vkJ5UOFJXfviTY8Xm+P1eXFAn/6r4iavRrGybznYbl3gaiSQLTCweUmywciPA/f
yyW3efZ2tJjxXU35Ufs8m1ooITEkU6bUGSCdokarKNdfSTYvHZJBQt1NQFQMsAySvdn9tyamHS1D
taBVM6xqwKx3Mmh3DZhKCY3g6skOPd39alTzAiPw68CFRqeGeQ7JUsXy33V2wiS/56/SeV5oKSdB
2Cn7zUo+zJ8ZDzJHqH4e8FCmprIPKBoJvNb/DAlay2+FMuq6RoZlJ7oIgg8rK+nTjvqhOtg7Z/lG
c67PZhPEFvTVttbEGJrV7CNSGMXFAKiQh5ZE3oYwQCR0g1unK7QjxMnLEW0LYiv4vn1vVVD1q1D3
XaQaZc7UfJuIehmewLMj2FjFGI9dMW1FPGqr8i5HhamLCNMpxQwNZ+TtKWuvpT0Bq+H+MWSCG6IL
s3JzpOuK4FRFXTXzhREBrHLk3JjfQ+5PVBcswnFzkZAk+WpF1kL7owAtR4ATbeBNWwOTXP5y7I6G
Jt6GR5PVXfksJKHaWb8zIkkrq7qPGGEG6RR8QNn58ZtjUsskbS+kaWHrW7kZAuKWUh471BQPEDNZ
UQmjYOMthWMDqRR38HAANxb4+rZlNP25z/fV1+31ZFoC+YGhiRpLLvMdjk91kHpwXjCT/CDQWvP2
PVJ6vs8Z+r+nTxZc0/D84P9J227V2LK5fWv3osKifqu6m5Ccx6r7t7VyUO3qQwwmUsBYjIfUQfTA
BLT/y+zoCTHPvcbh1de9Mh7TQ4cHJjDnb3itE6TpojYdpDEI/XIJqkEked0YySdohntln0Em6n01
vwiLphkLK+3/dLKqEdDVRuiWC+HczTgiSy0o+/NRWGkXFHDWRHTeI4EVA/dJFiljno5Bxh7NGT8D
tx0/VTgRf+5oB/dyNf/U1RxI407F7XS4Ny+FjYw2A+r3vP8XwLKVXUgCJR7z0RZDvJx6MtzKfG4C
VWVSQ1JTj8HnPTp2LjrLruZaKnJ4SR41YBICWgbMleHmxrbgXyWytHdqxVoWOEHM2WO8gKibB8SF
Z+lwjoRLTibTy2PzjhS4m4TlGI2iKhOQoLuksKEITo643UR05GJRpit3JviQ66cx35VmsRBiBs7k
3ik/NTtoGsaDCbCszOASMhGlepT4TnSWp6AIvR7iHgVfQbLKAb+h4ZNZncDkMo8G1HeS+kqvkc6m
+mQqlHDz6sMWkcp8/wOhIoXzbKtJDH+smbHXSafIOWBvQlFpU/ffJATRVXxiL+LdIMd+ljnyTNVw
thdVOPjYt6TJR/+iw0Wa7kj78lkqCb/9nLUqQEc8tcjgplN/kPQSeFr2UhUxzMaeZXhNDenAknhm
952LIdpl50u2XfGCbby8bbE+jE47bClnIUBYY6plFuH+QCXETHogVdmEXp8yAt/oKOSfuDdyF3pY
fEkuMcjdD3is17xhfWfIpQlqwW30ExymkMH3n0Fdn2LTnvkhvZmkG4GaFtP2t0T7uu9M9GnZBbaU
i0ONVD41hGfxOrDH7dD6JPLifMDyjoGkgeFbR9JMPUNuW7DE3izdLQDyZvPyUcJxqnKkopUkbF6/
e5I7bPne6N2q85z+typ5TlIDBJZhzTK7wHu4RsaT5yQN3k3KI/VKCMpUnCxpSEPhu6scDVHgknfZ
jTFbotMucLT2WiUv41oMcn5pyQvO2O5L3NsuUuntlP0TD1pCQe+mno7yzzW+Mp8QHjH6yl1OWP3h
5WtHW/3gdcWkaw3M8CIanrE6wl3gUl41oRnxjBQLXjnIojC3hHC6PS2l5Z+pZZaHW/OFteSZ7J46
wJDgaheOQRQ9MjKKrYceR4h+4KN42J/U6HNOVWhr8GIug/mYTOrHX4JEM4d57bXNUeRHcUpBOs06
q5gJ4EsJA6wanVSHf4IupUzJqvh9f6P9fCv38w5JZJ0prnYgnOS7nE/2EXtkG2zMu3DHPe13nmeF
KknxQ4nnikoDGdSCynsbxXihQYsPkoFivgRDZjo/Ex9mlMMdov7FHdhYyUqbfB4txD2JihHBIBUm
/0t/7HYAlWmsDsTtab7eCpNSVjREHnVjKZzFCVS1LZgP93mxwypeCfANQ5QHhOU499aoHkqDqTJL
R40O4pleYBjPsM5q/M8smtGgpKwn3HIyH51lD5MSjuiRa/HrNLx/feWptNgBZI/HiqOdySDNl2/T
OkuzLMhDtc/hMxGfiDEm+iKIdr9CnB0z6TISwrLiRsRHwP8d0wZ/140izdvrUP+W3dynDEJYP8w/
Cl+xhefAvFWj2a4nt4VnCpXrMNKx8iwKd5ikN2CL/80EX1khRSgQdUFshfXfWNCMdClvT83cOKlO
1sbgqx4QgVCGgjYt5gyHN4TDLNb4X9CMliAFvILMx1EcnchET/Vg8ZeyAyvf57yU84QkKm6gzqju
igRNY33EtfBmQqfJRaikMyGLd+6DwwAlY/C08T/EBOatkE/ANW5SS9rIT/qsJhqBHE1bEisqSbVZ
HCk865IDsqckH1cgE4cN2QVvXpkeAXYdInaIVlUcStC172gQ0VQWg0e075vxKH59oak8f1WH2kUu
ZSyNJdWnE35wO0nGq/7CNsLGdyHEDwKeWQH/Pd1JlV7qnAiSEY33Ebb9WKqukRzKFrGoNY++B1Pu
gOi1TxXp+5XTGFk8DkpbLThywPwgAGhoMx3ChtBa3SC7kaJytdVVaDNn6xTlvhnE4uHf6hLdMOnW
LlWct8xMjzyDXmWyIHT41NhPbEuelDkJJtNHMkp3zzuXSFrV7Scn6eqqyKMhMgeQYQ/x3SmZC0oC
xOGEaHrC+WKiNXapR2Uppg2+7YEt5G9SXlea3Nfj6p0XDMVGh2jgtxHtKQavwMvMGmdSDO2Necyj
fx1mwSWUWvxR+DPqyuXiD0UDjknXeeOUzl6t6LNl1t9XZKkAAJLKFWrenDofI8+gWKLwlHUMYgwj
U0BKwUBqaJUFOjR/YX0U5Cht94KkPdnWjjYfIr5yzOB7Fo9SBpUqDAzKSgCMwumNa08bb30f9hMd
/2Md+kCNJ/N2p+bjQKCHD3cgq6oL4O+O2M0gHYdE4GJ7qt1kUBugfV44/Y/b5jXoVMMm2NiUIA5s
zjXz5wuGCrlErj8OMauD29hd9ZNuF2DueXmOIi2VRM+54d8M4s+l6w4QBRSmHMRlVD4639RC9jn7
oK+PWiXgV89ngYcsQZqA/xGoqf6DgYyXfwyDE/AXMe+cOHwRZsQEdp9tD+7MP/gY+LBKIINNJTdm
fD2nGdLlbBpL2vwYOWYyrJCFtX896WFy/o2LFzPs53atp79LPeeHpGljzuuz4yN9Jplv+wBu4EE5
/pfCdQoWLo0upxUK8FOHDOg+ndXpyhFRXSXF+GLGwCcL36xmdNB2jtFF45jSLcOtDnG8nLpVre9C
VbdjJECQ5/ViCJ9klufzj4J9tylKxDbVga6sa3ILEIdYg0HyizRmD68yQ110t+vbu+Ipc0XZlOhN
Dfu6IDBIEpOaHkhfgALXEXzeQE84biEhE4teZrFbSQAYyyEYh5gySj6V0y+Mu0SMdcNd9LBiP4Vr
HAE1xIba8wS0g9Niq3HU4F7Sq3sj+51gwU+RlfN4lzZUq8ZqeRsPN4Q3ADfcXKI6eTgz5Mbms28E
yrX85i/iL/sXZN9l0Hk+I/wW392t0cjnlWOHIm2tWYxPXMuRFYxWWShQyMbdlqRALKgtLHVBQog0
HMDosOjoSIMFh8OIpDecZ5thxeqm9bUCppK3zJv2/w2QB8YaH+5qcj5HDNGZDHWSan3wm8PvhCoL
4NY6FTvLBrmLo6vrjpkIPg5sVKnG8EY3i32fXsLs3YCMw//bX2xz878Hm7Q7FjYbcafS1eZ2liJz
/+2ItBune/0Xb6WPwkQ8o6qwtaFBbKgG/f8a8jxyCO+SXIP0+8fp7jNjc1joMWEsbRggCRKGQ2dq
q3Ln+wfHtNl7bIns0JsUd50hjWTTRAh7yMKENkMyVC8E4AlNNo8KTAK/jrnMRP6xRYruCuHK1403
NgSAxJqy05K6mK1vztxQfwj8mGJ4surVkz5Vi3nmL3I38n9XfL+RhF80mNl1jMqzqsLQQqdzyJ/e
zjOvlyG2Y2uwnKGTHDftwCh6rIc7Tz2ZWxAhQA8FFdrslyQt40fLJz7uF5O67Tx2/E4z9+jceG1V
Py571VPkvaPsthD4yUQyZodI7Y8TL5i5HC3mPluy+/vYdjBtn+ND1mpoT2g95WktGOBZr7snIbxw
FeenAsefBFiaMJ70UdnlsJZ0gTncvcyEF/6EPR69jF+mTZ1O6s08hKTS7RdRCmJGmAcWnajfFsoU
PPtPPU9qs3E+X6t28QxxeepHZU6hZYtLinp9Q3n4ztUUDXRhj+3FnTLwqBdXT+2CcfsQmCb1lG/Q
QnipVvEQQRZSa4jA7MphT0Qoel3NWJcuhSkyAIY+caYe2AC6P53hJ5n9glcc0R/K8XTayToYi1KJ
+MvIEhLsrTiSbMUTngZ7+54RukNZJIRt490dbcJH7qiaWn6ufid3N3xOkJ2Rksy6dLU01lwS6fxM
BzlgYAbSUP3blTirRXXo4bxeps+HMahaeturVm3sl2mk1GjDyuwXMDKAwmIR1YRfxpcdgeE3j+3O
vT3yIMcdteT15jGBco+u9GnrlVVYf+/2+il+xjP4rDfrWlRoCAKbHrUX+zDUUzmCtWrddj/HbgW3
pzs/zm+6b6TIkgE6LzUNq3jZXI4raNRMqOvlBzAR2tQ8dbush1CPYzkCxHPhVB/HTcgEbCVbjnJS
xiw9JTrlbfFLWWat2/6N55/zpmAb5gPh8V5/o85rpqPav6WylLN67iR3BC1koxXSoV6giWT94Fhr
qFHw99/bWT6i7edrF8IkOTYspjNV1MPVvWwO6MjSP/KhKuf/NISIFfmFVNGVkZ6K8+IdKnFEkbf+
pIzbfPosyWMoIEZmEOvX/yhBl+Rgn92cU9vNC+C8h0ADc90F/L3spUgrXf5/b9IpGCGkw/j9pChF
AHQ8y3LCjQ+ElmRcAHoIPAUliijfI1D1yaUZaWreHMofpAOV7slPtjUxrJAvtHm2ts8Wql5W1I/1
ixaq4QZBnG6foujop6xuQ1FiRxh0CVl5M++LAeqsM2IqwCd9Nd03NO5/qqsoTGJHquzInnIzt2iE
bqAL2bXc6PYUiylHxxVmnV8i3eOHdwIdwu92qkVaZKU0wotAVaWqWlVZ4pSo9UYxHbUb33Ka7TPS
nlZdIdtGN8tqfPSpaH/bqsbkY8M1F8y1kIlvrt9D4iR9ublGqWGp2PR2aKaKwVgej/7J9H05/6/A
MjS6WWoZ1b9vsKcMaZvfyoOxB3zjwO5aawpSlP8Wc9NBv4WwOGWkkRALJ2+mfUJL8S6/T+8G0+Zd
XqMugkA/950PeMPJ+Wf4eMhD4NpwXxs6PAdJINIA2DGoMHMFJg+3TVJunxFztUnwnN6sWSTipnFX
ZJ3zHYk6eQ9zaVrdJouTfuXMQ8IeiP45vRcms2GsGBW/q3BN9Pnz88i1cUPHhgLnzujKmBVf6Y2O
Z/YUdyY+ZtV6diDg/tJYkKSQVUw54geIGu9tDElTR/q0HUCIwBIUnLYZcE/12Z7C7QmQlVJMP0A4
vX7ZBSDie8rZn6cPRlRGGtsRENNu/83rCVxwhRD74ZHlK9VnRCkXQ2Y2YnThiIAtI9E5iE+sZy7A
4tDNvB+GU+1zEHZenRDv87kR4etajDXgNdNZlE3Uk7w2x7oP41oF+Xsp5WD1e/AQjXd2gSURWeSM
VlVkYrRHyj14VjiOmMEFyYsnNrWms0cg4V4S64yGRz0MEkz3RzuCUvAKMcl0Xwu50lejWXhpKoDI
7mqsYATj1ow5xj6e2PYfp6BIu04f8oTcb7Lx/gIIx4hSQeu7ee1VQ9JQq6OxWKffTz3wTn2DmDNv
L72sfyEp8rarCgzPjpi1H4gFwRcFGQb5iO/3UcYPJbufjtqDlXDDqRPefTAwfGJ6AVV8GK4ur0C1
D/bN+4cZoLTmnFTrc0X6tFkRTBcSBIecRPVy+7IvAQ8KWWRaTpt9580BxMh1szcdldzwJfPJKFeW
tYYah8NiPbCHeIuXi23Ey9P9X5+HJ4Cu24d4UK4CJd0k3RSQ2lTqp0J5uUlV99suEhq3VrCp85xm
TNpIgIhs3xm8p60brh7eSYapT/qYyDFtb32Mg/mlI8j7fOL6yEwslt0UWoOk7adRRQqTac0zuubf
Yoz5J34Rc0QbwDCT+ukCnE1UpcQUCQQ0HGkrl1WBSI6xbKTdatLe5OEE06LknVyuFgVrDWiVyb8M
lwKCGid7897XgoV1ZD+bqNpxBDsEh6DOtD1kRRtzokmGSdkxvQyVcTI9T1kqvRQX4GW8lPG/bkvc
bYS2RDmWqQe+k8UoYA20MI7ssnebgc9UNMEYvMVMEncfWV8Mdgt2cahUuEgpxkAtk3vdG1zMq2eK
s4fTUFUkULDMsL7pCk8Q15klwt1m2ZdTajYfOviHAr8miVhFAyJlKwBG6cGNBY9ixq8nrwxgkZLO
4zeDTuWp01dTj/HeLXlWcZOlqawDGL6GkgEpUCdVoy1qgtW26dSZpE9HCsd8Se97mWW2uDMZLScE
qo/7NcuFSzFqR1tzxTZ2vP+oUwapXU/2kShsVzLxCbG0Mz5Dhd+MNb+IxZne4n7/EzEfdgKTLUJ1
HJUGlYuXaL32Fx/g7SAt9rbzPPQR5A8pUn0PtUtXQVXNdyqYdXqQVkaFRqMVFG3CJGXRoLO/fg6I
SDYAdiudpMto4eWyf0lWxNs/6jfkXloJdWBtAbF66Bp6VcQXxQ38fdwQzGCaIk4HEonYOfinSmkT
m0hlFfyRDbAPIo5Qt/3rrshetVys7sWToBgH1/+sYaFw4QfpYXTBLM1NX43TWluwyxT0GA/n70dZ
hVwLX68vqg4jmz8MOJN6vS2K7fCPnqCgsrfzzaV3oeiWYgUXS+y4yimIOOv5l/WQ5mid3JzpDgu+
42I/BtG6tNA3Di/M7X9JilR0n+XAPgtlmEomlGhEmmzLOs/qwmfZ1Jne1jJ3/Juo1sD4N+X3WQiw
D5MF1ByyzLozViJ4h8XpJptg+tHHab2rm3o7nVtGDTeA6uRXqTfxDBay3kQVPc3HDwP3clkU7s7J
7go7GtOJn8Gn0ttKievxDroiaVByIIsVd7Yc7ZRE1hA/DA2QYPVEqQS5VICgFyjo7/WpbbLN/z0Q
o/xi8RxjqFsaQwgDEjjwTBOn7VAzURs0/TvPkP8CLpF9cnt0m1PDe9MOnwpcVIQjmHxplANs26h+
O4o1vGwSUFeQ6zi06gVyAEcS74jlwOY9TUXQ8+TVOL/mKXveH5kDLdzyyoCjFyHcsjCX3zcTE0np
IWWlxSKWcO5mq+UOkwif8HOBrihVKoFfXsmfUsZyExM1UVS1mhCI0c4kBXz1yvX1FWIf+PIiZLrm
tfgitSAC2+Yy2s+lDerUSfWv//ZPcd98nUFGt8/tnO8k5fiuTQ0NUBR+bqWvUXaJbuMNddZON0wL
9j6J51uEU3Rb6Wifwp6fMoojOgSpcG+r1vv4O2pyKfiA58roDscpMgLr48Hc5QEfbCSTRokIghr/
e9fI7/8sfmyX2QG9BeaaBhz8bCg0b1eviI7/yadrVqBNnKDm2Dbit3z++ulSXOd0ki6IXu7sb/qK
+vmf1jeQagH09RoPm2LP/qlQnUMlZj7ZtPCtM40E+NktlWHBXkClkTlEJTOktiC+9+FN6mS05j78
Xj/uNuxaEJGIqXWxaUL5YYX2SWi96cqamPxQQUBNt51OQBhvXi/SkKr++DAy+dBPuqJV64MVGCKM
Q3lCP3bRstP4dF4DaKOHuBrN77dmUuB32y2QkxsGcWX1ocZzlOSuzkPYCPKbg51OuvY5Ky3ko16s
9SdJ7cEjRLpWzWSm4I+5vgctaXDK2oKelH/8G4KEPlGKxo+aKQGkoKvOJMw4+eNDLU4In9vm3n9o
kN3H9oYkTx31u4iemPksV7Y95wcDWuD4tKAaBhITXXZqdZFEpMeKAcfTsV6M7ztu16jnclxzL/Ff
G9U5lQjd7AJL8kfSRW+P0a4Yxjm51UHg4aCAjF6F8R/q5qqhcPHg5V/xH13asV6Io3TA+4apaSnx
HbekAn3DN7ExfW3QEFgXswOZ+VDk0f2fE3oia0vzWu4vlvxHaOfNenzK7C7T9H7oPSd/gyMJNJqR
UgjG25cB7PfYxVtUIWSVdqzROYHe2iyHKMk8nw+b9qNcSxrxa1buPeylk9NF3/a7p6G7VaXpM9oq
CLuer+fxriLX0mAk9rg5x5RsCV9Y3o83QqMhrK4IvLSsmbxDg4960G4dbjZt56CfMeqA0VnkYhbF
kKpOuQJYfb0hKWwBIcu/j0onMXakyg85nUktRnbijKiNiMHwn7KZ50//TwjIABfh+T7X+q+IQNB4
YxZPGltbUpEkndD2UdgyR53w4eI/H1SHNkeNXcSyONLi40Zi0VN19zRdXLlUEcQ79E3r8nSLRekl
5EfkGx6tIu5H4YahBDUBMVAoFOrneNwxe5RcxP6EjvnUBCPx314zC2BePscn0Ozj3JsbLezFChhs
PIAUGTO+f8C0IJU19dL2RGxe32e/P6l+B5pdF8Dy1lCVGAJxMdUKWz0VIVjPvg/RzjTtyxF9SjBi
NQ3hgEJWUilk9k4fO34sKKW43Cx/M48A4gYn3yy56YjjD4i329mCEIzJovPLEcCj3fHwWO6z9EVc
DOr8gQkoXGep2iUNkJpOabKw5Z7y0nvHcMpojWSOsD8QKfN5XSyG7GyzF00+JTwihY6q/pa3zggf
S1CnjE/ERPPeeK92l9XMQlqIS36Oia8jkEChcFRKiXC+oFiLUO1PsoQIAMUD+lfdTYYPbXKA4ZoZ
cPIEZcHLASfK5hU8g7cLkOkxkDEgLPsXhx8MCbeNzItEAxY2Uw3VJD1dL6pVTUvA3U6rkzcoYWcz
Wdii2Ahf+WeD1+f2h6y8GEvtZIqccdu6sr9V/QcGB8ltwmro8tr7kgIRP8UY10d1zYr7MgeX72Q6
G+Gb74tfBOoXBHDjAQNmn5a7XWM5ppOS+N5m+DaalrNAa7FKVl9+IOsisi/RrAKOTmscphGchQKm
W11MA9KO7silgNng1NFMSP48+ouJLWW3PmqeBr5v0lkJq6mbQda9RK++X2cdhEJaIMfAeauE6tX8
3v3IxGDviOaMCgxEjd8JrAnAmroXnh8/1R2oxFQ03Vw+8ED8i/z9OmyCa9h4VCwKE/Gr/aZ0PNWP
6GDB2FVbvwj5YKPJVCsVFNphszg86xH2+xlmLE22AAUrLzR0ELQ0S0jdCo6jr85VrqDhh1qLgGGF
bdE+pTESok3Gnp3cAkN10cHmSRMo5eiV4KixnOxGiTHf8ucGfq43Z7OZ458dKKvi+6QgSE387qPU
QJe8GRNTkJ+KNEwgMTyLhS7SRBufUX/UVIPrxyyuMUiG3v7ynrsZ0JxD2EkbvCg19I54jKrYNe/+
CVrFLuhDMElZR9AMUc5oPx2JiFqFHlbIUokz+JRJ/9cMq98AlCHSKH1LX4LSRDYBsS5rEIMgI0c4
EAfWUFqvs8f1UlC7CSWihKJbsENCoFKrywmedrEdizLHQnvHX2IFxl0opYtnmJgM1C2THWUB7mDg
0cHebjSUuoKaSrwdJPUWEZI8wfSkLBsfglv/IzbkVgc35KY2InImEwkqY/Kvqd6/VrjADhg2B2cr
pCiX+2KWwksP/E6m7wZHz/BaQiDAHc/dmxacOjgBmOUw8MoSeOkna+HV5mzHTS8GWM0tsKdn8sjo
DIzevWLZKHoDvAhl4sMegprOKsLfA590cSpiQW3ryPclLaCPqe9O6pHxmbTgG37k/rruvzPDBcu9
hs135dEijbpChmEzjnEa6cf8JQ5I0s8uE3anHNI57qAzCHs5wAaIrR8NDPveH5Tgmxviq7YWLd6S
MP9YbZgZAT3h8WKxGaoEWoPy2T2CBuwv1t1rskTMp+5BArC8YvEgdqfXoOzvmJnSqLKCWaqtvaXF
EyJZgfD+L0R6SBwkZFwxxAyhC9cuvtzDKrmFVHPBWCOs2DaxgcKbkkPp6nURrTOqT3hq5gkOU7E3
WSabXbIhzru8oo/k2uDxMqjRqFQ+4nKX8BIfJc4Dr4Pc8xxEz4eH54UBR3ZiODdYPAL971/bPVfq
iLSakPyLg6Sg/R5SXGbMCAS1OY4dcTuXvL0F4RW5MY1cq850EkJqa/l6Q0zqkmcvfJhrBulX2p4O
Et85VemUNG3kntuWASBZQQXfohekfJZKo2J+/FZGmxVFCiFJUtG3QD1dLXuQWz+Tle/DD9o2yE3K
+zhObBwpWPckhtRXfD8tftym9SS8qJzVwNj4W6frNmJRacs1tjFhkKCxQCAwlZflBj2jXKPCorAA
7+9avfdYzuwytkfB5iFD3nqEnJno7/Wn8WGKPvbu97setHWJug15cHQKfICAwt6GaMpoqaVLSYDg
ULNtRbB+5wBjLwm4Sj2wyu562OCfAH4SQWSXv4z4pL2OoeTGA8O333B5FGPnTXN9qBb8iiy8sHs9
tE3J+BEkjcJ9Ayo+eOvZEIrmzAGLfyFOrAa9G7G5lU46Lu5M7kdjbuuak2oAjsuv98+1BtSoU3Kc
q+1dtLkMJmPYP6XmTRvF2ApWDv8dIpmOb3fGquQHvHo7eshgeK644Hq5rrC3k84Ddp+xYXikqyLF
74vxbfprfFPgXpXX9eR5es6g6tdhKwOreRpG9BiIw6ovhb8/YqV/zVXccsLeNu+ZF7gs58nlGFSm
0DWktjcBnuSA0Ou/pW1i2hKCMgKjn6mY3jvUH6Bos+rDpKmBI5YVxgO86rqXML7fMM0cF4LVHD7l
s8oe5P37ujsUKAqF3HBUHLYRo3XgDsYY+Ki0gnwR2Am6zB5uQOpScsoDE0Bfh82voTVoRTOSGuFz
kX1XzZ8TG1BFneG9hUu96bRxybp3q3nVMgkt8+ejfv/nb5VLjrbggf9TrRhFHWx8706zqJVaTZ2x
TQhOI1YvFSwU4EnJVsU9g9foQg5zbTQWFwhnlVmvu7+4emsfXJyd15yHEgswwfxQD4uTv5pT/PPn
jfnWnPoJo8Gj+qTbiwtL/hUmyKVVDNQE378QpI8pm5Cf/vkoJWB1ydUR74Kk3zxEaICTPxQNLqIe
T+w/LBLVjUHyaP68QjeXIbVQN2K2cNSfHYZBtwZicwHPw6p1xrIYuTZdrE83AfyV81wyVBW74XGS
V4q6OAreZcEKlj4IAjWAU5iu6QZtODToEfvC1JshrEpGqxZTwO9pJOuS2bRGwpUHCpJT7NCna8+q
yvuJ8cz57ZgRMU2WksgX2SRNe0nJd0V7VwvN9PRAl9MN4J4MS2SDEkuFWGU1BfHHLrv7/cSRh6Xt
QjEujbYEyniWBXVGDbX7tDpE1YcIEQaMJbnQT3fqTzYTHcgVx3yBKB+p9fk+tqtI6K/IfwqiCVbI
BtqOeWacPohYbnD8SYwmuHco+ilvPHbO1t1alNreWjxJTeIp121VOwyJIb3r4kbmF2IcrkJO2MhR
dSBbU7rXnSYSHJyo+QbaZ27bjGcMrt2qnV5f+GRukyiC3uwGiFBV/tYs+ZIHPOoPNgjljkBYrTVw
VsAlkMpSE8diYSmQRwEaRMLVEbNwdi2+xaP3FSsCKfea/86Rn7rFhOX8qZzGCmHQsPVUm4+lk3w9
FTMrGx2MAJ5jRFG3s+T9+3KXOqvRKTkS8SHoxbbvJFHScyspRwfwJpvWtcx0RjIFBc/EuO+37X9h
pk52q1FaB5mb+PmShvS5le/KQfDP8Qoyk+jQtfwpbyqeYor9GCyMsrpCPY6UA/FLFugOFCueCoxX
MDu1BFs7M7KPQhs9AVrBl6FLd7ch7D8d6uRw/hdVXU971fz3EEXs81HwVCDLlRgnn9rDdfdJwvu/
wLk4hEvcVDaietyke8Gd4fcfT/e9SJCiOU/1wk86/WYrtDZcRZiQEaQ/mOf1xEoM/vL4xL9pNfHo
7xXkCifFZ5ZO27kFQPsTNNS+5OjTOgU1xyvHbYCi56Po+XiIjCp2LaW+J/sn15CzQVDZuyjbJerc
U+iJEahVdtPZqCBj1jf0NE+JkpXO/iEb7jnYdyWYUhKYknTuJsn/LD/7AAYFwrAj3k9QvElsUVUP
3fKYqHU3yKNY6lrknsxza5r9Q4T37vX596lHlu1AJ8FDMxKov6brdUi1BiioYKb9nh1nXdNnYrF0
PDSA8NN95r/nVcf/xBa3575mXjOTXks6/fFILRwkteoK0NIBRcd/iuYz2zcmRDMpvqePlyCzvjY1
Xf4uiPYgOQtJYZUHCxsO5aPK6ZYp4+MGnY2JcO6GePlF4KBjvERY497zpxeSQrdeiqeO+i6X7R25
qVVKGchzCkspZKvWLD/TxkQnQVA/NFuIB5/OepLYfy+DTyxyb+ZJiKk2fVpyEQotzUd+R0M+6cEh
4rjdPR+lIhDztE0FoN0rOm0u0vBw6diXuOYrVyR3AZlig/A5ENOR3WuOIwTQVgeFitSlRFYoSOFg
AQn9xgTbRNbvrwyT+3ValQIfkGmtm69TBFVS7Nj1HkdHlEioIuoJ2AaVlKUNJAwXd8KzGQyO5efK
xLcUZk/bn0fmdrgsRwbQMWkRiUBTASsYW2rLK7s/2ulbc+D+Rg4XlMarUAjtdF+L1GNlcYgL3FyS
oEkC1riA1CtWVYhYbwcBuZJBXZ3kmuEj0yAcpCoWtgdlB/uUjIB1CIY+hnedkjy9dZJ4tWnaYpfC
ZoayoufO71Q8rWvT6Jidh658tDe7/Lae5d8reQwie/Fk1P/6VT1GcGhBRvr3cr6jIgRtlidg2tAU
BGhypDjAfxcvz9HEla4cPWc6rMDLVb7CdUOZbj+mnGXpYy8X+5tefGDwputz4tu+6lu8eSaOmXSi
XEvSSQNlhnbdDRS42EI1Fh3n8c31iAtTRDHLcorQHUnLZNmEqSnTF9y0fRwWbMY+3UGghijoX/0m
LAdV5njyBXFavSyNp5kbaH5LFfkZWQj9jFt18Ricy/1H2xPZzeKf0OuTBejbrHRjvRAdzFTX7TFV
ZiEXB4yfqeMcHUCI2Eg6D1dWxfY3y9GhJLMrRAH4Xsb4EdYcih3H34oeUznQ1JzljQE4DdLPIQ3g
yz/zK6m11tPkItWxrHm81UAVzjwCOvLfv3sQluEctqDhLOfQhUB8L00/wwteBfIlN8KpRnHbpGxa
057otLewXOb7URd3TdKhFjWfHm+w34jPTE5Wvzh0B44QkkhdC/H8sfcYxy5STn9JliQ+duw4Q1KV
tKfAARBz2+Iq2ebn8316VBiynPMTkXHtbZNFzN0IQf7tZe6XpDRj/dl/guo3OtSDq1kmvpKqP6jv
R8stijvSgkE8hK3rh8yWRRkToJxXg4AdkN3PIsUO59YYC6WYVtVl6EJoWI7aHGbIyJu62ei7KASL
RBg08N5v7gHRhOzFrj54oCedb1QXDUFa+vVsgR8l0O2GNtL+JpsYOw01shwiDvVH8qnVOB67DdGj
XYCZr5/BJmcD9hJZ/OGs/1m4hi6xCk9jLA3FQ1oAiceM0MZrmMz/9seECnYhbGko5ZxUwfE2vpbb
e99D9kRwI8R8Q56KkbVDqaSZQROXqbHT1nBej8WP61xl0F7MaJBoI0j1tzdy8Zm1NFJq6n1eyT9s
GUyjyTeIVUECNipDerCn05dnetmD8R4wbHHMDekUO8kojwDvZg2+j9Lm27UWqEkCzRTLZCnLKina
4RMjXXnk+JBlmjtCumBE5Vs3yt6qKzNBCMGFPZyhWaTTV+Otf6OpriomZp2MLbMildgq5ld4YkbR
aqeVMCl3hAlOjNS0yUd9egiAuvSAw+I15LWZ4qlRaQXZ10OCJsMy8vTVCQK42iIQkwZdC9unLtuR
pfNVMm/pk15yevIHGebgKBWTyfTTNMMWkj2tX8xnSRQ57gnCSRM2rx07YaXlWugXqJELs+IxBZv1
EPx3y3HMD9Dtg8o8t2Ye0Ty7IpGUWEQMwwZUcQs7lK4tV4AhKxTuGbXVJAMXmHUQTQQMFCEMGWCx
r5BhO9q8CERHrV3ZMJJWokNRySDVo3H3hyZ+Isfzjxq+5bN8ipD7ZGPJdtYJTLGtNxZL3h1otb2s
P8Tiymfs0K+hBafq+Ul0h8tacG9tmDKvsIjE38KN0kiuBWLA0jtzJlOL0KSGbZE7Js5YJbKlWFy+
XM4LZMhkH6nO2MZZWgqBPdC32Ro+bEZZYC6pfE62XKCBjVn/zjTN3d05lUTGCD4oYeKD4fDlhyGy
DB1Z/YEdWqo9gH4CwghWMRnRSbl3FK2FArt4VI72//9t61Gbf3+OkZL6JXRdBVk1pPxz9v51UOWI
pXOSGyyzirXkfSE4cC4XlNVYi23QLFAhFUWnJsr4Knc4jH3zHapp0W8NmzQ3pu9+iQBMFGtNMxHd
jWQ4RwDxOlDKvufdUDZawMFfGuoouiTI8DWpgA3Rb94C4znXcLUFMtqQ/T+KgZL/S0oHXuV1OFxz
/L3aXVutaqRrJF8eXCpyczaKCLLiHz6AWPRxigj0YvoYEYBP9akX0qPg9wsx5T4IdxDAjg4eP2mn
1IyKgUse5U/6XayzdAJRUapV5k/TqQpt0GdEa/JbfCPx83mobyy1kUYI3RC7djDNu2E6ATVQSavn
O8ftCkTCpKeQmJfIAKujzt6sI+ZN0v3zcIxDKZUqFl4AISUOG5fS+qYRLWlgp6q/7NKVAtPVVbyE
uXZnviPYSIrihdDKaEtqOIiNdQEyEJXx6Jwc/gnWdDkqpWfNiBPzlbQqaQjtIyN+chVhod5F6aKs
ogFqbJdeIlOWMdTDsvl06NPQs1c/c4MJqL4yaEqImRJBydxME4BLgNtynqerTlXexcMz0Qro7YaY
61P9GHL3RVEy8p25aM/qJKZArLNwjIet3DpL2WUdhWN41ukEtFldHYeTSuheCRZIcDKD2lvLbTvY
buzZlQrEKi2w+pno5hjFACq3521T/RIPyV/4Tds4n1P+FQ5DwTesXrofVAJn8xztnU/ZOzgaErRY
uNcJS5W1w4Z11ZIQYoDHdPOUo/9M4LbXY7b0XlVFcnFGBlocU3aPSKqhElc4Ro4F+enOh4BrxYVV
3z+jq9G77m2+1EyWvf/fdeiH++yUNR5BIRpb6oHEdkbQiZykJUljVPomsJyOLAy2aBC0Va+LpqoQ
DPqKuq8yhs1sK8rbAYVRrJHOYVr4czgkMPo/m4tlAxunnIo+hPIjI7TsSLq6NfgwzywvlpTsy8KP
VetkP8r1/RETWlrFCYychT+zVLhvsViSOuz66syBl2KbI38Gz68wwzivGRUyI37Ux+nF5A+4TFcC
x2NOXIEs84kxOKplWmHZsJ0dG+ediiCdTu2Z+cX0rxGwuY4hJlo/h//y3ZbDMRUmmHEjIdXlzWCm
8ONbsGHi5JO7TQaOKkyirh3C3QrcE3t92gTPtJNq+NyN1qJ1R2rJdpnhk9qfEeYS57lLym6VGXJ9
qP/XpK0nJ1r3l3646e1azc/KNTOCnRhRzjVmk3EZNUMg8Oakh6m3LPiBUeYY3KMUT7d99MCgNCcE
NHZ6PaxVbIwj5G1lon3/N5HRq1n9hJEbg8fZyEB3Z49sXGisl+t8B25evhhK7ThWAaZVN/fEHbFk
3egB5Be92oo2DVxmuKjmaUxChhWW2DfB3ADGxhulBPgMtJDb8eDwz5je9tbL7eUodz5X7jJeXnOc
12QXETbEDGWInyELULGHwjvUJ4lxXMBEB3IsyzXiOScDW37gDPV8OMBHHHXx6L551UOOzTu0t/az
b7YAXtk1aIFkEXJNQP0x6KRB9gUmWURtyrIX/Pv2hsr2q40uR947RWFsahdwRmvAsbzxtCMM5bex
aSiotEDc237XYDCJzzRZN5VKTZwN0IyI5HSe+vE1KMff+MYTykAlpdCIxjV1OYmET1W4WqKdvg5i
k6+P/3oSr7yPwpGGvsQdHb29Xv5PLeAQpHjqBKtpCK9VkmsH3b1auxQnuCKLoepTYEJi+MOtRNAa
JzKwxF1A9DBqxfgKrJmrF+imabaF1aoiJa01FEzUT5SCf0TaSbZN9y2/O+UkG/6Vwbhuse1ot1UE
beIhNjLgi/srafdbm9XYeitTMtvlm+28nL6YMAcU1Bi8Rt7beFYdreurcmY/1UkY8vY71T1WnbaA
EhxZ2mS7D13rWjK/c1+09upcyfF5iZIBUYpaI0DUejjZgU/q00sRNGzqdjJsMifhXNpnGbu0qKUJ
HzvioBkD0zNwB4o1Cf0DVbAypaa1e/Geb+sReLwV3YgTC1W7XnFHeBsWVkTBWtsDcxPy5AiG6Tkv
weFIN383OZYMfgi67HVLjttFBuB7XMXFxh3EIj390nfJVjxYURUFp6NWZ+n+IX9P0KBh5PhKyj6G
KL88/PnLWwANtnnNAIvG4EJTuArrf2td8cZYZ6P7b2qx/QDIriKSX14d9aI0BUcGELaykww+QeEh
2Gi/03th8s2pIPCstNTt9gBHdm7bShftM5JC+CkB4Wf3q1kSZyILkbhiZwu9wW4Tvg6OALGtj9Vn
2dOwW0ZkrwBNTt1eS6RccWFlmwcoNe+SaksWiU9l8i0fOkBVMyanZdsYm6R7kXOAHSzAMV/qbxgp
a7D+PbnEY2mn+axWvR0lWb6EXjh5rYXeH32Vd08zRFRb5dqaPz93w2uHAej3/YeGHETwxNhOSGlT
2+kaqSY2lgiSG9HqgCjP7+sVh4+NEWsfQJwrmw8vnpVzBVyy9TWTikr9ShKqD4HKLsVrc4oSFu26
t5X28OZ79gnuP3FXfF8ohg04UWiKD5lWo3GlXQqQ9xenupWAG8oH0+6dVqmnaH7fdWINvcSbDkig
fmafBud2LaUfIsZyUwqZHmLGnKIhQFrei2Xy5IalLts84re4mL/tUNb40gu+tJhC6E38Odl4PGO8
TCiI7VRzwuXDXD2+fZuMzhuzMFFk6nWe+0uadzfn9SfAd0aASF8jbEuZRx7HSMtJpgELBG1ZXqYM
EoBMkY9T6+SfrW5RXWjd3KWa9Baf6wkfpIBv84Y3zf0sdQuBWKnRz3B413ybfUWw+mQbwBhSv6/L
56Q+grZ60SSnDqu/vNAp7Kt2YI/NEpFduLV1VbMwILyoXWnuwa53G6+7orVEzZJtlE/iSCHGIXMi
48t98S7LCDkFr7fRQDI0Yd+TtOTHj76+FxiqtDb/OndKgOrntZe5racJIFh/mhGTX5bqzvmwJ05I
NFJ2XNdNhDZe9l4RXk6HbjLwOLZnKBebI/kC4WT8pD0noMfaEulePhYQ/j58jP5d70sW5REy13Al
eDGFuVq2bR5FCWKs/C5/qG+8RJNcR3jYvkBfWivNGTwoLNqqGSB3TNree3mfF8U9MWSADyroUVjt
LAOcgGSYmb5UQHujCCBoTJHfSxM1l99JssWEQAiX8ZBQQHQm4ykaTsWOEEOGKGVFXJArLqSfVsTn
s7qBE/MlKxZsEPAwNJN3CH6e+0qSVfBfphNTUjiAcPYQGZvzII3xeopOVRKShAhK0cyoKfUofD5S
ubJ0JO/9pkvuyqOXyzNIf+GneXemYxbiJMX61CdOPesIpsW066pxEP4Eq0HxIPgNmfJd2xezOej7
IZtBUe2E9ixRwWGiP/gsoGOcK31/uIjgKlpr6kUt0W4h1JhPwuW5QtAVOPNhMDeKhavMUijob3Ov
qDw5EfHl7qR2QoGgV1YBlKMjRPauuk4/fWavZMCETNW7+ZWBHiJJ851C1GRXSQdMYeliL6WdvyQc
dXOUE5+H8/9GQVAIHc+kMDKXLkl36XdI/vpqh6KSH77El04Bg7vHyMBkUim7pYTvREREzskxVoND
dTW56GZ8OL+R5axf6C9Zgh77XOt/P3tIxG9YPDVlbzvnkv0J1M4Zj6L3MuOC27LSji4E+7IYqnxe
JdVuUO/NEs9KZyM9xBGQSjNzNQYExii70qczbde6oq/v+u/xKMipyYwePIUzADmV+2BoTNtknnUr
by/bqHU0/pSTdVjQnnJj229UE+zSsSqnB5h63PiqsNh3PDgkcz1MvqeAOgr0EczuJPs+WltJT9TA
syCiiwRS5QqDQnwU+4/FrpzTraPjjWfQDjNEfj339pKVIODKuJ8UtaPxc2PlfWgATT6tOzZ1SVO6
bMsFdAEfS79L7CuoPq08W4/QJHgLbBof6e0M/8o7T+nO91R8quL6t9sejJfhrVntZWLcjhO/w18E
Pm/vlMrcd5XQazq0UyBWY1eRQa+C3nyHgbzisF11LJjdKYavYfTqzgOq26NSgdWwMkccMbNCQ+pO
N0aIotS/JlixH0NlhXaZTV6v6ls0RYI7617lxg6gkwvQ43t35cwfORBF5EZiSuMJlERCoQttRLU0
gVs9mSVEnzrfFcF0NSL7qXsRO9jhbzpnROplcqL9usn9T/00IO16S5+4mv6tWZkl38XqimKSc+NE
mPS4IF5KRqkRANKDsnZjr8yS0ltsJwLuywzl0mXr+x1BGw+LM7dkwKcoIw+45YZesv7bX2A6Vh/p
2KT3rhTmOPXrJ+ACxaq0j/3t+k8qPtC3OJoGbFnVXtrx1/vogTJg7pg+MNrlGVVnu6J5FkhWnopZ
BRI3H2o5jdsL8rOYT5t7uKecw8ZLJTXNQ9LXkXxvlfNcpMSo+hqaF9w7M19EXYNi0s71aWOW12JN
ICzYV8o7rpH6U+OPgcMHKh72RUCDgfyjQ9XMna/IxyGhicC4M1JmFtp70HbW9sHTiOoc7iMTgr69
9BL1/RCNLdvVGOJWmr1PfKbEGWfQznDAeWj/c82+WyMgapiDDesSZXMzELYO7Z9YFmnQcfv/pDyS
ea/BvYYuNLZL+RP2ooZqRj4q7PFB/v+eGEPBgtxMLzGPb2c7p6lvF1pCQGye/x0K5JZgFtqYhYV4
NCM9mc4AKwtPB41XqDZ71M8+6HpYdWaqQsxp/JOikciqPihHHFFCgKVsYHgzerlyjE13nbZ/RsBH
Q2v1QyjGReLdtxk6Jlz2KapzmULy1V8M5bzqG2hwtZIgAbaYcRO1SVU1J0e7PJ3RGYwL/1SEFYE5
VJv1/fF0RHUZs677NW7jfngWlkQobbqkJ05xUziuAC7Eo5wjxf/d+7uiBF+clRPN0DS5YiOXSKb1
HvojLTVZfgahIeePv76nhE5LHbAAtJ+wZV4KBI0eyXLU39/llP2fV21RxkHtT5eSmR7uEz+F9N0x
FV3W8ijAz2ALeiVHp9FSY0/19+4mGTP4MtNnaV9aC9OOIdQCcDxoWuTZ6cA9H5rllzS68Z4nWnPI
XFhjxn1WKHYXLx/aeuYH8WEukF3XzT3jhiqCt5JhOVjyyzOVltC8aqa2EZtdwpANSdWKO3GUqmsO
97lKBzMDksTnXUU78GW7wDn5/pSmwgaZEPKHYckPnzzPxKBmZkM8iTvwlB7m7qo7OfU3TFhDxjgw
Ti7iQvLAgtSdfkykvWMO7ZwqO5s2lrQTwjQLUQY6sjxL7slPb7TcA1Cis2n9qFJJEXv53PKfiR7R
/LugimKPysTqaMTo85jr8N7EpV2qZQ0Mh9juPpy9X9zmbJpjFCiy3N0VC0mQW13n2cABkWv+RNb3
iFwpatXHyQn+PdmldbvMDBmGFnLp2bdzVqi9u2INR/IupgMWprN5y1+3eisnhje8OsMBR7fMGLLz
3KU59MerujVns6p6YtSiuf2co+h8nRfSfiPNtrvXKHxDCem3iJMAgP3HvKujvtVvFGhXwJk8KByY
YHf/h9WlTCbtF6xyQzLix2U+Zqe8qFSYs4/ZqUSq2D2fdFNekDqxcplrQV+lQcvGaCXwcmh4k2rt
CUuSMPLPVX1SRe5qMrZCTAM1iLugftl/PNKjvErzC+Yn41/h5Be6WpzIZluTzD20dgoai+HMgWH5
tTkEnKy/7A71fSnc3PPu7LqLkmY0WJeE3I2/IxQ/yI4mZW/yGTN6NIxmETd7fj1nh0QoiaozoM+t
Pfw097zhFn0gTgaN6x5Prx0yT3aXc337rKGEcVKy3B0I/L3OZecE+RZxT0w53zK3IyweZu19NQNO
5iU7TDfjS5cCNtZlMSq446juduU0KVzWXeRuK6yWOaG+TH5B839Yfgjt+U5nfBRPfwlbNgJIBm+s
uEqHL5NPl9VMnsyoFxqHEgpCVMRTB3GFx8IZVukJzdTVtGNPf2rO0hi/PHHpIXOTbCCmCf1JQ/v9
0LH8AFUR75dG9tl2nacuDWjtbsTwM7ITJoT0NKm+nF2uTYMX3QNJCo169F4++i/N/E/yBw1smV2j
YTCf6dPpm/745o6eQjdem7Ny26tNwAYHsQk9tE9wh5pUU5ysHMByGjcAC/lYgfTItFbBB04uENgE
EH1UyQJfbuVZLYUKFAFsA/czvA0mBZoM0kqTeIXYfNItoal+4E/fqt2ehuDJcasGaQvUENDZT0b5
dIytA+rq6yMa2LYAWKbG1m36HZZyl3aiOLlVyC4WVUIxaabo7envjEEVzoVmNK2tlQdYsmSDISrL
YUnU1QBk7aCyYwateBtyd9lHG2bLsIiOKJ3K9mRYBdDgYvoj0i9GADd9w5QXxEXmxopPyjyjNrdA
k8ra5RPIBp3VDElSZI+/qgoOfLHBYW2KwjlhHJhV76MADMuYf43uGchUEExQNqO/NG4iBoX6FGnQ
+ng/6104iUMOjipbtPL+DzvadBcATIVLdhFOW4U1+xPfo+IVXpT+sTWQy1EYhjv0buB/r5L4c1gE
6FdF18Fiy6I9qUVfcYQeRkxOn/1gEtF6dwbJsapRDP8N5RjK/9eTRsTKi3deOGhT1YwDhHEBv+Y8
FJXjkJGUjgP/Ipxy/RKT590zOmuvzX3RdrMGY2ccK5cbPQeip88vqSL4kaEXWkku86SNfKE5sWWY
UPByTe5BYX6DYGX0a+C3iYzeTCrN5y0ApbB2fO8wybaJw43URD25Qb3EYlZjeLeXIwL6wK7SDUSx
KLUNN6BswMzS2A8bwmAHy0IZPvA85k6sWN03co3Cvk/mjKCrQqXogT4YlkZaPDozYyf/lXuRijti
78UUZmJU3RK1oUx4FtGXeJ4TZjBfPtGIEDkpnT8TqACcZo4i1trRI0wuZmUVpqPdO2f7D5rkZgdE
DqFqjupoVOHN9D2Qp6GhbU1Mu7FftpH2+ECEA3LdW01xgtP/3OQcEjEkfI/DiuqV+Jxcu9YG+8eI
TB6cnCm9W0pIzgljZ8vvCF+KocasDcH1Gj2bI2/JjXC6hC1f0Dy4bQtm2BSQ58L6pf245h03HQfm
rqc+NjSbCewIw7F5H20Xj8KcMAut8r3hFQH9IJo8HR85R84YMo4jq8S33YoD30h4hQdsXqsw6sAW
R9QwIGRzOm3GKNn2Qma4Lac2syBo8yVy8fZViaVlDs2OO5m/XAly4U8yrKM40nZ7SpclYMZoETTM
DjXCgewwVd8Lo93m/9R9vBKsRN2OqN7+VTkAeTdVYzXqSBk8W8RwMXb+BIaOxV1bgiKFzlR5bx5W
wVIJHjOWHIYTBa/LHDydg7dQCNX/G2qwuF9e7JP+Y38CBryC1OHrzLEUeJ5yinPtnSHzjiuQClZp
knIuy19GGApu5HWw3+Ui7Xv5wHl3PVe5Xtr1eOVmCeDWD0jA29coFjXnzD3WaLKuRbaxtkZmqbcd
eLPCFeQEH4+5+XLFOHTIh03nQt6/z+ZoIc3mj/wGmjltdrFfBmtCweoJuomK4NV5GDqWpu/VPP/u
cRto1nG2JDxoUDxrSrkpamspALncDv8q7fTaum7pg9eNIxjbt0w+i27oAdsbi42YhQXEyAo2Q7qM
CctIiIG1GVQ7+g+IkxJf+9b+4iPokZCD7lDMKN2UwEci3tziARB+CjAe1zeiKyj5DU+mqWBLCrbt
Z9ruFdi0OlDFThVNcOswzeLnBaHZVYNEh3HhGQO30SghfULmXEOohJAfs/7cWQiGlLYgIXr0DmYy
6UTVZYkSWjVh+UCyBizlkzTSN1opFSsUdfKUBHUm5rczatDbQlEYZONoexC7mpvOZDCf4/Q/mnps
AXlZDl4p9ZvU35He+OXfNv1h7EWyAJwDrJoInLMze0ZlQODaUvlkHEkxZyw1T3lbagQgqSE61w4C
J4HMkCJbPy1ElUYtDTpi4yuJWfVNk9We2yUTcgSY6gVxWFS7wP5oNOPcJDVcnyUwi4vM/UiO1mhv
hqW0q/mRgmghrXo2FuYvpZVH9kPrXhMC4Fek33DxAyVndBUi5/dUK8frDc20ePjsQgg4sQMf/nbv
nFCq3ui6UEoNE8qjKy37mmoThpaq13nL6dawy+jO2I9/s4GOmke3RF8s5h9jd5wwFC6M9l6fO0Hk
B84LV767razc0pO9y1vPUPNSiYPlXcumC189eihRcswhm8kDIwKyAB6E9hL1akC9alNfu+j3A+0l
zIWbIA298gdSY42opg6wU5WYpNhgpmHeRX5CoN/+qDdzGopELC1WeAk+Ap74JjdJ5TwjgSq+7H66
6pLyG0o0N0H2amIkDGv/pmYqmslfghLYppLamJWyR8oTuZ49Gyuaj4ktiSrSePZ5TR/LYKqcLhB1
37oYhis3BZZJUqFI7jb+muICwz6Ut01T+JwXUDAepLXBkky2qf5jXC86uR5ClK6mR6M6TklIKzy/
H+EAS9nbDp/AfDewBgDs8HMlhISEx8bq92E9XZZHt50djwSwcBxuEHcBWcWb4Qn+jimBsI7OInAU
7pJPTwfBD9s2LGXi5RJpgdGXXGDo/pu4OmXvBxL6Ip9RkwIOD0GiZXb1M1AcfS3OlbS+FJZbypIy
US2OhdthpQu4G/cgd47+BzfzXcWzs3dbRJPljESFEKi7XpFCB6DxrnxRSdKCxBVbQMXRIKwgsdjp
MFC0c+BtBerWQ0JZ/n0MBkXj98eubawZLgkmQJqotL/0+bBNdvkjiUMrxlZpjMLnVMoKE9ox1bZT
UClO+HwxD26Dr3iSiLrstzxOOOuPaSgXke2NfS100CZkE+TWAphCMqLVOSnhr4Jwnz+eMuGxBfEw
XrrJRHdlGb68ZHO91sU275sDNZkaU/sk+6+yfjqGx0EoK3FBMXVHBXkfUv3+4JcICOP+vXet39E3
FsIQ8INvKOcxiNFyFGAlqXId73h33FZX74L+QNjPitMHp4JNo+drhISFV/sN0nHDg+Olai/DLsDL
Oue/4tWlLuc17ri5OYSMkHBI9fKsPFeSRYfFL6NBdceZaZnt/6omLfnm6X4fPMJ0bXapknjIVeB9
FodXDSfczuIRmMXDs1nTA03i08FVsVz/EJA2rxK5bovXv3Nm94iOCR8TkUVXnarJBY7kH4E6YDcT
2IcdUQA5VLpa9j8J9q+pDTdmqzRq7Hd6XL9uaJNHfQEhqZ9KXwS5r4maGPXzra3xZK4QId98QILM
niX+8Q5dhqOxrwLWTcpLtOOX2Qmh9jVoL/bZz5SPJEjDNtm6ZARNHxIYZuG8CTEj0mhbqFPcyvby
1uMpVO3ppOqKcdktOzci9vHTC1NYlqlmOwNLp/bscvPoiEB81HQoSaAm1OwSMKZYk+Aa2PYDZ/Mt
eMxOgn17+ZkGu7fvondcv7JHycESRgpXDFF20nSUG59YdZEzi7ZHttwnrvPoHZugK9aiN2/xVn1r
DhavPoPVZSp8xITN8i7x7lpQG5KV2AyV7chBzg1L0bVNdUTOS6H4IN0pvi4ua73O26yJheFGzOwg
+7ZjfxXzoJyU8zUqmjIDMGDVVbH3gq3Lg9Zxj3Ri/XcYxDNoijdQVeENfy47rRE8eXK6XAfBbqB2
hYXxGO80xH6C5X5Ni91t/tXMlsuukTWlV0hFQzZhf2RrG0P8UJgu5AX8KZCYMk8k3aOVlAFegPVe
XVTEE9KEe2uBxF8rTtboVIKAgLR7nkUpf9ydrgZ8LUljHSP3hXWmjpLlbcuEAX9c/xVmgsHP9wre
OiKrQxLknzj5C3a5VoogApZARs59WPErPqA5YK036ATLX8LIsabPdS5P4RDQubcz08wdVyWiCrFh
VliKHhWZR4QVg+Kipos/O9uKE+IVY89emq/Cug9PconHh5IdCN+rGlMhj0uCWkQCBhYAxPR3gcDF
PVZ40yuJ0BmLjrzFRFK80OXwZOQZes+VLe8fwslbrMoTxZ5Ko/T9fo7N6FvrxEoNsQOVftmxsz76
+1OrhW3h9zJBzpBCwE1cZggqR8ar/LsUTvwEoZjxELcR2mMHCcwwCu4VNvcjRFWq593qaBaMIss6
yq1XAEXIS0CsyLKD5QCWSaa1LghTDRH1pTUa7lJ3uCFF/r5ptEvqUGgM5HLLrlDblWb9dwko7BZn
uVtFaED0s7Xds2U/KgKywzGLBrs3GXn9GyAZKLwdB9eWRdMC9nMPKAziGzVb2FKfKpu+75DTuWaH
sSLM1XD/TDOypAIkdDBgLPg28pGwzw6LHTksvTJSzdGi++pwXirszBSeHaPoQFZ0eJk3gSJLFam9
Cto2opGOkVjE1Mmw6JyTH2ee/z1t/W4LzvMrRN/lHE//zugNXYQ2t0uilR7i9K2xhL9PyNlwgwPU
pWqAFzV8H7X6QsHr4ihu2uIxa60UxBDs5NvCFUeNbLr+Z4t8+4ZhaZ6uOeeg1i7TVChMIpi7/Sbi
Orw0nfjejsEf5I9uB0xpd0oCYxbCUmFaKLwxSlQj81A71XqLUKgjfjHSb1uSicvEKZs6KkU4mf7P
T09oncYw+J3FiqKhytErMIJzgr513W3qEjky/7voX23NkI9x7syPKcBG1pW7oQuKTh6oyO+GVzmS
x/LkJsUOoZy8kZr6NLAmlQIh05srl85jHmoJpjBiC9/O5cnTQybrOP1iidaS/qtcao7gClcY6XJW
CxrMhZW10lMNpom7c5EFu4MKnoicx68LikSUmg8mQFOaVZdmkuMytmMzyX2ucd8woVVeY4TFj75d
h9Nd9kzlAT5Dl80kfJHndq/92Bsa3wpzfFNTYwMWjiKHzmKJ7E2tOgUPSSKH3k6nlLM+r82OfX3c
6KHxvc2bo4FwgXlB09Nn1em3d2PVZ5Gamh+JkY7qRQI8rfTR18NJb6lxNR1IQ/2bKmBZr+2jme3q
Z7Vx1zbzi4Wu8eq0+UFtO6iwfotS6i+qos+Tlk1bPIuj/ggqX7491oa32Mr3240tplM17wo4ZBpT
7WEoWtelYMhUxiTzu1W/rPj6BQ2uQLpJMT850O4K2x+3YovcarV1BVP2WXCudAwrH2v45apxS5i0
LBgRO1dV0rnHWzlA+WVaPjUCiKSzkEcap71TEI9ueY60w2sNE7rB6kRzG5PA5mEl6ldvMmPCw/qG
EynQoGuRrEK0+u3zXz6k+MJgImFsksM7RVYFCpPwMrNeOnWelXIN5C+70L+lUnxpkY1uBFGJOOQK
RbVn1/JkC94UVkrifQ0y8FZgUihuxHgvXHrqINtirfvAgQ1wRAAPNm1CZrFThhwaHp/oaj8e2Vgw
AJYHO5XaYqXQsg/R6ZOEtzHbHniXWPeUYFFx6ApO63k/mC7wrB2LgjC5WLsoM15jbUw8GNp/taJQ
FFsoPtKAZnzcErAnUW+wGhnbKwJIHhyn+hMIQrpxxo2z6ZPeRhTN/oIU/GwmExZPxQfctCQRxgcd
45pZcOESH6q98nwtwU64AbTtM6/0rsKKSCl8bgSzF3RoKBjfNIpSPHLAhrPpzygbORgdIgcb5+dr
wyxL2ZAnMzoUJgTwnGz/5cah5cA+9p1B7VSCAMcx/f1b33ehml/RrsWHmh9N7w5or9Ti1MZDg/5U
hIfrJ/V96qr28EzKpOYDiH77SNELlaS6jwqFfx1TXrgEUd99kJzsD0/tnwQt6f/l69Ifg+ckIYle
xq107T1ZuyshPkQIAatMtRsnADi3mwJ+4zcGuGkBFHL0OB7X/9sonswIF7OezcHoInxyYi5k5Kwz
7Kc9oEEgEDAiKbhMqQe8eAFzs7CgPsQmF669HcSf2oz5si9yhCUI2+8v16j1cXfSpl6aNhIXS3Eu
D009jv8DuUHNkBNruRWX1NZfYmn+Mmcwi7S5S0fd8rpDneSs4A/itj+dgmU+tuEW1+p1p5885yPZ
AoGNcJa8LMwcW0nY+z/xUUbeN+7yy0+nUuNJocsivWilU06vOgD3cl8LntcXO85S2mI2yL4URkGO
1hQ7Jn2eg0KmXjP7B6pDEGdnWndCaQuIiNazPXBdZ/a1jlMUAbfQ+AUfV7XQbfo79xPJjzF4s88n
PMjZMvgqJeRDly7GM8kX/rovrf0aBYGhOo7XRx1A3q2aWY7MeqGLCB7R3SisQMcd3slqaLXoReYi
SD4YUYTvELAoBsfJuRC+86bEcWZNAns9bHw+Jpy/FOTpasKz1DmzKfg4qpXrg30Tc+BHpd/y+9Rl
LR+V2Uh/mJTlvh4n7HeG7OTioHG8SfGc6ThVtECtSeyzBVFE9NhJzzXPMnqgQHTvkarCrJ0FOUc0
gOjvZ/FkSuzpWGANfn8J2G51ajbs9/0Q1v+gp7zmi5uRae8RFu13ReSkjLnV8QlDMxYSaApbt0Gf
bQwyvfSQsqHxDoboDtoLUey5pQCKkDAfUNImWdG9PlciblzVL3GePrMw1JqBTy4UfVGdvykyifen
a4ik35ahuDktuwGtJS3Wb53CVk+X+GcH9FUzAEiEGT4igqSJMvxuXk0/JLmmEaMjyObkyf0UL9fa
Un38BwO+VQedxaKfpLdAh/uAdOYVlMLySC2IXM//EYkYrHcG1EDyNpqgb+NNsTcm9uf8Cptz2EsE
DzTp46IKn9HAoGvRq4066TELOegkvlTjWES9Z7euX8tHlr2q4b6w9YNgdOzUwM4FtlotPN7xTl0g
7S6mcNHjmMzguX3quWoZ/ZXwXcf/th8cP1W7UIKekGUYFDwm1ZHw23AAyDoondbscNrlGYeOyEhk
YA4ezRmMN/kulEowFChacJCZw46CZxZp4FLtt23+/3Nx9H6Btyh68+VlYbW9e3EEbASrWa/5C46D
WTh3x1hOTUoOJdoyxLYaAQCJO2U8exMgPYUnUlJd90LgGGHUMq3m1tNMgJfUMz93uJtBe8uTGwnV
+WjRuUmgyNLQmiSY4p0GTnwXYRm7DHbxd5ICGcxggxH4M74V+m8dUtKYCT8sfHLIFbBEtvnNG1OK
Fvq4dDuyVym/cU1/h0QQUWkE8BLLnE345j6t6VyQJ6MpMwICt+F+9c7O8uGEWMPfLHTZHAIo+nx0
5Sfcc4hPTRvdhqhVOVNygT8M+vQQSHc6qhZfbEvDRpxo4iA/VaUASoeMf3H6T5MMYnGJd52y7XQY
1acQ7HtUPOCrlPiNQakZRUwriwyKsfGeacRObt+ZQivyxcC1IWocEsj4h7fHXtGVIF+YnV4KphZC
dk/JQNiyHrw8sqtHlU4X0XIfhO5mURkYcgPidiBtz5Fn/3JieXJLxHMmoyO9lq5LnEJmWevnWhAD
hDF2vcWX6SMypWpz8p4kUfsPLL7IsoY4skkd6lOgqM/LKEBLBEyVgTqLTRubMI3itPv/hokflomU
oNOW7kk1i8vpvqsXZ2vEqxwnOAod3xZBALDAzrzh5Kj3mn17Crdc+bvwxRjKynn6K9RzTMtZPIJ5
KkxDyVuYjEoTJR73EeoV2SrWmXPbucdsNpR6sK9MV6vdMVqPTuw8Sl1NXom0Kera+Ph2go0EH8d3
XeZ4WFqrnJyMzdWFZ2OGp+Uo6YM81GkTsValo6U/nPhHW6p0mu1J7c360q4CqrSv2lSohqArGexo
EJZcGmTGwCBAAy9Y8kH3V6+ebHJ34QeOzsL0wGfHzqLYE94Ync7tsA9uV4Xum2YH6JAXHiGfBss3
MJ8RYceT88Kb493YMeFlgpglwjIBTzQj9YnwyLfq/r5defkgBnRe6uPd+Dzdtow+qV6WZhHh/PdJ
mPQocXPgoik1XO0ycOA1gJK9DFm2PuTc5flyjKTcYaK++Wpg8aPsLwol6/qudKI5SAC6KtJHaopA
noGIjiEVj4BVEctf3mn81MOVuPqkrYIZHRaOfKNQOl+rdM+IDGNOimaUOxj881Orx7as7bgT3AEX
SBtD0qaRxOar/7fII8HGcVFVf0r/fsr/dPmqtstUvEdfX2v74egTbtAWzLhH+bXVKg9gC4FYuqOk
jx4HsknvHfJ436gWi/zdcxkHZRDEB1FFlvYnt+xDEFQAGIXqOs5DgBNUxIbj7++YVcDgTk9+L2MH
ur2l2i64xu63C38DnCbWpNiJdJULRUN3mDSGONv++JRcuAsTyu4/bVeDf9OjYkC5DJLz1Au1B2pi
Vkir/u/+1Q+7AekD+1E5fA7Bv+/ULmQcgTYpPhSFDPoINfRn1CkCr7zu84LhfulzWIy2gM6vLy2Z
LhV8z/xO8K0Kn/d6L1zrzBfJ8rkyAMVaQ+GU53alI4Uzspd3VrSs5EG98FAEnkgBWfBuHcsnQ+oz
WlysENQIA3EphZ9ZaCAS71OTtwLMRNGx9WKQXLu2RPfhYlMziazNDLGeqmHqFC7r22JmXduu+TID
8OAmiOaqYq6QATvrAZL0RRfIJwN6VtBJaHj8kfUkSbD+vRC8w6OSeT8rkoQFzSzLFIx9yKZDoLTM
iBYh4dZc44HUFFQijsqFg0ysXlXUkkwl+3VsXxrLOhDP3bNFLwzoUAwPsWVPiVPvnNy9x8wlguwe
ip/7OVMJHNzVXpXmL9+HR72DGnM9qyPZmtzHNyhWLgPYTLCDu8k4wvlDiwWuN8nK7DdhDwk2oSt3
UHYnGj5MsESrBtrclyI0icrYVfRlH0DkbCwiIngxaV01nRgkyfBaGtcy0aNT15Ymdqg+myhxb0a+
VOM/Ou62JIaEMdWrLKBPJlZk3te7A8bsWxD0GZ210ZavGODenUf+LsgoMYBb2jzrpgjYEn458siw
T07Yx8ENWk70jolsqwJyQr1kMZRMzxNYa/m04l/Ao8MlHKZZwYQvnwJma9Uv3EUXwe8e4o67YmZY
Zd/qT7xoVQ5lXGDNJVWG4lvfLzxpkasQ349hnrCnny4IP0UmZ1YoH+ezPzfaqq568WpwzRn4xraa
OECFauXmu2EtCIU8tEh0FeOey+aYYwgHtcD1xXR4WuhbgVr27atDmufnGojFYKupjmGKca9FmZ1k
jMiOuZU1gbGMDBKwrG3v7/0dhXRI+1KEXgoUCRGGXpKRJdzBmLD9JPb94q5kCXGuzRW8TsTTR5YP
U8+EeT5vSizezXf1XdMQO6Lz1Nvs35Wv39ms24xFJuJiKuNaOXSAqgeYkxKXu79et1cjFxwY/TbC
VmEOsFEy6ZCb1uH5PgKyG426+Gvw9F5imGqyDMPFI6WoSmENg5dsDsSK8AKVWA5+d/ptg3GjvU+z
/jpIikC4zo4zLO+OY+GU6yEAmvEvy+E5d6hZ5GdytZXq5XnHJ8nAeZvtIRMrpeDu9KkfV8NkO0FS
Gh1mBbvXy/o8e8a8cj0wqsrcbG1sPZ5GC/7cxtypqFqrkmNx7Aw2j3njz0m92cZS6LbrOFjJFhz5
wgjoqiekxZ+B0Shztd0fK4bKvWvxoN0XBXTKFy22l3ctAie0+NI6sAAt5ac5z6HFEXQfrR4ciqHL
j4deMh2G+2jK7n7c3R9Z9sL064i+0S5DOdQZx+DZzNTokkOy2XepQJn9zkEB7zoaYw+0H0nzJ3LE
1cmrvC0HJhJGoEyKvrsSsQqJmg7HMqbyWGeBz/JMPNM3ukpnsuM5gylOi9dazZ9Z4RbkjhLVmr/1
uNBNt1wX9UwhnS/GnAm+kHmMU+0VFIRUqmASkp8bMrteQ+SGew0ECQTURu/4ZxwBPjpK0JPZVHhg
aVDr8c5WOoQ1kLhN3h0NRVsohkr07dnpbuqGC3BRg6bUlMVca571m7B64e/5fmYwxFrcUx84+EW9
OFDq1FLSPSP0zAMOExvTrjiS/pQLlqYJlKfq2uv45EnvpQoHjrLzV75C49rocVeWjX8UkVXxd6fH
wsUr3peduX9d6LNwuDUt2OfIppRInA2G9G5psY1YkrcwNsyrj9mkIdLrjfgT5MtLdPQDjzl6937G
dxV6/+7qqUVP/ZQfLsDJkTJFtar64xhfxlc7ESz47wqKQJxrvrUMlfv7O9kDYXiXFPxk0hE2M084
uYX2xgkv4Nbh+SDverR/yXs3vxwqxbWGFlEOIhDi+Ril6ZYTgJyyXI8H7DoG6OiVVqTCNxCafrAi
XRpwz4D+e5oYJ+aGym5AV3LqzAWsVCTFJsGJKGx1vjRF32/d7bYmZMF4IQ3GtpfPHF776IyjA6wa
rA4Q/ri1+LA1WXqsh+fghcScZI9F7jZvMsGu019wNhZH68GyOqefmqLWw+SsBb3b9BfMfy/KiC69
cbm4ouTA4CczETObVTy/C+A/Ix2YzHFRWZkTUjMIUtPUqwfPCKtcXhkWyQ3M65Li0kW0FgSgPCCm
hEeqZNcZXNFX6rqJbiJFFNLUjvtnhwEcR5ChMQzdHFqX/B353s6W/PZpShKRjdJ8ei3ktkgo0s2J
L4cQk5SF9mHIzczym3UVAyoMVlZB0Gve7WVNyvzjwweXFv1BO3Yl/NgzIkhlQLJCJqf5L/fuXROa
XLs4ox4yclBRbqrzbWyzqhSnbsDEkytq0c5MwN5KfxaKxOfJyKGtyJLXhdmsL/yi3zVN0pGSqhgA
1lyOu1oxUuOLbJxmXA4QsTEJo0BywjQsAwlFDzab+w47lFeO+SxAyhvGSJY0ecjOQxOZ4GNYci2Q
/4961Mub6MN8B8qPEG2wpPvqufV5dRK6wq7DLW2Vqtp2zLqFpUAtl2LwjK925lVnG8QlcSAxaZlf
o9+2MMJPrx4MmL/1f1/BP5DUq+x28A40NORFBMiR6BYXpC0krmv+6Adg0ZAJK+fdLlIMNnfZYfoe
95bPbVItaKAh5Ajuvxy62DUT37JY2m1r5eCZqoujw0dD63V2A2znCMemIljLm75/v0gpANYX4038
Lh7OEwP+wKxf3JH09KmSUYfWux+eMcGMAsxZDYzq+NOt9tfbf8xTAmeQDm7a9/uFykqdnMgbTcQY
RUee36YwiZxvaRJhcF/r/bcbemGuQC8G5uwJcfK48WkPRmG7MRdbPfcEHoJNiWP5/BUZMQNJ8FP+
UYXa7QVpCwYi2pJG5Ku6bI0KurXx7aUDrp7787bV4EbLMxpqx8mokDPGAyUzWOYRDeqAD2ec8afh
HFZTg2iqyvzCouEwKzPZg9cfjO9odoGYV8eZD8B6f8boWAHh1rE+2eOs0kqeFak9mJgtjPqAtk75
+Om90b+OOwdsEgZa0JlQe3vqXn/XGqh8sbR8N/hGsAgLMcfVirBRXERVRwtvZ2oz0CrOEh8OSHyY
gkxuxwAkxffD3w/VJSf2AHdoYs8I2axVrdGhk1L5WffupmpECQIm98SWMppUypaaHwXYHOUA1ba2
z+iH0eZlJiqdG2qWi7WMDKC1z14bchhA1BeFqYC8Z+HS2IOLVO//hMdIrJ84DZdo+2RR6jHq1mKL
Fu5kuTlQxMgpLjPP0YZ1OqzjInC5dfo8OZa4rJ02xWqJm0bxOjnxrTfNgRcJlPYd5lNsk4LKkupy
nd+67thbmpf4M/8shZjaODQnHqiay9WZgzazv4kL3Zz+nUA7FTSe94hCGgHry0VBcl//RPArfjCG
bFE0MGxQsL3IfRckAf2iU9e2uJIhWPE3FCBPi5kXK73l8bbvGQcgW8Zg0QmvG6DhViGo2dmar+VE
tkTg4aGxtnFEGTJiS6a2UCPvyTs+Mx9AhkEKlD1rnyHvDQ8vjc8dC1juFbX1ENwQ1Lmpg4BExVoT
43hSykEM7h2M1jo+YCmn7ExfUHj8V/cdvUTRtZdU8oxi0KF/Ph/+jsKFe1A+XIuE0hoZtbxJWLUz
JjYfxAiJlxEnDDN4UFTz2RAHgGQVGuov+Y649xwI9XvalbKXsOgdz6uBGOPIATPkp7HY+4qR7Y8C
zyonGimncPmg6ggrpB3iX4pIdRuyrkubRa/izrN5/+/bnokjzhDH74gYhiu6/Z4vkB1vYXwb1sqd
kxBDKn4KDK4KXswf0gtr/AWnzmRJXnc8xE9yzmsJ9fjRevIdB8/tHNy4HCVNPYMfkJjvTRs7qzvk
QiKjFjzwTXDG/49LUKuaA11gCy7S5ZTa7foeseOG/ch7/BrgQ7jou0r9aJ1P+Jd5GIpChAkA5F0j
Y0lsDfUh1U5kYr6u9b6XVJb1ezUYoAm15B/Qyu8uzEps+z9FIJRU2ul1uZiXF5a87IVuztB8hs61
f94unRtKW23oq/3WlGwYRZgUpdPyL0+Eh6UcY3CfLd1DS0CsBkPQk+Kf88wEwxAqkGpQi1WmTzOM
AzY6fClN71Y6dGB0DhpdBj/lpvE7P87YDefUxVrSXTSIrF+pn8c9KdCeOgprKEgVi0tpQGTTwtFN
sfO05DPUvqVGNjiwkLVo9GckY2XRZzdEujeI40UMNHgzCj5Uthlk9KDGZrTlXP0/oExUL8BDe9yC
I8UEFz3FwIDUUkR9AHM/IiratdHjUD0P+PCXwNToweLQDLfnFOv+uojWf8O0vIKZIWs1GAp2cwXe
mFPrKsnKF5uX0S/FVpBLjdBWYkhjM/RXbYhobjk7adfcZoDO5NV6q5cU2+BHIAd1+TqP7wpCVFBN
VshqyA0fLeFWN3XUFqtDSpKIeqF4L5NWusH+rOuhUrj0MeRa3pk1Hf9N+O4ZO6K/0Bn/ABtkD8A+
4vW7A0i7xZKjky67hFgz9FYgxTuskMvYdOPGO94WkpYguF22lmfdg7Ub9rULooYT0YF/zSHZDQxB
dm0gmGA1ciLGIp8ZCCy4ES0TkmLGMHKptYx1XEf1cWfyJ0S1wZp78PZTYcwO2fvbXKlIJgSpi/Ca
ZSqkTs1KTHip4nToB4N84A5/cEjRJGQErJI2YAAYMZxTHYJUi9S7XalSL3k5sApSuaGRoZhYWHNe
lSnsQ/6AG65EmybbAV5REiclID4SVC2Lgb4aNWDPd5cR98GiSUSmqMxh0XLhoZTyWE1UH3b9E1L1
4t2wX9LL+7AEOG9++my1mNBuAGgQ9u+5RBpY10WjuPvMe2oy9A6SNZEsi5TQJfo683Ukkrm1Qwcc
SXTsN1+h+MiIhopzVWgZ0xTaYTu1gsG6bLTHoc5PfOSbtj0iqeDcy5Pk+AYjNbpN7rAfjxp4IxRf
qrRDurCt/lt/rl+1FdJ/XDoEIpZF6hUPr+OyyW+kPz/flLy84t24czwkBrKTHosKmov3dF123VSc
9rFarX65k2JAmD8ADiU/pLEMdTuiAU0WrqIQf2HtmC9NLmm2zaoHN+T/a443w4TQK+if1QTytD+H
AdcmmTVzDaIJ6PopCKsDpeldZxnv9tkUALU7lE9uVzDNK0XBhJ0zOiKwCf2j8l8xz6wjABXXg/as
OmH5HGqjpmTbSaEwyu/lLTyGqxlEqF7DmjJmqjl/eMv2HJ2iDhm4GJAFB8F0KP37MAirY7cmYTnl
bqb+hICexh0khEXGCNp5NiUGEqq8Qr7/+yUVrzMZRHi6WnZ0CCDjCmCUfOCFAHY8pdeEaAC3CU9G
Y4oSrOWhRlZWs23KSDSVidZyDehi8VTCFdb6A0vqSfHIdRehwd73n+cBWdBzNMZaBy/o/a9PA985
TYn2BbuzI+dl5sX9hgIZhvsGOaDvlMcGN7qY6AM9GQ5yk3j0reclkCnKBqmcPYBwVVBaLYroPZXu
TZn2d/qZve3hlBYb2+wOK9l3Fqw2gQercY/C703WTcicZY3cn0ngAsQCJzk/CBtbmasEzwPoim78
jOGoIduW8mS+qvb647Rn3Lums7i9vfM5ln6jC8DcN4IFmnZc1arhLXFJPihuZsFozwnoLKMTtSNu
gzKa2asOLcj2wvsStyicPiamdSR/YA8QK2bP2sBpk/JNGrp7opeHJth2G99gUNa1RyoenF1Y8+TB
88wl/Pvx6jThSVsZJr7Xy848YuWWsohYx6UCHYkITLY7JA3ps8m4abHazaIZpSf/gvL0Mo7BnqvU
g6w7YtAF+iaXVTKCJQkivGoxjm5J8+LzV0RHQ/vPQkPOyevlWzNfI2AXNBERfKSc8IQpJY72aTPc
igTmQOL0K0Y4TF9OlCJjt7PZ0TQLrZy2cmis7ZpsGt5knWRyEmr8s0jf8A+laYxK/53RR16VOcOn
N37NrRvd2ndLLghpE1OWMOFGuAWT913rITlXps5nXNQ4yqQeAM54aHIAe0Z5VYl2/0zZoFLCjpqO
IUvAeyRHrReNxwAeQL/1ls7JpSP+kmPEI+v6G5uMSVRcVKBiFp3ya2xyQ9Dg/lX39ojlO3HiJpFU
WT1pwlfPBTjrkZt7K9f8gWzh+lF2cPy6r1UE1RZPA9MuxtrEzoXWOroBH6cbrzV4fkQh+FpLSXQQ
QId+5Fd+ooIM7lB0OVY91hwBOOMJ87b0hWLAdEYeXspoHrvTgsN7vRfsepJggOcjzMHQOsbFEPih
HxOfSiA13RR/iCMvORuYiUZT4Fj5FSEXr7siADUjdRnmKijbWZXFF2IdY1XocD0RE8sF3xY1oOW+
Hj+wyPllcrhd4kz9c+YUnd+1ialjYmfnPrts2qGW9s0DtvyQlcpkICn8FXCYjXtcpDp/tXzwNOhs
eMVvLPj+/9qwWuJKd7xr8BH/GMeK0ZuPaW8rnQYkGrdGsNvnjn+0UTeeEmSqfTZzm95edI10mmyy
OXsjl3ey19EpOwi8DEBIgQOvlqrPwOQjwq5jCReW1NtPFXq4MkOt2L3DONNYIXMFNoOxf+BAlrrh
tOvD9J979QTpG1L1YY9Yx770st2SXh1c3/2AiVF9W0r13ra/CjTlZq68OuEq2ZiCGN2zEZupvfw9
GIZHtYQAFDMFSz1BwC+e4xz5pzNS+GzDlrCYyO9H7KuNvfHWiyS+Rjb413/yldKgj0Qwohymyx+m
V/+cxAXnUCNYRIqGwbaRt+h0EOZAI+TLotjQbDcG+2isCSMC8/ftRggQTug0rngodjLq3QiKSd3O
Ah5MbdTBQkWRRyoZNyg+pHLvHsFUOl4p/xGPOd3jx7VD9Sx+gphso16G3fiYhJSgDHI6Su7oLx/r
UDTGJ0HANxluL9/AUSLBU5nmZbvkVBcyKzv+sblcKba8sN/CGgpd7RB8oWptTS3QOCwrxEIS0Sgt
YSw9RmxpdGVI7Pcz9mxMEztNCKxRZtKxBCMaJaylUGVxnT0vLYLzBCC4IBvgaROiaEjM/YAJQHIV
rgX2FUxSFQQIZHlesSx5S5WyAksKT4hIz/Fl2kdU9YGYC7d8DKFCPYi/YGwEWZFyvDLvl5Ao2jj+
G3srXcjO0ypHLOZHtCW4nEf3rq70Ao429gycXJhxPZdj/LUriTAeezJ5nA/nzPGFGC6byheoR+fw
m8YpGqF3LdQfx0zXov6FqIJ1dKj9vykYHMCKRa4iZimcu/I7Pn75e8QrCL7u/qtITVdwnTpKozsV
qSsgWJmdV45aLb2v+Rmn2ZB89RGZP2jzmW1OaU6hjS6SeBo5DcG1c8f/BU/iwa1mzzrcXTFf+b9D
jGrjNtu4oc2XzE10XwrGAl8F+PO6oVcDlhfzydVFy9y6T4YwLlcjZw9blCKcfYnxCu8oHK5bZMM9
VaUFz5QGh/4grpIkro47J6p5I3DPW+wMynl8MZMG0IAASOLHg+QCBMqvfvbrcpe5eOaTAr7zGAG6
WGaJTGjgzRoo5viTdLXwoP85DajbhPLbM7tZuZGhHIyoMTl2ylxab1D9CCDXBoE/jeOlTQ37ocxV
GUrQAM6jnF6GRBu7ssaBCXdEwgtDs1NBdrvquYxKJnLy6uNZY+RyQuo7ggnpUMXSfFts2FfDT+dt
NxTAfZ1WXTmQA8dZHDlDm7thAdF+y23ZhNzHaZI8bJe6iQvss+ScwlqF9WRaEeEqqgQQ2HSJZk8G
Nj3yROU9F5eMG6ZZ+N7ybMDi3m2Vc3HVJFfgYCMy85TvEgSUan03AmLf0gFMLWgVHPewkk/S9JjE
E0dMQKAQ378RtFNHwP43THmONJ71fF23ANBAc31G2IAgarFXBDlMmSgI8RvJftWEee+IETIj27Vq
W7V92a1NMiFR+jbwF8XqOE8CKafIl3GmEt7EDcv5U3XbqvyD8KYNoZdUUyOyLrfNQRkM2re2kWlV
KXe3whW+T80svuHdSeKNKlI+Whub08BLi85I5fbBUqD8kjonuHX0gqp2PoeS4RRsG6YWAomC/0yd
/uiMblovQE9WQHVN3c0vEDCgyUAJNRz32XMuGHKNeGkjyOxAJsDxcwMn7DvKjR9+VpNNYAScdfGo
R9HkhQgDUgtzfexR/taj43hXHAMfvYjtkmxv6OY6G43LQcIsFtcRgeWYCVyTNcnf67LB48xfWUt7
+dk39V/FsN5bEm1MYsTptitptzAEus5Kd1bhjw5yhVDxDCeH834wAwzIIeOutWDb1T7odR8WRfn2
/IYP0ZEf01nvE2LDLo9L+89/xj7dpb2E2x+awhcSN6MGbmv0IMcnO/2XlZsVLH+3L7FDD9u09m4s
7CMYivEIJoEiXJS9hwyAr4IA5C9Szs+IsVc0l4wN0ylx3ju4Nf+VX1Mqq+SZYMAxXpysydxPH17y
QzQlL0xFTaAyyyEdME0bHcaV7lV2u5PE3g4knnvlMxru/4UhSE6TsHnxG6EHr4xl7opteh57x2Ug
lEqKaGHzXhSS94V+P+8pqKf3daj/Eou5AxyK58CuXppk4TzmvevdqkObPfL7YLPj6+otk8/TejJ/
okb28fi5sPApLOS28GKk3ujRL1h11cMjn27kKVSNervFUmmT5vpPvB82BWf78Lc6wsoNdl2Yh77C
tRsJ/zNQD7/e8xXHQ3iiurY+62eFAYegtEPLfjgAesIClMwOdn1oiEaatNCwn4nn8J2UG0s2UtH3
RnwBFkFM8y4VvYhc5khY3cqrw9BgZIrdXkqTOye68HogxZRe0R4cHzabmp5AUcxyeuEvbJ3MKxWf
kCW8/5tV5oWZflIzOFOzzwOP2Sg9Rgfvu2D9zdtb+YqpMOF9Te1dQHhIO6g9WST/YkRv7KWUkbak
fIxrhqRjggnVrzjUnyU1oxb74tw7LLqZ0S+4AUjWjOdb8LzxrdB96aalcoVvaXPaZEOe2SVQa2Td
ukuKa/DYnWbCbPRvY/I9uaChVr2BfIf3LUAkpPp8vVzWjC7jofW7hG3xcqBnJk+ESj/fD4eZCHit
tK8RZJWcJ7RerStfSI8JLtwIDLqIgRr0jiENatpStb1MzGtHONr9uDj0WtvS2it+eKmRSowhLFHq
cN81/uVIf1O0Cajzv6zAKhmEFpoJbqfns1HGGTF7T2fhfv5GXrdLZf03f0XQbh4ILrV8HkIUaKNS
ZF2otc47uqftzlbl1F2kvR2uxk7wat9AIcWCuFdEbZmXiqH8X5qJLK30c5/nJXWhXr+RxiSftHE/
NHHoqX4Fv96vm7Ro60Np6YylMXVfHWToJXSUhy/DS9BqMKMgi7FCECp2sHJFn5TV4xIb+CWY37H9
MedZHyGcF8bBXxdlFzKMvrYtrd+dmHiQMoMTkaKCE6uAuVvIcR8+79kNRknVDpOHfa+o4hO6rBIY
iCmgp15hzsHlxPqODJL9Hl9HY78Twh/NIpdKAuyoX0W7Ebcjg/h4PPwAOLaLdN0Av2Mo1tJRZOJc
/xty5Bpj22/bjxz0ofuHa/o0wmvXrYrM9knoa9AbxC1lFqSmKpUDKJb7OqD3L1R0FZDD+D/E4pUY
JbrsRI9Qt7T4B1cns/+NZ37uMhutq36CsrxRxGzciMuuDA8SkTjFj7bBe2G8UGhLq6+CCF6al41X
QG4oy6jDXDSYJFlUYBB6zC5EjTQQKNV3Rb9FuPfxQBidI2Z6RNgGmiiIORtmKTg0YfRyHbNqiLoP
GsoPFvCKX+gaULOAbdZcEUVWhghDhfYs2q+LIStb2yxJKPuSbwXMiS9vROsdHUiQ+QXjSc+v42gN
iB/f4ypLhGRMt0rurtPT12HhxmIdluE1WnuljsNecq+Z84Up9anKvHyrvKe1fX/ms+CmrTaWBGWF
ddObPzAX+dDRVHxlsUONJUydAqiJWT2VR2aH0qveqaYO6DDVhXsLjFJPeTOdtLGfXyTkdoeroxd/
+4HnhhpGJFjOop88uEck3fjl4s5zSJEu4/wzgBuxJUc12efwlEsn0i4XZYqfV7x0JoMBsU0DRvRN
AQvxzvB/m37Irre/aWvabqzuuMw+8BKlFa7OqTSA2OLBPYif/kwrxCV1C9diiHpHJZ7v90+A2ptQ
CWIKZpEwz9qATKaa8l3Yay3pQ6DOoPi4yD3jpW6ulrWYRCaKUTj3Eli57mN8Nwk6WDM4HoWuzTfz
iUPLdEI0DVnaX5DTZhcIYqH8Evi4LAx88Wihvgn28cci3JopxrzcP+YbvsGh8mm0tfYZBmQwQUv8
1YBw+6DoaaZ26AW7HxnXGlXxZKPHGRR3yjBCkxBOsQMTsUXeR21EDSBLGHH9p25IL7x5aN+vrDM4
DkoJK5iNVEyA2P9XuQ3bRAJTebc9E4D4Bc4si3uSbmg7Cllp7EytcfdaB8APyPBc8uMD5tsUZVFg
pn2gFaM9rNelHzt6jz/ueadOKJw8+4kU1gGKj8n+fCM0P4QEd9gOeged3YHL+Mx4N9Pac58obD8s
G5bQEU714UENZpAxD70AuTzv9d+t/2ZWURhvKGmsUVdq5eikhdR4b2WXpxPGc9jf0FgQiKYT0EnC
kQHVRFSZzVm+VBNnbqymwnktDpnTd3BkPoPXg2RjgSBhTX979VwSVzjALZIz1CDJwfARtoG4moLG
wpprg9GYILiwJPRhop4gxsxdD8ycU6Ap76nmwoWbKx/ySLbpVhh3FhGvvGXsR2PqJUUCu4Lcqb8F
RCBhfinNDPjBRIIZU3FOR1pD0ZIZDWdBysG45NJtPbNPmfoyv+DwTXfhN24UbljZSDTIVSH+Q3jz
HLlOwal0v/6SSLe2dqxagbjI9KiuHllzHcLfwdLx2g82XXgZUF+3PtvxvoctXVY1FHV9qUXsvLBc
/BcmA8K9sABT5AvRNug6/C0MZugDmyL2Gd0QrAAwjiJQdi79CnVmmsym7cSnN5QSGK3rfORN2stV
s8gjSfYtyvA8macQp7FnsXCmXlUGEfRs2UL4yXl61aNYM2rIcdzEeahT/cKXcxIE5vgsEZJtGa0A
Z0asC2A0Pg+LPmU/atuy11tW8rM5RJDH3Q4j7s9bLoUUKVgYmDhg+yR2v4ffaMbB8gqohVYzIJ2v
GOxarMEeLqtDk0q98re7F3HMV4A4MjJhAC+dvl9LB28BG2F0WnIB3ybRM0h+StR15R6BPR7TWgHA
sGAU41GmAHbIZ12oKVngC2aBbwuqNYm1s3gnaO4KfrsdNF7yMHOeCx9Y+KJAR/TlhuS0be+Lt4oZ
gwOaFVP2nbA0OWuafGeftM7e/JMW5RaUhKKFgeESN6Q1yZwsdsYjVydMcxj0FqOJyPaBwTCdEarv
XEHtTVwWIpNH1kQnpvq8jBARbV9fDmmUYOhKyWxPhlnEtTOyY8Ki0S+SKilK+e0jJtPWBERHYnf4
5A/NeCi1d9XZ+54q+MFbxqXlRmXnx1h5gKhs7A37tbr9BYaa/guTP6K/q2/CM+N2m2VQ83n0Eil+
U+94e6SCTGCPEiXNK4Qi8QpB5s3pf3gEHjSAiagsvJ66PEDvFEmBXCXMwpdL1vJJkWpifbAjxwh6
PT+AlEDLnmRd0Mjivpeb40PqDIc9YFzkUPznzdQ+i9B6uUGyCc5xR9U/PT7Rt/I/n85mZzYxqlv6
drEquR4W75hUnaaxhDKnkhz58Zb65m46uFALXp/R1tN53eLS39c1BPVnRnrXe+QP44+ix6N2t/LC
+THeI/Om84a2/x1ULCK+2dt5u1xJUCNpvfLRqAPYLE5R2RA4xg+ROwzGT2gWj7VKmBs4lU+rqr4h
5vmoHotr9P4YZHGfvZGIfbR2g9WhP7FmYX2Ti9OqlTW/EyORJ5I/gfDCP5N0zdFK20QIN2B7kQBy
ZgHWlc17ft3UnQNUVLzmZt2Dx2z7sfzTCRz3JNH3UPHU8KUn77WwNUp/S4dUChm/aifwBufhuGYI
RZ0rEQwTZfhP/v/LBHoRTBz6vUpxBLEp0JiAWrVYQIhQowWlzaJXsg8rnZsOfx1Xhp+0pBNetP8V
XASB67sVn7nz0JJaisg2KUg3JFOhfA2b3NfZ5+8Qb5QcbL0LGJSGnDiTV9gpd3VBMBGWD6cp4vkM
B3+9MnGcA7JRnX50tBj8cmG+ViLJ5JAjVfj1QG6B0XccLM4XrRMI6r1MQEKdxeCFuym4F/8jnez8
ZPiNjMB6wt5W1kWXt8x01bb7lCD8gUnqWV3khDpj9nfcv7KpPm3jMQpNkAN+QBO+1cAYx/z0WvQr
9tVbFVU9pek+r0sw4sG1+5mGgNEtqjUQ3xqodcls0n8JKJ4HG+AJab/aJQ06jd3QGAEPhUSAWPom
TDCQ7tLkki3T81BzAXEHUwECNzaJlbt4bFiaJgojd696ostwPK6yQ+P3ICPW4ODdeSNW3+LKZB//
5Ff5hxnVTB+RxAFuxDg3c3FP4qqrOSs1susujjKW8ZA5jR3EPHwK2QZJ71l2x/94kJFgmOuQDsO+
V+H6NnaafrL0F0BkHNZoZRGpcyCaY76E7Qx1hkYSmVS5Rf9EWR3GIOvBufQ1OvoMIreUJhdVtZRx
demlaksiWHfE/Gib+iCCWpCREbwFfz9F2qCur+0SK1I+gnNFKxC6oFznJN/QD8AS9gAF8bF1Ojor
Efhybt2AgBtRC54DR+clXKTsYiaGz8l8enkaUkyq/W2TtNhKqOiGARaNoa6M5fQ6SNqfcLlDA3Jx
nSoG1m8N01BaOGNYGuTQvv+huIBlu6HWOu7kGE0kaK+hq07AoKDiA8F3cY+kDrpa8J9mS4v+MSXO
YBaJ/qiADeG36frVzu4NnGy2qN2y5yFND3nRKB+tN8Y2e7SKacj9s910gqt6Lg4Le0MqGjlCIcsw
dZA1vYY1R7uK/ZaKqGspfEoGaP6DZfUTODOTY7rQ2BH8jsARgm5vXxQnU8F416LDE3o7YLasyfJt
zTVweWIY9Htm2Gf6ZAvIQRsInWBOTa/l7BrbWKxWSJHxwlueAlmvuyIQJPvrNaEFzpCSGd7JqoDQ
wl+EWMgWKenssA9JRExr2vGLOLA4mNN2a3z80/VOp9jfWdTKgTUSctyQyr/IQLXdZqsK4jyddvs7
+saum0h+3GrN3uVFJSmMm91qW2f5e/bTtbdjeA8iZpnjKcHn/31vjWDoi5/7ROP5Ag2ZWiKd3ZcH
+KsTT4FTktRjK3arcwvrwntjEYeW6IogVxhE9EXBQFKlsCNp8MODHOCRp1+fc45GDMOEoG2i9gwi
lEpbL9dBjsd928TuL3OT7IsZLyT9CrigEYRR/0I1dP5D06uY3PRD5aXbveIM0Kk8ADHY8FVat2fV
bCZvRqZ5aXylHtVB23pezIrwKl3tznH58BYmLl5OU57FlyskxZ4nTmoanjodaX/DvK9PX2/zf1pd
B3HaHKCFlaJqw1hyC0mxackF/T4CzYjhKlvjNp46cnV/G3+GxoAMSDHvaT6B0EQOO0VKqwVYzn9Q
iR+M7b2G/TsHtqsyfPrr4kIudFZ+tK/seBR3N2WSkyCkTKRC1+siCVNPVhK5YWsChfrAhZxoSnve
9l5ow6KlcevTJh/4eZs34SyIswIdn6AjLtA4HqjX3xiqjO9Qo7oVeRmgNaLZpLLlajSL1D9uOWsM
s7NFxy81sIC6/UWVUGaZJbEg0dg6a7ryKIdQyztD/J06/i+MLWwz8tcyhcruUUI10qOz8G5KEhZ2
efBv6nVIvY2ybMg7SugkmWvsKVK9DHMttBUB04akyrNT7eSXnFimbo56yiiehf1Y54dfzvPbDdO9
C7xnI3iQbwSSHgVxdXqfTbHU9VU8XnhfqBW1BekUgC6WalwpwT2cvuSkEKdTLk1fboB49DgENTvm
y8uwQNbN0yTPlIGFkrWx/PFcFQDal2GmXXWPdhhP6Bd9MPmKJyXD2wHekcTCH/ACN1sd5eBSvpUT
XL52D/M23HMwOGAHTDd5LP87edp/YMz86/1OeYRuGnEurjzSUBGpZr9ZIR77el6isSxyHwEMVcCC
k9FQu88er/K1rnwBoH3ejGiq/8sHb16zsI1IjAW7wLip4JbkZa9RdPk3p8csq4d32cS85WIx7jBP
VMyDZ+W09n3KjzjfHqpCnM6ZJn62wFmVLJak0vv3UbQMoUD7KBQs+kx7BP+s4w6RAx8r0bVzGDFw
6FMeLMu5keqrC0sKrB/9C3t/14GfG1hRngWiL52v5smeSIe07xJ5x6kjNgHl9nceYFiZ9GGS2D7P
SfkntUjcPq4P/zKFCmA21pJxgf/h0KUtInf5/9C9AweuX3OtcJKElm9wn07ZjzF+9JZjb5fJIPvC
EJAjOROesoaxl6ZQlCjH74/eX0FrjcZdMJ1/2JBRlAZfq3v1lnZCjGyn0wCrOQgTU4+gGeBGpD6N
OrTKLNtqE0oSCd7dPY4T4xNaPHVF+sIHWoTQTGCSkHOWslt9GYotptDgtB9jS5c+SlfZ+GZ6xwxH
h7zpHGv+TOls6sINqhwZygWsuHm6/dfZ/Zkj8K6evzBOJ6xdEKGW93G7iM0TEPyXUA2hnHSGmup3
YiDjnADMhkF0A6Cx7LhToDzlvQ39dX+2l7vpVkNzzBVKMIzscpzrtQOH4qzRllCxfj19euzrdBMk
54qkNhiJ36Ox8br4VAI/jpsqhgT8w96I85IC7PVs8OTaGiZSyZ4H2F26WKx7zkUwZsQ3lnIULHNw
VGuwnSYxG+EIgtUcpXmWpTsNrF1YyfG1VWWmg9fNgTsbAwTY8BpxJM7bRORsAz6eb1Z9k8j57z2b
UiZrWI68T0q+33RFFfEY1oxiBU4G4b84DUkANeVGJJsYCN+Y/+HkV6PV88IqtU/UyNiS5zq2Eii7
wHmIlqpYTPRckcxsPBVKQHSOJWhXfynXpiz3UnD7ark7SWNqF7SZ/zcNorZ3UzMnck8ogFmSkqAs
uVx8j6WvqdiU2y9YVZP1egAfbuNbWC5dkhhT2BQBm1A1oKthroCbKSBxigSyy5XQDQcoXro0dSs2
lPks5OJVnrJVKp13E8i7XLfgn1lrBeSOZ00BCGx1JLVFo8iNLxnYnzqt5r92idpzP/OnNEsc+3Ai
2aQn6XIf9UP2Crcp15PcvrjckBJC2QuOWowXb25bmXlTI3OdqSIMqSgY8z3B68pYjwaek9oAlBUh
x1AooCHIR5/2nD4Jc0n3o5ylq38yaCnBnD8Dg+zWucLdHt/IhLZYsaV8usPeUDOMa5mPaFsOX8PM
X/jfByFyUhD2cW8s7M9xIsnSBG+URjIC9W7BHuxCSPpoMYdcZLeKu3hsetLx9EPNOxCwwHoHNb7N
kOjO7glPqlYLP7soTSO66uFNzSUcRB0YnRHapYZsDiQWe+leDyw9aUk9zo9PZ6DeJ5AoNsXXTPTd
qLMxetLk2GWaKPHiF1n5OlanTsq+RzTpwqdRx7D7pqIS65hxCwQdCNFUXFHLy86Mf8HtHIxb77VR
On1igv6yZlEZ3nIc1zKnpSi+f8NyDgN/qAu4V1Uokx9GNPoe57W9NyThkCac65EvnOAdhVvmUsVV
F0Ow18hpgl5Ewhzi+MyeUgJQKsZneZaxOBR+aF87Ez8eiDpM7rgfSphtOz2myQ566zODgwQ60TPA
Sk7URWKb1xHdEdtTGOo69F8L+QcgTF8dBRxE30u8xb9JQOytvxh26JPabqVTtCtjhHYbhtYoxHV3
A8C4O46rHwik0nz2Tl/dUj32WKRknSKiYLAwqWLgGsPZ//bFEcumbc6h+B80DBNmbNETHYu/DzRE
S0GCMANQXm7v8GRIac7eyl5jtiT5sqpOj69zFcCrybzXcnGKokmNknw92gMplQnyu7mKW3fuimR/
BSodIdy+MoVz/SKiA21/Iw22Fpp/QrzyxGRIUugFbJad3qDqwo1feHF70sS7CyXYxEgQf1BjlBMa
jLte4awikyURd2naFDcReFEK3x9kG3RQ7Z7cS/uCYRUeXk3mIh30nqOIWL4HbJSNfIloam9Tlqg/
0lOq32Bj1ErEN9ntyB8Uc+J54k4ZKMZc2HqzCjd6EINU4eQRZ4BI+hmIWozbPHQdg10tGa0O5kQm
XGWzLfyknSOiNbW/YRBqDx+fN1xN+RsyiYCxIwdarurDVMOz90ZeK6/2lj0HIuxVTdVpfk+5A79V
QgzHPxzSwajNeVCRntBv2JrcKkJBIaSqal9Rp5A+I9z0GIdfmRA/K48TfY98cjVUbbwfjdrbxkr0
B5GMQN3rL6Z6Nacb/9LZRGK2koNyQN29d4H7aocqbjhqTratjUBITC2G3/sYdOetPeMgY4dZDgND
R58ucCSHpWC/HDyapgdmIO9le30YsJkAnadfKHuGDksKqtZWFdHrRpzGY9J7yFe72EtaUSG3EsHN
ZRXMnTnSBJixefy6l5Gtoq2g/K4t8fuK10aCZjaJ8SPrfL9iZe79owrYdob1OP/zpbRo5blk0fu5
r4KdCGQsXhV0GsTVbuucjc9simLwqgPEPOggPZIcq36z4hwke4Tblh+TQFGp57bJ2HgY1zxo6Ht9
Ac9dapY4M37KgVavUYSYYFXYVRA4Um2SL5LAcMNvwF8eXlTOf2jLumvCYwgwxu7RUzLPuEx8Cdjy
SPlsv09eUYZ8uAiiRjMTbYl16W95wgx6CIrNqk1dQK3FPNnmyXNEIRNktdfIfbtummyC5SCXmHof
BIVqVdxVsKifRddGpczNNvlJfT94h+boW4jyb/AH5V3gXIJGA6XLWVdGrGQ9wzstfRlSSsKUKqBY
PynUcvNJWaDZdjklLRtMkeIAHBndDB01WrWjuNvj+/XuTzcc+Bxx+Wofa1SdHmT0jWg043lo0tNu
kL3kKbq0V/sk4ZsXIttxqfDVhcO5BOCKBJCbqcJv+nD8iznDkwCk8XGOPrDiZ+tSDo9HTs6KyPaI
IV5Sd/G8X/tUwEbIv2Y09GgOiPW1YwURQf6fGBhbtV3/e29LBH1twvPmcqkyAwZBFqEy/8v6hkLs
6tvpXz6n+rejfGUWs91fz4wHKKZdBnBxrHnoBdE2s04W4pDMn9BHsZ0GzJLilQUgHqChj5drDM2M
WzmvFyThVgSA81LZGTtVDgu9oaCJsEl8jSklfHsiXMDRlJPP70m266Kz/h+uhTvTTU1gEcO3EmNO
wKF7r8c62MA19yp9hBq/z9gOg2FYNTIpWnILsuM9rYni1YaUJseH0PAqf5pvc7/U01FrHMeCeOOC
aXtvpLY1A+VI+RwlnYC+iTU9xDtye0h6l9zIjKoUDVukaG98k+9du7a3wPr6YCLwUMnILdnTvabx
8HM+BSnfCAJr/SqMKXLA0vgDg8Z/etBF6ryyFIRUltqxBV/RwFDULwmmbU4O1U8Hz4DPsbwqXTMt
iqwYohjBY4YsfToBVHgXtCmvexeiewdPCbDQ2cnkZLxWwcQCn2CaZ3DzDB3hnl9YRZvXAdP9l4hT
HrQX5JFOHPHEq5U3OU901yuitJ0GxNYtpYhXy4wLb6IPmqyPg2EDuCE5gsLhIT2LMa3C5LdNmKqN
psboIpn+9wT7k09C4vsmEOG2BqW42XdTLZ9T28kKRj/LC11/AE8lW5spfNM+1KW2EA4S6djJYQTo
I2QuY4oib9ld+G6h8rnhBk/6ASq3iiBKoLUsxSlYS5xEKebLK8RCZZ6TXDI8Cm8Abdl8a+38Ui7m
w4gA6FHPuIFiA6Jqrsnv8A8awjUFlDsg1fix80FEpXXg6hXdV8ouJ7dn7qNssy1DVXq/IwI94aZU
RSA/Fznv5PDCVTOQO9FlZWcRW3xjP3JG41MdrASXui8RiQKojFpbk2irqswPP2G0yItq8+xLXUTi
7dsu8n4kfjz6fmgokYkKLzS2rnNJyQT5tIeq8coXJoJQr4vs5anKu6R74x+H3ramImG05O5W85JM
SIB/iGcM9NZESJzZIF+yxdiM2aqRVDuyZ3JCci1dv7PJAtHATw849RggynV+sXbv3i/Ri1KXUsOw
dVL0dmt1v8B/JUT5ju5XTDxgE5ddU6+2Ff7XHyDaaomALkbNY1p6GR/crNryIOmRI0VNdhRDpn+e
iJarQRcEWpJTZlfOoMDHgLQacqPaoqIHB0QUthY7lbZBMHhhWTaTemR87K9dKQitohT9sT2xCTzA
2cP7bkywaR6qmtIbIFQtVOIXx5kzEuO3xg9lRJckeEl5f1RurmvLeGS3sZofJIvaHvMM740BVzoU
QHQz1rlIQvxt+kOytJtGXJxCa2HDUFP1GQMwm9cqbmI2DLWUAdVdXY8OjC6+B9N68FQZPPorMpDa
e51nC0Yf9EOXSoO4rwW7KdIQTeoxehAOIx50saFlFW7CD80v5WiSFPfGLE297thMof3y1XTCvxIC
oCo01gVwGkgr7klrHyDBhdU84cLZh5+lDgKwPm/GrgTCwA0w1RZteSyq4YjlYDUT3/vmcRAa88eh
Oi2DnAMFQzSMn6zpDSuhgRt4KoBVWPSX7y9evYXUO6zA12wtFxD8XjQ/8X7g8ooiHJhdEUBTp0aq
UfcLEzBQLi96Z3eI/hQhwYbW7faovgqWrURk69mHy504RoOoTZ2xF9Dhs4+L204nd8/r4vSKLxxp
WYp9WcbfZN9IuD2ScZFvt5Zvhu73xKFWrAuIhjYvi7to4Aagc6tG1cGMiJLPrFX8WtujxsO48Kc2
++BBLnkj7wYCr5Q9H7FXZQnGOlUpbHfxk8Wq/gLaJ0qNvpULtew4QNQ2wfimKIUlvyX0qrzVqXAp
SzauQ/34lf8SDhva2ohl0TxEYcJIMGd6HeHc2fiKxx1CYuZze46F4Ou9UYOCcow6tnpJo9oyjkrR
1YHOsODJLBpv5NCwowi8TksejECo6dOVo25bEQ+UiwP2xzp24LpHV0KDXcNk2LL3B8y9p6NHT234
e3hQeUBdng9ZoGuC6tHR3tw6Q26xfcos26AqTSLIy5t3WHbv6SBwNxTHc3oNCdjdmfrGi/UZ6YXY
JLT3YkX+Ms1brtFqyZFQSj+QzTCG2MzT6QDXQU16AwaFlYHvMPkLhsef56ywCNIXbONHPfjlbTtI
5gRkHsqWVdWL07P6/8oidiG/3ZTnIG+SIi8gSg0OkTzMksVgaY2KnODgnA4QjO5LGiyu9AEuiSHE
l3RW3bokOA2rMRjZxgZer8OSfAywzV0O/2rgj32ZvNeVh8/a0n9IbbvMdSMv3G6wCP6AkiGasAWR
TorzI9IMIooaXjHh5NwuqHJMIc8sDaf0h7NB6fenav+7V2NazJDxFOCd25gNkFUQQFAL526YPedl
fota3f+4P6IPJvvCE78pYgpEhgKAf8hmh0RS0anCVR2XUvRKR7Ybj8KLNipT2JDvVbVv9MySfiun
WBHt6eP2U+8SvNnoNnAz1z6EBZjCcuAGbeOtq0bkMSF08BAmOna9BerZSrSJ0jCJcUxMO/mDhEqU
qXjZ5fwmQGQ/AwV8wLLYcPuaSPpPldg3UVdSbtcX1HiX3coks4PqJXSa6KsLGFaS8Gvt0MRRXOqh
cmwLxCef4tIb8HxQrghrFvQznl5q/4oiO9tXTnan4FWyJKi/jf41LeqU67n07f88ucPc5ghZRToH
TtcRYJfm7l/w92pjN0IYdGf6h9FJknPuGcyXqEV/tKFaKL2vhyzmHoKut3ym1JXrQ53ekurYKolh
loGtivgT4kzgN6JI2kAlKV+rEay8f75OODDfTfUCiLaKgyFFGoQfwLmmKddlbPm5/3s67Hrg1Snf
dlhDNZcDzNlSxaTw+/ss04Wd/eFjUmNERQA+W3yacVUvvrJ6yQ7JTMNjxjF7oHUwTlGpURiaBiVD
8GY2Uu/W2mWr4Hl0xFGWNxrwlQjcVp8yOp3vP9eMp93cxEsRJWXk8GH9ZJIFimrAIbj00WF+Sy02
qPGSKEebO8i2yKaZKYbxNjC+eZkUuzV+zyGmNwtSwJWgmv30q5XBe5cYhcIkyh1p+8Ql0BUVoXeJ
LhDC5ndR0IeEQ5qxfhYYYsgLoTNTxhB4pUx5UL9GRzSnZjmfPrWAZbc3cRL5WTzpWpNDaTI4dtN3
GWjai6QUEET/yukWAVAdaFgm4EHVZW4zG0V/btpzXWq67PH2Z7QeAUeeRdiRF97NF9Mzb9MdRJVg
ts/Rq/tZcX11kTNz0JtnJ+YeNPiXCNRzC81Rz4c+NLLadgNlF30jNwZxER62uIwjdNS83cJl63pB
XCjDgo/jOIcDvWou1//eVXW+/teGmFRqIUXMYAJ64oK2XDEx91b4VauXNDQbQvBj0AuNXpnemWP7
JxkoWpqXgmEMhDkb9od/nSYjoEfyKdF08FIRx+34LUP68OBa1EGaK+bfcu2aLyTX/VqO7QLLFDfE
o7XufVFMM6XP4T084UpdnqHYHr7tlWAMfLj2+Y77mTFGyCUiN4Egk+CUIJk+SXFqzxv/VZj7zns+
QA50yifV1sBeh1UHLVoIvQwdl7jJ8hk+iI5+NXpjeVuaEMc6iO8y5N52kXgh/jQPNl6Lg+eRDOBC
qFPZnmqF9ggrbc/rbEN1rcSwJA704C5TMlB1VDu+ItRFffGPtEiSxfOqkLpaIZXUkY/B4nIqCAlB
eGydUslr7JGCkNc4+cpMOMgVK/H3nhWrT5ScLMBtF3N8sboUylmbWRlBLmLdXDibSPpSgkWKEolb
yE6aPZlj1WfudK4p1OURMDyK5jDlXQ/oPM0IIB18K+VN3b9FsIcDU/Z8fw5QSId5/8Hp1AoApJrX
MRiBLDigY1eks4WzYevy0WbugJcx8j4cesUP6bkE0VjCoxEEd17iZYqKh47zW1AugefY1bAs3Gh+
8AU4jPPVJMzI+301CIo10HoapDOvyF96FmmT0qH/Cp32kOq44X75ywaXzclf87PUHfBtVo0UhZnn
pC0SWM5MtQcNyc7DjF3tP50L/EyUKyrdSCVy8RHsO3qf68lX0tE70nnTHT3weHPEVHA7cQ0Gl55s
DEJkDbwbCDJ/r5KziTfLam6//SzpAcXBabHRZvSca8V6mAUIvSb8DIhR1rPMAjG1B0AxlX04mpZe
gfYWBDQsliOajB2tPp9jSUuTASMtuY631RLMMMSr1818SSRuq+fGEH/P1My89m4C9KXmgj2qqKVw
aN7ZnXN8fVvtKgjuExknRZ2/nscTPRwIqyrw+l2Z6F2eegYC/qOzbNhS9iapzJDyrVeTBJFEDW9M
i14Fu5wG0T2s4h0zfUdddBbV5wavnkz4jflPe4bTvWGh/r6J+FrISkM+O+nomTHAsIZqlBw3O+sB
BEleFwsmuaZ+o4DD2A4SFkP7bb/hl4Z5MZXya8Ga8qgf4lVz5JzYz4NhhwHE4yVd1LTB6wzU6H3c
ms7XgtKMwl0aL92os6zbeRrcq96BFLkl+UBsWeJaabNUoQz9Xqo+Pj4bDFoTSOMaWTuczGGaXUiq
Hg0OKiIvQ7m3REjlgZIb8/Bzvxgma41LZojBn4W3a+uFloR7tlp0X/bdp3LrrnO95DPwLvr0MrqC
LPIuZC19a+aFlhKs+tA+bX/2Y80a29yczFTJzyHfjIlecsepsrVQb5mnQ7MFZJV4OLReBFGVAad+
V4AYaHE2pEsBFSnfECegsdL/OcvYiBp6hO9UitMFzwufVxtwhMXF2yhUzb8onj9CAko4z0a9vO+H
BQaZsbA0RGZ322xtJtz7oqR3vHdEIXIYsuBPUXYcEdHT+yXo7AH9igZLbYxlld72G6ALQxDQwXr0
6dCEnTu6wfxavy3WXqmx7pCU9urgIe3LEiidhRIMuXApqQgUF4TVpDrXYNfHyYyg0lbyPoFD+1mF
TmIvt/ay63NDzwsxVY/3QeXuQmFCwnHT9SkqX3Q+Hb/MvipM9mrzXzYzINaDuldtbwudyczrV8kc
G/TS/nqFsy7fcDKVu+u2asQ2Qab2qeEXaKtVHHIPOuRF1LERYRG38+BgfhnBoj65V/O4LuuOwaaI
tXfi/lRRRI55lyQmjhZiwowzbQVgOAsKPPQ1N3nIDSu5yZSmMKfu7WtmVwJuvLlVYwmfxo86q3S/
ihqpARrZCW/ENn1xlMm9BoRxs6KNqrjtkPDNGwmn0DIGiS6ejOxqNJNGw+x1H60gd1RDSgOPAeXm
mI30TfnrnCzam8M1ESvK8lFhnMviMAQ+q3pPcFsi3QOGt/9M3+BcAkwCqpGHEUljDdOQpdysoiEw
kBz6TB7uHak+OTPO+gbiqbY5gj/tfQuTv7GZF3Fc5B4/oqhFYoaHP6mWjfkT5zqunwRrrx7dCbAj
cxnq5IxI054UlW7aOfAB93SXcSbHvBIhfWQ29JUdox5X62/8Vxbem+pdM32wXc4DBeN9wxOc6D9j
JS20PEKNScCz825rX+uZLl3cVRWweLHTGDI5JG3UoZlm1UIW8Ftbb4PckoyTvGBl84+YNPXTeCQo
lLLFCGkG3Q35tauOBtVHu1zF035GKLvwxaesJxD83koQPTYUKBytxJKH+LIfe2aiVaKnZF2J45kT
QYWMLhOG3OpAvTTGkaDv9Ka1omdeem+aiAgVU9gu0ddVovPpQXWwUCqD5TotpYjs4qN7aN0Fp+Gw
yuB3Ca8d/xiX2RQd5ezyq4rlKnD6c0coct4nvwpMFbH8gSKYTrP7Hk/TFp5LUuEjOeLA8mDgsUXx
7rqm9ReuFJOOOVm2k2f1f76Wd9Hxl4z9qpe0rHgKzDaIJmtRs5W6frLxC2o4ExBjnc+3jiQTUUXk
stAepeg08ORJQZ/AwN8BUpbW+2uNijdPsyz/945D7gS5qMTSXRLM5UTuZZoYt6MZ23vC4ySR27dV
f78K22O907TjUCAQFUDMuYn//pCA0hU8wspYmfrM49oEHo1+xwjXKrYki279NPmJg3b3SldFAqMX
XAb6J7Wxp25TPWOSElNE5uWF0onE0VFuBJ4X5MT/aHross3r0ARmFtVgdX/AH15Tex9TuYR6xbGK
1JbuqPhd4okmf6+77rhn6KvDj1mtuUeN3BseyhHTAty0bRp/Q9sODqw47CiZ9aRQwtqbRYhvU+w/
ScJ4NXnIPqls0osF3wZ3/hgfGKpL26FeG796VkY860EhTS+0yE7hf9ZJjkRSuOnalvKN7jiVQLtW
tZUh+Qyi7sGyvD+A1/j6fTtrOaLoJ+txiwVkk5pZJzYsipSJVpdTPUiUw0XfjUTgp+Nr0AGNgo+U
90QkUiaNw03ImIL8IOorng4F4/RtnSJ+2oW9EjLSYexsyOXE7rD65g8yi0NSUztdX0FSyabdywMU
1W5ztNQ9YNNQXthn0ogrfXbmqJ5BEG5lNl1JzQaKJLykGhVRj1SGMmM7OKlK27sy8BQbH7zlFaKN
+/c26A18KpQoGkoQJTGII3e2VnFTUxShr8tlJeACO6MamKSZiirsa5ahro3pE3L+nIds9O4Ej1Nf
D7Bpxw9ialz5DFkC2yMXRJOXx+G8x/gya2oKKT+xDzNUvM4USzeyPSF11m5/bpUqd8E+sCzE9We4
tBqfzCMNULstTmNj/LW+74MP+nrjFGHTUkPISPl55c9atvZ9y1dedifPFJyr05wkCNiYt4GDcKZ/
mI9tf7LmoVfeToFRe5ckFoeckHyc/HhsnHdwls4Ookcg71/BOpPLTsQ7Xv5GJd3RlaTw8LLhuHh6
2fC9cxKQ/3jRugcIe2wkJQzNoCYvDz+dA8l+FgNile7nc8IZDGlsjI8ss5Cjbpji0AKPGZ0o1zcq
tNlMsDXFP0JqjLz3KRG+hh60gqtg72c3IC/IN4OKZlAAHwRHiNB1fNiPwBwmdiFg8NlTOzaNQL/g
7ukLwpnFaEkfzTQLMO0PWm7IkTAe/UtChlfphixCrQG71e1G+9I2HqH79bKadwSD8YWLzdDnHKhl
EM5MIGoC1lmbX86bSKum5nFr4S+BwdA3B6HnlIuxhTJdSe7gkTpck4eRgjxXIhM6kRI3zmTnQ36g
4zJBvkZkznWL8/lvikS0q6Z1MXq5+vxby0XF9lXubsUjFo9N9euKihPMno02kfFhhGqy8C99I2fB
9q7qZE/lZEyjzUokgwVTXPGHz/WwpT6/TnNpSpMzeRhST8qJS0wwNoP6OpNTifusECdxmeFLkGAj
NXJ6kvbtzeu9fZUKNjsvemYD17ufwk4xYiVpxPiVdPI//OLtrw79y5KgtPG7gHM3xZvEquG2Q0RM
RMv95/Q2u0uBU7XjsOE0bVc4oZLThxKhgLhxVnZQNl9wCjwIpdQAkvFbj2LmbXGNle8AXa9DpYOU
zldXle45p3sIdyjWP/8VRkwWb1lnYon8ge+EAmOXR+omfLNoSHv0yrkuC0i0toUcLbQ4FopyHJ4i
FAyh+QVyDJFDbhkxzsqe00I7JJMg6FOL0BIdnaSCgSDsqfTnwHHS5V8jGvn28VD8KFbNI4XzVF3U
BLJskFESCgYPG7+09IdLkE/KVL/CWdUX5gA74gIU3mWY8dpCZq1dCFkQhXlinczt902Ymn7mYd9H
QtOC+gps5oCLzOzhwjwTFuIiLmG95ZqrjIj9yPQvVsfcgw9j+0DvCH0xtLY3hPEIGU3ZD8ooL3j3
5TRHL395577TJ5nc3rQh29lSN/EHL+06z6vGekDLtwBDQ6SP3lMFZ7BKbfh9YoOwR1cj++5tI2iE
o4Pw6NnqQgdDlukIqldPalbJN5CmTZBD/zY1E/DimFyuG3EooeUQlD4/N/e7Jfdt5QIiGTjowOsA
9leAQJHOyrMhR8Evx5SX2NpNPy+FUFmwg6qxB7HnxNe0wRdD0YHODNGHCYtQpLd/XCTkby9WzGOG
X/ZqRvB39SwZLi/ORiz2ojFsV+PUzx9gAJqxLs2X7dpG97m04KJflyvVHs0Xm35cP1L7nH0YTDvf
rQobkUlbxriC9E+oO6le+MjNQYC4mPHlr7jtNMLbtjAhs5e5KEZ0rnuZk1CHjZjKW06wuLq7rLSQ
BGkqRx9w4xiuyawHAF6W2HZt1M4ZeCda48qtwH5BIhAdZEX1/g4UzRHjVQIP5d7Mr9iLbjHT/lUX
YIkeeFKyT4W0bGqEPNG3uSH8lpEbYZMY+CMxEU68zEMqq1SPYTejS8y89S+QWRSo5u79wyG881gA
B9qQ5oB0amFK1TgSL+fPJKSFhkyXU2FTSgN2uI1SuJ7JcKgaXSqE2qRDDfh+Xkv2n43lhPOBWeS6
0qfrZ6gxejTJveVM6sYz70AFQNQQlZop/r+BLIISAUWax59OQLrPKwWF8FqPOCDovEAsFjgE0osI
h3xcw082fUw0n6+E2NkkdEBrsqg+uCPgemn4vKF5XuOU0f0cDV9QVkPLlyIktzXqCYQ7kFxNTqAg
uOmWXfT7/Y1PUxvKsVEKX0EJX+03WEKYVxQoOB1yIyWRfJQFTWaEIDmABVOE/vprZ6oyciIGQVdy
V4lgxQT6j3F0KkPqAqcffRopdKnPIxOn769y2vFi2Aiff86sOEDZmgp4IF9bO/E249iGmpl44mu2
t4qjPEQyWStnoxQA2Jb3CXVdybCVm0Wz8aW1G1W60CVVMGzMC4SDaBLTabh8YZZZfnLx7DDVhOHk
KUZk+72c4rdaUc+8dGigACwfaGiP+PVQLXgLH0dwdREF5nS2nXoYVGTVR7EQ8qsmwUHB4eQNbdXs
h4ipBq5OO1Ll5Ep+Q307691i51PkXKlMS14ElFPTjaeyNnTvrJRrh9P8U4kT9X11QzDmfAKKXYlu
jlGq2fqB2kOlqpTI3s+XCy5dZxHGdKHL56C4kg1dbfix7lLMpatv+F3IMMo9kmPYskth70bV6bZe
Zjil/CoGVNDHrE06i58/F6j5E7Q6mihVSp+tTKLW9slsIznNm5bYDVbvhorzjz3N/rhXcKZ4zoYu
nruwfR7qmnuyCzIVosRN6XI6VELIPAQs9vIS8TpXZgm56mjk2pIrB9yZmP+CWj2s7Jk3PpW8sEaM
vZp1vk1mE+UCpgsygPTvIfvU+ExnK7OQ4I5IkcrZAFyo6Eat6BQLWjGHG9DdMIn747i1VT8yY5P0
EPNI98Z2w6oRqsP1a5Y8espI6muIMIeWWzwtckeUBVWXKJxJb/Ft4CBC1cWcvMIoNhV34kho5k45
IlikVzy60v8jVx5+j6MbtRDpcVFOGTDRlm6TDM4l3LuBPtrraKkEwkr3U/KEe7by9mM+nFknKcEb
bg6QZJWCZdotHdhyyFfwFUTRqY7CwC6z7g9IzJwRX6UZfo5Fk5/lRbI830RzTTdHUT24Yt1YdaIN
6NyeuNocCYgbG/59JoB+c6dbpHzOnH8/nrrZgzRmSP8UL4hc9apGkTh9PxKh60hytiuxmXklN332
K/8Ssyytij0PQtcQKDdt6sTHdC6NLi+nhNFEfoz+HQo4BqH6o9aA0ibqepzcGN5L0spt9OshM3D+
ffb9M5MzMpqWMbD1+h7bxPDAInzlZSpd5V0RV+Te3vjkgipFRGTzbqYcc19XG/l/fTvhaMwYUQuZ
84gGljNFsKQL021/ReTufYu2nSyHOS/4PEakUy8Ia03OSr/sSqhu3CWgNIFuvnI+9OKffZvfeTYi
x8v8jDlXCT/4kGgd59DqFV6h6gkbROnMO93HdZ0Uba17/vuDKaTCHb5d5LOAcxZ8eIxV/Q+5wT/S
7sercK2Aj8u/bq7+lVYGU9C8GbS+Yo3szFJBlwwMT8iuD8v+znPso+D9kUof3DCBuInEiXORYOjl
fOb8YBmodMCA4aUDXBcxc4ZdBYzqaFsUzWVkH5Y2vyoGyn+ROIzFvrN689gTOASaXXHsSRzcD6XW
e/I+WVeJ2nlNY5Xir7LXk7P5c8islRjpF0np1MnC9WFEMiUe+3DYRSwSqA/VRt1qv2KObRI3m0PS
H9ufd6/U8jydiZ6mAKbykQcmeAU/Y5CJtnMiAe6qElHJHMEKpnMn0VlgYw1VuQnySnrR+rFsjhWT
g6HkvI9O37nlJdM/Wmep8SlnHv4BTBFSXjE/fHJlybKxksXOxh/IkR9jUUCpFXy/qWSNlIe/FI2P
rK4I2SmceI5E8T5dzLXONj2+tfJTfsERPy89uSCaJuel5XWhzmdiq++mGzfsDEotuUE2ERemvosN
OfTFYYL2Bfn0zS0ieOjvxVphBkLpxP2W3rrFX7CEBy+SrsYdHW8/95xDDlcHiQ+PBJj4dnDCPwzp
C9U4cKl/vFm5KmNFGWUtJw1cH2JnStKRshQz+i68U8XtCPhdhY8H7O+cSpo7MF2/+KRaIpTENrQN
rmkXrNPRWHiIsdrkfRk5ho7FFjgrwgFuzDokbD+LjGFpX4deqFjnhSgu70geB1tkzqyfyybOFUUi
2Z6NIeI0J8wvSNWhLZ71PwruAna4mPbgpsORJyE+FGlq21NXKYsgmTNl9LPtqeZcN24i0ij8BOJ5
bj+wtlTDVE1dDm1BLKvswuIdyyzDT9EdtfVXXHMKQWGqPD3/5PbVmOzgAkfmAg8j97y0xi9jh7YA
PnCC24ZFa1WyEjdoAvrOajh3bq8+ZZgQQyfO/W63ZlkFnCbeypBjJq3O+yDhcmh2sdZE0kzxHBnU
EbnGnlXu28uFfiQKm0E6jR6tjUsHv58P0Q3+pUYez5WIcKmeG44fVPnxs16gc5/W41lMGzJoL/Nj
vX5fr3txFtVmcA+o2hXwdr9qONP1KQXAw2md/ofJmSZfaT8l1NL+D4nKGv4lEswybcJEyBGcmvEO
nNl/G6JVsDvV/82aeTD+uV6whPp8dkMIoZuYknu1gfy8/VQnVXNpBoEf16qQaNcE7p6IE2OV23XW
VsfptcOLJ4TBn2IXo0HnQHIDvlcrCy9JzPaYnZwqLdUe+QPrpvwjSoGeB++l3XFu5kPVD3ysi9jr
Pa0jdnyKRYi3SZql1pHCEsOxZEJAJ9MgfY3+jujyD4xofhi653DjIhKlt8j9qzcTjuyZl3K6KX5q
lInjUdWn+udCfRXGKQRwtyxEOJhnqNTRa8Et/wHP5wMj2CnwtX+l4SL99vfriGis/B5l1Ty+o3MD
TNbzyd/b6W/oDEnZIdTTxcWgcsGQjwCgPVyL3OkGFxixvn3R/lCjnuamVHowhgt9aOmej4EQKrkB
L4Fr34WN4u2zr1GK/6uZTjnjwhk/gAm4jVmpLkmNzwGjnKdq3ZzJX5ySFnXpnXDxOhn70oKjt0kN
tDIvREpdnpjXMUoutbZXoBkaOkDfodsiO7sgvI6s3bIa1H5W1GB34D09u93GhNie2pLCtBtf5EFb
gzwjczviGSrvNKPJoxjWyZM+cdqbH5Wr6X7uea0z2pn4FnOlVnhEAgT4zeYFLT/BKqJXGSRQ8j9/
3gZ4KMCGjknsg0l45PcBZWUE7OtqyIX36gAdTJS8xhNMlqnCONFFOFZlcpgPudrgnYx5MPsSbKbn
cSGPzZZouS3PTE5YfGjYWdD2V1ZK8xmlPK79ykgf53wL109wZJvPTYuQ5GoE3fhPIL+LQkXgkABH
UTJ4cad7zx4z35jnew70bFhm8RO2YX6iaOZlfP2uiIfXYVQqMJALJHZx5Xbr8ieaLtUEltKlHPxM
s1lepmL0mKRqTM9XJompW+hhzuHF1Fz6s0cJWv6o6/wqzZ79OwALhGqcijiZZo+q8QM3vVah2BHx
N0eeE6WTeCqbX8LYnguDbh38x3yw3lhJ2tjaR5i/07Y50oN2wF97tkqPE0NME4Fau9vHMHP0BS6w
gKEFYtrBX+Xfns2nnJbnOcLzaZ3UxNd80uFfWbesLcnOO4wBgPOsmIpdl1erT41xyX6gI4gdsWDd
KpjBldmA1nBI6+QDiJGC6obznxQ/VSiqBvyrl6j0pLk25SNCMjNb39MvHEGYNHGkHGjZpXHNkP/2
PRXZTU970k4ip33EX2nB4Lv/kfrGjRzdT3ADTijDi4Sm60ZGWBculOvsurcIwb0rnXu2XNGmZ68T
nEtiUt7cgyFl+XVmg7esB5gaTeHya040JdhUYT0B4VQ0fdr3F48apHTT6WYwU9d/DNwVha5CS5e4
9oSjNZrb+/hSdW4ap3UPAprJifaliRzhy7oqlQ2hwwq8Bs9V9dxGFekA5d0gxCu6Nh636E2K44ty
+YVziQaTUNjSUDA2YLnJNXNo+heGIlYffybAnGEeB3h8z39W5tTqbYdYfZw1Ocf6yGaOCkNLcwtA
hZ959Z2onz5m47c7DWwX0277uD280ybuSfiB6vggYQg4WDRdZYPIGR2uUT1fdKg/CjnqP5qCiIS+
PePBAGFKwGlh4475tN0t6DjtEWZ508Mlj3JCE0tjLQWuucRxt/H8nyvuf2pDdF72yE5ERzfnfpOp
g2Zu8TqF+Nh6dyXh1fr8OKXPYuOFSIikK6WdT+FmdEQsVJOdz02nT5zDHhIB/1MJlzZfSwWFba/H
/FzQhvC4U9c723pmCZWQ441rxYR7EhmpoFjT0zCLAtUt+4NIdca+7Impqikp1pDmDPycvAsKLgLw
yRywpZDcBLqp
`protect end_protected
