`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZT7+RCzMGpoBYSuObDu7GHIWP4wbG2z0+NZPy5ctMvSzcpDtYTeVa9Rt2jwWGft47o5EJP3ckUaz
ga/PA8jA7w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nez6Bl347nb6+rwYEAGUgNCAGAzNmFU5MeAC9+3K2UzYt8qxPFrJ/SFJLhvmq05ak2WdPG0DC6DY
KQm2he2dsLt5QsRiFYmj2xAL1KdqCGiHsVFY+u/PuU8GEcfn2GTMt2pBI+06udHlKRy3Gt2+icT+
Rzwp56VKG96Z/MuGTf4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bJ23shOZkE3PVggRHLeGJ2PbG8xrPMkBPZCJ8ZYfdCaWhZ4ZYd1C1zb43X+ojqULL2oHyUgAMgSj
ecIJtiACC+HQhYS9ZAedcNObDtyg4oslk+vfdk+TM2FZF2Etrw/yAEbq1f/PH0Kn+mbNEo33Zwe5
Rm8FZ1wDWOyOXh016tcp0RwCvdj2XR1Kw/zAigz9XUFsy0aJtcUXIJIlKcvvsjSATgFtlJhxEDo0
pnsWRjWP0UYdXkfmSQNXFz8qVRQRGSAtue/7tEuKBK7i+2io/Fn8ReAkkGJiWskeE9nOr9dx+4DE
9tfPWFjj0ZgyCy6JPKhTrEZyje87nH/0x9mcFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dilSTjuujT5h2DrLDbS/v0rUBHgSqc1odhqH2k0dTfIZcb7N2jGBdTrXFekiehlmoGDjU9sGGdlh
yFg/bT9j8pTdVb3lIkuOyMiLP0CoFYVl1z2IegKN7b9yFR+7EZbxn0N/B1ycLjS4ssnQq+SGbWl2
k2N7LLrQtkLu5td7xjU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pVPXt9t5C8qS/9IP6M6Y37REfDMW0SGfG45oP1DNSuCggimX25Htte0JNMgNJo8ar+6qTjWsopD4
IXOQzxTzbzczkdAIs6+pl9RpNOeJpa0bvybm+uwfWb8+Rcnz3NLflVxnmjLM1ayKKYARNVh7gQb9
C4SQt1FdooQ2JWlTXbp3V2aZpvw5F49u06L9Z5ayEEDdOQE/HQgnVfIryQKYB8stQTSh++L7A6Hi
fnnwsPjJQ2SynIHMSopYLmrhF02KU9HJ3WVKZ+nUrhCKV9djJvyWE9gZFn3X/nfyIkmo23lpYTgC
rYvCI0W4K/uiiwV05xGsCFhMYz37LiZv5/YMUw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4016)
`protect data_block
6Wo5rjfCVuPcU2g0iGcqP9tvT8tu0bB2joNIAOyeYj7XhN9i3gnhamfxv0DpYtwkP51HLRtLcsSX
ILx9f6y/6E1soWPaenpfUF8Elhc6vIelGxvGb5wfpvwx+Q2/Yt7L3tLerLAqWAvcyjL8wuiPP+Dm
6g1PmsO44zatHkhb8wUiIrWFqZatHA7yD8ynK9s4w+Y1bVgD7UI4ZsmPpnrtWc48Lpify74Rb1ke
The1G4ZPU4rsUFD6LefSHhsfu8wNDmMilPhnQoYIJ1uqdtk/KP0n2xa2TFMC9jhEGhPCQKvbIDS0
Lx2an9qEHrbTN3O+3Ao2/WXABJ1CkOfaksrrs3P3TyUUkMa958JAfvPwgr+4cDcCcIa/jlWLJFas
9eDbmG9IQE6UWYk0fMF/Iw3f0HFKVs74SPHR+0IXOTGoTTN4Xge1qD/G/75WFbxxeCq3nqJQXkhb
eh0raNjcMvfi6HacS3SCdQdGG8XgCHXtXKREW9N9yLpjQgkvYVaMlY2rYCD1lMITAvRNkhXmimMr
n9jFLRjbZEGSNoVAUEaL93RqCphJBlIScELR51MJHoWZw/MgoHvrJGvHMxMcc7DcdHtgpmIM9m+x
bjd/6uAsRrloWWeJOR+FsGiAyYI5i0K4TObv49NU8mkWKGIeCw1f5hHF0Zh8yCxPqRnNQ9J1Ns4P
hVnXwqmrHkuiFZz4P8UULY5tTwdChi25f//cFcNfrGqO/yNJsAqizy/rWgdNSI5AL6U3vVK8bK78
ykFnqmgE9Q9SFAfbfkB2J58n2E9nPUrPvgtNPEb991PZ0s+4Z3RIZZJ7ihXwBRnkMJRHmx2DWoY6
3Vs88TYoJtzKRUUd0FKnipBsYZzvHFSe/yKEUYwnw4mV1UisVw8qZ4vuyg/L38CSu/v8b5ndUYYR
ikygo4k7m3Y/PkJpz1B+zVSwyxFWu3hELvcWBD2sAXF0YsVLbp8kwach/tSGcE4ZC36Mb1MkjoiG
rkmjgrWfbPFmpPNnYjA4fL7dnFkOmMCJ7xn1jrsvwk8/2/xcw99VypFSXzy7hWEM7wTndPs2AwB+
emGXLPMcbjGISs5ZJf7wc/x9tI/HmHc95/qY8foqfNIxooF3jxMK5xlLoiwR01UD02HzBYidCXlA
CLhK4ZqRbIP7/GGORmawMvlWC/+GRo5fiJChNnEYbd/8yKpHD5ifzZTgdI0ROpnxDJnSOEJ/JZpx
ypOGn3OFHd2l615AYapfVp77rDDucoJOkSEN3Lzw82xhq79SsGzXSzzKH7IwPs/ozy458iEDicKh
IN0800aFvt2dl1umRfkDDLGo36/4pXZLJXnS42PM9KOrPOlwY64o5p4ggeaWEFlz1ZIHpiFDO6t/
bWkqkdGpe8UG3xBE+jY9/ce5jZacn+4Xx8foGhiaqL3YfiuJcr1sbyUSx+aCN3gD+4UN9iPwKbKj
VdLlWFJgr258+OhLG1eis3HybVY9yRueYrNxvfnuetpRVrQSFLXSa4GUs9Uws/fvYfUKRY/YrdfE
PV49jyIwnfIGmVg05pgFe+fvYhtuQpwLkvv5RJrV//Vg8FdcGnzCBirLdntmnooKbO66BIFIH0cw
s8ihj9SRUYP+jGljycY20vRPKzNTPlu67F9u1gwfIVBjYhXkGYsA8Q2JGKzJdHCbJmW7hhhfRClI
9+1SAs4Rg5ewQg++fp6l+0lxNX967MR03wgB/9/SpNKGZILR42J6qokqj0vOEoqBWD/AnpAVt8Ox
OiY/SWvUecIVf0Vti3iu4m2quCgWYPQg0hJwHcStjppOiPrsA6XoOQmc1KvrDjfJykV6QOoJb6ib
W5Hx02okqmnogyp0mNHndHVd5kztXOH98jN6jaWqajk96T/qEa27bXPfSsxhoCbLoFDAFzbQrVzm
9QpTDV/Hx6fK8OUhpzJene4xqhAYtM2tFHoi9hDLxiLBs01c55drhzxsJCjPYHqEzpXlPdsJc6d6
+vNtzEDO/p2dSRX+Q6Xswnvp8giqpOkwb6ifh0/l1bBRZOgzvXLOFp7CMNoqcOUBvD2Y8HTaYWFQ
rPtuOyOPB39FcrE19mmWNxTCJWznyhai40pl9bSLB50ilpTge31TrBmp8FKNqOh+/9EwMhDUDEP1
V9+DCLYLSRamFboIGg28Da1Z5+Pt03YJ08yXqqqXtoOHsBe0t9U6BrwwU6QTll0ORRbPNBPD0Bd7
2Cnt0xCk6JOCVSmv3GSREfrFjzK2k0ea2weTqG9nsDg2VnlL88upUNGhqrTIzH6N8RZzG8dDZKqT
yaDWXE7KdKvLOXBP0gwSjMzpSSpTupKdAtH0XGSopAlo6O2TNmtwcgn3PuSRvfmWP4nu88H6weOY
MurGmfFaJa9uOwOYkEJ5WL0ERUVrqnq0nYsylAsSBrh+nM+IUF6NI9x4s+yQf6XVcZwGN21qA7sq
14FbxOh3vFzxAMdctirP84z38MYNounjcl6KxpQshESRvYXO4eAjNEo6tASVGnwoDN3l/Rrb/lgU
2UOKEr1huVyx4hKjctl0/gl870+crOJewWHFa8W0KYNv5stLTFOZzUJ+huwQSq2L7auP240N4yZm
UOkisqu3PWwDpLLq7gxZ+K2iRoFbO6z2jx5c0eRWTqmntcJgd6UuZ2AAwlNRubIu+m9F1DG1cYt5
TFGnskVP9fVE8m66adkJd61y7X0wZnU7IXUY+FjxWEVXF+Jd0o19udQeU7X4dRvUzU7p1YRwSLhN
5tu0uN+Vt5PuNS9S24O7BdohbenGEjewjf0/mbNoxZbVyTy68FvV6wVenMQoYfvVQGeso+hUJ8z7
cgyiHTZWEnwOzCHpRDLtMrVi/9MiseRXNgGyk3jk4UmvW70ZmAS0YjxBskkz/Bf8XlP/bNKSQpDa
uBUdsuievjzE0ZEKJ74f6EaJ1iQBg6+DnvtBQB4RZchtrpNLm7Fegg3qeXY6dMysgnTIuXmI4YVU
cj9R1eSb2vNXPPT1Lyasxzao086XKRQ96ejDmv6ePiQaDYefzwV6MfPreNgPQrltaloQa4yjuoPW
7vUdlJetlwcDsv9NnMw9FoXjPLB6XMjKn2YTiZn1cdHbjp3masuKXPwqG35zc3lKJlLw4h0nwmRr
RGOgytpbyHWLpbzYRHprcvqqx2pxWwg/BHvzborJooZgIbs7/OC1VniQMMnf+STcldBo9DIxwIZ2
ZR0IX3tJEHGoIoYzw+OHIna5TdzpU8EhRWUR3PMUDR9A15edg7ZYUhA71elxT0bYuIOBVM9ettgT
0GyATB8mPD5qGPQ8uUml2EZuMD62/5WaGBB+XKrFAc9Pob/0GbW4HbftVtF0O8WaUiIfyqKpqgDR
nOtyi2kmNm0chc0NPvq/ULTqeQsxfgHERzwTXh8dQ5MP/8/cXUbEzy+gwxeN6J5ucpcGUpJUSbXU
wVYO6EzplcydNwsBWt62KOWhjNejqK5siCP/PLFD5FRRbUpIoEAggAvsW2UNaI5iICzLXpL0GduY
5H+DHCvw9668DfyVvPiiZ7Cd7xvD98+ewJZZhsPs1qP+rrMsZmpApq1wIHNnE8abfUq8RBeNVuI5
xyPhzr9Vdkn9pzyJBMbWPHmvrCLpITGSCnsBuOoH3EKJHa7WP/NqaKe6NSVRiZh32dJYN1dspIO6
NBMN++b+lJK0+dWumzNpSmJBUldj4c3UJEqcFeCLmjv3NLLw1wU3QMZ503yEerD8xWbpENPSrUeU
UNO6KJkw5lLJrxSphgyNI0hf9V17n9+sNX6gxmwZhFtnCUeEVg07YnUcg/GrdUuOWh1B/E/6QGlf
fCn88TWYQOrQvy8vwEhqH7A4a/Avg+cHvP+wndHEvKLR5yt2408o20a6TAn45Da33k0Tr0U3XmQ4
DWjJ+9QrNDgE7xV8BM9hWfcO6WAb2IR58dn1Xy6fWzDvMNWsx5miVYD19XbkugNKMmHtn1uOS3UK
hP2Co6MHoFFP5ED0l/1XHxYHQ9bKEEwYNYTU1bJSkFIjrFQEDLxqI50HtfnTM5tgrTMWPGbM3D5G
kP7XrTlBA7/c5BdZnk89DMcXM5dIWrr/mMjYJ/l9XVXpwrKSjs+xmJHt1zrKJPoB0SLQFqYcECfY
q0jGqw83PsmDYkeXdSC4npUVzxMswz81Diw3JFz+nrFQYYbQHQecsxpaQtWzOWRhGJ2KmhvvJ/SJ
xaXy2XvdKVAE+mZXRIk9vmUFBaULcj7Th98Te85xCiDBrDPPHNkDlPWCVW6vyagWuye4wlrVTPbt
Tuqq7KHolYkZQWqtIYPkooanML5h6IRg/J2oz1ughg65JduYhbBYLjaaYJd5K6SMKStMTHdWCXr0
Zbb4i+71VVral70iVEPnThkP130Lo24QptN7qQym+btP0r/F3i7RBn2sTJOTjQeh6izFqB2rCgyo
Z+LY4HB6aYEUH6YVWPRFHE1ZOrQ5vOFi4u8/GTIWXTu09MRXluh3y1B40zxqPToMuZ3XIchGI1sm
X/PP0OfIcEIMaP2fB9iNTfoYCJ9VVX8oxY/Cu7NRVEMi3Lou5LLw4ISKu2TcJKv4PdJaucOzzgbY
qh8l5vcAlxgGzbIYkwqUGkXSaUJI5ofZhHzdJBcAN3MiH3nox+rjyxfAIYks27Rk+tk2koFlZnr3
cOe4ZsNsXBHqFSUAE0MNSX5rtC34+axxc+uXRsgBaEhW94GGHIR5qb0KeRp+SO7kBfQBwQKp5WPd
cbgyS+3/+rVBNtYzYTTcyruM8SQZKHE6OdszL+4/BUvvpps7U6CVTHLt4Nbg4H5qRvXpnfhYffa8
Z0Fxs83L+e3x323yh/XD4RCvOyFSrLEKWfvbJwV5NZyto+bs3Cv+lPv3HW4XST535b/oNTixANB5
+KWD+Jyn/8OHHgVormjYCJELa2IIteZ1ZMFxQVvbyMiyJZbCitKms5azjK9YWl6p8qAEKTBlfR/X
bGJzcKCMzK2VmuO0RGGeQZferKp9WQlQ4TQWbF+BpYDXtgEbyP0yNi2laiaiNgNItOgdxW0/tBGB
DAYUcgyu8XLKTrNC70lh/KWEwwhWWL64/mnkAtCw7yLR9D3ElDDJEPqqg8/oPtsP0UEdQs4Sm2Z5
l+01AuxtdcikfQo2BEFGrf7t0+/LS7ofhMXXfNXFPPwof0v5oazNTSLuATijfIO+LKzvjo8k7ddH
MEeqd06Wh06VuFTWabH98mJM/0Bj5vig3gyXPoc9f7wpEO8QLk62m7HfSjGSFwZwqiDxPaVeiL+5
8n7IB8bCi36leTL6kVrd9g/EK7RV9H7fzOSmG+2vWWEvnxnQMaNhIpabtfqmr3E6IjFfEQAWN9nt
DxgHhXY2vc/cLag/HjUoplng6m261RMgtng=
`protect end_protected
